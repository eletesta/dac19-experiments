// Benchmark "mapping" written by ABC on Mon Nov 19 13:13:48 2018

module mapping ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128;
  wire n387, n389, n390, n391, n393, n394, n395, n396, n398, n399, n400,
    n401, n403, n404, n405, n407, n408, n409, n410, n411, n412, n413, n414,
    n416, n417, n418, n420, n421, n422, n423, n424, n425, n426, n427, n429,
    n430, n431, n433, n434, n435, n436, n437, n438, n439, n440, n442, n443,
    n444, n446, n447, n448, n449, n450, n451, n452, n454, n455, n456, n458,
    n459, n460, n461, n462, n463, n464, n465, n467, n468, n469, n471, n472,
    n473, n474, n475, n476, n477, n478, n480, n481, n482, n484, n485, n486,
    n487, n488, n489, n490, n491, n493, n494, n495, n497, n498, n499, n500,
    n501, n502, n503, n504, n506, n507, n508, n510, n511, n512, n513, n514,
    n515, n516, n518, n519, n520, n522, n523, n524, n525, n526, n527, n528,
    n529, n531, n532, n533, n535, n536, n537, n538, n539, n540, n541, n542,
    n544, n545, n546, n548, n549, n550, n551, n552, n553, n554, n555, n557,
    n558, n559, n561, n562, n563, n564, n565, n566, n567, n568, n570, n571,
    n572, n574, n575, n576, n577, n578, n579, n580, n582, n583, n584, n586,
    n587, n588, n589, n590, n591, n592, n593, n595, n596, n597, n599, n600,
    n601, n602, n603, n604, n605, n606, n608, n609, n610, n612, n613, n614,
    n615, n616, n617, n618, n619, n621, n622, n623, n625, n626, n627, n628,
    n629, n630, n631, n632, n634, n635, n636, n638, n639, n640, n641, n642,
    n643, n644, n646, n647, n648, n650, n651, n652, n653, n654, n655, n656,
    n657, n659, n660, n661, n663, n664, n665, n666, n667, n668, n669, n670,
    n672, n673, n674, n676, n677, n678, n679, n680, n681, n682, n683, n685,
    n686, n687, n689, n690, n691, n692, n693, n694, n695, n696, n698, n699,
    n700, n702, n703, n704, n705, n706, n707, n708, n710, n711, n712, n714,
    n715, n716, n717, n718, n719, n720, n721, n723, n724, n725, n727, n728,
    n729, n730, n731, n732, n733, n734, n736, n737, n738, n740, n741, n742,
    n743, n744, n745, n746, n747, n749, n750, n751, n753, n754, n755, n756,
    n757, n758, n759, n760, n762, n763, n764, n766, n767, n768, n769, n770,
    n771, n772, n774, n775, n776, n778, n779, n780, n781, n782, n783, n784,
    n785, n787, n788, n789, n791, n792, n793, n794, n795, n796, n797, n798,
    n800, n801, n802, n804, n805, n806, n807, n808, n809, n810, n811, n813,
    n814, n815, n817, n818, n819, n820, n821, n822, n823, n824, n826, n827,
    n828, n830, n831, n832, n833, n834, n835, n836, n838, n839, n840, n842,
    n843, n844, n845, n846, n847, n848, n849, n851, n852, n853, n855, n856,
    n857, n858, n859, n860, n861, n862, n864, n865, n866, n868, n869, n870,
    n871, n872, n873, n874, n875, n877, n878, n879, n881, n882, n883, n884,
    n885, n886, n887, n888, n890, n891, n892, n894, n895, n896, n897, n898,
    n899, n900, n902, n903, n904, n906, n907, n908, n909, n910, n911, n912,
    n913, n915, n916, n917, n919, n920, n921, n922, n923, n924, n925, n926,
    n928, n929, n930, n932, n933, n934, n935, n936, n937, n938, n939, n941,
    n942, n943, n945, n946, n947, n948, n949, n950, n951, n952, n954, n955,
    n956, n958, n959, n960, n961, n962, n963, n964, n966, n967, n968, n970,
    n971, n972, n973, n974, n975, n976, n978, n979, n980, n981, n983, n984,
    n985, n986, n987, n989, n990, n991, n992, n994, n995, n996, n997, n998,
    n1000, n1001, n1002, n1003, n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1014, n1015, n1016, n1017, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1028, n1029, n1030, n1031, n1033, n1034,
    n1035, n1036, n1037, n1038, n1039, n1040, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1050, n1051, n1052, n1053, n1055, n1056, n1057,
    n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1076, n1077, n1078, n1080, n1081,
    n1082, n1083, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
    n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1102, n1103, n1104,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1114, n1115, n1116,
    n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1126, n1127, n1128,
    n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1138, n1139, n1140,
    n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1150, n1151, n1152,
    n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1162, n1163, n1164,
    n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1174, n1175, n1176,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1186, n1187, n1188,
    n1190;
  assign n387 = pi000 & pi128;
  assign po000 = ~pi000 ^ ~pi128;
  assign n389 = ~pi001 & ~pi129;
  assign n390 = pi001 ^ ~pi129;
  assign n391 = ~n387 & ~n390;
  assign po001 = n387 ^ ~n390;
  assign n393 = ~n391 & ~n389;
  assign n394 = ~pi002 & ~pi130;
  assign n395 = pi002 ^ ~pi130;
  assign n396 = ~n393 & ~n395;
  assign po002 = n393 ^ ~n395;
  assign n398 = ~n396 & ~n394;
  assign n399 = pi003 & pi131;
  assign n400 = pi003 ^ ~pi131;
  assign n401 = n398 & ~n400;
  assign po003 = ~n398 ^ n400;
  assign n403 = ~n401 & ~n399;
  assign n404 = ~pi004 & ~pi132;
  assign n405 = pi004 ^ ~pi132;
  assign po004 = ~n403 ^ ~n405;
  assign n407 = ~n400 & ~n405;
  assign n408 = n398 & n407;
  assign n409 = ~n399 & ~n405;
  assign n410 = ~n409 & ~n404;
  assign n411 = ~n408 & ~n410;
  assign n412 = pi005 & pi133;
  assign n413 = pi005 ^ ~pi133;
  assign n414 = ~n411 & ~n413;
  assign po005 = ~n411 ^ ~n413;
  assign n416 = ~n414 & ~n412;
  assign n417 = ~pi006 & ~pi134;
  assign n418 = pi006 ^ ~pi134;
  assign po006 = ~n416 ^ ~n418;
  assign n420 = ~n413 & ~n418;
  assign n421 = ~n411 & n420;
  assign n422 = ~n412 & ~n418;
  assign n423 = ~n422 & ~n417;
  assign n424 = ~n421 & ~n423;
  assign n425 = pi007 & pi135;
  assign n426 = pi007 ^ ~pi135;
  assign n427 = ~n424 & ~n426;
  assign po007 = ~n424 ^ ~n426;
  assign n429 = ~n427 & ~n425;
  assign n430 = ~pi008 & ~pi136;
  assign n431 = pi008 ^ ~pi136;
  assign po008 = ~n429 ^ ~n431;
  assign n433 = ~n426 & ~n431;
  assign n434 = ~n424 & n433;
  assign n435 = ~n425 & ~n431;
  assign n436 = ~n435 & ~n430;
  assign n437 = ~n434 & ~n436;
  assign n438 = pi009 & pi137;
  assign n439 = pi009 ^ ~pi137;
  assign n440 = ~n437 & ~n439;
  assign po009 = ~n437 ^ ~n439;
  assign n442 = ~n440 & ~n438;
  assign n443 = ~pi010 & ~pi138;
  assign n444 = pi010 ^ ~pi138;
  assign po010 = ~n442 ^ ~n444;
  assign n446 = n440 & ~n444;
  assign n447 = ~n438 & ~n444;
  assign n448 = ~n447 & ~n443;
  assign n449 = ~n446 & ~n448;
  assign n450 = pi011 & pi139;
  assign n451 = pi011 ^ ~pi139;
  assign n452 = ~n449 & ~n451;
  assign po011 = ~n449 ^ ~n451;
  assign n454 = ~n452 & ~n450;
  assign n455 = ~pi012 & ~pi140;
  assign n456 = pi012 ^ ~pi140;
  assign po012 = n454 ^ n456;
  assign n458 = ~n451 & ~n456;
  assign n459 = ~n449 & n458;
  assign n460 = ~n450 & ~n456;
  assign n461 = ~n460 & ~n455;
  assign n462 = ~n459 & ~n461;
  assign n463 = pi013 & pi141;
  assign n464 = pi013 ^ ~pi141;
  assign n465 = ~n462 & ~n464;
  assign po013 = ~n462 ^ ~n464;
  assign n467 = ~n465 & ~n463;
  assign n468 = ~pi014 & ~pi142;
  assign n469 = pi014 ^ ~pi142;
  assign po014 = ~n467 ^ ~n469;
  assign n471 = ~n464 & ~n469;
  assign n472 = ~n462 & n471;
  assign n473 = ~n463 & ~n469;
  assign n474 = ~n473 & ~n468;
  assign n475 = ~n472 & ~n474;
  assign n476 = pi015 & pi143;
  assign n477 = pi015 ^ ~pi143;
  assign n478 = ~n475 & ~n477;
  assign po015 = ~n475 ^ ~n477;
  assign n480 = ~n478 & ~n476;
  assign n481 = ~pi016 & ~pi144;
  assign n482 = pi016 ^ ~pi144;
  assign po016 = ~n480 ^ ~n482;
  assign n484 = ~n477 & ~n482;
  assign n485 = ~n475 & n484;
  assign n486 = ~n476 & ~n482;
  assign n487 = ~n486 & ~n481;
  assign n488 = ~n485 & ~n487;
  assign n489 = pi017 & pi145;
  assign n490 = pi017 ^ ~pi145;
  assign n491 = ~n488 & ~n490;
  assign po017 = ~n488 ^ ~n490;
  assign n493 = ~n491 & ~n489;
  assign n494 = ~pi018 & ~pi146;
  assign n495 = pi018 ^ ~pi146;
  assign po018 = ~n493 ^ ~n495;
  assign n497 = ~n490 & ~n495;
  assign n498 = ~n488 & n497;
  assign n499 = ~n489 & ~n495;
  assign n500 = ~n499 & ~n494;
  assign n501 = ~n498 & ~n500;
  assign n502 = pi019 & pi147;
  assign n503 = pi019 ^ ~pi147;
  assign n504 = ~n501 & ~n503;
  assign po019 = ~n501 ^ ~n503;
  assign n506 = ~n504 & ~n502;
  assign n507 = ~pi020 & ~pi148;
  assign n508 = pi020 ^ ~pi148;
  assign po020 = ~n506 ^ ~n508;
  assign n510 = n504 & ~n508;
  assign n511 = ~n502 & ~n508;
  assign n512 = ~n511 & ~n507;
  assign n513 = ~n510 & ~n512;
  assign n514 = pi021 & pi149;
  assign n515 = pi021 ^ ~pi149;
  assign n516 = ~n513 & ~n515;
  assign po021 = ~n513 ^ ~n515;
  assign n518 = ~n516 & ~n514;
  assign n519 = ~pi022 & ~pi150;
  assign n520 = pi022 ^ ~pi150;
  assign po022 = n518 ^ n520;
  assign n522 = ~n515 & ~n520;
  assign n523 = ~n513 & n522;
  assign n524 = ~n514 & ~n520;
  assign n525 = ~n524 & ~n519;
  assign n526 = ~n523 & ~n525;
  assign n527 = pi023 & pi151;
  assign n528 = pi023 ^ ~pi151;
  assign n529 = ~n526 & ~n528;
  assign po023 = ~n526 ^ ~n528;
  assign n531 = ~n529 & ~n527;
  assign n532 = ~pi024 & ~pi152;
  assign n533 = pi024 ^ ~pi152;
  assign po024 = ~n531 ^ ~n533;
  assign n535 = ~n528 & ~n533;
  assign n536 = ~n526 & n535;
  assign n537 = ~n527 & ~n533;
  assign n538 = ~n537 & ~n532;
  assign n539 = ~n536 & ~n538;
  assign n540 = pi025 & pi153;
  assign n541 = pi025 ^ ~pi153;
  assign n542 = ~n539 & ~n541;
  assign po025 = ~n539 ^ ~n541;
  assign n544 = ~n542 & ~n540;
  assign n545 = ~pi026 & ~pi154;
  assign n546 = pi026 ^ ~pi154;
  assign po026 = ~n544 ^ ~n546;
  assign n548 = ~n541 & ~n546;
  assign n549 = ~n539 & n548;
  assign n550 = ~n540 & ~n546;
  assign n551 = ~n550 & ~n545;
  assign n552 = ~n549 & ~n551;
  assign n553 = pi027 & pi155;
  assign n554 = pi027 ^ ~pi155;
  assign n555 = ~n552 & ~n554;
  assign po027 = ~n552 ^ ~n554;
  assign n557 = ~n555 & ~n553;
  assign n558 = ~pi028 & ~pi156;
  assign n559 = pi028 ^ ~pi156;
  assign po028 = ~n557 ^ ~n559;
  assign n561 = ~n554 & ~n559;
  assign n562 = ~n552 & n561;
  assign n563 = ~n553 & ~n559;
  assign n564 = ~n563 & ~n558;
  assign n565 = ~n562 & ~n564;
  assign n566 = pi029 & pi157;
  assign n567 = pi029 ^ ~pi157;
  assign n568 = ~n565 & ~n567;
  assign po029 = ~n565 ^ ~n567;
  assign n570 = ~n568 & ~n566;
  assign n571 = ~pi030 & ~pi158;
  assign n572 = pi030 ^ ~pi158;
  assign po030 = ~n570 ^ ~n572;
  assign n574 = n568 & ~n572;
  assign n575 = ~n566 & ~n572;
  assign n576 = ~n575 & ~n571;
  assign n577 = ~n574 & ~n576;
  assign n578 = pi031 & pi159;
  assign n579 = pi031 ^ ~pi159;
  assign n580 = ~n577 & ~n579;
  assign po031 = ~n577 ^ ~n579;
  assign n582 = ~n580 & ~n578;
  assign n583 = ~pi032 & ~pi160;
  assign n584 = pi032 ^ ~pi160;
  assign po032 = n582 ^ n584;
  assign n586 = ~n579 & ~n584;
  assign n587 = ~n577 & n586;
  assign n588 = ~n578 & ~n584;
  assign n589 = ~n588 & ~n583;
  assign n590 = ~n587 & ~n589;
  assign n591 = pi033 & pi161;
  assign n592 = pi033 ^ ~pi161;
  assign n593 = ~n590 & ~n592;
  assign po033 = ~n590 ^ ~n592;
  assign n595 = ~n593 & ~n591;
  assign n596 = ~pi034 & ~pi162;
  assign n597 = pi034 ^ ~pi162;
  assign po034 = ~n595 ^ ~n597;
  assign n599 = ~n592 & ~n597;
  assign n600 = ~n590 & n599;
  assign n601 = ~n591 & ~n597;
  assign n602 = ~n601 & ~n596;
  assign n603 = ~n600 & ~n602;
  assign n604 = pi035 & pi163;
  assign n605 = pi035 ^ ~pi163;
  assign n606 = ~n603 & ~n605;
  assign po035 = ~n603 ^ ~n605;
  assign n608 = ~n606 & ~n604;
  assign n609 = ~pi036 & ~pi164;
  assign n610 = pi036 ^ ~pi164;
  assign po036 = ~n608 ^ ~n610;
  assign n612 = ~n605 & ~n610;
  assign n613 = ~n603 & n612;
  assign n614 = ~n604 & ~n610;
  assign n615 = ~n614 & ~n609;
  assign n616 = ~n613 & ~n615;
  assign n617 = pi037 & pi165;
  assign n618 = pi037 ^ ~pi165;
  assign n619 = ~n616 & ~n618;
  assign po037 = ~n616 ^ ~n618;
  assign n621 = ~n619 & ~n617;
  assign n622 = ~pi038 & ~pi166;
  assign n623 = pi038 ^ ~pi166;
  assign po038 = ~n621 ^ ~n623;
  assign n625 = ~n618 & ~n623;
  assign n626 = ~n616 & n625;
  assign n627 = ~n617 & ~n623;
  assign n628 = ~n627 & ~n622;
  assign n629 = ~n626 & ~n628;
  assign n630 = pi039 & pi167;
  assign n631 = pi039 ^ ~pi167;
  assign n632 = ~n629 & ~n631;
  assign po039 = ~n629 ^ ~n631;
  assign n634 = ~n632 & ~n630;
  assign n635 = ~pi040 & ~pi168;
  assign n636 = pi040 ^ ~pi168;
  assign po040 = ~n634 ^ ~n636;
  assign n638 = n632 & ~n636;
  assign n639 = ~n630 & ~n636;
  assign n640 = ~n639 & ~n635;
  assign n641 = ~n638 & ~n640;
  assign n642 = pi041 & pi169;
  assign n643 = pi041 ^ ~pi169;
  assign n644 = ~n641 & ~n643;
  assign po041 = ~n641 ^ ~n643;
  assign n646 = ~n644 & ~n642;
  assign n647 = ~pi042 & ~pi170;
  assign n648 = pi042 ^ ~pi170;
  assign po042 = n646 ^ n648;
  assign n650 = ~n643 & ~n648;
  assign n651 = ~n641 & n650;
  assign n652 = ~n642 & ~n648;
  assign n653 = ~n652 & ~n647;
  assign n654 = ~n651 & ~n653;
  assign n655 = pi043 & pi171;
  assign n656 = pi043 ^ ~pi171;
  assign n657 = ~n654 & ~n656;
  assign po043 = ~n654 ^ ~n656;
  assign n659 = ~n657 & ~n655;
  assign n660 = ~pi044 & ~pi172;
  assign n661 = pi044 ^ ~pi172;
  assign po044 = ~n659 ^ ~n661;
  assign n663 = ~n656 & ~n661;
  assign n664 = ~n654 & n663;
  assign n665 = ~n655 & ~n661;
  assign n666 = ~n665 & ~n660;
  assign n667 = ~n664 & ~n666;
  assign n668 = pi045 & pi173;
  assign n669 = pi045 ^ ~pi173;
  assign n670 = ~n667 & ~n669;
  assign po045 = ~n667 ^ ~n669;
  assign n672 = ~n670 & ~n668;
  assign n673 = ~pi046 & ~pi174;
  assign n674 = pi046 ^ ~pi174;
  assign po046 = ~n672 ^ ~n674;
  assign n676 = ~n669 & ~n674;
  assign n677 = ~n667 & n676;
  assign n678 = ~n668 & ~n674;
  assign n679 = ~n678 & ~n673;
  assign n680 = ~n677 & ~n679;
  assign n681 = pi047 & pi175;
  assign n682 = pi047 ^ ~pi175;
  assign n683 = ~n680 & ~n682;
  assign po047 = ~n680 ^ ~n682;
  assign n685 = ~n683 & ~n681;
  assign n686 = ~pi048 & ~pi176;
  assign n687 = pi048 ^ ~pi176;
  assign po048 = ~n685 ^ ~n687;
  assign n689 = ~n682 & ~n687;
  assign n690 = ~n680 & n689;
  assign n691 = ~n681 & ~n687;
  assign n692 = ~n691 & ~n686;
  assign n693 = ~n690 & ~n692;
  assign n694 = pi049 & pi177;
  assign n695 = pi049 ^ ~pi177;
  assign n696 = ~n693 & ~n695;
  assign po049 = ~n693 ^ ~n695;
  assign n698 = ~n696 & ~n694;
  assign n699 = ~pi050 & ~pi178;
  assign n700 = pi050 ^ ~pi178;
  assign po050 = ~n698 ^ ~n700;
  assign n702 = n696 & ~n700;
  assign n703 = ~n694 & ~n700;
  assign n704 = ~n703 & ~n699;
  assign n705 = ~n702 & ~n704;
  assign n706 = pi051 & pi179;
  assign n707 = pi051 ^ ~pi179;
  assign n708 = ~n705 & ~n707;
  assign po051 = ~n705 ^ ~n707;
  assign n710 = ~n708 & ~n706;
  assign n711 = ~pi052 & ~pi180;
  assign n712 = pi052 ^ ~pi180;
  assign po052 = n710 ^ n712;
  assign n714 = ~n707 & ~n712;
  assign n715 = ~n705 & n714;
  assign n716 = ~n706 & ~n712;
  assign n717 = ~n716 & ~n711;
  assign n718 = ~n715 & ~n717;
  assign n719 = pi053 & pi181;
  assign n720 = pi053 ^ ~pi181;
  assign n721 = ~n718 & ~n720;
  assign po053 = ~n718 ^ ~n720;
  assign n723 = ~n721 & ~n719;
  assign n724 = ~pi054 & ~pi182;
  assign n725 = pi054 ^ ~pi182;
  assign po054 = ~n723 ^ ~n725;
  assign n727 = ~n720 & ~n725;
  assign n728 = ~n718 & n727;
  assign n729 = ~n719 & ~n725;
  assign n730 = ~n729 & ~n724;
  assign n731 = ~n728 & ~n730;
  assign n732 = pi055 & pi183;
  assign n733 = pi055 ^ ~pi183;
  assign n734 = ~n731 & ~n733;
  assign po055 = ~n731 ^ ~n733;
  assign n736 = ~n734 & ~n732;
  assign n737 = ~pi056 & ~pi184;
  assign n738 = pi056 ^ ~pi184;
  assign po056 = ~n736 ^ ~n738;
  assign n740 = ~n733 & ~n738;
  assign n741 = ~n731 & n740;
  assign n742 = ~n732 & ~n738;
  assign n743 = ~n742 & ~n737;
  assign n744 = ~n741 & ~n743;
  assign n745 = pi057 & pi185;
  assign n746 = pi057 ^ ~pi185;
  assign n747 = ~n744 & ~n746;
  assign po057 = ~n744 ^ ~n746;
  assign n749 = ~n747 & ~n745;
  assign n750 = ~pi058 & ~pi186;
  assign n751 = pi058 ^ ~pi186;
  assign po058 = ~n749 ^ ~n751;
  assign n753 = ~n746 & ~n751;
  assign n754 = ~n744 & n753;
  assign n755 = ~n745 & ~n751;
  assign n756 = ~n755 & ~n750;
  assign n757 = ~n754 & ~n756;
  assign n758 = pi059 & pi187;
  assign n759 = pi059 ^ ~pi187;
  assign n760 = ~n757 & ~n759;
  assign po059 = ~n757 ^ ~n759;
  assign n762 = ~n760 & ~n758;
  assign n763 = ~pi060 & ~pi188;
  assign n764 = pi060 ^ ~pi188;
  assign po060 = ~n762 ^ ~n764;
  assign n766 = n760 & ~n764;
  assign n767 = ~n758 & ~n764;
  assign n768 = ~n767 & ~n763;
  assign n769 = ~n766 & ~n768;
  assign n770 = pi061 & pi189;
  assign n771 = pi061 ^ ~pi189;
  assign n772 = ~n769 & ~n771;
  assign po061 = ~n769 ^ ~n771;
  assign n774 = ~n772 & ~n770;
  assign n775 = ~pi062 & ~pi190;
  assign n776 = pi062 ^ ~pi190;
  assign po062 = n774 ^ n776;
  assign n778 = ~n771 & ~n776;
  assign n779 = ~n769 & n778;
  assign n780 = ~n770 & ~n776;
  assign n781 = ~n780 & ~n775;
  assign n782 = ~n779 & ~n781;
  assign n783 = pi063 & pi191;
  assign n784 = pi063 ^ ~pi191;
  assign n785 = ~n782 & ~n784;
  assign po063 = ~n782 ^ ~n784;
  assign n787 = ~n785 & ~n783;
  assign n788 = ~pi064 & ~pi192;
  assign n789 = pi064 ^ ~pi192;
  assign po064 = ~n787 ^ ~n789;
  assign n791 = ~n784 & ~n789;
  assign n792 = ~n782 & n791;
  assign n793 = ~n783 & ~n789;
  assign n794 = ~n793 & ~n788;
  assign n795 = ~n792 & ~n794;
  assign n796 = pi065 & pi193;
  assign n797 = pi065 ^ ~pi193;
  assign n798 = ~n795 & ~n797;
  assign po065 = ~n795 ^ ~n797;
  assign n800 = ~n798 & ~n796;
  assign n801 = ~pi066 & ~pi194;
  assign n802 = pi066 ^ ~pi194;
  assign po066 = ~n800 ^ ~n802;
  assign n804 = ~n797 & ~n802;
  assign n805 = ~n795 & n804;
  assign n806 = ~n796 & ~n802;
  assign n807 = ~n806 & ~n801;
  assign n808 = ~n805 & ~n807;
  assign n809 = pi067 & pi195;
  assign n810 = pi067 ^ ~pi195;
  assign n811 = ~n808 & ~n810;
  assign po067 = ~n808 ^ ~n810;
  assign n813 = ~n811 & ~n809;
  assign n814 = ~pi068 & ~pi196;
  assign n815 = pi068 ^ ~pi196;
  assign po068 = ~n813 ^ ~n815;
  assign n817 = ~n810 & ~n815;
  assign n818 = ~n808 & n817;
  assign n819 = ~n809 & ~n815;
  assign n820 = ~n819 & ~n814;
  assign n821 = ~n818 & ~n820;
  assign n822 = pi069 & pi197;
  assign n823 = pi069 ^ ~pi197;
  assign n824 = ~n821 & ~n823;
  assign po069 = ~n821 ^ ~n823;
  assign n826 = ~n824 & ~n822;
  assign n827 = ~pi070 & ~pi198;
  assign n828 = pi070 ^ ~pi198;
  assign po070 = ~n826 ^ ~n828;
  assign n830 = n824 & ~n828;
  assign n831 = ~n822 & ~n828;
  assign n832 = ~n831 & ~n827;
  assign n833 = ~n830 & ~n832;
  assign n834 = pi071 & pi199;
  assign n835 = pi071 ^ ~pi199;
  assign n836 = ~n833 & ~n835;
  assign po071 = ~n833 ^ ~n835;
  assign n838 = ~n836 & ~n834;
  assign n839 = ~pi072 & ~pi200;
  assign n840 = pi072 ^ ~pi200;
  assign po072 = n838 ^ n840;
  assign n842 = ~n835 & ~n840;
  assign n843 = ~n833 & n842;
  assign n844 = ~n834 & ~n840;
  assign n845 = ~n844 & ~n839;
  assign n846 = ~n843 & ~n845;
  assign n847 = pi073 & pi201;
  assign n848 = pi073 ^ ~pi201;
  assign n849 = ~n846 & ~n848;
  assign po073 = ~n846 ^ ~n848;
  assign n851 = ~n849 & ~n847;
  assign n852 = ~pi074 & ~pi202;
  assign n853 = pi074 ^ ~pi202;
  assign po074 = ~n851 ^ ~n853;
  assign n855 = ~n848 & ~n853;
  assign n856 = ~n846 & n855;
  assign n857 = ~n847 & ~n853;
  assign n858 = ~n857 & ~n852;
  assign n859 = ~n856 & ~n858;
  assign n860 = pi075 & pi203;
  assign n861 = pi075 ^ ~pi203;
  assign n862 = ~n859 & ~n861;
  assign po075 = ~n859 ^ ~n861;
  assign n864 = ~n862 & ~n860;
  assign n865 = ~pi076 & ~pi204;
  assign n866 = pi076 ^ ~pi204;
  assign po076 = ~n864 ^ ~n866;
  assign n868 = ~n861 & ~n866;
  assign n869 = ~n859 & n868;
  assign n870 = ~n860 & ~n866;
  assign n871 = ~n870 & ~n865;
  assign n872 = ~n869 & ~n871;
  assign n873 = pi077 & pi205;
  assign n874 = pi077 ^ ~pi205;
  assign n875 = ~n872 & ~n874;
  assign po077 = ~n872 ^ ~n874;
  assign n877 = ~n875 & ~n873;
  assign n878 = ~pi078 & ~pi206;
  assign n879 = pi078 ^ ~pi206;
  assign po078 = ~n877 ^ ~n879;
  assign n881 = ~n874 & ~n879;
  assign n882 = ~n872 & n881;
  assign n883 = ~n873 & ~n879;
  assign n884 = ~n883 & ~n878;
  assign n885 = ~n882 & ~n884;
  assign n886 = pi079 & pi207;
  assign n887 = pi079 ^ ~pi207;
  assign n888 = ~n885 & ~n887;
  assign po079 = ~n885 ^ ~n887;
  assign n890 = ~n888 & ~n886;
  assign n891 = ~pi080 & ~pi208;
  assign n892 = pi080 ^ ~pi208;
  assign po080 = ~n890 ^ ~n892;
  assign n894 = n888 & ~n892;
  assign n895 = ~n886 & ~n892;
  assign n896 = ~n895 & ~n891;
  assign n897 = ~n894 & ~n896;
  assign n898 = pi081 & pi209;
  assign n899 = pi081 ^ ~pi209;
  assign n900 = ~n897 & ~n899;
  assign po081 = ~n897 ^ ~n899;
  assign n902 = ~n900 & ~n898;
  assign n903 = ~pi082 & ~pi210;
  assign n904 = pi082 ^ ~pi210;
  assign po082 = n902 ^ n904;
  assign n906 = ~n899 & ~n904;
  assign n907 = ~n897 & n906;
  assign n908 = ~n898 & ~n904;
  assign n909 = ~n908 & ~n903;
  assign n910 = ~n907 & ~n909;
  assign n911 = pi083 & pi211;
  assign n912 = pi083 ^ ~pi211;
  assign n913 = ~n910 & ~n912;
  assign po083 = ~n910 ^ ~n912;
  assign n915 = ~n913 & ~n911;
  assign n916 = ~pi084 & ~pi212;
  assign n917 = pi084 ^ ~pi212;
  assign po084 = ~n915 ^ ~n917;
  assign n919 = ~n912 & ~n917;
  assign n920 = ~n910 & n919;
  assign n921 = ~n911 & ~n917;
  assign n922 = ~n921 & ~n916;
  assign n923 = ~n920 & ~n922;
  assign n924 = pi085 & pi213;
  assign n925 = pi085 ^ ~pi213;
  assign n926 = ~n923 & ~n925;
  assign po085 = ~n923 ^ ~n925;
  assign n928 = ~n926 & ~n924;
  assign n929 = ~pi086 & ~pi214;
  assign n930 = pi086 ^ ~pi214;
  assign po086 = ~n928 ^ ~n930;
  assign n932 = ~n925 & ~n930;
  assign n933 = ~n923 & n932;
  assign n934 = ~n924 & ~n930;
  assign n935 = ~n934 & ~n929;
  assign n936 = ~n933 & ~n935;
  assign n937 = pi087 & pi215;
  assign n938 = pi087 ^ ~pi215;
  assign n939 = ~n936 & ~n938;
  assign po087 = ~n936 ^ ~n938;
  assign n941 = ~n939 & ~n937;
  assign n942 = ~pi088 & ~pi216;
  assign n943 = pi088 ^ ~pi216;
  assign po088 = ~n941 ^ ~n943;
  assign n945 = ~n938 & ~n943;
  assign n946 = ~n936 & n945;
  assign n947 = ~n937 & ~n943;
  assign n948 = ~n947 & ~n942;
  assign n949 = ~n946 & ~n948;
  assign n950 = pi089 & pi217;
  assign n951 = pi089 ^ ~pi217;
  assign n952 = ~n949 & ~n951;
  assign po089 = ~n949 ^ ~n951;
  assign n954 = ~n952 & ~n950;
  assign n955 = ~pi090 & ~pi218;
  assign n956 = pi090 ^ ~pi218;
  assign po090 = ~n954 ^ ~n956;
  assign n958 = n952 & ~n956;
  assign n959 = ~n950 & ~n956;
  assign n960 = ~n959 & ~n955;
  assign n961 = ~n958 & ~n960;
  assign n962 = pi091 & pi219;
  assign n963 = pi091 ^ ~pi219;
  assign n964 = ~n961 & ~n963;
  assign po091 = ~n961 ^ ~n963;
  assign n966 = ~n964 & ~n962;
  assign n967 = ~pi092 & ~pi220;
  assign n968 = pi092 ^ ~pi220;
  assign po092 = ~n966 ^ ~n968;
  assign n970 = n964 & ~n968;
  assign n971 = ~n962 & ~n968;
  assign n972 = ~n971 & ~n967;
  assign n973 = ~n970 & ~n972;
  assign n974 = pi093 & pi221;
  assign n975 = pi093 ^ ~pi221;
  assign n976 = ~n973 & ~n975;
  assign po093 = ~n973 ^ ~n975;
  assign n978 = ~n976 & ~n974;
  assign n979 = pi094 & pi222;
  assign n980 = ~pi094 & ~pi222;
  assign n981 = pi094 ^ ~pi222;
  assign po094 = ~n978 ^ ~n981;
  assign n983 = pi095 & pi223;
  assign n984 = pi095 ^ ~pi223;
  assign n985 = ~n978 & ~n980;
  assign n986 = ~n985 & ~n979;
  assign n987 = ~n986 & ~n984;
  assign po095 = ~n986 ^ ~n984;
  assign n989 = ~n987 & ~n983;
  assign n990 = ~n989 & pi224;
  assign n991 = n989 & ~pi224;
  assign n992 = pi096 ^ pi224;
  assign po096 = n989 ^ ~n992;
  assign n994 = pi097 & pi225;
  assign n995 = ~pi097 & ~pi225;
  assign n996 = pi097 ^ ~pi225;
  assign n997 = ~n991 & pi096;
  assign n998 = ~n997 & ~n990;
  assign po097 = ~n998 ^ ~n996;
  assign n1000 = ~pi098 & ~pi226;
  assign n1001 = pi098 ^ ~pi226;
  assign n1002 = ~n998 & ~n995;
  assign n1003 = ~n1002 & ~n994;
  assign po098 = ~n1003 ^ ~n1001;
  assign n1005 = ~n996 & ~n1001;
  assign n1006 = ~n998 & n1005;
  assign n1007 = ~n994 & ~n1001;
  assign n1008 = ~n1007 & ~n1000;
  assign n1009 = ~n1006 & ~n1008;
  assign n1010 = pi099 & pi227;
  assign n1011 = ~pi099 & ~pi227;
  assign n1012 = pi099 ^ ~pi227;
  assign po099 = n1009 ^ n1012;
  assign n1014 = ~pi100 & ~pi228;
  assign n1015 = pi100 ^ ~pi228;
  assign n1016 = ~n1009 & ~n1011;
  assign n1017 = ~n1016 & ~n1010;
  assign po100 = ~n1017 ^ ~n1015;
  assign n1019 = ~n1012 & ~n1015;
  assign n1020 = ~n1009 & n1019;
  assign n1021 = ~n1010 & ~n1015;
  assign n1022 = ~n1021 & ~n1014;
  assign n1023 = ~n1020 & ~n1022;
  assign n1024 = pi101 & pi229;
  assign n1025 = ~pi101 & ~pi229;
  assign n1026 = pi101 ^ ~pi229;
  assign po101 = n1023 ^ n1026;
  assign n1028 = ~pi102 & ~pi230;
  assign n1029 = pi102 ^ ~pi230;
  assign n1030 = ~n1023 & ~n1025;
  assign n1031 = ~n1030 & ~n1024;
  assign po102 = ~n1031 ^ ~n1029;
  assign n1033 = ~n1026 & ~n1029;
  assign n1034 = ~n1023 & n1033;
  assign n1035 = ~n1024 & ~n1029;
  assign n1036 = ~n1035 & ~n1028;
  assign n1037 = ~n1034 & ~n1036;
  assign n1038 = ~n1037 & pi231;
  assign n1039 = n1037 & ~pi231;
  assign n1040 = pi103 ^ pi231;
  assign po103 = n1037 ^ ~n1040;
  assign n1042 = ~pi104 & ~pi232;
  assign n1043 = pi104 & pi232;
  assign n1044 = pi104 ^ ~pi232;
  assign n1045 = ~n1039 & pi103;
  assign n1046 = ~n1045 & ~n1038;
  assign n1047 = ~n1046 & ~n1042;
  assign n1048 = ~n1047 & ~n1043;
  assign po104 = ~n1046 ^ ~n1044;
  assign n1050 = ~pi105 & ~pi233;
  assign n1051 = pi105 & pi233;
  assign n1052 = pi105 ^ ~pi233;
  assign n1053 = n1048 & ~n1051;
  assign po105 = ~n1048 ^ ~n1052;
  assign n1055 = ~pi106 & ~pi234;
  assign n1056 = pi106 ^ ~pi234;
  assign n1057 = ~n1053 & ~n1050;
  assign po106 = n1057 ^ ~n1056;
  assign n1059 = ~n1052 & ~n1056;
  assign n1060 = ~n1048 & n1059;
  assign n1061 = ~n1051 & ~n1056;
  assign n1062 = ~n1061 & ~n1055;
  assign n1063 = ~n1060 & ~n1062;
  assign n1064 = ~n1063 & pi235;
  assign n1065 = n1063 & ~pi235;
  assign n1066 = pi107 ^ pi235;
  assign po107 = n1063 ^ ~n1066;
  assign n1068 = pi108 & pi236;
  assign n1069 = ~pi108 & ~pi236;
  assign n1070 = pi108 ^ ~pi236;
  assign n1071 = ~n1065 & pi107;
  assign n1072 = ~n1071 & ~n1064;
  assign n1073 = ~n1072 & ~n1069;
  assign n1074 = ~n1073 & ~n1068;
  assign po108 = ~n1072 ^ ~n1070;
  assign n1076 = pi109 & pi237;
  assign n1077 = ~pi109 & ~pi237;
  assign n1078 = pi109 ^ ~pi237;
  assign po109 = ~n1074 ^ ~n1078;
  assign n1080 = ~pi110 & ~pi238;
  assign n1081 = pi110 ^ ~pi238;
  assign n1082 = ~n1074 & ~n1077;
  assign n1083 = ~n1082 & ~n1076;
  assign po110 = ~n1083 ^ ~n1081;
  assign n1085 = ~n1078 & ~n1081;
  assign n1086 = ~n1074 & n1085;
  assign n1087 = ~n1076 & ~n1081;
  assign n1088 = ~n1087 & ~n1080;
  assign n1089 = ~n1086 & ~n1088;
  assign n1090 = pi111 & pi239;
  assign n1091 = ~pi111 & ~pi239;
  assign n1092 = pi111 ^ ~pi239;
  assign po111 = n1089 ^ n1092;
  assign n1094 = ~n1089 & ~n1091;
  assign n1095 = ~n1094 & ~n1090;
  assign n1096 = pi112 & pi240;
  assign n1097 = ~pi112 & ~pi240;
  assign n1098 = n1095 & ~n1096;
  assign n1099 = ~n1098 & ~n1097;
  assign n1100 = pi112 ^ ~pi240;
  assign po112 = n1095 ^ n1100;
  assign n1102 = ~n1099 & ~pi241;
  assign n1103 = n1099 & pi241;
  assign n1104 = pi113 ^ pi241;
  assign po113 = ~n1099 ^ ~n1104;
  assign n1106 = ~n1103 & ~pi113;
  assign n1107 = ~n1106 & ~n1102;
  assign n1108 = ~pi114 & ~pi242;
  assign n1109 = pi114 & pi242;
  assign n1110 = ~n1107 & ~n1109;
  assign n1111 = ~n1110 & ~n1108;
  assign n1112 = pi114 ^ ~pi242;
  assign po114 = n1107 ^ ~n1112;
  assign n1114 = ~n1111 & ~pi243;
  assign n1115 = n1111 & pi243;
  assign n1116 = pi115 ^ pi243;
  assign po115 = ~n1111 ^ ~n1116;
  assign n1118 = ~n1115 & ~pi115;
  assign n1119 = ~n1118 & ~n1114;
  assign n1120 = pi116 & pi244;
  assign n1121 = ~pi116 & ~pi244;
  assign n1122 = ~n1119 & ~n1120;
  assign n1123 = ~n1122 & ~n1121;
  assign n1124 = pi116 ^ ~pi244;
  assign po116 = n1119 ^ ~n1124;
  assign n1126 = ~n1123 & ~pi245;
  assign n1127 = n1123 & pi245;
  assign n1128 = pi117 ^ pi245;
  assign po117 = ~n1123 ^ ~n1128;
  assign n1130 = ~n1127 & ~pi117;
  assign n1131 = ~n1130 & ~n1126;
  assign n1132 = pi118 & pi246;
  assign n1133 = ~pi118 & ~pi246;
  assign n1134 = ~n1131 & ~n1132;
  assign n1135 = ~n1134 & ~n1133;
  assign n1136 = pi118 ^ ~pi246;
  assign po118 = n1131 ^ ~n1136;
  assign n1138 = ~n1135 & ~pi247;
  assign n1139 = n1135 & pi247;
  assign n1140 = pi119 ^ pi247;
  assign po119 = ~n1135 ^ ~n1140;
  assign n1142 = ~n1139 & ~pi119;
  assign n1143 = ~n1142 & ~n1138;
  assign n1144 = pi120 & pi248;
  assign n1145 = ~pi120 & ~pi248;
  assign n1146 = ~n1143 & ~n1144;
  assign n1147 = ~n1146 & ~n1145;
  assign n1148 = pi120 ^ ~pi248;
  assign po120 = n1143 ^ ~n1148;
  assign n1150 = ~n1147 & ~pi249;
  assign n1151 = n1147 & pi249;
  assign n1152 = pi121 ^ pi249;
  assign po121 = ~n1147 ^ ~n1152;
  assign n1154 = ~n1151 & ~pi121;
  assign n1155 = ~n1154 & ~n1150;
  assign n1156 = pi122 & pi250;
  assign n1157 = ~pi122 & ~pi250;
  assign n1158 = ~n1155 & ~n1156;
  assign n1159 = ~n1158 & ~n1157;
  assign n1160 = pi122 ^ ~pi250;
  assign po122 = n1155 ^ ~n1160;
  assign n1162 = ~n1159 & ~pi251;
  assign n1163 = n1159 & pi251;
  assign n1164 = pi123 ^ pi251;
  assign po123 = ~n1159 ^ ~n1164;
  assign n1166 = ~n1163 & ~pi123;
  assign n1167 = ~n1166 & ~n1162;
  assign n1168 = pi124 & pi252;
  assign n1169 = ~pi124 & ~pi252;
  assign n1170 = ~n1167 & ~n1168;
  assign n1171 = ~n1170 & ~n1169;
  assign n1172 = pi124 ^ ~pi252;
  assign po124 = n1167 ^ ~n1172;
  assign n1174 = ~n1171 & ~pi253;
  assign n1175 = n1171 & pi253;
  assign n1176 = pi125 ^ pi253;
  assign po125 = ~n1171 ^ ~n1176;
  assign n1178 = ~n1175 & ~pi125;
  assign n1179 = ~n1178 & ~n1174;
  assign n1180 = pi126 & pi254;
  assign n1181 = ~pi126 & ~pi254;
  assign n1182 = ~n1179 & ~n1180;
  assign n1183 = ~n1182 & ~n1181;
  assign n1184 = pi126 ^ ~pi254;
  assign po126 = n1179 ^ ~n1184;
  assign n1186 = pi127 & pi255;
  assign n1187 = ~pi127 & ~pi255;
  assign n1188 = pi127 ^ ~pi255;
  assign po127 = n1183 ^ ~n1188;
  assign n1190 = n1183 & ~n1187;
  assign po128 = n1190 | n1186;
endmodule


