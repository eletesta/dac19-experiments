module top(n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438);
  input n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63;
  output n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438;
  wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405;
  assign n406 = n0 ^ n32;
  assign n373 = n5 & n37;
  assign n336 = n4 & n36;
  assign n340 = n10 & n42;
  assign n366 = n14 & n46;
  assign n341 = n24 & n56;
  assign n342 = n8 & n40;
  assign n343 = n1 & n33;
  assign n348 = n7 & n39;
  assign n349 = n28 & n60;
  assign n350 = n19 & n51;
  assign n351 = n2 & n34;
  assign n364 = n30 & n62;
  assign n352 = n13 & n45;
  assign n353 = n18 & n50;
  assign n355 = n11 & n43;
  assign n356 = n3 & n35;
  assign n359 = n16 & n48;
  assign n357 = n31 & n63;
  assign n358 = n27 & n59;
  assign n360 = n15 & n47;
  assign n361 = n17 & n49;
  assign n363 = n9 & n41;
  assign n278 = n32 & n0;
  assign n362 = n29 & n61;
  assign n365 = n6 & n38;
  assign n354 = n25 & n57;
  assign n367 = n20 & n52;
  assign n331 = n22 & n54;
  assign n371 = n21 & n53;
  assign n372 = n12 & n44;
  assign n339 = n23 & n55;
  assign n368 = n26 & n58;
  assign n398 = ~n56;
  assign n314 = ~n3;
  assign n346 = ~n40;
  assign n378 = ~n62;
  assign n389 = ~n6;
  assign n401 = ~n28;
  assign n377 = ~n10;
  assign n391 = ~n13;
  assign n335 = ~n27;
  assign n387 = ~n7;
  assign n399 = ~n24;
  assign n327 = ~n54;
  assign n315 = ~n36;
  assign n332 = ~n52;
  assign n380 = ~n50;
  assign n404 = ~n57;
  assign n323 = ~n31;
  assign n317 = ~n55;
  assign n381 = ~n18;
  assign n400 = ~n60;
  assign n322 = ~n5;
  assign n395 = ~n14;
  assign n402 = ~n47;
  assign n347 = ~n8;
  assign n385 = ~n19;
  assign n374 = ~n53;
  assign n330 = ~n29;
  assign n382 = ~n1;
  assign n344 = ~n34;
  assign n333 = ~n20;
  assign n321 = ~n37;
  assign n390 = ~n45;
  assign n338 = ~n11;
  assign n376 = ~n42;
  assign n370 = ~n12;
  assign n388 = ~n38;
  assign n318 = ~n23;
  assign n392 = ~n41;
  assign n329 = ~n61;
  assign n403 = ~n15;
  assign n396 = ~n48;
  assign n320 = ~n26;
  assign n337 = ~n43;
  assign n334 = ~n59;
  assign n393 = ~n9;
  assign n319 = ~n58;
  assign n326 = ~n17;
  assign n369 = ~n44;
  assign n375 = ~n21;
  assign n325 = ~n49;
  assign n397 = ~n16;
  assign n405 = ~n25;
  assign n384 = ~n51;
  assign n316 = ~n4;
  assign n345 = ~n2;
  assign n386 = ~n39;
  assign n394 = ~n46;
  assign n313 = ~n35;
  assign n328 = ~n22;
  assign n324 = ~n63;
  assign n383 = ~n33;
  assign n379 = ~n30;
  assign n282 = n313 & n314;
  assign n283 = n315 & n316;
  assign n284 = n317 & n318;
  assign n299 = n319 & n320;
  assign n285 = n321 & n322;
  assign n286 = n323 & n324;
  assign n288 = n325 & n326;
  assign n289 = n327 & n328;
  assign n290 = n329 & n330;
  assign n130 = ~n331;
  assign n287 = n332 & n333;
  assign n292 = n334 & n335;
  assign n256 = ~n336;
  assign n293 = n337 & n338;
  assign n123 = ~n339;
  assign n214 = ~n340;
  assign n116 = ~n341;
  assign n228 = ~n342;
  assign n276 = ~n343;
  assign n310 = n344 & n345;
  assign n300 = n346 & n347;
  assign n235 = ~n348;
  assign n88 = ~n349;
  assign n151 = ~n350;
  assign n270 = ~n351;
  assign n193 = ~n352;
  assign n158 = ~n353;
  assign n109 = ~n354;
  assign n207 = ~n355;
  assign n263 = ~n356;
  assign n66 = ~n357;
  assign n95 = ~n358;
  assign n172 = ~n359;
  assign n179 = ~n360;
  assign n165 = ~n361;
  assign n81 = ~n362;
  assign n221 = ~n363;
  assign n74 = ~n364;
  assign n242 = ~n365;
  assign n186 = ~n366;
  assign n144 = ~n367;
  assign n102 = ~n368;
  assign n301 = n369 & n370;
  assign n137 = ~n371;
  assign n200 = ~n372;
  assign n249 = ~n373;
  assign n298 = n374 & n375;
  assign n296 = n376 & n377;
  assign n291 = n378 & n379;
  assign n297 = n380 & n381;
  assign n306 = n382 & n383;
  assign n294 = n384 & n385;
  assign n295 = n386 & n387;
  assign n302 = n388 & n389;
  assign n303 = n390 & n391;
  assign n304 = n392 & n393;
  assign n305 = n394 & n395;
  assign n307 = n396 & n397;
  assign n308 = n398 & n399;
  assign n309 = n400 & n401;
  assign n311 = n402 & n403;
  assign n312 = n404 & n405;
  assign n266 = ~n282;
  assign n259 = ~n283;
  assign n126 = ~n284;
  assign n252 = ~n285;
  assign n69 = ~n286;
  assign n147 = ~n287;
  assign n168 = ~n288;
  assign n133 = ~n289;
  assign n84 = ~n290;
  assign n77 = ~n291;
  assign n98 = ~n292;
  assign n210 = ~n293;
  assign n154 = ~n294;
  assign n238 = ~n295;
  assign n217 = ~n296;
  assign n161 = ~n297;
  assign n140 = ~n298;
  assign n105 = ~n299;
  assign n231 = ~n300;
  assign n203 = ~n301;
  assign n245 = ~n302;
  assign n196 = ~n303;
  assign n224 = ~n304;
  assign n189 = ~n305;
  assign n281 = ~n306;
  assign n175 = ~n307;
  assign n119 = ~n308;
  assign n91 = ~n309;
  assign n273 = ~n310;
  assign n182 = ~n311;
  assign n112 = ~n312;
  assign n277 = n281 & n276;
  assign n279 = n69 & n66;
  assign n280 = n281 & n278;
  assign n407 = n277 ^ n278;
  assign n71 = ~n279;
  assign n275 = ~n280;
  assign n274 = n275 & n276;
  assign n271 = ~n274;
  assign n268 = n2 ^ n271;
  assign n272 = n271 & n273;
  assign n408 = n34 ^ n268;
  assign n269 = ~n272;
  assign n267 = n269 & n270;
  assign n264 = ~n267;
  assign n261 = n3 ^ n264;
  assign n265 = n264 & n266;
  assign n409 = n35 ^ n261;
  assign n262 = ~n265;
  assign n260 = n262 & n263;
  assign n257 = ~n260;
  assign n253 = n4 ^ n257;
  assign n258 = n257 & n259;
  assign n410 = n36 ^ n253;
  assign n255 = ~n258;
  assign n254 = n255 & n256;
  assign n250 = ~n254;
  assign n247 = n5 ^ n250;
  assign n251 = n250 & n252;
  assign n411 = n37 ^ n247;
  assign n248 = ~n251;
  assign n246 = n248 & n249;
  assign n243 = ~n246;
  assign n239 = n6 ^ n243;
  assign n244 = n243 & n245;
  assign n412 = n38 ^ n239;
  assign n241 = ~n244;
  assign n240 = n241 & n242;
  assign n236 = ~n240;
  assign n233 = n7 ^ n236;
  assign n237 = n236 & n238;
  assign n413 = n39 ^ n233;
  assign n234 = ~n237;
  assign n232 = n234 & n235;
  assign n229 = ~n232;
  assign n226 = n8 ^ n229;
  assign n230 = n229 & n231;
  assign n414 = n40 ^ n226;
  assign n227 = ~n230;
  assign n225 = n227 & n228;
  assign n222 = ~n225;
  assign n219 = n9 ^ n222;
  assign n223 = n222 & n224;
  assign n415 = n41 ^ n219;
  assign n220 = ~n223;
  assign n218 = n220 & n221;
  assign n215 = ~n218;
  assign n212 = n10 ^ n215;
  assign n216 = n215 & n217;
  assign n416 = n42 ^ n212;
  assign n213 = ~n216;
  assign n211 = n213 & n214;
  assign n208 = ~n211;
  assign n205 = n11 ^ n208;
  assign n209 = n208 & n210;
  assign n417 = n43 ^ n205;
  assign n206 = ~n209;
  assign n204 = n206 & n207;
  assign n201 = ~n204;
  assign n198 = n12 ^ n201;
  assign n202 = n201 & n203;
  assign n418 = n44 ^ n198;
  assign n199 = ~n202;
  assign n197 = n199 & n200;
  assign n195 = ~n197;
  assign n190 = n13 ^ n195;
  assign n194 = n195 & n196;
  assign n419 = n45 ^ n190;
  assign n192 = ~n194;
  assign n191 = n192 & n193;
  assign n187 = ~n191;
  assign n183 = n14 ^ n187;
  assign n188 = n187 & n189;
  assign n420 = n46 ^ n183;
  assign n185 = ~n188;
  assign n184 = n185 & n186;
  assign n180 = ~n184;
  assign n177 = n15 ^ n180;
  assign n181 = n180 & n182;
  assign n421 = n47 ^ n177;
  assign n178 = ~n181;
  assign n176 = n178 & n179;
  assign n173 = ~n176;
  assign n170 = n48 ^ n173;
  assign n174 = n173 & n175;
  assign n422 = n16 ^ n170;
  assign n171 = ~n174;
  assign n169 = n171 & n172;
  assign n166 = ~n169;
  assign n163 = n17 ^ n166;
  assign n167 = n166 & n168;
  assign n423 = n49 ^ n163;
  assign n164 = ~n167;
  assign n162 = n164 & n165;
  assign n159 = ~n162;
  assign n156 = n18 ^ n159;
  assign n160 = n159 & n161;
  assign n424 = n50 ^ n156;
  assign n157 = ~n160;
  assign n155 = n157 & n158;
  assign n152 = ~n155;
  assign n149 = n19 ^ n152;
  assign n153 = n152 & n154;
  assign n425 = n51 ^ n149;
  assign n150 = ~n153;
  assign n148 = n150 & n151;
  assign n145 = ~n148;
  assign n141 = n20 ^ n145;
  assign n146 = n145 & n147;
  assign n426 = n52 ^ n141;
  assign n143 = ~n146;
  assign n142 = n143 & n144;
  assign n138 = ~n142;
  assign n135 = n53 ^ n138;
  assign n139 = n138 & n140;
  assign n427 = n21 ^ n135;
  assign n136 = ~n139;
  assign n134 = n136 & n137;
  assign n132 = ~n134;
  assign n127 = n22 ^ n132;
  assign n131 = n132 & n133;
  assign n428 = n54 ^ n127;
  assign n129 = ~n131;
  assign n128 = n129 & n130;
  assign n124 = ~n128;
  assign n121 = n23 ^ n124;
  assign n125 = n124 & n126;
  assign n429 = n55 ^ n121;
  assign n122 = ~n125;
  assign n120 = n122 & n123;
  assign n117 = ~n120;
  assign n114 = n24 ^ n117;
  assign n118 = n117 & n119;
  assign n430 = n56 ^ n114;
  assign n115 = ~n118;
  assign n113 = n115 & n116;
  assign n110 = ~n113;
  assign n107 = n25 ^ n110;
  assign n111 = n110 & n112;
  assign n431 = n57 ^ n107;
  assign n108 = ~n111;
  assign n106 = n108 & n109;
  assign n103 = ~n106;
  assign n100 = n26 ^ n103;
  assign n104 = n103 & n105;
  assign n432 = n58 ^ n100;
  assign n101 = ~n104;
  assign n99 = n101 & n102;
  assign n96 = ~n99;
  assign n93 = n59 ^ n96;
  assign n97 = n96 & n98;
  assign n433 = n27 ^ n93;
  assign n94 = ~n97;
  assign n92 = n94 & n95;
  assign n89 = ~n92;
  assign n86 = n28 ^ n89;
  assign n90 = n89 & n91;
  assign n434 = n60 ^ n86;
  assign n87 = ~n90;
  assign n85 = n87 & n88;
  assign n83 = ~n85;
  assign n79 = n61 ^ n83;
  assign n82 = n83 & n84;
  assign n435 = n29 ^ n79;
  assign n80 = ~n82;
  assign n78 = n80 & n81;
  assign n76 = ~n78;
  assign n72 = n30 ^ n76;
  assign n75 = n76 & n77;
  assign n436 = n62 ^ n72;
  assign n73 = ~n75;
  assign n70 = n73 & n74;
  assign n437 = n70 ^ n71;
  assign n68 = ~n70;
  assign n67 = n68 & n69;
  assign n65 = ~n67;
  assign n64 = n65 & n66;
  assign n438 = ~n64;
endmodule
