module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32;
  wire n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248;
  assign n65 = x32 ^ x0;
  assign n67 = x0 & x32;
  assign n66 = x33 ^ x1;
  assign n68 = n67 ^ n66;
  assign n69 = x1 & x33;
  assign n70 = ~x1 & ~x33;
  assign n71 = n67 & ~n70;
  assign n72 = ~n69 & ~n71;
  assign n73 = n72 ^ x2;
  assign n74 = n73 ^ x34;
  assign n75 = x34 ^ x2;
  assign n76 = n72 ^ x34;
  assign n77 = n75 & n76;
  assign n78 = n77 ^ x2;
  assign n79 = n78 ^ x3;
  assign n80 = n79 ^ x35;
  assign n81 = x35 ^ x3;
  assign n82 = n78 ^ x35;
  assign n83 = n81 & ~n82;
  assign n84 = n83 ^ x3;
  assign n85 = n84 ^ x4;
  assign n86 = n85 ^ x36;
  assign n87 = x36 ^ x4;
  assign n88 = n84 ^ x36;
  assign n89 = n87 & ~n88;
  assign n90 = n89 ^ x4;
  assign n91 = n90 ^ x5;
  assign n92 = n91 ^ x37;
  assign n93 = x37 ^ x5;
  assign n94 = n90 ^ x37;
  assign n95 = n93 & ~n94;
  assign n96 = n95 ^ x5;
  assign n97 = n96 ^ x6;
  assign n98 = n97 ^ x38;
  assign n99 = x38 ^ x6;
  assign n100 = n96 ^ x38;
  assign n101 = n99 & ~n100;
  assign n102 = n101 ^ x6;
  assign n103 = n102 ^ x7;
  assign n104 = n103 ^ x39;
  assign n105 = x39 ^ x7;
  assign n106 = n102 ^ x39;
  assign n107 = n105 & ~n106;
  assign n108 = n107 ^ x7;
  assign n109 = n108 ^ x8;
  assign n110 = n109 ^ x40;
  assign n111 = x40 ^ x8;
  assign n112 = n108 ^ x40;
  assign n113 = n111 & ~n112;
  assign n114 = n113 ^ x8;
  assign n115 = n114 ^ x9;
  assign n116 = n115 ^ x41;
  assign n117 = x41 ^ x9;
  assign n118 = n114 ^ x41;
  assign n119 = n117 & ~n118;
  assign n120 = n119 ^ x9;
  assign n121 = n120 ^ x10;
  assign n122 = n121 ^ x42;
  assign n123 = x42 ^ x10;
  assign n124 = n120 ^ x42;
  assign n125 = n123 & ~n124;
  assign n126 = n125 ^ x10;
  assign n127 = n126 ^ x11;
  assign n128 = n127 ^ x43;
  assign n129 = x43 ^ x11;
  assign n130 = n126 ^ x43;
  assign n131 = n129 & ~n130;
  assign n132 = n131 ^ x11;
  assign n133 = n132 ^ x12;
  assign n134 = n133 ^ x44;
  assign n135 = x44 ^ x12;
  assign n136 = n132 ^ x44;
  assign n137 = n135 & ~n136;
  assign n138 = n137 ^ x12;
  assign n139 = n138 ^ x13;
  assign n140 = n139 ^ x45;
  assign n141 = x45 ^ x13;
  assign n142 = n138 ^ x45;
  assign n143 = n141 & ~n142;
  assign n144 = n143 ^ x13;
  assign n145 = n144 ^ x14;
  assign n146 = n145 ^ x46;
  assign n147 = x46 ^ x14;
  assign n148 = n144 ^ x46;
  assign n149 = n147 & ~n148;
  assign n150 = n149 ^ x14;
  assign n151 = n150 ^ x15;
  assign n152 = n151 ^ x47;
  assign n153 = x47 ^ x15;
  assign n154 = n150 ^ x47;
  assign n155 = n153 & ~n154;
  assign n156 = n155 ^ x15;
  assign n157 = n156 ^ x48;
  assign n158 = n157 ^ x16;
  assign n159 = x48 ^ x16;
  assign n160 = ~n157 & n159;
  assign n161 = n160 ^ x16;
  assign n162 = n161 ^ x17;
  assign n163 = n162 ^ x49;
  assign n164 = x49 ^ x17;
  assign n165 = n161 ^ x49;
  assign n166 = n164 & ~n165;
  assign n167 = n166 ^ x17;
  assign n168 = n167 ^ x18;
  assign n169 = n168 ^ x50;
  assign n170 = x50 ^ x18;
  assign n171 = n167 ^ x50;
  assign n172 = n170 & ~n171;
  assign n173 = n172 ^ x18;
  assign n174 = n173 ^ x19;
  assign n175 = n174 ^ x51;
  assign n176 = x51 ^ x19;
  assign n177 = n173 ^ x51;
  assign n178 = n176 & ~n177;
  assign n179 = n178 ^ x19;
  assign n180 = n179 ^ x20;
  assign n181 = n180 ^ x52;
  assign n182 = x52 ^ x20;
  assign n183 = n179 ^ x52;
  assign n184 = n182 & ~n183;
  assign n185 = n184 ^ x20;
  assign n186 = n185 ^ x53;
  assign n187 = n186 ^ x21;
  assign n188 = x53 ^ x21;
  assign n189 = ~n186 & n188;
  assign n190 = n189 ^ x21;
  assign n191 = n190 ^ x22;
  assign n192 = n191 ^ x54;
  assign n193 = x54 ^ x22;
  assign n194 = n190 ^ x54;
  assign n195 = n193 & ~n194;
  assign n196 = n195 ^ x22;
  assign n197 = n196 ^ x23;
  assign n198 = n197 ^ x55;
  assign n199 = x55 ^ x23;
  assign n200 = n196 ^ x55;
  assign n201 = n199 & ~n200;
  assign n202 = n201 ^ x23;
  assign n203 = n202 ^ x24;
  assign n204 = n203 ^ x56;
  assign n205 = x56 ^ x24;
  assign n206 = n202 ^ x56;
  assign n207 = n205 & ~n206;
  assign n208 = n207 ^ x24;
  assign n209 = n208 ^ x25;
  assign n210 = n209 ^ x57;
  assign n211 = x57 ^ x25;
  assign n212 = n208 ^ x57;
  assign n213 = n211 & ~n212;
  assign n214 = n213 ^ x25;
  assign n215 = n214 ^ x26;
  assign n216 = n215 ^ x58;
  assign n217 = x58 ^ x26;
  assign n218 = n214 ^ x58;
  assign n219 = n217 & ~n218;
  assign n220 = n219 ^ x26;
  assign n221 = n220 ^ x59;
  assign n222 = n221 ^ x27;
  assign n223 = x59 ^ x27;
  assign n224 = ~n221 & n223;
  assign n225 = n224 ^ x27;
  assign n226 = n225 ^ x28;
  assign n227 = n226 ^ x60;
  assign n228 = x60 ^ x28;
  assign n229 = n225 ^ x60;
  assign n230 = n228 & ~n229;
  assign n231 = n230 ^ x28;
  assign n232 = n231 ^ x61;
  assign n233 = n232 ^ x29;
  assign n234 = x61 ^ x29;
  assign n235 = ~n232 & n234;
  assign n236 = n235 ^ x29;
  assign n237 = n236 ^ x30;
  assign n238 = n237 ^ x62;
  assign n240 = x62 ^ x30;
  assign n241 = n236 ^ x62;
  assign n242 = n240 & ~n241;
  assign n243 = n242 ^ x30;
  assign n239 = x63 ^ x31;
  assign n244 = n243 ^ n239;
  assign n245 = x31 & x63;
  assign n246 = ~x31 & ~x63;
  assign n247 = n243 & ~n246;
  assign n248 = ~n245 & ~n247;
  assign y0 = n65;
  assign y1 = n68;
  assign y2 = ~n74;
  assign y3 = n80;
  assign y4 = n86;
  assign y5 = n92;
  assign y6 = n98;
  assign y7 = n104;
  assign y8 = n110;
  assign y9 = n116;
  assign y10 = n122;
  assign y11 = n128;
  assign y12 = n134;
  assign y13 = n140;
  assign y14 = n146;
  assign y15 = n152;
  assign y16 = n158;
  assign y17 = n163;
  assign y18 = n169;
  assign y19 = n175;
  assign y20 = n181;
  assign y21 = n187;
  assign y22 = n192;
  assign y23 = n198;
  assign y24 = n204;
  assign y25 = n210;
  assign y26 = n216;
  assign y27 = n222;
  assign y28 = n227;
  assign y29 = n233;
  assign y30 = n238;
  assign y31 = n244;
  assign y32 = ~n248;
endmodule
