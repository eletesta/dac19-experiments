module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63;
  wire n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579;
  assign n65 = x0 & x32;
  assign n71 = x33 & ~n65;
  assign n68 = ~x32 & x33;
  assign n69 = ~x0 & n68;
  assign n66 = x33 ^ x1;
  assign n67 = x32 & n66;
  assign n70 = n69 ^ n67;
  assign n72 = n71 ^ n70;
  assign n77 = x33 ^ x2;
  assign n78 = x32 & n77;
  assign n76 = ~x1 & n68;
  assign n79 = n78 ^ n76;
  assign n74 = x34 ^ x33;
  assign n75 = x0 & n74;
  assign n80 = n79 ^ n75;
  assign n73 = n70 & n71;
  assign n81 = n80 ^ n73;
  assign n105 = n75 ^ n73;
  assign n106 = ~n80 & n105;
  assign n107 = n106 ^ n73;
  assign n99 = x33 ^ x0;
  assign n100 = ~n74 & n99;
  assign n101 = n100 ^ x0;
  assign n102 = x35 & ~n101;
  assign n97 = ~x2 & n68;
  assign n95 = x33 ^ x3;
  assign n96 = x32 & n95;
  assign n98 = n97 ^ n96;
  assign n103 = n102 ^ n98;
  assign n82 = x35 & n74;
  assign n83 = ~x1 & n82;
  assign n84 = x35 ^ x34;
  assign n85 = ~n74 & n84;
  assign n86 = x35 & n85;
  assign n87 = ~x0 & n86;
  assign n88 = ~n83 & ~n87;
  assign n89 = ~x35 & n74;
  assign n90 = x1 & n89;
  assign n91 = ~x35 & n85;
  assign n92 = x0 & n91;
  assign n93 = ~n90 & ~n92;
  assign n94 = n88 & n93;
  assign n104 = n103 ^ n94;
  assign n108 = n107 ^ n104;
  assign n126 = n107 ^ n94;
  assign n127 = n104 & ~n126;
  assign n128 = n127 ^ n107;
  assign n121 = x33 ^ x4;
  assign n122 = x32 & n121;
  assign n120 = ~x3 & n68;
  assign n123 = n122 ^ n120;
  assign n112 = x2 & n89;
  assign n113 = x1 & n91;
  assign n114 = ~n112 & ~n113;
  assign n115 = ~x2 & n82;
  assign n116 = ~x1 & n86;
  assign n117 = ~n115 & ~n116;
  assign n118 = n114 & n117;
  assign n110 = x36 ^ x35;
  assign n111 = x0 & n110;
  assign n119 = n118 ^ n111;
  assign n124 = n123 ^ n119;
  assign n109 = n98 & n102;
  assign n125 = n124 ^ n109;
  assign n129 = n128 ^ n125;
  assign n166 = n128 ^ n109;
  assign n167 = n125 & n166;
  assign n168 = n167 ^ n128;
  assign n161 = n123 ^ n111;
  assign n162 = n123 ^ n118;
  assign n163 = n161 & n162;
  assign n164 = n163 ^ n111;
  assign n146 = x37 & n110;
  assign n147 = ~x1 & n146;
  assign n148 = x37 ^ x36;
  assign n149 = ~n110 & n148;
  assign n150 = x37 & n149;
  assign n151 = ~x0 & n150;
  assign n152 = ~n147 & ~n151;
  assign n153 = ~x37 & n110;
  assign n154 = x1 & n153;
  assign n155 = ~x37 & n149;
  assign n156 = x0 & n155;
  assign n157 = ~n154 & ~n156;
  assign n158 = n152 & n157;
  assign n139 = x3 & n89;
  assign n140 = x2 & n91;
  assign n141 = ~n139 & ~n140;
  assign n142 = ~x3 & n82;
  assign n143 = ~x2 & n86;
  assign n144 = ~n142 & ~n143;
  assign n145 = n141 & n144;
  assign n159 = n158 ^ n145;
  assign n134 = x35 ^ x0;
  assign n135 = ~n110 & n134;
  assign n136 = n135 ^ x0;
  assign n137 = x37 & ~n136;
  assign n132 = ~x4 & n68;
  assign n130 = x33 ^ x5;
  assign n131 = x32 & n130;
  assign n133 = n132 ^ n131;
  assign n138 = n137 ^ n133;
  assign n160 = n159 ^ n138;
  assign n165 = n164 ^ n160;
  assign n169 = n168 ^ n165;
  assign n199 = n168 ^ n160;
  assign n200 = ~n165 & n199;
  assign n201 = n200 ^ n168;
  assign n195 = n158 ^ n138;
  assign n196 = n159 & n195;
  assign n197 = n196 ^ n145;
  assign n192 = n133 & n137;
  assign n185 = ~x2 & n146;
  assign n186 = ~x1 & n150;
  assign n187 = ~n185 & ~n186;
  assign n188 = x2 & n153;
  assign n189 = x1 & n155;
  assign n190 = ~n188 & ~n189;
  assign n191 = n187 & n190;
  assign n193 = n192 ^ n191;
  assign n177 = ~x4 & n82;
  assign n178 = ~x3 & n86;
  assign n179 = ~n177 & ~n178;
  assign n180 = x4 & n89;
  assign n181 = x3 & n91;
  assign n182 = ~n180 & ~n181;
  assign n183 = n179 & n182;
  assign n173 = x33 ^ x6;
  assign n174 = x32 & n173;
  assign n172 = ~x5 & n68;
  assign n175 = n174 ^ n172;
  assign n170 = x38 ^ x37;
  assign n171 = x0 & n170;
  assign n176 = n175 ^ n171;
  assign n184 = n183 ^ n176;
  assign n194 = n193 ^ n184;
  assign n198 = n197 ^ n194;
  assign n202 = n201 ^ n198;
  assign n250 = n201 ^ n194;
  assign n251 = n198 & n250;
  assign n252 = n251 ^ n201;
  assign n246 = n192 ^ n184;
  assign n247 = ~n193 & n246;
  assign n248 = n247 ^ n191;
  assign n241 = n183 ^ n175;
  assign n242 = n176 & n241;
  assign n243 = n242 ^ n171;
  assign n236 = x37 ^ x0;
  assign n237 = ~n170 & n236;
  assign n238 = n237 ^ x0;
  assign n239 = x39 & ~n238;
  assign n234 = ~x6 & n68;
  assign n232 = x33 ^ x7;
  assign n233 = x32 & n232;
  assign n235 = n234 ^ n233;
  assign n240 = n239 ^ n235;
  assign n244 = n243 ^ n240;
  assign n223 = x5 & n89;
  assign n224 = x4 & n91;
  assign n225 = ~n223 & ~n224;
  assign n226 = ~x5 & n82;
  assign n227 = ~x4 & n86;
  assign n228 = ~n226 & ~n227;
  assign n229 = n225 & n228;
  assign n210 = x39 & n170;
  assign n211 = ~x1 & n210;
  assign n212 = x39 ^ x38;
  assign n213 = ~n170 & n212;
  assign n214 = x39 & n213;
  assign n215 = ~x0 & n214;
  assign n216 = ~n211 & ~n215;
  assign n217 = ~x39 & n170;
  assign n218 = x1 & n217;
  assign n219 = ~x39 & n213;
  assign n220 = x0 & n219;
  assign n221 = ~n218 & ~n220;
  assign n222 = n216 & n221;
  assign n230 = n229 ^ n222;
  assign n203 = x3 & n153;
  assign n204 = x2 & n155;
  assign n205 = ~n203 & ~n204;
  assign n206 = ~x3 & n146;
  assign n207 = ~x2 & n150;
  assign n208 = ~n206 & ~n207;
  assign n209 = n205 & n208;
  assign n231 = n230 ^ n209;
  assign n245 = n244 ^ n231;
  assign n249 = n248 ^ n245;
  assign n253 = n252 ^ n249;
  assign n297 = n252 ^ n245;
  assign n298 = ~n249 & ~n297;
  assign n299 = n298 ^ n252;
  assign n292 = n240 ^ n231;
  assign n293 = n243 ^ n231;
  assign n294 = ~n292 & n293;
  assign n295 = n294 ^ n240;
  assign n286 = n222 ^ n209;
  assign n287 = n229 ^ n209;
  assign n288 = n286 & ~n287;
  assign n289 = n288 ^ n222;
  assign n278 = ~x2 & n210;
  assign n279 = ~x1 & n214;
  assign n280 = ~n278 & ~n279;
  assign n281 = x2 & n217;
  assign n282 = x1 & n219;
  assign n283 = ~n281 & ~n282;
  assign n284 = n280 & n283;
  assign n274 = x33 ^ x8;
  assign n275 = x32 & n274;
  assign n273 = ~x7 & n68;
  assign n276 = n275 ^ n273;
  assign n271 = x40 ^ x39;
  assign n272 = x0 & n271;
  assign n277 = n276 ^ n272;
  assign n285 = n284 ^ n277;
  assign n290 = n289 ^ n285;
  assign n262 = ~x4 & n146;
  assign n263 = ~x3 & n150;
  assign n264 = ~n262 & ~n263;
  assign n265 = x4 & n153;
  assign n266 = x3 & n155;
  assign n267 = ~n265 & ~n266;
  assign n268 = n264 & n267;
  assign n255 = ~x6 & n82;
  assign n256 = ~x5 & n86;
  assign n257 = ~n255 & ~n256;
  assign n258 = x6 & n89;
  assign n259 = x5 & n91;
  assign n260 = ~n258 & ~n259;
  assign n261 = n257 & n260;
  assign n269 = n268 ^ n261;
  assign n254 = n235 & n239;
  assign n270 = n269 ^ n254;
  assign n291 = n290 ^ n270;
  assign n296 = n295 ^ n291;
  assign n300 = n299 ^ n296;
  assign n361 = n299 ^ n291;
  assign n362 = ~n296 & n361;
  assign n363 = n362 ^ n299;
  assign n356 = n285 ^ n270;
  assign n357 = n289 ^ n270;
  assign n358 = ~n356 & n357;
  assign n359 = n358 ^ n285;
  assign n351 = n268 ^ n254;
  assign n352 = n269 & n351;
  assign n353 = n352 ^ n261;
  assign n342 = ~x3 & n210;
  assign n343 = ~x2 & n214;
  assign n344 = ~n342 & ~n343;
  assign n345 = x3 & n217;
  assign n346 = x2 & n219;
  assign n347 = ~n345 & ~n346;
  assign n348 = n344 & n347;
  assign n329 = x41 & n271;
  assign n330 = ~x1 & n329;
  assign n331 = x41 ^ x40;
  assign n332 = ~n271 & n331;
  assign n333 = x41 & n332;
  assign n334 = ~x0 & n333;
  assign n335 = ~n330 & ~n334;
  assign n336 = ~x41 & n271;
  assign n337 = x1 & n336;
  assign n338 = ~x41 & n332;
  assign n339 = x0 & n338;
  assign n340 = ~n337 & ~n339;
  assign n341 = n335 & n340;
  assign n349 = n348 ^ n341;
  assign n327 = ~x8 & n68;
  assign n325 = x33 ^ x9;
  assign n326 = x32 & n325;
  assign n328 = n327 ^ n326;
  assign n350 = n349 ^ n328;
  assign n354 = n353 ^ n350;
  assign n321 = n284 ^ n276;
  assign n322 = n277 & n321;
  assign n323 = n322 ^ n272;
  assign n312 = ~x7 & n82;
  assign n313 = ~x6 & n86;
  assign n314 = ~n312 & ~n313;
  assign n315 = x7 & n89;
  assign n316 = x6 & n91;
  assign n317 = ~n315 & ~n316;
  assign n318 = n314 & n317;
  assign n308 = x39 ^ x0;
  assign n309 = ~n271 & n308;
  assign n310 = n309 ^ x0;
  assign n311 = x41 & ~n310;
  assign n319 = n318 ^ n311;
  assign n301 = x5 & n153;
  assign n302 = x4 & n155;
  assign n303 = ~n301 & ~n302;
  assign n304 = ~x5 & n146;
  assign n305 = ~x4 & n150;
  assign n306 = ~n304 & ~n305;
  assign n307 = n303 & n306;
  assign n320 = n319 ^ n307;
  assign n324 = n323 ^ n320;
  assign n355 = n354 ^ n324;
  assign n360 = n359 ^ n355;
  assign n364 = n363 ^ n360;
  assign n419 = n363 ^ n355;
  assign n420 = ~n360 & ~n419;
  assign n421 = n420 ^ n363;
  assign n414 = n350 ^ n324;
  assign n415 = n353 ^ n324;
  assign n416 = n414 & n415;
  assign n417 = n416 ^ n350;
  assign n409 = n323 ^ n319;
  assign n410 = n320 & n409;
  assign n411 = n410 ^ n307;
  assign n404 = x33 ^ x10;
  assign n405 = x32 & n404;
  assign n403 = ~x9 & n68;
  assign n406 = n405 ^ n403;
  assign n396 = ~x2 & n329;
  assign n397 = ~x1 & n333;
  assign n398 = ~n396 & ~n397;
  assign n399 = x2 & n336;
  assign n400 = x1 & n338;
  assign n401 = ~n399 & ~n400;
  assign n402 = n398 & n401;
  assign n407 = n406 ^ n402;
  assign n389 = ~x6 & n146;
  assign n390 = ~x5 & n150;
  assign n391 = ~n389 & ~n390;
  assign n392 = x6 & n153;
  assign n393 = x5 & n155;
  assign n394 = ~n392 & ~n393;
  assign n395 = n391 & n394;
  assign n408 = n407 ^ n395;
  assign n412 = n411 ^ n408;
  assign n384 = n341 ^ n328;
  assign n385 = ~n349 & ~n384;
  assign n386 = n385 ^ n328;
  assign n383 = n311 & ~n318;
  assign n387 = n386 ^ n383;
  assign n374 = ~x8 & n82;
  assign n375 = ~x7 & n86;
  assign n376 = ~n374 & ~n375;
  assign n377 = x8 & n89;
  assign n378 = x7 & n91;
  assign n379 = ~n377 & ~n378;
  assign n380 = n376 & n379;
  assign n372 = x42 ^ x41;
  assign n373 = x0 & n372;
  assign n381 = n380 ^ n373;
  assign n365 = x4 & n217;
  assign n366 = x3 & n219;
  assign n367 = ~n365 & ~n366;
  assign n368 = ~x4 & n210;
  assign n369 = ~x3 & n214;
  assign n370 = ~n368 & ~n369;
  assign n371 = n367 & n370;
  assign n382 = n381 ^ n371;
  assign n388 = n387 ^ n382;
  assign n413 = n412 ^ n388;
  assign n418 = n417 ^ n413;
  assign n422 = n421 ^ n418;
  assign n495 = n421 ^ n413;
  assign n496 = n418 & ~n495;
  assign n497 = n496 ^ n421;
  assign n490 = n408 ^ n388;
  assign n491 = n411 ^ n388;
  assign n492 = n490 & n491;
  assign n493 = n492 ^ n408;
  assign n486 = n383 ^ n382;
  assign n487 = ~n387 & n486;
  assign n488 = n487 ^ n382;
  assign n480 = n380 ^ n371;
  assign n481 = ~n381 & ~n480;
  assign n482 = n481 ^ n373;
  assign n477 = n402 ^ n395;
  assign n478 = ~n407 & ~n477;
  assign n479 = n478 ^ n406;
  assign n483 = n482 ^ n479;
  assign n468 = ~x3 & n329;
  assign n469 = ~x2 & n333;
  assign n470 = ~n468 & ~n469;
  assign n471 = x3 & n336;
  assign n472 = x2 & n338;
  assign n473 = ~n471 & ~n472;
  assign n474 = n470 & n473;
  assign n461 = ~x5 & n210;
  assign n462 = ~x4 & n214;
  assign n463 = ~n461 & ~n462;
  assign n464 = x5 & n217;
  assign n465 = x4 & n219;
  assign n466 = ~n464 & ~n465;
  assign n467 = n463 & n466;
  assign n475 = n474 ^ n467;
  assign n459 = ~x10 & n68;
  assign n457 = x33 ^ x11;
  assign n458 = x32 & n457;
  assign n460 = n459 ^ n458;
  assign n476 = n475 ^ n460;
  assign n484 = n483 ^ n476;
  assign n448 = x9 & n89;
  assign n449 = x8 & n91;
  assign n450 = ~n448 & ~n449;
  assign n451 = ~x9 & n82;
  assign n452 = ~x8 & n86;
  assign n453 = ~n451 & ~n452;
  assign n454 = n450 & n453;
  assign n444 = x41 ^ x0;
  assign n445 = ~n372 & n444;
  assign n446 = n445 ^ x0;
  assign n447 = x43 & ~n446;
  assign n455 = n454 ^ n447;
  assign n430 = ~x43 & n372;
  assign n431 = x1 & n430;
  assign n432 = x43 ^ x42;
  assign n433 = ~n372 & n432;
  assign n434 = ~x43 & n433;
  assign n435 = x0 & n434;
  assign n436 = ~n431 & ~n435;
  assign n437 = x43 & n372;
  assign n438 = ~x1 & n437;
  assign n439 = x43 & n433;
  assign n440 = ~x0 & n439;
  assign n441 = ~n438 & ~n440;
  assign n442 = n436 & n441;
  assign n423 = ~x7 & n146;
  assign n424 = ~x6 & n150;
  assign n425 = ~n423 & ~n424;
  assign n426 = x7 & n153;
  assign n427 = x6 & n155;
  assign n428 = ~n426 & ~n427;
  assign n429 = n425 & n428;
  assign n443 = n442 ^ n429;
  assign n456 = n455 ^ n443;
  assign n485 = n484 ^ n456;
  assign n489 = n488 ^ n485;
  assign n494 = n493 ^ n489;
  assign n498 = n497 ^ n494;
  assign n564 = n497 ^ n489;
  assign n565 = n494 & ~n564;
  assign n566 = n565 ^ n497;
  assign n560 = n488 ^ n484;
  assign n561 = ~n485 & ~n560;
  assign n562 = n561 ^ n456;
  assign n555 = n479 ^ n476;
  assign n556 = ~n483 & n555;
  assign n557 = n556 ^ n476;
  assign n551 = n467 ^ n460;
  assign n552 = ~n475 & ~n551;
  assign n553 = n552 ^ n460;
  assign n549 = n447 & ~n454;
  assign n542 = ~x8 & n146;
  assign n543 = ~x7 & n150;
  assign n544 = ~n542 & ~n543;
  assign n545 = x8 & n153;
  assign n546 = x7 & n155;
  assign n547 = ~n545 & ~n546;
  assign n548 = n544 & n547;
  assign n550 = n549 ^ n548;
  assign n554 = n553 ^ n550;
  assign n558 = n557 ^ n554;
  assign n538 = n455 ^ n442;
  assign n539 = n443 & ~n538;
  assign n540 = n539 ^ n429;
  assign n532 = x33 ^ x12;
  assign n533 = x32 & n532;
  assign n531 = ~x11 & n68;
  assign n534 = n533 ^ n531;
  assign n524 = ~x4 & n329;
  assign n525 = ~x3 & n333;
  assign n526 = ~n524 & ~n525;
  assign n527 = x4 & n336;
  assign n528 = x3 & n338;
  assign n529 = ~n527 & ~n528;
  assign n530 = n526 & n529;
  assign n535 = n534 ^ n530;
  assign n517 = x2 & n430;
  assign n518 = x1 & n434;
  assign n519 = ~n517 & ~n518;
  assign n520 = ~x2 & n437;
  assign n521 = ~x1 & n439;
  assign n522 = ~n520 & ~n521;
  assign n523 = n519 & n522;
  assign n536 = n535 ^ n523;
  assign n508 = x10 & n89;
  assign n509 = x9 & n91;
  assign n510 = ~n508 & ~n509;
  assign n511 = ~x10 & n82;
  assign n512 = ~x9 & n86;
  assign n513 = ~n511 & ~n512;
  assign n514 = n510 & n513;
  assign n506 = x44 ^ x43;
  assign n507 = x0 & n506;
  assign n515 = n514 ^ n507;
  assign n499 = ~x6 & n210;
  assign n500 = ~x5 & n214;
  assign n501 = ~n499 & ~n500;
  assign n502 = x6 & n217;
  assign n503 = x5 & n219;
  assign n504 = ~n502 & ~n503;
  assign n505 = n501 & n504;
  assign n516 = n515 ^ n505;
  assign n537 = n536 ^ n516;
  assign n541 = n540 ^ n537;
  assign n559 = n558 ^ n541;
  assign n563 = n562 ^ n559;
  assign n567 = n566 ^ n563;
  assign n652 = n566 ^ n559;
  assign n653 = n563 & n652;
  assign n654 = n653 ^ n566;
  assign n648 = n554 ^ n541;
  assign n649 = n558 & n648;
  assign n650 = n649 ^ n541;
  assign n643 = n540 ^ n536;
  assign n644 = n537 & n643;
  assign n645 = n644 ^ n516;
  assign n639 = n530 ^ n523;
  assign n640 = ~n535 & ~n639;
  assign n641 = n640 ^ n534;
  assign n634 = n507 ^ n505;
  assign n635 = n514 ^ n505;
  assign n636 = ~n634 & ~n635;
  assign n637 = n636 ^ n507;
  assign n629 = x43 ^ x0;
  assign n630 = ~n506 & n629;
  assign n631 = n630 ^ x0;
  assign n632 = x45 & ~n631;
  assign n627 = ~x12 & n68;
  assign n625 = x33 ^ x13;
  assign n626 = x32 & n625;
  assign n628 = n627 ^ n626;
  assign n633 = n632 ^ n628;
  assign n638 = n637 ^ n633;
  assign n642 = n641 ^ n638;
  assign n646 = n645 ^ n642;
  assign n621 = n553 ^ n549;
  assign n622 = ~n550 & ~n621;
  assign n623 = n622 ^ n548;
  assign n611 = x3 & n430;
  assign n612 = x2 & n434;
  assign n613 = ~n611 & ~n612;
  assign n614 = ~x3 & n437;
  assign n615 = ~x2 & n439;
  assign n616 = ~n614 & ~n615;
  assign n617 = n613 & n616;
  assign n604 = ~x9 & n146;
  assign n605 = ~x8 & n150;
  assign n606 = ~n604 & ~n605;
  assign n607 = x9 & n153;
  assign n608 = x8 & n155;
  assign n609 = ~n607 & ~n608;
  assign n610 = n606 & n609;
  assign n618 = n617 ^ n610;
  assign n591 = x45 & n506;
  assign n592 = ~x1 & n591;
  assign n593 = x45 ^ x44;
  assign n594 = ~n506 & n593;
  assign n595 = x45 & n594;
  assign n596 = ~x0 & n595;
  assign n597 = ~n592 & ~n596;
  assign n598 = ~x45 & n506;
  assign n599 = x1 & n598;
  assign n600 = ~x45 & n594;
  assign n601 = x0 & n600;
  assign n602 = ~n599 & ~n601;
  assign n603 = n597 & n602;
  assign n619 = n618 ^ n603;
  assign n582 = ~x11 & n82;
  assign n583 = ~x10 & n86;
  assign n584 = ~n582 & ~n583;
  assign n585 = x11 & n89;
  assign n586 = x10 & n91;
  assign n587 = ~n585 & ~n586;
  assign n588 = n584 & n587;
  assign n575 = x7 & n217;
  assign n576 = x6 & n219;
  assign n577 = ~n575 & ~n576;
  assign n578 = ~x7 & n210;
  assign n579 = ~x6 & n214;
  assign n580 = ~n578 & ~n579;
  assign n581 = n577 & n580;
  assign n589 = n588 ^ n581;
  assign n568 = x5 & n336;
  assign n569 = x4 & n338;
  assign n570 = ~n568 & ~n569;
  assign n571 = ~x5 & n329;
  assign n572 = ~x4 & n333;
  assign n573 = ~n571 & ~n572;
  assign n574 = n570 & n573;
  assign n590 = n589 ^ n574;
  assign n620 = n619 ^ n590;
  assign n624 = n623 ^ n620;
  assign n647 = n646 ^ n624;
  assign n651 = n650 ^ n647;
  assign n655 = n654 ^ n651;
  assign n733 = n654 ^ n647;
  assign n734 = ~n651 & ~n733;
  assign n735 = n734 ^ n654;
  assign n729 = n645 ^ n624;
  assign n730 = n646 & n729;
  assign n731 = n730 ^ n642;
  assign n725 = n623 ^ n619;
  assign n726 = n620 & ~n725;
  assign n727 = n726 ^ n590;
  assign n720 = n641 ^ n637;
  assign n721 = n638 & ~n720;
  assign n722 = n721 ^ n633;
  assign n710 = x2 & n598;
  assign n711 = x1 & n600;
  assign n712 = ~n710 & ~n711;
  assign n713 = ~x2 & n591;
  assign n714 = ~x1 & n595;
  assign n715 = ~n713 & ~n714;
  assign n716 = n712 & n715;
  assign n703 = x4 & n430;
  assign n704 = x3 & n434;
  assign n705 = ~n703 & ~n704;
  assign n706 = ~x4 & n437;
  assign n707 = ~x3 & n439;
  assign n708 = ~n706 & ~n707;
  assign n709 = n705 & n708;
  assign n717 = n716 ^ n709;
  assign n702 = n628 & n632;
  assign n718 = n717 ^ n702;
  assign n693 = ~x6 & n329;
  assign n694 = ~x5 & n333;
  assign n695 = ~n693 & ~n694;
  assign n696 = x6 & n336;
  assign n697 = x5 & n338;
  assign n698 = ~n696 & ~n697;
  assign n699 = n695 & n698;
  assign n686 = x8 & n217;
  assign n687 = x7 & n219;
  assign n688 = ~n686 & ~n687;
  assign n689 = ~x8 & n210;
  assign n690 = ~x7 & n214;
  assign n691 = ~n689 & ~n690;
  assign n692 = n688 & n691;
  assign n700 = n699 ^ n692;
  assign n679 = x10 & n153;
  assign n680 = x9 & n155;
  assign n681 = ~n679 & ~n680;
  assign n682 = ~x10 & n146;
  assign n683 = ~x9 & n150;
  assign n684 = ~n682 & ~n683;
  assign n685 = n681 & n684;
  assign n701 = n700 ^ n685;
  assign n719 = n718 ^ n701;
  assign n723 = n722 ^ n719;
  assign n674 = n617 ^ n603;
  assign n675 = n618 & ~n674;
  assign n676 = n675 ^ n610;
  assign n671 = n588 ^ n574;
  assign n672 = n589 & ~n671;
  assign n673 = n672 ^ n581;
  assign n677 = n676 ^ n673;
  assign n663 = ~x12 & n82;
  assign n664 = ~x11 & n86;
  assign n665 = ~n663 & ~n664;
  assign n666 = x12 & n89;
  assign n667 = x11 & n91;
  assign n668 = ~n666 & ~n667;
  assign n669 = n665 & n668;
  assign n659 = x33 ^ x14;
  assign n660 = x32 & n659;
  assign n658 = ~x13 & n68;
  assign n661 = n660 ^ n658;
  assign n656 = x46 ^ x45;
  assign n657 = x0 & n656;
  assign n662 = n661 ^ n657;
  assign n670 = n669 ^ n662;
  assign n678 = n677 ^ n670;
  assign n724 = n723 ^ n678;
  assign n728 = n727 ^ n724;
  assign n732 = n731 ^ n728;
  assign n736 = n735 ^ n732;
  assign n833 = n735 ^ n728;
  assign n834 = n732 & ~n833;
  assign n835 = n834 ^ n735;
  assign n829 = n727 ^ n723;
  assign n830 = n724 & ~n829;
  assign n831 = n830 ^ n678;
  assign n824 = n722 ^ n718;
  assign n825 = ~n719 & ~n824;
  assign n826 = n825 ^ n701;
  assign n818 = n692 ^ n685;
  assign n819 = n699 ^ n685;
  assign n820 = n818 & ~n819;
  assign n821 = n820 ^ n692;
  assign n809 = ~x11 & n146;
  assign n810 = ~x10 & n150;
  assign n811 = ~n809 & ~n810;
  assign n812 = x11 & n153;
  assign n813 = x10 & n155;
  assign n814 = ~n812 & ~n813;
  assign n815 = n811 & n814;
  assign n802 = ~x7 & n329;
  assign n803 = ~x6 & n333;
  assign n804 = ~n802 & ~n803;
  assign n805 = x7 & n336;
  assign n806 = x6 & n338;
  assign n807 = ~n805 & ~n806;
  assign n808 = n804 & n807;
  assign n816 = n815 ^ n808;
  assign n795 = x5 & n430;
  assign n796 = x4 & n434;
  assign n797 = ~n795 & ~n796;
  assign n798 = ~x5 & n437;
  assign n799 = ~x4 & n439;
  assign n800 = ~n798 & ~n799;
  assign n801 = n797 & n800;
  assign n817 = n816 ^ n801;
  assign n822 = n821 ^ n817;
  assign n780 = ~x47 & n656;
  assign n781 = x1 & n780;
  assign n782 = x47 ^ x46;
  assign n783 = ~n656 & n782;
  assign n784 = ~x47 & n783;
  assign n785 = x0 & n784;
  assign n786 = ~n781 & ~n785;
  assign n787 = x47 & n656;
  assign n788 = ~x1 & n787;
  assign n789 = x47 & n783;
  assign n790 = ~x0 & n789;
  assign n791 = ~n788 & ~n790;
  assign n792 = n786 & n791;
  assign n773 = ~x13 & n82;
  assign n774 = ~x12 & n86;
  assign n775 = ~n773 & ~n774;
  assign n776 = x13 & n89;
  assign n777 = x12 & n91;
  assign n778 = ~n776 & ~n777;
  assign n779 = n775 & n778;
  assign n793 = n792 ^ n779;
  assign n766 = x9 & n217;
  assign n767 = x8 & n219;
  assign n768 = ~n766 & ~n767;
  assign n769 = ~x9 & n210;
  assign n770 = ~x8 & n214;
  assign n771 = ~n769 & ~n770;
  assign n772 = n768 & n771;
  assign n794 = n793 ^ n772;
  assign n823 = n822 ^ n794;
  assign n827 = n826 ^ n823;
  assign n762 = n673 ^ n670;
  assign n763 = ~n677 & n762;
  assign n764 = n763 ^ n670;
  assign n758 = n716 ^ n702;
  assign n759 = n717 & n758;
  assign n760 = n759 ^ n709;
  assign n754 = n669 ^ n661;
  assign n755 = n662 & n754;
  assign n756 = n755 ^ n657;
  assign n748 = x45 ^ x0;
  assign n749 = ~n656 & n748;
  assign n750 = n749 ^ x0;
  assign n751 = x47 & ~n750;
  assign n746 = ~x14 & n68;
  assign n744 = x33 ^ x15;
  assign n745 = x32 & n744;
  assign n747 = n746 ^ n745;
  assign n752 = n751 ^ n747;
  assign n737 = ~x3 & n591;
  assign n738 = ~x2 & n595;
  assign n739 = ~n737 & ~n738;
  assign n740 = x3 & n598;
  assign n741 = x2 & n600;
  assign n742 = ~n740 & ~n741;
  assign n743 = n739 & n742;
  assign n753 = n752 ^ n743;
  assign n757 = n756 ^ n753;
  assign n761 = n760 ^ n757;
  assign n765 = n764 ^ n761;
  assign n828 = n827 ^ n765;
  assign n832 = n831 ^ n828;
  assign n836 = n835 ^ n832;
  assign n929 = n835 ^ n828;
  assign n930 = ~n832 & ~n929;
  assign n931 = n930 ^ n835;
  assign n924 = n823 ^ n765;
  assign n925 = n826 ^ n765;
  assign n926 = n924 & ~n925;
  assign n927 = n926 ^ n823;
  assign n919 = n764 ^ n760;
  assign n920 = n761 & ~n919;
  assign n921 = n920 ^ n757;
  assign n908 = ~x6 & n437;
  assign n909 = ~x5 & n439;
  assign n910 = ~n908 & ~n909;
  assign n911 = x6 & n430;
  assign n912 = x5 & n434;
  assign n913 = ~n911 & ~n912;
  assign n914 = n910 & n913;
  assign n901 = x12 & n153;
  assign n902 = x11 & n155;
  assign n903 = ~n901 & ~n902;
  assign n904 = ~x12 & n146;
  assign n905 = ~x11 & n150;
  assign n906 = ~n904 & ~n905;
  assign n907 = n903 & n906;
  assign n915 = n914 ^ n907;
  assign n894 = x4 & n598;
  assign n895 = x3 & n600;
  assign n896 = ~n894 & ~n895;
  assign n897 = ~x4 & n591;
  assign n898 = ~x3 & n595;
  assign n899 = ~n897 & ~n898;
  assign n900 = n896 & n899;
  assign n916 = n915 ^ n900;
  assign n886 = ~x14 & n82;
  assign n887 = ~x13 & n86;
  assign n888 = ~n886 & ~n887;
  assign n889 = x14 & n89;
  assign n890 = x13 & n91;
  assign n891 = ~n889 & ~n890;
  assign n892 = n888 & n891;
  assign n882 = x33 ^ x16;
  assign n883 = x32 & n882;
  assign n881 = ~x15 & n68;
  assign n884 = n883 ^ n881;
  assign n879 = x48 ^ x47;
  assign n880 = x0 & n879;
  assign n885 = n884 ^ n880;
  assign n893 = n892 ^ n885;
  assign n917 = n916 ^ n893;
  assign n870 = x10 & n217;
  assign n871 = x9 & n219;
  assign n872 = ~n870 & ~n871;
  assign n873 = ~x10 & n210;
  assign n874 = ~x9 & n214;
  assign n875 = ~n873 & ~n874;
  assign n876 = n872 & n875;
  assign n863 = ~x2 & n787;
  assign n864 = ~x1 & n789;
  assign n865 = ~n863 & ~n864;
  assign n866 = x2 & n780;
  assign n867 = x1 & n784;
  assign n868 = ~n866 & ~n867;
  assign n869 = n865 & n868;
  assign n877 = n876 ^ n869;
  assign n856 = x8 & n336;
  assign n857 = x7 & n338;
  assign n858 = ~n856 & ~n857;
  assign n859 = ~x8 & n329;
  assign n860 = ~x7 & n333;
  assign n861 = ~n859 & ~n860;
  assign n862 = n858 & n861;
  assign n878 = n877 ^ n862;
  assign n918 = n917 ^ n878;
  assign n922 = n921 ^ n918;
  assign n851 = n817 ^ n794;
  assign n852 = n821 ^ n794;
  assign n853 = n851 & ~n852;
  assign n854 = n853 ^ n817;
  assign n847 = n756 ^ n752;
  assign n848 = ~n753 & ~n847;
  assign n849 = n848 ^ n743;
  assign n842 = n808 ^ n801;
  assign n843 = n815 ^ n801;
  assign n844 = n842 & ~n843;
  assign n845 = n844 ^ n808;
  assign n838 = n792 ^ n772;
  assign n839 = n793 & ~n838;
  assign n840 = n839 ^ n779;
  assign n837 = n747 & n751;
  assign n841 = n840 ^ n837;
  assign n846 = n845 ^ n841;
  assign n850 = n849 ^ n846;
  assign n855 = n854 ^ n850;
  assign n923 = n922 ^ n855;
  assign n928 = n927 ^ n923;
  assign n932 = n931 ^ n928;
  assign n1041 = n931 ^ n923;
  assign n1042 = n928 & n1041;
  assign n1043 = n1042 ^ n931;
  assign n1036 = n918 ^ n855;
  assign n1037 = n921 ^ n855;
  assign n1038 = ~n1036 & n1037;
  assign n1039 = n1038 ^ n918;
  assign n1031 = n854 ^ n849;
  assign n1032 = ~n850 & ~n1031;
  assign n1033 = n1032 ^ n846;
  assign n1020 = ~x11 & n210;
  assign n1021 = ~x10 & n214;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = x11 & n217;
  assign n1024 = x10 & n219;
  assign n1025 = ~n1023 & ~n1024;
  assign n1026 = n1022 & n1025;
  assign n1013 = ~x3 & n787;
  assign n1014 = ~x2 & n789;
  assign n1015 = ~n1013 & ~n1014;
  assign n1016 = x3 & n780;
  assign n1017 = x2 & n784;
  assign n1018 = ~n1016 & ~n1017;
  assign n1019 = n1015 & n1018;
  assign n1027 = n1026 ^ n1019;
  assign n1000 = x49 & n879;
  assign n1001 = ~x1 & n1000;
  assign n1002 = x49 ^ x48;
  assign n1003 = ~n879 & n1002;
  assign n1004 = x49 & n1003;
  assign n1005 = ~x0 & n1004;
  assign n1006 = ~n1001 & ~n1005;
  assign n1007 = ~x49 & n879;
  assign n1008 = x1 & n1007;
  assign n1009 = ~x49 & n1003;
  assign n1010 = x0 & n1009;
  assign n1011 = ~n1008 & ~n1010;
  assign n1012 = n1006 & n1011;
  assign n1028 = n1027 ^ n1012;
  assign n991 = x9 & n336;
  assign n992 = x8 & n338;
  assign n993 = ~n991 & ~n992;
  assign n994 = ~x9 & n329;
  assign n995 = ~x8 & n333;
  assign n996 = ~n994 & ~n995;
  assign n997 = n993 & n996;
  assign n984 = x15 & n89;
  assign n985 = x14 & n91;
  assign n986 = ~n984 & ~n985;
  assign n987 = ~x15 & n82;
  assign n988 = ~x14 & n86;
  assign n989 = ~n987 & ~n988;
  assign n990 = n986 & n989;
  assign n998 = n997 ^ n990;
  assign n977 = ~x13 & n146;
  assign n978 = ~x12 & n150;
  assign n979 = ~n977 & ~n978;
  assign n980 = x13 & n153;
  assign n981 = x12 & n155;
  assign n982 = ~n980 & ~n981;
  assign n983 = n979 & n982;
  assign n999 = n998 ^ n983;
  assign n1029 = n1028 ^ n999;
  assign n968 = ~x7 & n437;
  assign n969 = ~x6 & n439;
  assign n970 = ~n968 & ~n969;
  assign n971 = x7 & n430;
  assign n972 = x6 & n434;
  assign n973 = ~n971 & ~n972;
  assign n974 = n970 & n973;
  assign n961 = x5 & n598;
  assign n962 = x4 & n600;
  assign n963 = ~n961 & ~n962;
  assign n964 = ~x5 & n591;
  assign n965 = ~x4 & n595;
  assign n966 = ~n964 & ~n965;
  assign n967 = n963 & n966;
  assign n975 = n974 ^ n967;
  assign n956 = x47 ^ x0;
  assign n957 = ~n879 & n956;
  assign n958 = n957 ^ x0;
  assign n959 = x49 & ~n958;
  assign n954 = ~x16 & n68;
  assign n952 = x33 ^ x17;
  assign n953 = x32 & n952;
  assign n955 = n954 ^ n953;
  assign n960 = n959 ^ n955;
  assign n976 = n975 ^ n960;
  assign n1030 = n1029 ^ n976;
  assign n1034 = n1033 ^ n1030;
  assign n948 = n916 ^ n878;
  assign n949 = n917 & ~n948;
  assign n950 = n949 ^ n893;
  assign n944 = n845 ^ n840;
  assign n945 = ~n841 & ~n944;
  assign n946 = n945 ^ n837;
  assign n940 = n876 ^ n862;
  assign n941 = n877 & ~n940;
  assign n942 = n941 ^ n869;
  assign n936 = n907 ^ n900;
  assign n937 = ~n915 & n936;
  assign n938 = n937 ^ n900;
  assign n933 = n892 ^ n884;
  assign n934 = n885 & n933;
  assign n935 = n934 ^ n880;
  assign n939 = n938 ^ n935;
  assign n943 = n942 ^ n939;
  assign n947 = n946 ^ n943;
  assign n951 = n950 ^ n947;
  assign n1035 = n1034 ^ n951;
  assign n1040 = n1039 ^ n1035;
  assign n1044 = n1043 ^ n1040;
  assign n1147 = n1043 ^ n1035;
  assign n1148 = ~n1040 & ~n1147;
  assign n1149 = n1148 ^ n1043;
  assign n1142 = n1030 ^ n951;
  assign n1143 = n1033 ^ n951;
  assign n1144 = ~n1142 & n1143;
  assign n1145 = n1144 ^ n1030;
  assign n1137 = n950 ^ n943;
  assign n1138 = ~n947 & ~n1137;
  assign n1139 = n1138 ^ n950;
  assign n1132 = n974 ^ n960;
  assign n1133 = n975 & n1132;
  assign n1134 = n1133 ^ n967;
  assign n1123 = x2 & n1007;
  assign n1124 = x1 & n1009;
  assign n1125 = ~n1123 & ~n1124;
  assign n1126 = ~x2 & n1000;
  assign n1127 = ~x1 & n1004;
  assign n1128 = ~n1126 & ~n1127;
  assign n1129 = n1125 & n1128;
  assign n1116 = x4 & n780;
  assign n1117 = x3 & n784;
  assign n1118 = ~n1116 & ~n1117;
  assign n1119 = ~x4 & n787;
  assign n1120 = ~x3 & n789;
  assign n1121 = ~n1119 & ~n1120;
  assign n1122 = n1118 & n1121;
  assign n1130 = n1129 ^ n1122;
  assign n1109 = ~x16 & n82;
  assign n1110 = ~x15 & n86;
  assign n1111 = ~n1109 & ~n1110;
  assign n1112 = x16 & n89;
  assign n1113 = x15 & n91;
  assign n1114 = ~n1112 & ~n1113;
  assign n1115 = n1111 & n1114;
  assign n1131 = n1130 ^ n1115;
  assign n1135 = n1134 ^ n1131;
  assign n1105 = n1019 ^ n1012;
  assign n1106 = ~n1027 & n1105;
  assign n1107 = n1106 ^ n1012;
  assign n1103 = n955 & n959;
  assign n1096 = x6 & n598;
  assign n1097 = x5 & n600;
  assign n1098 = ~n1096 & ~n1097;
  assign n1099 = ~x6 & n591;
  assign n1100 = ~x5 & n595;
  assign n1101 = ~n1099 & ~n1100;
  assign n1102 = n1098 & n1101;
  assign n1104 = n1103 ^ n1102;
  assign n1108 = n1107 ^ n1104;
  assign n1136 = n1135 ^ n1108;
  assign n1140 = n1139 ^ n1136;
  assign n1091 = n942 ^ n938;
  assign n1092 = ~n939 & ~n1091;
  assign n1093 = n1092 ^ n935;
  assign n1088 = n999 ^ n976;
  assign n1089 = ~n1029 & ~n1088;
  assign n1090 = n1089 ^ n976;
  assign n1094 = n1093 ^ n1090;
  assign n1083 = n997 ^ n983;
  assign n1084 = n998 & ~n1083;
  assign n1085 = n1084 ^ n990;
  assign n1074 = ~x14 & n146;
  assign n1075 = ~x13 & n150;
  assign n1076 = ~n1074 & ~n1075;
  assign n1077 = x14 & n153;
  assign n1078 = x13 & n155;
  assign n1079 = ~n1077 & ~n1078;
  assign n1080 = n1076 & n1079;
  assign n1067 = ~x10 & n329;
  assign n1068 = ~x9 & n333;
  assign n1069 = ~n1067 & ~n1068;
  assign n1070 = x10 & n336;
  assign n1071 = x9 & n338;
  assign n1072 = ~n1070 & ~n1071;
  assign n1073 = n1069 & n1072;
  assign n1081 = n1080 ^ n1073;
  assign n1060 = ~x8 & n437;
  assign n1061 = ~x7 & n439;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = x8 & n430;
  assign n1064 = x7 & n434;
  assign n1065 = ~n1063 & ~n1064;
  assign n1066 = n1062 & n1065;
  assign n1082 = n1081 ^ n1066;
  assign n1086 = n1085 ^ n1082;
  assign n1052 = ~x12 & n210;
  assign n1053 = ~x11 & n214;
  assign n1054 = ~n1052 & ~n1053;
  assign n1055 = x12 & n217;
  assign n1056 = x11 & n219;
  assign n1057 = ~n1055 & ~n1056;
  assign n1058 = n1054 & n1057;
  assign n1048 = x33 ^ x18;
  assign n1049 = x32 & n1048;
  assign n1047 = ~x17 & n68;
  assign n1050 = n1049 ^ n1047;
  assign n1045 = x50 ^ x49;
  assign n1046 = x0 & n1045;
  assign n1051 = n1050 ^ n1046;
  assign n1059 = n1058 ^ n1051;
  assign n1087 = n1086 ^ n1059;
  assign n1095 = n1094 ^ n1087;
  assign n1141 = n1140 ^ n1095;
  assign n1146 = n1145 ^ n1141;
  assign n1150 = n1149 ^ n1146;
  assign n1271 = n1149 ^ n1141;
  assign n1272 = ~n1146 & n1271;
  assign n1273 = n1272 ^ n1149;
  assign n1266 = n1136 ^ n1095;
  assign n1267 = n1139 ^ n1095;
  assign n1268 = ~n1266 & ~n1267;
  assign n1269 = n1268 ^ n1136;
  assign n1261 = n1090 ^ n1087;
  assign n1262 = ~n1094 & ~n1261;
  assign n1263 = n1262 ^ n1087;
  assign n1256 = n1107 ^ n1103;
  assign n1257 = ~n1104 & n1256;
  assign n1258 = n1257 ^ n1102;
  assign n1247 = x17 & n89;
  assign n1248 = x16 & n91;
  assign n1249 = ~n1247 & ~n1248;
  assign n1250 = ~x17 & n82;
  assign n1251 = ~x16 & n86;
  assign n1252 = ~n1250 & ~n1251;
  assign n1253 = n1249 & n1252;
  assign n1234 = ~x51 & n1045;
  assign n1235 = x1 & n1234;
  assign n1236 = x51 ^ x50;
  assign n1237 = ~n1045 & n1236;
  assign n1238 = ~x51 & n1237;
  assign n1239 = x0 & n1238;
  assign n1240 = ~n1235 & ~n1239;
  assign n1241 = x51 & n1045;
  assign n1242 = ~x1 & n1241;
  assign n1243 = x51 & n1237;
  assign n1244 = ~x0 & n1243;
  assign n1245 = ~n1242 & ~n1244;
  assign n1246 = n1240 & n1245;
  assign n1254 = n1253 ^ n1246;
  assign n1227 = x11 & n336;
  assign n1228 = x10 & n338;
  assign n1229 = ~n1227 & ~n1228;
  assign n1230 = ~x11 & n329;
  assign n1231 = ~x10 & n333;
  assign n1232 = ~n1230 & ~n1231;
  assign n1233 = n1229 & n1232;
  assign n1255 = n1254 ^ n1233;
  assign n1259 = n1258 ^ n1255;
  assign n1223 = n1122 ^ n1115;
  assign n1224 = ~n1130 & n1223;
  assign n1225 = n1224 ^ n1115;
  assign n1219 = n1058 ^ n1050;
  assign n1220 = n1051 & n1219;
  assign n1221 = n1220 ^ n1046;
  assign n1214 = x49 ^ x0;
  assign n1215 = ~n1045 & n1214;
  assign n1216 = n1215 ^ x0;
  assign n1217 = x51 & ~n1216;
  assign n1212 = ~x18 & n68;
  assign n1210 = x33 ^ x19;
  assign n1211 = x32 & n1210;
  assign n1213 = n1212 ^ n1211;
  assign n1218 = n1217 ^ n1213;
  assign n1222 = n1221 ^ n1218;
  assign n1226 = n1225 ^ n1222;
  assign n1260 = n1259 ^ n1226;
  assign n1264 = n1263 ^ n1260;
  assign n1206 = n1134 ^ n1108;
  assign n1207 = n1135 & n1206;
  assign n1208 = n1207 ^ n1131;
  assign n1202 = n1082 ^ n1059;
  assign n1203 = ~n1086 & n1202;
  assign n1204 = n1203 ^ n1059;
  assign n1197 = n1073 ^ n1066;
  assign n1198 = ~n1081 & n1197;
  assign n1199 = n1198 ^ n1066;
  assign n1188 = ~x9 & n437;
  assign n1189 = ~x8 & n439;
  assign n1190 = ~n1188 & ~n1189;
  assign n1191 = x9 & n430;
  assign n1192 = x8 & n434;
  assign n1193 = ~n1191 & ~n1192;
  assign n1194 = n1190 & n1193;
  assign n1181 = ~x15 & n146;
  assign n1182 = ~x14 & n150;
  assign n1183 = ~n1181 & ~n1182;
  assign n1184 = x15 & n153;
  assign n1185 = x14 & n155;
  assign n1186 = ~n1184 & ~n1185;
  assign n1187 = n1183 & n1186;
  assign n1195 = n1194 ^ n1187;
  assign n1174 = ~x7 & n591;
  assign n1175 = ~x6 & n595;
  assign n1176 = ~n1174 & ~n1175;
  assign n1177 = x7 & n598;
  assign n1178 = x6 & n600;
  assign n1179 = ~n1177 & ~n1178;
  assign n1180 = n1176 & n1179;
  assign n1196 = n1195 ^ n1180;
  assign n1200 = n1199 ^ n1196;
  assign n1165 = x5 & n780;
  assign n1166 = x4 & n784;
  assign n1167 = ~n1165 & ~n1166;
  assign n1168 = ~x5 & n787;
  assign n1169 = ~x4 & n789;
  assign n1170 = ~n1168 & ~n1169;
  assign n1171 = n1167 & n1170;
  assign n1158 = x13 & n217;
  assign n1159 = x12 & n219;
  assign n1160 = ~n1158 & ~n1159;
  assign n1161 = ~x13 & n210;
  assign n1162 = ~x12 & n214;
  assign n1163 = ~n1161 & ~n1162;
  assign n1164 = n1160 & n1163;
  assign n1172 = n1171 ^ n1164;
  assign n1151 = ~x3 & n1000;
  assign n1152 = ~x2 & n1004;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = x3 & n1007;
  assign n1155 = x2 & n1009;
  assign n1156 = ~n1154 & ~n1155;
  assign n1157 = n1153 & n1156;
  assign n1173 = n1172 ^ n1157;
  assign n1201 = n1200 ^ n1173;
  assign n1205 = n1204 ^ n1201;
  assign n1209 = n1208 ^ n1205;
  assign n1265 = n1264 ^ n1209;
  assign n1270 = n1269 ^ n1265;
  assign n1274 = n1273 ^ n1270;
  assign n1392 = n1273 ^ n1265;
  assign n1393 = n1270 & ~n1392;
  assign n1394 = n1393 ^ n1273;
  assign n1387 = n1260 ^ n1209;
  assign n1388 = n1263 ^ n1209;
  assign n1389 = n1387 & ~n1388;
  assign n1390 = n1389 ^ n1260;
  assign n1381 = n1208 ^ n1201;
  assign n1382 = n1208 ^ n1204;
  assign n1383 = n1381 & ~n1382;
  assign n1384 = n1383 ^ n1201;
  assign n1377 = n1255 ^ n1226;
  assign n1378 = n1258 ^ n1226;
  assign n1379 = n1377 & ~n1378;
  assign n1380 = n1379 ^ n1255;
  assign n1385 = n1384 ^ n1380;
  assign n1371 = n1196 ^ n1173;
  assign n1372 = n1199 ^ n1173;
  assign n1373 = n1371 & ~n1372;
  assign n1374 = n1373 ^ n1196;
  assign n1367 = n1225 ^ n1221;
  assign n1368 = n1222 & n1367;
  assign n1369 = n1368 ^ n1218;
  assign n1358 = ~x8 & n591;
  assign n1359 = ~x7 & n595;
  assign n1360 = ~n1358 & ~n1359;
  assign n1361 = x8 & n598;
  assign n1362 = x7 & n600;
  assign n1363 = ~n1361 & ~n1362;
  assign n1364 = n1360 & n1363;
  assign n1351 = ~x10 & n437;
  assign n1352 = ~x9 & n439;
  assign n1353 = ~n1351 & ~n1352;
  assign n1354 = x10 & n430;
  assign n1355 = x9 & n434;
  assign n1356 = ~n1354 & ~n1355;
  assign n1357 = n1353 & n1356;
  assign n1365 = n1364 ^ n1357;
  assign n1350 = n1213 & n1217;
  assign n1366 = n1365 ^ n1350;
  assign n1370 = n1369 ^ n1366;
  assign n1375 = n1374 ^ n1370;
  assign n1345 = n1246 ^ n1233;
  assign n1346 = ~n1254 & n1345;
  assign n1347 = n1346 ^ n1233;
  assign n1341 = n1171 ^ n1157;
  assign n1342 = n1172 & ~n1341;
  assign n1343 = n1342 ^ n1164;
  assign n1338 = n1194 ^ n1180;
  assign n1339 = n1195 & ~n1338;
  assign n1340 = n1339 ^ n1187;
  assign n1344 = n1343 ^ n1340;
  assign n1348 = n1347 ^ n1344;
  assign n1327 = ~x6 & n787;
  assign n1328 = ~x5 & n789;
  assign n1329 = ~n1327 & ~n1328;
  assign n1330 = x6 & n780;
  assign n1331 = x5 & n784;
  assign n1332 = ~n1330 & ~n1331;
  assign n1333 = n1329 & n1332;
  assign n1320 = ~x4 & n1000;
  assign n1321 = ~x3 & n1004;
  assign n1322 = ~n1320 & ~n1321;
  assign n1323 = x4 & n1007;
  assign n1324 = x3 & n1009;
  assign n1325 = ~n1323 & ~n1324;
  assign n1326 = n1322 & n1325;
  assign n1334 = n1333 ^ n1326;
  assign n1313 = ~x18 & n82;
  assign n1314 = ~x17 & n86;
  assign n1315 = ~n1313 & ~n1314;
  assign n1316 = x18 & n89;
  assign n1317 = x17 & n91;
  assign n1318 = ~n1316 & ~n1317;
  assign n1319 = n1315 & n1318;
  assign n1335 = n1334 ^ n1319;
  assign n1305 = ~x14 & n210;
  assign n1306 = ~x13 & n214;
  assign n1307 = ~n1305 & ~n1306;
  assign n1308 = x14 & n217;
  assign n1309 = x13 & n219;
  assign n1310 = ~n1308 & ~n1309;
  assign n1311 = n1307 & n1310;
  assign n1301 = x33 ^ x20;
  assign n1302 = x32 & n1301;
  assign n1300 = ~x19 & n68;
  assign n1303 = n1302 ^ n1300;
  assign n1298 = x52 ^ x51;
  assign n1299 = x0 & n1298;
  assign n1304 = n1303 ^ n1299;
  assign n1312 = n1311 ^ n1304;
  assign n1336 = n1335 ^ n1312;
  assign n1289 = ~x12 & n329;
  assign n1290 = ~x11 & n333;
  assign n1291 = ~n1289 & ~n1290;
  assign n1292 = x12 & n336;
  assign n1293 = x11 & n338;
  assign n1294 = ~n1292 & ~n1293;
  assign n1295 = n1291 & n1294;
  assign n1282 = ~x2 & n1241;
  assign n1283 = ~x1 & n1243;
  assign n1284 = ~n1282 & ~n1283;
  assign n1285 = x2 & n1234;
  assign n1286 = x1 & n1238;
  assign n1287 = ~n1285 & ~n1286;
  assign n1288 = n1284 & n1287;
  assign n1296 = n1295 ^ n1288;
  assign n1275 = x16 & n153;
  assign n1276 = x15 & n155;
  assign n1277 = ~n1275 & ~n1276;
  assign n1278 = ~x16 & n146;
  assign n1279 = ~x15 & n150;
  assign n1280 = ~n1278 & ~n1279;
  assign n1281 = n1277 & n1280;
  assign n1297 = n1296 ^ n1281;
  assign n1337 = n1336 ^ n1297;
  assign n1349 = n1348 ^ n1337;
  assign n1376 = n1375 ^ n1349;
  assign n1386 = n1385 ^ n1376;
  assign n1391 = n1390 ^ n1386;
  assign n1395 = n1394 ^ n1391;
  assign n1529 = n1394 ^ n1386;
  assign n1530 = ~n1391 & ~n1529;
  assign n1531 = n1530 ^ n1394;
  assign n1525 = n1380 ^ n1376;
  assign n1526 = ~n1385 & n1525;
  assign n1527 = n1526 ^ n1376;
  assign n1521 = n1375 ^ n1348;
  assign n1522 = n1349 & ~n1521;
  assign n1523 = n1522 ^ n1337;
  assign n1516 = n1374 ^ n1366;
  assign n1517 = n1374 ^ n1369;
  assign n1518 = ~n1516 & n1517;
  assign n1519 = n1518 ^ n1366;
  assign n1510 = n1347 ^ n1343;
  assign n1511 = n1344 & ~n1510;
  assign n1512 = n1511 ^ n1340;
  assign n1505 = n1326 ^ n1319;
  assign n1506 = n1333 ^ n1319;
  assign n1507 = n1505 & ~n1506;
  assign n1508 = n1507 ^ n1326;
  assign n1496 = x19 & n89;
  assign n1497 = x18 & n91;
  assign n1498 = ~n1496 & ~n1497;
  assign n1499 = ~x19 & n82;
  assign n1500 = ~x18 & n86;
  assign n1501 = ~n1499 & ~n1500;
  assign n1502 = n1498 & n1501;
  assign n1492 = x51 ^ x0;
  assign n1493 = ~n1298 & n1492;
  assign n1494 = n1493 ^ x0;
  assign n1495 = x53 & ~n1494;
  assign n1503 = n1502 ^ n1495;
  assign n1485 = x9 & n598;
  assign n1486 = x8 & n600;
  assign n1487 = ~n1485 & ~n1486;
  assign n1488 = ~x9 & n591;
  assign n1489 = ~x8 & n595;
  assign n1490 = ~n1488 & ~n1489;
  assign n1491 = n1487 & n1490;
  assign n1504 = n1503 ^ n1491;
  assign n1509 = n1508 ^ n1504;
  assign n1513 = n1512 ^ n1509;
  assign n1480 = n1295 ^ n1281;
  assign n1481 = n1296 & ~n1480;
  assign n1482 = n1481 ^ n1288;
  assign n1477 = n1311 ^ n1303;
  assign n1478 = n1304 & n1477;
  assign n1479 = n1478 ^ n1299;
  assign n1483 = n1482 ^ n1479;
  assign n1472 = x33 ^ x21;
  assign n1473 = x32 & n1472;
  assign n1471 = ~x20 & n68;
  assign n1474 = n1473 ^ n1471;
  assign n1464 = ~x17 & n146;
  assign n1465 = ~x16 & n150;
  assign n1466 = ~n1464 & ~n1465;
  assign n1467 = x17 & n153;
  assign n1468 = x16 & n155;
  assign n1469 = ~n1467 & ~n1468;
  assign n1470 = n1466 & n1469;
  assign n1475 = n1474 ^ n1470;
  assign n1457 = ~x11 & n437;
  assign n1458 = ~x10 & n439;
  assign n1459 = ~n1457 & ~n1458;
  assign n1460 = x11 & n430;
  assign n1461 = x10 & n434;
  assign n1462 = ~n1460 & ~n1461;
  assign n1463 = n1459 & n1462;
  assign n1476 = n1475 ^ n1463;
  assign n1484 = n1483 ^ n1476;
  assign n1514 = n1513 ^ n1484;
  assign n1453 = n1335 ^ n1297;
  assign n1454 = n1336 & ~n1453;
  assign n1455 = n1454 ^ n1312;
  assign n1449 = n1364 ^ n1350;
  assign n1450 = n1365 & n1449;
  assign n1451 = n1450 ^ n1357;
  assign n1439 = ~x15 & n210;
  assign n1440 = ~x14 & n214;
  assign n1441 = ~n1439 & ~n1440;
  assign n1442 = x15 & n217;
  assign n1443 = x14 & n219;
  assign n1444 = ~n1442 & ~n1443;
  assign n1445 = n1441 & n1444;
  assign n1432 = x7 & n780;
  assign n1433 = x6 & n784;
  assign n1434 = ~n1432 & ~n1433;
  assign n1435 = ~x7 & n787;
  assign n1436 = ~x6 & n789;
  assign n1437 = ~n1435 & ~n1436;
  assign n1438 = n1434 & n1437;
  assign n1446 = n1445 ^ n1438;
  assign n1425 = ~x5 & n1000;
  assign n1426 = ~x4 & n1004;
  assign n1427 = ~n1425 & ~n1426;
  assign n1428 = x5 & n1007;
  assign n1429 = x4 & n1009;
  assign n1430 = ~n1428 & ~n1429;
  assign n1431 = n1427 & n1430;
  assign n1447 = n1446 ^ n1431;
  assign n1416 = x3 & n1234;
  assign n1417 = x2 & n1238;
  assign n1418 = ~n1416 & ~n1417;
  assign n1419 = ~x3 & n1241;
  assign n1420 = ~x2 & n1243;
  assign n1421 = ~n1419 & ~n1420;
  assign n1422 = n1418 & n1421;
  assign n1409 = ~x13 & n329;
  assign n1410 = ~x12 & n333;
  assign n1411 = ~n1409 & ~n1410;
  assign n1412 = x13 & n336;
  assign n1413 = x12 & n338;
  assign n1414 = ~n1412 & ~n1413;
  assign n1415 = n1411 & n1414;
  assign n1423 = n1422 ^ n1415;
  assign n1396 = x53 & n1298;
  assign n1397 = ~x1 & n1396;
  assign n1398 = x53 ^ x52;
  assign n1399 = ~n1298 & n1398;
  assign n1400 = x53 & n1399;
  assign n1401 = ~x0 & n1400;
  assign n1402 = ~n1397 & ~n1401;
  assign n1403 = ~x53 & n1298;
  assign n1404 = x1 & n1403;
  assign n1405 = ~x53 & n1399;
  assign n1406 = x0 & n1405;
  assign n1407 = ~n1404 & ~n1406;
  assign n1408 = n1402 & n1407;
  assign n1424 = n1423 ^ n1408;
  assign n1448 = n1447 ^ n1424;
  assign n1452 = n1451 ^ n1448;
  assign n1456 = n1455 ^ n1452;
  assign n1515 = n1514 ^ n1456;
  assign n1520 = n1519 ^ n1515;
  assign n1524 = n1523 ^ n1520;
  assign n1528 = n1527 ^ n1524;
  assign n1532 = n1531 ^ n1528;
  assign n1660 = n1531 ^ n1524;
  assign n1661 = n1528 & n1660;
  assign n1662 = n1661 ^ n1531;
  assign n1655 = n1523 ^ n1515;
  assign n1656 = n1523 ^ n1519;
  assign n1657 = n1655 & n1656;
  assign n1658 = n1657 ^ n1515;
  assign n1651 = n1514 ^ n1452;
  assign n1652 = n1456 & ~n1651;
  assign n1653 = n1652 ^ n1455;
  assign n1645 = n1509 ^ n1484;
  assign n1646 = n1512 ^ n1484;
  assign n1647 = n1645 & ~n1646;
  assign n1648 = n1647 ^ n1509;
  assign n1640 = n1508 ^ n1503;
  assign n1641 = n1504 & ~n1640;
  assign n1642 = n1641 ^ n1491;
  assign n1630 = x2 & n1403;
  assign n1631 = x1 & n1405;
  assign n1632 = ~n1630 & ~n1631;
  assign n1633 = ~x2 & n1396;
  assign n1634 = ~x1 & n1400;
  assign n1635 = ~n1633 & ~n1634;
  assign n1636 = n1632 & n1635;
  assign n1623 = x4 & n1234;
  assign n1624 = x3 & n1238;
  assign n1625 = ~n1623 & ~n1624;
  assign n1626 = ~x4 & n1241;
  assign n1627 = ~x3 & n1243;
  assign n1628 = ~n1626 & ~n1627;
  assign n1629 = n1625 & n1628;
  assign n1637 = n1636 ^ n1629;
  assign n1621 = ~x21 & n68;
  assign n1619 = x33 ^ x22;
  assign n1620 = x32 & n1619;
  assign n1622 = n1621 ^ n1620;
  assign n1638 = n1637 ^ n1622;
  assign n1610 = x20 & n89;
  assign n1611 = x19 & n91;
  assign n1612 = ~n1610 & ~n1611;
  assign n1613 = ~x20 & n82;
  assign n1614 = ~x19 & n86;
  assign n1615 = ~n1613 & ~n1614;
  assign n1616 = n1612 & n1615;
  assign n1608 = x54 ^ x53;
  assign n1609 = x0 & n1608;
  assign n1617 = n1616 ^ n1609;
  assign n1601 = ~x16 & n210;
  assign n1602 = ~x15 & n214;
  assign n1603 = ~n1601 & ~n1602;
  assign n1604 = x16 & n217;
  assign n1605 = x15 & n219;
  assign n1606 = ~n1604 & ~n1605;
  assign n1607 = n1603 & n1606;
  assign n1618 = n1617 ^ n1607;
  assign n1639 = n1638 ^ n1618;
  assign n1643 = n1642 ^ n1639;
  assign n1596 = n1445 ^ n1431;
  assign n1597 = n1446 & ~n1596;
  assign n1598 = n1597 ^ n1438;
  assign n1587 = ~x12 & n437;
  assign n1588 = ~x11 & n439;
  assign n1589 = ~n1587 & ~n1588;
  assign n1590 = x12 & n430;
  assign n1591 = x11 & n434;
  assign n1592 = ~n1590 & ~n1591;
  assign n1593 = n1589 & n1592;
  assign n1580 = ~x18 & n146;
  assign n1581 = ~x17 & n150;
  assign n1582 = ~n1580 & ~n1581;
  assign n1583 = x18 & n153;
  assign n1584 = x17 & n155;
  assign n1585 = ~n1583 & ~n1584;
  assign n1586 = n1582 & n1585;
  assign n1594 = n1593 ^ n1586;
  assign n1573 = ~x10 & n591;
  assign n1574 = ~x9 & n595;
  assign n1575 = ~n1573 & ~n1574;
  assign n1576 = x10 & n598;
  assign n1577 = x9 & n600;
  assign n1578 = ~n1576 & ~n1577;
  assign n1579 = n1575 & n1578;
  assign n1595 = n1594 ^ n1579;
  assign n1599 = n1598 ^ n1595;
  assign n1564 = ~x6 & n1000;
  assign n1565 = ~x5 & n1004;
  assign n1566 = ~n1564 & ~n1565;
  assign n1567 = x6 & n1007;
  assign n1568 = x5 & n1009;
  assign n1569 = ~n1567 & ~n1568;
  assign n1570 = n1566 & n1569;
  assign n1557 = x8 & n780;
  assign n1558 = x7 & n784;
  assign n1559 = ~n1557 & ~n1558;
  assign n1560 = ~x8 & n787;
  assign n1561 = ~x7 & n789;
  assign n1562 = ~n1560 & ~n1561;
  assign n1563 = n1559 & n1562;
  assign n1571 = n1570 ^ n1563;
  assign n1550 = x14 & n336;
  assign n1551 = x13 & n338;
  assign n1552 = ~n1550 & ~n1551;
  assign n1553 = ~x14 & n329;
  assign n1554 = ~x13 & n333;
  assign n1555 = ~n1553 & ~n1554;
  assign n1556 = n1552 & n1555;
  assign n1572 = n1571 ^ n1556;
  assign n1600 = n1599 ^ n1572;
  assign n1644 = n1643 ^ n1600;
  assign n1649 = n1648 ^ n1644;
  assign n1546 = n1451 ^ n1447;
  assign n1547 = n1448 & ~n1546;
  assign n1548 = n1547 ^ n1424;
  assign n1542 = n1479 ^ n1476;
  assign n1543 = n1483 & n1542;
  assign n1544 = n1543 ^ n1476;
  assign n1538 = n1415 ^ n1408;
  assign n1539 = ~n1423 & n1538;
  assign n1540 = n1539 ^ n1408;
  assign n1534 = n1470 ^ n1463;
  assign n1535 = ~n1475 & ~n1534;
  assign n1536 = n1535 ^ n1474;
  assign n1533 = n1495 & ~n1502;
  assign n1537 = n1536 ^ n1533;
  assign n1541 = n1540 ^ n1537;
  assign n1545 = n1544 ^ n1541;
  assign n1549 = n1548 ^ n1545;
  assign n1650 = n1649 ^ n1549;
  assign n1654 = n1653 ^ n1650;
  assign n1659 = n1658 ^ n1654;
  assign n1663 = n1662 ^ n1659;
  assign n1809 = n1662 ^ n1654;
  assign n1810 = n1659 & n1809;
  assign n1811 = n1810 ^ n1662;
  assign n1805 = n1653 ^ n1649;
  assign n1806 = ~n1650 & ~n1805;
  assign n1807 = n1806 ^ n1549;
  assign n1800 = n1648 ^ n1643;
  assign n1801 = n1644 & ~n1800;
  assign n1802 = n1801 ^ n1600;
  assign n1797 = n1548 ^ n1544;
  assign n1798 = ~n1545 & n1797;
  assign n1799 = n1798 ^ n1541;
  assign n1803 = n1802 ^ n1799;
  assign n1792 = n1642 ^ n1638;
  assign n1793 = n1639 & n1792;
  assign n1794 = n1793 ^ n1618;
  assign n1788 = n1540 ^ n1536;
  assign n1789 = n1537 & n1788;
  assign n1790 = n1789 ^ n1533;
  assign n1778 = x9 & n780;
  assign n1779 = x8 & n784;
  assign n1780 = ~n1778 & ~n1779;
  assign n1781 = ~x9 & n787;
  assign n1782 = ~x8 & n789;
  assign n1783 = ~n1781 & ~n1782;
  assign n1784 = n1780 & n1783;
  assign n1771 = ~x17 & n210;
  assign n1772 = ~x16 & n214;
  assign n1773 = ~n1771 & ~n1772;
  assign n1774 = x17 & n217;
  assign n1775 = x16 & n219;
  assign n1776 = ~n1774 & ~n1775;
  assign n1777 = n1773 & n1776;
  assign n1785 = n1784 ^ n1777;
  assign n1764 = ~x7 & n1000;
  assign n1765 = ~x6 & n1004;
  assign n1766 = ~n1764 & ~n1765;
  assign n1767 = x7 & n1007;
  assign n1768 = x6 & n1009;
  assign n1769 = ~n1767 & ~n1768;
  assign n1770 = n1766 & n1769;
  assign n1786 = n1785 ^ n1770;
  assign n1755 = ~x21 & n82;
  assign n1756 = ~x20 & n86;
  assign n1757 = ~n1755 & ~n1756;
  assign n1758 = x21 & n89;
  assign n1759 = x20 & n91;
  assign n1760 = ~n1758 & ~n1759;
  assign n1761 = n1757 & n1760;
  assign n1751 = x53 ^ x0;
  assign n1752 = ~n1608 & n1751;
  assign n1753 = n1752 ^ x0;
  assign n1754 = x55 & ~n1753;
  assign n1762 = n1761 ^ n1754;
  assign n1743 = ~x11 & n591;
  assign n1744 = ~x10 & n595;
  assign n1745 = ~n1743 & ~n1744;
  assign n1746 = x11 & n598;
  assign n1747 = x10 & n600;
  assign n1748 = ~n1746 & ~n1747;
  assign n1749 = n1745 & n1748;
  assign n1736 = ~x13 & n437;
  assign n1737 = ~x12 & n439;
  assign n1738 = ~n1736 & ~n1737;
  assign n1739 = x13 & n430;
  assign n1740 = x12 & n434;
  assign n1741 = ~n1739 & ~n1740;
  assign n1742 = n1738 & n1741;
  assign n1750 = n1749 ^ n1742;
  assign n1763 = n1762 ^ n1750;
  assign n1787 = n1786 ^ n1763;
  assign n1791 = n1790 ^ n1787;
  assign n1795 = n1794 ^ n1791;
  assign n1730 = n1595 ^ n1572;
  assign n1731 = n1598 ^ n1572;
  assign n1732 = n1730 & ~n1731;
  assign n1733 = n1732 ^ n1595;
  assign n1725 = n1609 ^ n1607;
  assign n1726 = n1616 ^ n1607;
  assign n1727 = ~n1725 & ~n1726;
  assign n1728 = n1727 ^ n1609;
  assign n1721 = n1629 ^ n1622;
  assign n1722 = ~n1637 & ~n1721;
  assign n1723 = n1722 ^ n1622;
  assign n1718 = n1593 ^ n1579;
  assign n1719 = n1594 & ~n1718;
  assign n1720 = n1719 ^ n1586;
  assign n1724 = n1723 ^ n1720;
  assign n1729 = n1728 ^ n1724;
  assign n1734 = n1733 ^ n1729;
  assign n1713 = n1563 ^ n1556;
  assign n1714 = ~n1571 & n1713;
  assign n1715 = n1714 ^ n1556;
  assign n1708 = x33 ^ x23;
  assign n1709 = x32 & n1708;
  assign n1707 = ~x22 & n68;
  assign n1710 = n1709 ^ n1707;
  assign n1700 = x19 & n153;
  assign n1701 = x18 & n155;
  assign n1702 = ~n1700 & ~n1701;
  assign n1703 = ~x19 & n146;
  assign n1704 = ~x18 & n150;
  assign n1705 = ~n1703 & ~n1704;
  assign n1706 = n1702 & n1705;
  assign n1711 = n1710 ^ n1706;
  assign n1687 = x55 & n1608;
  assign n1688 = ~x1 & n1687;
  assign n1689 = x55 ^ x54;
  assign n1690 = ~n1608 & n1689;
  assign n1691 = x55 & n1690;
  assign n1692 = ~x0 & n1691;
  assign n1693 = ~n1688 & ~n1692;
  assign n1694 = ~x55 & n1608;
  assign n1695 = x1 & n1694;
  assign n1696 = ~x55 & n1690;
  assign n1697 = x0 & n1696;
  assign n1698 = ~n1695 & ~n1697;
  assign n1699 = n1693 & n1698;
  assign n1712 = n1711 ^ n1699;
  assign n1716 = n1715 ^ n1712;
  assign n1678 = x5 & n1234;
  assign n1679 = x4 & n1238;
  assign n1680 = ~n1678 & ~n1679;
  assign n1681 = ~x5 & n1241;
  assign n1682 = ~x4 & n1243;
  assign n1683 = ~n1681 & ~n1682;
  assign n1684 = n1680 & n1683;
  assign n1671 = x15 & n336;
  assign n1672 = x14 & n338;
  assign n1673 = ~n1671 & ~n1672;
  assign n1674 = ~x15 & n329;
  assign n1675 = ~x14 & n333;
  assign n1676 = ~n1674 & ~n1675;
  assign n1677 = n1673 & n1676;
  assign n1685 = n1684 ^ n1677;
  assign n1664 = ~x3 & n1396;
  assign n1665 = ~x2 & n1400;
  assign n1666 = ~n1664 & ~n1665;
  assign n1667 = x3 & n1403;
  assign n1668 = x2 & n1405;
  assign n1669 = ~n1667 & ~n1668;
  assign n1670 = n1666 & n1669;
  assign n1686 = n1685 ^ n1670;
  assign n1717 = n1716 ^ n1686;
  assign n1735 = n1734 ^ n1717;
  assign n1796 = n1795 ^ n1735;
  assign n1804 = n1803 ^ n1796;
  assign n1808 = n1807 ^ n1804;
  assign n1812 = n1811 ^ n1808;
  assign n1951 = n1811 ^ n1804;
  assign n1952 = ~n1808 & n1951;
  assign n1953 = n1952 ^ n1811;
  assign n1947 = n1799 ^ n1796;
  assign n1948 = ~n1803 & ~n1947;
  assign n1949 = n1948 ^ n1796;
  assign n1942 = n1791 ^ n1735;
  assign n1943 = n1794 ^ n1735;
  assign n1944 = n1942 & ~n1943;
  assign n1945 = n1944 ^ n1791;
  assign n1937 = n1729 ^ n1717;
  assign n1938 = ~n1734 & ~n1937;
  assign n1939 = n1938 ^ n1717;
  assign n1933 = n1790 ^ n1786;
  assign n1934 = n1787 & n1933;
  assign n1935 = n1934 ^ n1763;
  assign n1928 = n1728 ^ n1720;
  assign n1929 = n1724 & ~n1928;
  assign n1930 = n1929 ^ n1728;
  assign n1925 = n1762 ^ n1749;
  assign n1926 = n1750 & ~n1925;
  assign n1927 = n1926 ^ n1742;
  assign n1931 = n1930 ^ n1927;
  assign n1921 = n1677 ^ n1670;
  assign n1922 = ~n1685 & n1921;
  assign n1923 = n1922 ^ n1670;
  assign n1919 = n1754 & ~n1761;
  assign n1912 = ~x12 & n591;
  assign n1913 = ~x11 & n595;
  assign n1914 = ~n1912 & ~n1913;
  assign n1915 = x12 & n598;
  assign n1916 = x11 & n600;
  assign n1917 = ~n1915 & ~n1916;
  assign n1918 = n1914 & n1917;
  assign n1920 = n1919 ^ n1918;
  assign n1924 = n1923 ^ n1920;
  assign n1932 = n1931 ^ n1924;
  assign n1936 = n1935 ^ n1932;
  assign n1940 = n1939 ^ n1936;
  assign n1907 = n1712 ^ n1686;
  assign n1908 = n1716 & ~n1907;
  assign n1909 = n1908 ^ n1686;
  assign n1902 = n1777 ^ n1770;
  assign n1903 = ~n1785 & n1902;
  assign n1904 = n1903 ^ n1770;
  assign n1899 = n1706 ^ n1699;
  assign n1900 = ~n1711 & ~n1899;
  assign n1901 = n1900 ^ n1710;
  assign n1905 = n1904 ^ n1901;
  assign n1890 = ~x20 & n146;
  assign n1891 = ~x19 & n150;
  assign n1892 = ~n1890 & ~n1891;
  assign n1893 = x20 & n153;
  assign n1894 = x19 & n155;
  assign n1895 = ~n1893 & ~n1894;
  assign n1896 = n1892 & n1895;
  assign n1883 = ~x2 & n1687;
  assign n1884 = ~x1 & n1691;
  assign n1885 = ~n1883 & ~n1884;
  assign n1886 = x2 & n1694;
  assign n1887 = x1 & n1696;
  assign n1888 = ~n1886 & ~n1887;
  assign n1889 = n1885 & n1888;
  assign n1897 = n1896 ^ n1889;
  assign n1876 = ~x14 & n437;
  assign n1877 = ~x13 & n439;
  assign n1878 = ~n1876 & ~n1877;
  assign n1879 = x14 & n430;
  assign n1880 = x13 & n434;
  assign n1881 = ~n1879 & ~n1880;
  assign n1882 = n1878 & n1881;
  assign n1898 = n1897 ^ n1882;
  assign n1906 = n1905 ^ n1898;
  assign n1910 = n1909 ^ n1906;
  assign n1865 = ~x4 & n1396;
  assign n1866 = ~x3 & n1400;
  assign n1867 = ~n1865 & ~n1866;
  assign n1868 = x4 & n1403;
  assign n1869 = x3 & n1405;
  assign n1870 = ~n1868 & ~n1869;
  assign n1871 = n1867 & n1870;
  assign n1858 = ~x6 & n1241;
  assign n1859 = ~x5 & n1243;
  assign n1860 = ~n1858 & ~n1859;
  assign n1861 = x6 & n1234;
  assign n1862 = x5 & n1238;
  assign n1863 = ~n1861 & ~n1862;
  assign n1864 = n1860 & n1863;
  assign n1872 = n1871 ^ n1864;
  assign n1856 = ~x23 & n68;
  assign n1854 = x33 ^ x24;
  assign n1855 = x32 & n1854;
  assign n1857 = n1856 ^ n1855;
  assign n1873 = n1872 ^ n1857;
  assign n1845 = ~x22 & n82;
  assign n1846 = ~x21 & n86;
  assign n1847 = ~n1845 & ~n1846;
  assign n1848 = x22 & n89;
  assign n1849 = x21 & n91;
  assign n1850 = ~n1848 & ~n1849;
  assign n1851 = n1847 & n1850;
  assign n1843 = x56 ^ x55;
  assign n1844 = x0 & n1843;
  assign n1852 = n1851 ^ n1844;
  assign n1836 = ~x18 & n210;
  assign n1837 = ~x17 & n214;
  assign n1838 = ~n1836 & ~n1837;
  assign n1839 = x18 & n217;
  assign n1840 = x17 & n219;
  assign n1841 = ~n1839 & ~n1840;
  assign n1842 = n1838 & n1841;
  assign n1853 = n1852 ^ n1842;
  assign n1874 = n1873 ^ n1853;
  assign n1827 = x10 & n780;
  assign n1828 = x9 & n784;
  assign n1829 = ~n1827 & ~n1828;
  assign n1830 = ~x10 & n787;
  assign n1831 = ~x9 & n789;
  assign n1832 = ~n1830 & ~n1831;
  assign n1833 = n1829 & n1832;
  assign n1820 = x8 & n1007;
  assign n1821 = x7 & n1009;
  assign n1822 = ~n1820 & ~n1821;
  assign n1823 = ~x8 & n1000;
  assign n1824 = ~x7 & n1004;
  assign n1825 = ~n1823 & ~n1824;
  assign n1826 = n1822 & n1825;
  assign n1834 = n1833 ^ n1826;
  assign n1813 = ~x16 & n329;
  assign n1814 = ~x15 & n333;
  assign n1815 = ~n1813 & ~n1814;
  assign n1816 = x16 & n336;
  assign n1817 = x15 & n338;
  assign n1818 = ~n1816 & ~n1817;
  assign n1819 = n1815 & n1818;
  assign n1835 = n1834 ^ n1819;
  assign n1875 = n1874 ^ n1835;
  assign n1911 = n1910 ^ n1875;
  assign n1941 = n1940 ^ n1911;
  assign n1946 = n1945 ^ n1941;
  assign n1950 = n1949 ^ n1946;
  assign n1954 = n1953 ^ n1950;
  assign n2114 = n1953 ^ n1946;
  assign n2115 = ~n1950 & n2114;
  assign n2116 = n2115 ^ n1953;
  assign n2110 = n1945 ^ n1940;
  assign n2111 = n1941 & ~n2110;
  assign n2112 = n2111 ^ n1911;
  assign n2105 = n1939 ^ n1935;
  assign n2106 = n1936 & n2105;
  assign n2107 = n2106 ^ n1932;
  assign n2100 = n1901 ^ n1898;
  assign n2101 = n1905 & ~n2100;
  assign n2102 = n2101 ^ n1898;
  assign n2096 = n1864 ^ n1857;
  assign n2097 = ~n1872 & ~n2096;
  assign n2098 = n2097 ^ n1857;
  assign n2091 = n1826 ^ n1819;
  assign n2092 = n1833 ^ n1819;
  assign n2093 = n2091 & ~n2092;
  assign n2094 = n2093 ^ n1826;
  assign n2083 = x23 & n89;
  assign n2084 = x22 & n91;
  assign n2085 = ~n2083 & ~n2084;
  assign n2086 = ~x23 & n82;
  assign n2087 = ~x22 & n86;
  assign n2088 = ~n2086 & ~n2087;
  assign n2089 = n2085 & n2088;
  assign n2079 = x55 ^ x0;
  assign n2080 = ~n1843 & n2079;
  assign n2081 = n2080 ^ x0;
  assign n2082 = x57 & ~n2081;
  assign n2090 = n2089 ^ n2082;
  assign n2095 = n2094 ^ n2090;
  assign n2099 = n2098 ^ n2095;
  assign n2103 = n2102 ^ n2099;
  assign n2068 = x7 & n1234;
  assign n2069 = x6 & n1238;
  assign n2070 = ~n2068 & ~n2069;
  assign n2071 = ~x7 & n1241;
  assign n2072 = ~x6 & n1243;
  assign n2073 = ~n2071 & ~n2072;
  assign n2074 = n2070 & n2073;
  assign n2061 = ~x17 & n329;
  assign n2062 = ~x16 & n333;
  assign n2063 = ~n2061 & ~n2062;
  assign n2064 = x17 & n336;
  assign n2065 = x16 & n338;
  assign n2066 = ~n2064 & ~n2065;
  assign n2067 = n2063 & n2066;
  assign n2075 = n2074 ^ n2067;
  assign n2054 = x5 & n1403;
  assign n2055 = x4 & n1405;
  assign n2056 = ~n2054 & ~n2055;
  assign n2057 = ~x5 & n1396;
  assign n2058 = ~x4 & n1400;
  assign n2059 = ~n2057 & ~n2058;
  assign n2060 = n2056 & n2059;
  assign n2076 = n2075 ^ n2060;
  assign n2045 = ~x11 & n787;
  assign n2046 = ~x10 & n789;
  assign n2047 = ~n2045 & ~n2046;
  assign n2048 = x11 & n780;
  assign n2049 = x10 & n784;
  assign n2050 = ~n2048 & ~n2049;
  assign n2051 = n2047 & n2050;
  assign n2038 = ~x19 & n210;
  assign n2039 = ~x18 & n214;
  assign n2040 = ~n2038 & ~n2039;
  assign n2041 = x19 & n217;
  assign n2042 = x18 & n219;
  assign n2043 = ~n2041 & ~n2042;
  assign n2044 = n2040 & n2043;
  assign n2052 = n2051 ^ n2044;
  assign n2031 = ~x9 & n1000;
  assign n2032 = ~x8 & n1004;
  assign n2033 = ~n2031 & ~n2032;
  assign n2034 = x9 & n1007;
  assign n2035 = x8 & n1009;
  assign n2036 = ~n2034 & ~n2035;
  assign n2037 = n2033 & n2036;
  assign n2053 = n2052 ^ n2037;
  assign n2077 = n2076 ^ n2053;
  assign n2026 = x33 ^ x25;
  assign n2027 = x32 & n2026;
  assign n2025 = ~x24 & n68;
  assign n2028 = n2027 ^ n2025;
  assign n2018 = x15 & n430;
  assign n2019 = x14 & n434;
  assign n2020 = ~n2018 & ~n2019;
  assign n2021 = ~x15 & n437;
  assign n2022 = ~x14 & n439;
  assign n2023 = ~n2021 & ~n2022;
  assign n2024 = n2020 & n2023;
  assign n2029 = n2028 ^ n2024;
  assign n2011 = x3 & n1694;
  assign n2012 = x2 & n1696;
  assign n2013 = ~n2011 & ~n2012;
  assign n2014 = ~x3 & n1687;
  assign n2015 = ~x2 & n1691;
  assign n2016 = ~n2014 & ~n2015;
  assign n2017 = n2013 & n2016;
  assign n2030 = n2029 ^ n2017;
  assign n2078 = n2077 ^ n2030;
  assign n2104 = n2103 ^ n2078;
  assign n2108 = n2107 ^ n2104;
  assign n2005 = n1927 ^ n1924;
  assign n2006 = n1930 ^ n1924;
  assign n2007 = ~n2005 & ~n2006;
  assign n2008 = n2007 ^ n1927;
  assign n2002 = n1906 ^ n1875;
  assign n2003 = n1910 & ~n2002;
  assign n2004 = n2003 ^ n1875;
  assign n2009 = n2008 ^ n2004;
  assign n1997 = n1853 ^ n1835;
  assign n1998 = n1873 ^ n1835;
  assign n1999 = ~n1997 & n1998;
  assign n2000 = n1999 ^ n1853;
  assign n1993 = n1923 ^ n1919;
  assign n1994 = ~n1920 & n1993;
  assign n1995 = n1994 ^ n1918;
  assign n1987 = n1889 ^ n1882;
  assign n1988 = n1896 ^ n1882;
  assign n1989 = n1987 & ~n1988;
  assign n1990 = n1989 ^ n1889;
  assign n1984 = n1851 ^ n1842;
  assign n1985 = ~n1852 & ~n1984;
  assign n1986 = n1985 ^ n1844;
  assign n1991 = n1990 ^ n1986;
  assign n1975 = ~x21 & n146;
  assign n1976 = ~x20 & n150;
  assign n1977 = ~n1975 & ~n1976;
  assign n1978 = x21 & n153;
  assign n1979 = x20 & n155;
  assign n1980 = ~n1978 & ~n1979;
  assign n1981 = n1977 & n1980;
  assign n1962 = x57 & n1843;
  assign n1963 = ~x1 & n1962;
  assign n1964 = x57 ^ x56;
  assign n1965 = ~n1843 & n1964;
  assign n1966 = x57 & n1965;
  assign n1967 = ~x0 & n1966;
  assign n1968 = ~n1963 & ~n1967;
  assign n1969 = ~x57 & n1843;
  assign n1970 = x1 & n1969;
  assign n1971 = ~x57 & n1965;
  assign n1972 = x0 & n1971;
  assign n1973 = ~n1970 & ~n1972;
  assign n1974 = n1968 & n1973;
  assign n1982 = n1981 ^ n1974;
  assign n1955 = ~x13 & n591;
  assign n1956 = ~x12 & n595;
  assign n1957 = ~n1955 & ~n1956;
  assign n1958 = x13 & n598;
  assign n1959 = x12 & n600;
  assign n1960 = ~n1958 & ~n1959;
  assign n1961 = n1957 & n1960;
  assign n1983 = n1982 ^ n1961;
  assign n1992 = n1991 ^ n1983;
  assign n1996 = n1995 ^ n1992;
  assign n2001 = n2000 ^ n1996;
  assign n2010 = n2009 ^ n2001;
  assign n2109 = n2108 ^ n2010;
  assign n2113 = n2112 ^ n2109;
  assign n2117 = n2116 ^ n2113;
  assign n2271 = n2116 ^ n2109;
  assign n2272 = n2113 & ~n2271;
  assign n2273 = n2272 ^ n2116;
  assign n2266 = n2104 ^ n2010;
  assign n2267 = n2107 ^ n2010;
  assign n2268 = n2266 & ~n2267;
  assign n2269 = n2268 ^ n2104;
  assign n2261 = n2004 ^ n2001;
  assign n2262 = ~n2009 & n2261;
  assign n2263 = n2262 ^ n2001;
  assign n2254 = n2028 ^ n2017;
  assign n2255 = n2024 ^ n2017;
  assign n2256 = ~n2254 & ~n2255;
  assign n2257 = n2256 ^ n2028;
  assign n2249 = n2067 ^ n2060;
  assign n2250 = n2074 ^ n2060;
  assign n2251 = n2249 & ~n2250;
  assign n2252 = n2251 ^ n2067;
  assign n2246 = n2051 ^ n2037;
  assign n2247 = n2052 & ~n2246;
  assign n2248 = n2247 ^ n2044;
  assign n2253 = n2252 ^ n2248;
  assign n2258 = n2257 ^ n2253;
  assign n2243 = n2082 & ~n2089;
  assign n2235 = ~x14 & n591;
  assign n2236 = ~x13 & n595;
  assign n2237 = ~n2235 & ~n2236;
  assign n2238 = x14 & n598;
  assign n2239 = x13 & n600;
  assign n2240 = ~n2238 & ~n2239;
  assign n2241 = n2237 & n2240;
  assign n2228 = x22 & n153;
  assign n2229 = x21 & n155;
  assign n2230 = ~n2228 & ~n2229;
  assign n2231 = ~x22 & n146;
  assign n2232 = ~x21 & n150;
  assign n2233 = ~n2231 & ~n2232;
  assign n2234 = n2230 & n2233;
  assign n2242 = n2241 ^ n2234;
  assign n2244 = n2243 ^ n2242;
  assign n2218 = ~x16 & n437;
  assign n2219 = ~x15 & n439;
  assign n2220 = ~n2218 & ~n2219;
  assign n2221 = x16 & n430;
  assign n2222 = x15 & n434;
  assign n2223 = ~n2221 & ~n2222;
  assign n2224 = n2220 & n2223;
  assign n2211 = ~x4 & n1687;
  assign n2212 = ~x3 & n1691;
  assign n2213 = ~n2211 & ~n2212;
  assign n2214 = x4 & n1694;
  assign n2215 = x3 & n1696;
  assign n2216 = ~n2214 & ~n2215;
  assign n2217 = n2213 & n2216;
  assign n2225 = n2224 ^ n2217;
  assign n2204 = ~x2 & n1962;
  assign n2205 = ~x1 & n1966;
  assign n2206 = ~n2204 & ~n2205;
  assign n2207 = x2 & n1969;
  assign n2208 = x1 & n1971;
  assign n2209 = ~n2207 & ~n2208;
  assign n2210 = n2206 & n2209;
  assign n2226 = n2225 ^ n2210;
  assign n2195 = x12 & n780;
  assign n2196 = x11 & n784;
  assign n2197 = ~n2195 & ~n2196;
  assign n2198 = ~x12 & n787;
  assign n2199 = ~x11 & n789;
  assign n2200 = ~n2198 & ~n2199;
  assign n2201 = n2197 & n2200;
  assign n2188 = x10 & n1007;
  assign n2189 = x9 & n1009;
  assign n2190 = ~n2188 & ~n2189;
  assign n2191 = ~x10 & n1000;
  assign n2192 = ~x9 & n1004;
  assign n2193 = ~n2191 & ~n2192;
  assign n2194 = n2190 & n2193;
  assign n2202 = n2201 ^ n2194;
  assign n2181 = ~x18 & n329;
  assign n2182 = ~x17 & n333;
  assign n2183 = ~n2181 & ~n2182;
  assign n2184 = x18 & n336;
  assign n2185 = x17 & n338;
  assign n2186 = ~n2184 & ~n2185;
  assign n2187 = n2183 & n2186;
  assign n2203 = n2202 ^ n2187;
  assign n2227 = n2226 ^ n2203;
  assign n2245 = n2244 ^ n2227;
  assign n2259 = n2258 ^ n2245;
  assign n2176 = n1981 ^ n1961;
  assign n2177 = n1982 & ~n2176;
  assign n2178 = n2177 ^ n1974;
  assign n2167 = ~x24 & n82;
  assign n2168 = ~x23 & n86;
  assign n2169 = ~n2167 & ~n2168;
  assign n2170 = x24 & n89;
  assign n2171 = x23 & n91;
  assign n2172 = ~n2170 & ~n2171;
  assign n2173 = n2169 & n2172;
  assign n2165 = x58 ^ x57;
  assign n2166 = x0 & n2165;
  assign n2174 = n2173 ^ n2166;
  assign n2158 = ~x20 & n210;
  assign n2159 = ~x19 & n214;
  assign n2160 = ~n2158 & ~n2159;
  assign n2161 = x20 & n217;
  assign n2162 = x19 & n219;
  assign n2163 = ~n2161 & ~n2162;
  assign n2164 = n2160 & n2163;
  assign n2175 = n2174 ^ n2164;
  assign n2179 = n2178 ^ n2175;
  assign n2149 = ~x8 & n1241;
  assign n2150 = ~x7 & n1243;
  assign n2151 = ~n2149 & ~n2150;
  assign n2152 = x8 & n1234;
  assign n2153 = x7 & n1238;
  assign n2154 = ~n2152 & ~n2153;
  assign n2155 = n2151 & n2154;
  assign n2142 = ~x6 & n1396;
  assign n2143 = ~x5 & n1400;
  assign n2144 = ~n2142 & ~n2143;
  assign n2145 = x6 & n1403;
  assign n2146 = x5 & n1405;
  assign n2147 = ~n2145 & ~n2146;
  assign n2148 = n2144 & n2147;
  assign n2156 = n2155 ^ n2148;
  assign n2140 = ~x25 & n68;
  assign n2138 = x33 ^ x26;
  assign n2139 = x32 & n2138;
  assign n2141 = n2140 ^ n2139;
  assign n2157 = n2156 ^ n2141;
  assign n2180 = n2179 ^ n2157;
  assign n2260 = n2259 ^ n2180;
  assign n2264 = n2263 ^ n2260;
  assign n2134 = n2099 ^ n2078;
  assign n2135 = n2103 & n2134;
  assign n2136 = n2135 ^ n2078;
  assign n2129 = n2000 ^ n1992;
  assign n2130 = n2000 ^ n1995;
  assign n2131 = n2129 & n2130;
  assign n2132 = n2131 ^ n1992;
  assign n2125 = n2076 ^ n2030;
  assign n2126 = n2077 & n2125;
  assign n2127 = n2126 ^ n2053;
  assign n2121 = n1986 ^ n1983;
  assign n2122 = n1991 & ~n2121;
  assign n2123 = n2122 ^ n1983;
  assign n2118 = n2098 ^ n2094;
  assign n2119 = n2095 & n2118;
  assign n2120 = n2119 ^ n2090;
  assign n2124 = n2123 ^ n2120;
  assign n2128 = n2127 ^ n2124;
  assign n2133 = n2132 ^ n2128;
  assign n2137 = n2136 ^ n2133;
  assign n2265 = n2264 ^ n2137;
  assign n2270 = n2269 ^ n2265;
  assign n2274 = n2273 ^ n2270;
  assign n2445 = n2273 ^ n2265;
  assign n2446 = ~n2270 & ~n2445;
  assign n2447 = n2446 ^ n2273;
  assign n2440 = n2260 ^ n2137;
  assign n2441 = n2263 ^ n2137;
  assign n2442 = n2440 & ~n2441;
  assign n2443 = n2442 ^ n2260;
  assign n2435 = n2136 ^ n2132;
  assign n2436 = ~n2133 & ~n2435;
  assign n2437 = n2436 ^ n2128;
  assign n2430 = n2244 ^ n2226;
  assign n2431 = n2227 & n2430;
  assign n2432 = n2431 ^ n2203;
  assign n2419 = x23 & n153;
  assign n2420 = x22 & n155;
  assign n2421 = ~n2419 & ~n2420;
  assign n2422 = ~x23 & n146;
  assign n2423 = ~x22 & n150;
  assign n2424 = ~n2422 & ~n2423;
  assign n2425 = n2421 & n2424;
  assign n2412 = x3 & n1969;
  assign n2413 = x2 & n1971;
  assign n2414 = ~n2412 & ~n2413;
  assign n2415 = ~x3 & n1962;
  assign n2416 = ~x2 & n1966;
  assign n2417 = ~n2415 & ~n2416;
  assign n2418 = n2414 & n2417;
  assign n2426 = n2425 ^ n2418;
  assign n2399 = ~x59 & n2165;
  assign n2400 = x1 & n2399;
  assign n2401 = x59 ^ x58;
  assign n2402 = ~n2165 & n2401;
  assign n2403 = ~x59 & n2402;
  assign n2404 = x0 & n2403;
  assign n2405 = ~n2400 & ~n2404;
  assign n2406 = x59 & n2165;
  assign n2407 = ~x1 & n2406;
  assign n2408 = x59 & n2402;
  assign n2409 = ~x0 & n2408;
  assign n2410 = ~n2407 & ~n2409;
  assign n2411 = n2405 & n2410;
  assign n2427 = n2426 ^ n2411;
  assign n2390 = ~x13 & n787;
  assign n2391 = ~x12 & n789;
  assign n2392 = ~n2390 & ~n2391;
  assign n2393 = x13 & n780;
  assign n2394 = x12 & n784;
  assign n2395 = ~n2393 & ~n2394;
  assign n2396 = n2392 & n2395;
  assign n2383 = x21 & n217;
  assign n2384 = x20 & n219;
  assign n2385 = ~n2383 & ~n2384;
  assign n2386 = ~x21 & n210;
  assign n2387 = ~x20 & n214;
  assign n2388 = ~n2386 & ~n2387;
  assign n2389 = n2385 & n2388;
  assign n2397 = n2396 ^ n2389;
  assign n2376 = ~x11 & n1000;
  assign n2377 = ~x10 & n1004;
  assign n2378 = ~n2376 & ~n2377;
  assign n2379 = x11 & n1007;
  assign n2380 = x10 & n1009;
  assign n2381 = ~n2379 & ~n2380;
  assign n2382 = n2378 & n2381;
  assign n2398 = n2397 ^ n2382;
  assign n2428 = n2427 ^ n2398;
  assign n2371 = x33 ^ x27;
  assign n2372 = x32 & n2371;
  assign n2370 = ~x26 & n68;
  assign n2373 = n2372 ^ n2370;
  assign n2363 = ~x17 & n437;
  assign n2364 = ~x16 & n439;
  assign n2365 = ~n2363 & ~n2364;
  assign n2366 = x17 & n430;
  assign n2367 = x16 & n434;
  assign n2368 = ~n2366 & ~n2367;
  assign n2369 = n2365 & n2368;
  assign n2374 = n2373 ^ n2369;
  assign n2356 = ~x5 & n1687;
  assign n2357 = ~x4 & n1691;
  assign n2358 = ~n2356 & ~n2357;
  assign n2359 = x5 & n1694;
  assign n2360 = x4 & n1696;
  assign n2361 = ~n2359 & ~n2360;
  assign n2362 = n2358 & n2361;
  assign n2375 = n2374 ^ n2362;
  assign n2429 = n2428 ^ n2375;
  assign n2433 = n2432 ^ n2429;
  assign n2351 = n2243 ^ n2241;
  assign n2352 = n2242 & n2351;
  assign n2353 = n2352 ^ n2234;
  assign n2342 = ~x9 & n1241;
  assign n2343 = ~x8 & n1243;
  assign n2344 = ~n2342 & ~n2343;
  assign n2345 = x9 & n1234;
  assign n2346 = x8 & n1238;
  assign n2347 = ~n2345 & ~n2346;
  assign n2348 = n2344 & n2347;
  assign n2335 = x19 & n336;
  assign n2336 = x18 & n338;
  assign n2337 = ~n2335 & ~n2336;
  assign n2338 = ~x19 & n329;
  assign n2339 = ~x18 & n333;
  assign n2340 = ~n2338 & ~n2339;
  assign n2341 = n2337 & n2340;
  assign n2349 = n2348 ^ n2341;
  assign n2328 = ~x7 & n1396;
  assign n2329 = ~x6 & n1400;
  assign n2330 = ~n2328 & ~n2329;
  assign n2331 = x7 & n1403;
  assign n2332 = x6 & n1405;
  assign n2333 = ~n2331 & ~n2332;
  assign n2334 = n2330 & n2333;
  assign n2350 = n2349 ^ n2334;
  assign n2354 = n2353 ^ n2350;
  assign n2324 = n2173 ^ n2164;
  assign n2325 = ~n2174 & ~n2324;
  assign n2326 = n2325 ^ n2166;
  assign n2315 = ~x25 & n82;
  assign n2316 = ~x24 & n86;
  assign n2317 = ~n2315 & ~n2316;
  assign n2318 = x25 & n89;
  assign n2319 = x24 & n91;
  assign n2320 = ~n2318 & ~n2319;
  assign n2321 = n2317 & n2320;
  assign n2311 = x57 ^ x0;
  assign n2312 = ~n2165 & n2311;
  assign n2313 = n2312 ^ x0;
  assign n2314 = x59 & ~n2313;
  assign n2322 = n2321 ^ n2314;
  assign n2304 = x15 & n598;
  assign n2305 = x14 & n600;
  assign n2306 = ~n2304 & ~n2305;
  assign n2307 = ~x15 & n591;
  assign n2308 = ~x14 & n595;
  assign n2309 = ~n2307 & ~n2308;
  assign n2310 = n2306 & n2309;
  assign n2323 = n2322 ^ n2310;
  assign n2327 = n2326 ^ n2323;
  assign n2355 = n2354 ^ n2327;
  assign n2434 = n2433 ^ n2355;
  assign n2438 = n2437 ^ n2434;
  assign n2299 = n2127 ^ n2120;
  assign n2300 = ~n2124 & n2299;
  assign n2301 = n2300 ^ n2127;
  assign n2295 = n2245 ^ n2180;
  assign n2296 = n2258 ^ n2180;
  assign n2297 = ~n2295 & n2296;
  assign n2298 = n2297 ^ n2245;
  assign n2302 = n2301 ^ n2298;
  assign n2290 = n2257 ^ n2252;
  assign n2291 = n2253 & n2290;
  assign n2292 = n2291 ^ n2248;
  assign n2287 = n2175 ^ n2157;
  assign n2288 = n2179 & n2287;
  assign n2289 = n2288 ^ n2157;
  assign n2293 = n2292 ^ n2289;
  assign n2283 = n2224 ^ n2210;
  assign n2284 = n2225 & ~n2283;
  assign n2285 = n2284 ^ n2217;
  assign n2279 = n2148 ^ n2141;
  assign n2280 = ~n2156 & ~n2279;
  assign n2281 = n2280 ^ n2141;
  assign n2275 = n2194 ^ n2187;
  assign n2276 = n2201 ^ n2187;
  assign n2277 = n2275 & ~n2276;
  assign n2278 = n2277 ^ n2194;
  assign n2282 = n2281 ^ n2278;
  assign n2286 = n2285 ^ n2282;
  assign n2294 = n2293 ^ n2286;
  assign n2303 = n2302 ^ n2294;
  assign n2439 = n2438 ^ n2303;
  assign n2444 = n2443 ^ n2439;
  assign n2448 = n2447 ^ n2444;
  assign n2613 = n2447 ^ n2439;
  assign n2614 = n2444 & n2613;
  assign n2615 = n2614 ^ n2447;
  assign n2608 = n2434 ^ n2303;
  assign n2609 = n2437 ^ n2303;
  assign n2610 = ~n2608 & n2609;
  assign n2611 = n2610 ^ n2434;
  assign n2602 = n2298 ^ n2294;
  assign n2603 = n2301 ^ n2294;
  assign n2604 = ~n2602 & ~n2603;
  assign n2605 = n2604 ^ n2298;
  assign n2598 = n2289 ^ n2286;
  assign n2599 = n2293 & n2598;
  assign n2600 = n2599 ^ n2286;
  assign n2594 = n2353 ^ n2327;
  assign n2595 = n2354 & n2594;
  assign n2596 = n2595 ^ n2350;
  assign n2583 = ~x2 & n2406;
  assign n2584 = ~x1 & n2408;
  assign n2585 = ~n2583 & ~n2584;
  assign n2586 = x2 & n2399;
  assign n2587 = x1 & n2403;
  assign n2588 = ~n2586 & ~n2587;
  assign n2589 = n2585 & n2588;
  assign n2576 = x24 & n153;
  assign n2577 = x23 & n155;
  assign n2578 = ~n2576 & ~n2577;
  assign n2579 = ~x24 & n146;
  assign n2580 = ~x23 & n150;
  assign n2581 = ~n2579 & ~n2580;
  assign n2582 = n2578 & n2581;
  assign n2590 = n2589 ^ n2582;
  assign n2569 = ~x16 & n591;
  assign n2570 = ~x15 & n595;
  assign n2571 = ~n2569 & ~n2570;
  assign n2572 = x16 & n598;
  assign n2573 = x15 & n600;
  assign n2574 = ~n2572 & ~n2573;
  assign n2575 = n2571 & n2574;
  assign n2591 = n2590 ^ n2575;
  assign n2560 = ~x26 & n82;
  assign n2561 = ~x25 & n86;
  assign n2562 = ~n2560 & ~n2561;
  assign n2563 = x26 & n89;
  assign n2564 = x25 & n91;
  assign n2565 = ~n2563 & ~n2564;
  assign n2566 = n2562 & n2565;
  assign n2558 = x60 ^ x59;
  assign n2559 = x0 & n2558;
  assign n2567 = n2566 ^ n2559;
  assign n2551 = x22 & n217;
  assign n2552 = x21 & n219;
  assign n2553 = ~n2551 & ~n2552;
  assign n2554 = ~x22 & n210;
  assign n2555 = ~x21 & n214;
  assign n2556 = ~n2554 & ~n2555;
  assign n2557 = n2553 & n2556;
  assign n2568 = n2567 ^ n2557;
  assign n2592 = n2591 ^ n2568;
  assign n2542 = x8 & n1403;
  assign n2543 = x7 & n1405;
  assign n2544 = ~n2542 & ~n2543;
  assign n2545 = ~x8 & n1396;
  assign n2546 = ~x7 & n1400;
  assign n2547 = ~n2545 & ~n2546;
  assign n2548 = n2544 & n2547;
  assign n2535 = x10 & n1234;
  assign n2536 = x9 & n1238;
  assign n2537 = ~n2535 & ~n2536;
  assign n2538 = ~x10 & n1241;
  assign n2539 = ~x9 & n1243;
  assign n2540 = ~n2538 & ~n2539;
  assign n2541 = n2537 & n2540;
  assign n2549 = n2548 ^ n2541;
  assign n2533 = ~x27 & n68;
  assign n2531 = x33 ^ x28;
  assign n2532 = x32 & n2531;
  assign n2534 = n2533 ^ n2532;
  assign n2550 = n2549 ^ n2534;
  assign n2593 = n2592 ^ n2550;
  assign n2597 = n2596 ^ n2593;
  assign n2601 = n2600 ^ n2597;
  assign n2606 = n2605 ^ n2601;
  assign n2526 = n2429 ^ n2355;
  assign n2527 = n2432 ^ n2355;
  assign n2528 = n2526 & n2527;
  assign n2529 = n2528 ^ n2429;
  assign n2521 = n2326 ^ n2322;
  assign n2522 = n2323 & n2521;
  assign n2523 = n2522 ^ n2310;
  assign n2517 = n2285 ^ n2278;
  assign n2518 = n2282 & n2517;
  assign n2519 = n2518 ^ n2285;
  assign n2508 = ~x6 & n1687;
  assign n2509 = ~x5 & n1691;
  assign n2510 = ~n2508 & ~n2509;
  assign n2511 = x6 & n1694;
  assign n2512 = x5 & n1696;
  assign n2513 = ~n2511 & ~n2512;
  assign n2514 = n2510 & n2513;
  assign n2501 = x18 & n430;
  assign n2502 = x17 & n434;
  assign n2503 = ~n2501 & ~n2502;
  assign n2504 = ~x18 & n437;
  assign n2505 = ~x17 & n439;
  assign n2506 = ~n2504 & ~n2505;
  assign n2507 = n2503 & n2506;
  assign n2515 = n2514 ^ n2507;
  assign n2494 = ~x4 & n1962;
  assign n2495 = ~x3 & n1966;
  assign n2496 = ~n2494 & ~n2495;
  assign n2497 = x4 & n1969;
  assign n2498 = x3 & n1971;
  assign n2499 = ~n2497 & ~n2498;
  assign n2500 = n2496 & n2499;
  assign n2516 = n2515 ^ n2500;
  assign n2520 = n2519 ^ n2516;
  assign n2524 = n2523 ^ n2520;
  assign n2490 = n2398 ^ n2375;
  assign n2491 = ~n2428 & ~n2490;
  assign n2492 = n2491 ^ n2375;
  assign n2485 = n2348 ^ n2334;
  assign n2486 = n2349 & ~n2485;
  assign n2487 = n2486 ^ n2341;
  assign n2481 = n2396 ^ n2382;
  assign n2482 = n2397 & ~n2481;
  assign n2483 = n2482 ^ n2389;
  assign n2480 = n2314 & ~n2321;
  assign n2484 = n2483 ^ n2480;
  assign n2488 = n2487 ^ n2484;
  assign n2475 = n2425 ^ n2411;
  assign n2476 = n2426 & ~n2475;
  assign n2477 = n2476 ^ n2418;
  assign n2472 = n2369 ^ n2362;
  assign n2473 = ~n2374 & ~n2472;
  assign n2474 = n2473 ^ n2373;
  assign n2478 = n2477 ^ n2474;
  assign n2463 = ~x12 & n1000;
  assign n2464 = ~x11 & n1004;
  assign n2465 = ~n2463 & ~n2464;
  assign n2466 = x12 & n1007;
  assign n2467 = x11 & n1009;
  assign n2468 = ~n2466 & ~n2467;
  assign n2469 = n2465 & n2468;
  assign n2456 = ~x14 & n787;
  assign n2457 = ~x13 & n789;
  assign n2458 = ~n2456 & ~n2457;
  assign n2459 = x14 & n780;
  assign n2460 = x13 & n784;
  assign n2461 = ~n2459 & ~n2460;
  assign n2462 = n2458 & n2461;
  assign n2470 = n2469 ^ n2462;
  assign n2449 = ~x20 & n329;
  assign n2450 = ~x19 & n333;
  assign n2451 = ~n2449 & ~n2450;
  assign n2452 = x20 & n336;
  assign n2453 = x19 & n338;
  assign n2454 = ~n2452 & ~n2453;
  assign n2455 = n2451 & n2454;
  assign n2471 = n2470 ^ n2455;
  assign n2479 = n2478 ^ n2471;
  assign n2489 = n2488 ^ n2479;
  assign n2493 = n2492 ^ n2489;
  assign n2525 = n2524 ^ n2493;
  assign n2530 = n2529 ^ n2525;
  assign n2607 = n2606 ^ n2530;
  assign n2612 = n2611 ^ n2607;
  assign n2616 = n2615 ^ n2612;
  assign n2799 = n2615 ^ n2607;
  assign n2800 = ~n2612 & ~n2799;
  assign n2801 = n2800 ^ n2615;
  assign n2795 = n2601 ^ n2530;
  assign n2796 = ~n2606 & ~n2795;
  assign n2797 = n2796 ^ n2530;
  assign n2790 = n2600 ^ n2596;
  assign n2791 = n2597 & n2790;
  assign n2792 = n2791 ^ n2593;
  assign n2787 = n2529 ^ n2524;
  assign n2788 = ~n2525 & n2787;
  assign n2789 = n2788 ^ n2493;
  assign n2793 = n2792 ^ n2789;
  assign n2782 = n2492 ^ n2479;
  assign n2783 = ~n2489 & n2782;
  assign n2784 = n2783 ^ n2492;
  assign n2777 = n2523 ^ n2516;
  assign n2778 = n2523 ^ n2519;
  assign n2779 = n2777 & ~n2778;
  assign n2780 = n2779 ^ n2516;
  assign n2766 = ~x21 & n329;
  assign n2767 = ~x20 & n333;
  assign n2768 = ~n2766 & ~n2767;
  assign n2769 = x21 & n336;
  assign n2770 = x20 & n338;
  assign n2771 = ~n2769 & ~n2770;
  assign n2772 = n2768 & n2771;
  assign n2759 = ~x13 & n1000;
  assign n2760 = ~x12 & n1004;
  assign n2761 = ~n2759 & ~n2760;
  assign n2762 = x13 & n1007;
  assign n2763 = x12 & n1009;
  assign n2764 = ~n2762 & ~n2763;
  assign n2765 = n2761 & n2764;
  assign n2773 = n2772 ^ n2765;
  assign n2752 = x11 & n1234;
  assign n2753 = x10 & n1238;
  assign n2754 = ~n2752 & ~n2753;
  assign n2755 = ~x11 & n1241;
  assign n2756 = ~x10 & n1243;
  assign n2757 = ~n2755 & ~n2756;
  assign n2758 = n2754 & n2757;
  assign n2774 = n2773 ^ n2758;
  assign n2743 = ~x5 & n1962;
  assign n2744 = ~x4 & n1966;
  assign n2745 = ~n2743 & ~n2744;
  assign n2746 = x5 & n1969;
  assign n2747 = x4 & n1971;
  assign n2748 = ~n2746 & ~n2747;
  assign n2749 = n2745 & n2748;
  assign n2736 = ~x7 & n1687;
  assign n2737 = ~x6 & n1691;
  assign n2738 = ~n2736 & ~n2737;
  assign n2739 = x7 & n1694;
  assign n2740 = x6 & n1696;
  assign n2741 = ~n2739 & ~n2740;
  assign n2742 = n2738 & n2741;
  assign n2750 = n2749 ^ n2742;
  assign n2729 = ~x17 & n591;
  assign n2730 = ~x16 & n595;
  assign n2731 = ~n2729 & ~n2730;
  assign n2732 = x17 & n598;
  assign n2733 = x16 & n600;
  assign n2734 = ~n2732 & ~n2733;
  assign n2735 = n2731 & n2734;
  assign n2751 = n2750 ^ n2735;
  assign n2775 = n2774 ^ n2751;
  assign n2720 = x25 & n153;
  assign n2721 = x24 & n155;
  assign n2722 = ~n2720 & ~n2721;
  assign n2723 = ~x25 & n146;
  assign n2724 = ~x24 & n150;
  assign n2725 = ~n2723 & ~n2724;
  assign n2726 = n2722 & n2725;
  assign n2713 = ~x9 & n1396;
  assign n2714 = ~x8 & n1400;
  assign n2715 = ~n2713 & ~n2714;
  assign n2716 = x9 & n1403;
  assign n2717 = x8 & n1405;
  assign n2718 = ~n2716 & ~n2717;
  assign n2719 = n2715 & n2718;
  assign n2727 = n2726 ^ n2719;
  assign n2706 = ~x19 & n437;
  assign n2707 = ~x18 & n439;
  assign n2708 = ~n2706 & ~n2707;
  assign n2709 = x19 & n430;
  assign n2710 = x18 & n434;
  assign n2711 = ~n2709 & ~n2710;
  assign n2712 = n2708 & n2711;
  assign n2728 = n2727 ^ n2712;
  assign n2776 = n2775 ^ n2728;
  assign n2781 = n2780 ^ n2776;
  assign n2785 = n2784 ^ n2781;
  assign n2700 = n2568 ^ n2550;
  assign n2701 = n2591 ^ n2550;
  assign n2702 = n2700 & n2701;
  assign n2703 = n2702 ^ n2568;
  assign n2696 = n2487 ^ n2483;
  assign n2697 = ~n2484 & ~n2696;
  assign n2698 = n2697 ^ n2480;
  assign n2681 = x61 & n2558;
  assign n2682 = ~x1 & n2681;
  assign n2683 = x61 ^ x60;
  assign n2684 = ~n2558 & n2683;
  assign n2685 = x61 & n2684;
  assign n2686 = ~x0 & n2685;
  assign n2687 = ~n2682 & ~n2686;
  assign n2688 = ~x61 & n2558;
  assign n2689 = x1 & n2688;
  assign n2690 = ~x61 & n2684;
  assign n2691 = x0 & n2690;
  assign n2692 = ~n2689 & ~n2691;
  assign n2693 = n2687 & n2692;
  assign n2674 = x3 & n2399;
  assign n2675 = x2 & n2403;
  assign n2676 = ~n2674 & ~n2675;
  assign n2677 = ~x3 & n2406;
  assign n2678 = ~x2 & n2408;
  assign n2679 = ~n2677 & ~n2678;
  assign n2680 = n2676 & n2679;
  assign n2694 = n2693 ^ n2680;
  assign n2670 = x33 ^ x29;
  assign n2671 = x32 & n2670;
  assign n2669 = ~x28 & n68;
  assign n2672 = n2671 ^ n2669;
  assign n2665 = x59 ^ x0;
  assign n2666 = ~n2558 & n2665;
  assign n2667 = n2666 ^ x0;
  assign n2668 = x61 & ~n2667;
  assign n2673 = n2672 ^ n2668;
  assign n2695 = n2694 ^ n2673;
  assign n2699 = n2698 ^ n2695;
  assign n2704 = n2703 ^ n2699;
  assign n2660 = n2474 ^ n2471;
  assign n2661 = n2478 & ~n2660;
  assign n2662 = n2661 ^ n2471;
  assign n2656 = n2469 ^ n2455;
  assign n2657 = n2470 & ~n2656;
  assign n2658 = n2657 ^ n2462;
  assign n2652 = n2541 ^ n2534;
  assign n2653 = ~n2549 & ~n2652;
  assign n2654 = n2653 ^ n2534;
  assign n2648 = n2559 ^ n2557;
  assign n2649 = n2566 ^ n2557;
  assign n2650 = ~n2648 & ~n2649;
  assign n2651 = n2650 ^ n2559;
  assign n2655 = n2654 ^ n2651;
  assign n2659 = n2658 ^ n2655;
  assign n2663 = n2662 ^ n2659;
  assign n2643 = n2582 ^ n2575;
  assign n2644 = ~n2590 & n2643;
  assign n2645 = n2644 ^ n2575;
  assign n2640 = n2507 ^ n2500;
  assign n2641 = ~n2515 & n2640;
  assign n2642 = n2641 ^ n2500;
  assign n2646 = n2645 ^ n2642;
  assign n2631 = ~x23 & n210;
  assign n2632 = ~x22 & n214;
  assign n2633 = ~n2631 & ~n2632;
  assign n2634 = x23 & n217;
  assign n2635 = x22 & n219;
  assign n2636 = ~n2634 & ~n2635;
  assign n2637 = n2633 & n2636;
  assign n2624 = x27 & n89;
  assign n2625 = x26 & n91;
  assign n2626 = ~n2624 & ~n2625;
  assign n2627 = ~x27 & n82;
  assign n2628 = ~x26 & n86;
  assign n2629 = ~n2627 & ~n2628;
  assign n2630 = n2626 & n2629;
  assign n2638 = n2637 ^ n2630;
  assign n2617 = ~x15 & n787;
  assign n2618 = ~x14 & n789;
  assign n2619 = ~n2617 & ~n2618;
  assign n2620 = x15 & n780;
  assign n2621 = x14 & n784;
  assign n2622 = ~n2620 & ~n2621;
  assign n2623 = n2619 & n2622;
  assign n2639 = n2638 ^ n2623;
  assign n2647 = n2646 ^ n2639;
  assign n2664 = n2663 ^ n2647;
  assign n2705 = n2704 ^ n2664;
  assign n2786 = n2785 ^ n2705;
  assign n2794 = n2793 ^ n2786;
  assign n2798 = n2797 ^ n2794;
  assign n2802 = n2801 ^ n2798;
  assign n2978 = n2801 ^ n2794;
  assign n2979 = n2798 & n2978;
  assign n2980 = n2979 ^ n2801;
  assign n2974 = n2789 ^ n2786;
  assign n2975 = n2793 & ~n2974;
  assign n2976 = n2975 ^ n2786;
  assign n2970 = n2785 ^ n2704;
  assign n2971 = ~n2705 & ~n2970;
  assign n2972 = n2971 ^ n2664;
  assign n2964 = n2784 ^ n2776;
  assign n2965 = n2784 ^ n2780;
  assign n2966 = ~n2964 & n2965;
  assign n2967 = n2966 ^ n2776;
  assign n2959 = n2751 ^ n2728;
  assign n2960 = ~n2775 & n2959;
  assign n2961 = n2960 ^ n2728;
  assign n2955 = n2658 ^ n2651;
  assign n2956 = ~n2655 & ~n2955;
  assign n2957 = n2956 ^ n2658;
  assign n2951 = n2637 ^ n2623;
  assign n2952 = n2638 & ~n2951;
  assign n2953 = n2952 ^ n2630;
  assign n2949 = n2668 & n2672;
  assign n2942 = ~x2 & n2681;
  assign n2943 = ~x1 & n2685;
  assign n2944 = ~n2942 & ~n2943;
  assign n2945 = x2 & n2688;
  assign n2946 = x1 & n2690;
  assign n2947 = ~n2945 & ~n2946;
  assign n2948 = n2944 & n2947;
  assign n2950 = n2949 ^ n2948;
  assign n2954 = n2953 ^ n2950;
  assign n2958 = n2957 ^ n2954;
  assign n2962 = n2961 ^ n2958;
  assign n2937 = n2642 ^ n2639;
  assign n2938 = ~n2646 & n2937;
  assign n2939 = n2938 ^ n2639;
  assign n2933 = n2749 ^ n2735;
  assign n2934 = n2750 & ~n2933;
  assign n2935 = n2934 ^ n2742;
  assign n2929 = n2772 ^ n2758;
  assign n2930 = n2773 & ~n2929;
  assign n2931 = n2930 ^ n2765;
  assign n2926 = n2726 ^ n2712;
  assign n2927 = n2727 & ~n2926;
  assign n2928 = n2927 ^ n2719;
  assign n2932 = n2931 ^ n2928;
  assign n2936 = n2935 ^ n2932;
  assign n2940 = n2939 ^ n2936;
  assign n2922 = n2693 ^ n2673;
  assign n2923 = n2694 & n2922;
  assign n2924 = n2923 ^ n2680;
  assign n2912 = ~x12 & n1241;
  assign n2913 = ~x11 & n1243;
  assign n2914 = ~n2912 & ~n2913;
  assign n2915 = x12 & n1234;
  assign n2916 = x11 & n1238;
  assign n2917 = ~n2915 & ~n2916;
  assign n2918 = n2914 & n2917;
  assign n2905 = ~x22 & n329;
  assign n2906 = ~x21 & n333;
  assign n2907 = ~n2905 & ~n2906;
  assign n2908 = x22 & n336;
  assign n2909 = x21 & n338;
  assign n2910 = ~n2908 & ~n2909;
  assign n2911 = n2907 & n2910;
  assign n2919 = n2918 ^ n2911;
  assign n2898 = ~x10 & n1396;
  assign n2899 = ~x9 & n1400;
  assign n2900 = ~n2898 & ~n2899;
  assign n2901 = x10 & n1403;
  assign n2902 = x9 & n1405;
  assign n2903 = ~n2901 & ~n2902;
  assign n2904 = n2900 & n2903;
  assign n2920 = n2919 ^ n2904;
  assign n2889 = ~x16 & n787;
  assign n2890 = ~x15 & n789;
  assign n2891 = ~n2889 & ~n2890;
  assign n2892 = x16 & n780;
  assign n2893 = x15 & n784;
  assign n2894 = ~n2892 & ~n2893;
  assign n2895 = n2891 & n2894;
  assign n2882 = x24 & n217;
  assign n2883 = x23 & n219;
  assign n2884 = ~n2882 & ~n2883;
  assign n2885 = ~x24 & n210;
  assign n2886 = ~x23 & n214;
  assign n2887 = ~n2885 & ~n2886;
  assign n2888 = n2884 & n2887;
  assign n2896 = n2895 ^ n2888;
  assign n2875 = ~x14 & n1000;
  assign n2876 = ~x13 & n1004;
  assign n2877 = ~n2875 & ~n2876;
  assign n2878 = x14 & n1007;
  assign n2879 = x13 & n1009;
  assign n2880 = ~n2878 & ~n2879;
  assign n2881 = n2877 & n2880;
  assign n2897 = n2896 ^ n2881;
  assign n2921 = n2920 ^ n2897;
  assign n2925 = n2924 ^ n2921;
  assign n2941 = n2940 ^ n2925;
  assign n2963 = n2962 ^ n2941;
  assign n2968 = n2967 ^ n2963;
  assign n2870 = n2703 ^ n2695;
  assign n2871 = n2703 ^ n2698;
  assign n2872 = n2870 & ~n2871;
  assign n2873 = n2872 ^ n2695;
  assign n2866 = n2659 ^ n2647;
  assign n2867 = ~n2663 & n2866;
  assign n2868 = n2867 ^ n2647;
  assign n2855 = ~x18 & n591;
  assign n2856 = ~x17 & n595;
  assign n2857 = ~n2855 & ~n2856;
  assign n2858 = x18 & n598;
  assign n2859 = x17 & n600;
  assign n2860 = ~n2858 & ~n2859;
  assign n2861 = n2857 & n2860;
  assign n2848 = ~x6 & n1962;
  assign n2849 = ~x5 & n1966;
  assign n2850 = ~n2848 & ~n2849;
  assign n2851 = x6 & n1969;
  assign n2852 = x5 & n1971;
  assign n2853 = ~n2851 & ~n2852;
  assign n2854 = n2850 & n2853;
  assign n2862 = n2861 ^ n2854;
  assign n2841 = x4 & n2399;
  assign n2842 = x3 & n2403;
  assign n2843 = ~n2841 & ~n2842;
  assign n2844 = ~x4 & n2406;
  assign n2845 = ~x3 & n2408;
  assign n2846 = ~n2844 & ~n2845;
  assign n2847 = n2843 & n2846;
  assign n2863 = n2862 ^ n2847;
  assign n2833 = ~x28 & n82;
  assign n2834 = ~x27 & n86;
  assign n2835 = ~n2833 & ~n2834;
  assign n2836 = x28 & n89;
  assign n2837 = x27 & n91;
  assign n2838 = ~n2836 & ~n2837;
  assign n2839 = n2835 & n2838;
  assign n2830 = x62 ^ x61;
  assign n2831 = x0 & n2830;
  assign n2828 = ~x29 & n68;
  assign n2826 = x33 ^ x30;
  assign n2827 = x32 & n2826;
  assign n2829 = n2828 ^ n2827;
  assign n2832 = n2831 ^ n2829;
  assign n2840 = n2839 ^ n2832;
  assign n2864 = n2863 ^ n2840;
  assign n2817 = ~x20 & n437;
  assign n2818 = ~x19 & n439;
  assign n2819 = ~n2817 & ~n2818;
  assign n2820 = x20 & n430;
  assign n2821 = x19 & n434;
  assign n2822 = ~n2820 & ~n2821;
  assign n2823 = n2819 & n2822;
  assign n2810 = ~x26 & n146;
  assign n2811 = ~x25 & n150;
  assign n2812 = ~n2810 & ~n2811;
  assign n2813 = x26 & n153;
  assign n2814 = x25 & n155;
  assign n2815 = ~n2813 & ~n2814;
  assign n2816 = n2812 & n2815;
  assign n2824 = n2823 ^ n2816;
  assign n2803 = x8 & n1694;
  assign n2804 = x7 & n1696;
  assign n2805 = ~n2803 & ~n2804;
  assign n2806 = ~x8 & n1687;
  assign n2807 = ~x7 & n1691;
  assign n2808 = ~n2806 & ~n2807;
  assign n2809 = n2805 & n2808;
  assign n2825 = n2824 ^ n2809;
  assign n2865 = n2864 ^ n2825;
  assign n2869 = n2868 ^ n2865;
  assign n2874 = n2873 ^ n2869;
  assign n2969 = n2968 ^ n2874;
  assign n2973 = n2972 ^ n2969;
  assign n2977 = n2976 ^ n2973;
  assign n2981 = n2980 ^ n2977;
  assign n3176 = n2980 ^ n2973;
  assign n3177 = ~n2977 & ~n3176;
  assign n3178 = n3177 ^ n2980;
  assign n3171 = n2972 ^ n2874;
  assign n3172 = n2972 ^ n2968;
  assign n3173 = ~n3171 & n3172;
  assign n3174 = n3173 ^ n2874;
  assign n3167 = n2967 ^ n2962;
  assign n3168 = ~n2963 & n3167;
  assign n3169 = n3168 ^ n2941;
  assign n3162 = n2873 ^ n2868;
  assign n3163 = n2869 & n3162;
  assign n3164 = n3163 ^ n2865;
  assign n3156 = n2924 ^ n2920;
  assign n3157 = n2921 & ~n3156;
  assign n3158 = n3157 ^ n2897;
  assign n3152 = n2840 ^ n2825;
  assign n3153 = n2863 ^ n2825;
  assign n3154 = n3152 & ~n3153;
  assign n3155 = n3154 ^ n2840;
  assign n3159 = n3158 ^ n3155;
  assign n3141 = x19 & n598;
  assign n3142 = x18 & n600;
  assign n3143 = ~n3141 & ~n3142;
  assign n3144 = ~x19 & n591;
  assign n3145 = ~x18 & n595;
  assign n3146 = ~n3144 & ~n3145;
  assign n3147 = n3143 & n3146;
  assign n3134 = ~x5 & n2406;
  assign n3135 = ~x4 & n2408;
  assign n3136 = ~n3134 & ~n3135;
  assign n3137 = x5 & n2399;
  assign n3138 = x4 & n2403;
  assign n3139 = ~n3137 & ~n3138;
  assign n3140 = n3136 & n3139;
  assign n3148 = n3147 ^ n3140;
  assign n3127 = ~x3 & n2681;
  assign n3128 = ~x2 & n2685;
  assign n3129 = ~n3127 & ~n3128;
  assign n3130 = x3 & n2688;
  assign n3131 = x2 & n2690;
  assign n3132 = ~n3130 & ~n3131;
  assign n3133 = n3129 & n3132;
  assign n3149 = n3148 ^ n3133;
  assign n3118 = ~x25 & n210;
  assign n3119 = ~x24 & n214;
  assign n3120 = ~n3118 & ~n3119;
  assign n3121 = x25 & n217;
  assign n3122 = x24 & n219;
  assign n3123 = ~n3121 & ~n3122;
  assign n3124 = n3120 & n3123;
  assign n3111 = ~x29 & n82;
  assign n3112 = ~x28 & n86;
  assign n3113 = ~n3111 & ~n3112;
  assign n3114 = x29 & n89;
  assign n3115 = x28 & n91;
  assign n3116 = ~n3114 & ~n3115;
  assign n3117 = n3113 & n3116;
  assign n3125 = n3124 ^ n3117;
  assign n3098 = x63 & n2830;
  assign n3099 = ~x1 & n3098;
  assign n3100 = x63 ^ x62;
  assign n3101 = ~n2830 & n3100;
  assign n3102 = x63 & n3101;
  assign n3103 = ~x0 & n3102;
  assign n3104 = ~n3099 & ~n3103;
  assign n3105 = ~x63 & n2830;
  assign n3106 = x1 & n3105;
  assign n3107 = ~x63 & n3101;
  assign n3108 = x0 & n3107;
  assign n3109 = ~n3106 & ~n3108;
  assign n3110 = n3104 & n3109;
  assign n3126 = n3125 ^ n3110;
  assign n3150 = n3149 ^ n3126;
  assign n3089 = x17 & n780;
  assign n3090 = x16 & n784;
  assign n3091 = ~n3089 & ~n3090;
  assign n3092 = ~x17 & n787;
  assign n3093 = ~x16 & n789;
  assign n3094 = ~n3092 & ~n3093;
  assign n3095 = n3091 & n3094;
  assign n3082 = ~x15 & n1000;
  assign n3083 = ~x14 & n1004;
  assign n3084 = ~n3082 & ~n3083;
  assign n3085 = x15 & n1007;
  assign n3086 = x14 & n1009;
  assign n3087 = ~n3085 & ~n3086;
  assign n3088 = n3084 & n3087;
  assign n3096 = n3095 ^ n3088;
  assign n3075 = ~x23 & n329;
  assign n3076 = ~x22 & n333;
  assign n3077 = ~n3075 & ~n3076;
  assign n3078 = x23 & n336;
  assign n3079 = x22 & n338;
  assign n3080 = ~n3078 & ~n3079;
  assign n3081 = n3077 & n3080;
  assign n3097 = n3096 ^ n3081;
  assign n3151 = n3150 ^ n3097;
  assign n3160 = n3159 ^ n3151;
  assign n3070 = n2953 ^ n2949;
  assign n3071 = ~n2950 & n3070;
  assign n3072 = n3071 ^ n2948;
  assign n3066 = n2861 ^ n2847;
  assign n3067 = n2862 & ~n3066;
  assign n3068 = n3067 ^ n2854;
  assign n3062 = n2823 ^ n2809;
  assign n3063 = n2824 & ~n3062;
  assign n3064 = n3063 ^ n2816;
  assign n3059 = n2918 ^ n2904;
  assign n3060 = n2919 & ~n3059;
  assign n3061 = n3060 ^ n2911;
  assign n3065 = n3064 ^ n3061;
  assign n3069 = n3068 ^ n3065;
  assign n3073 = n3072 ^ n3069;
  assign n3055 = n2895 ^ n2881;
  assign n3056 = n2896 & ~n3055;
  assign n3057 = n3056 ^ n2888;
  assign n3051 = n2839 ^ n2829;
  assign n3052 = n2832 & n3051;
  assign n3053 = n3052 ^ n2831;
  assign n3047 = x33 ^ x31;
  assign n3048 = x32 & n3047;
  assign n3046 = ~x30 & n68;
  assign n3049 = n3048 ^ n3046;
  assign n3042 = x61 ^ x0;
  assign n3043 = ~n2830 & n3042;
  assign n3044 = n3043 ^ x0;
  assign n3045 = x63 & ~n3044;
  assign n3050 = n3049 ^ n3045;
  assign n3054 = n3053 ^ n3050;
  assign n3058 = n3057 ^ n3054;
  assign n3074 = n3073 ^ n3058;
  assign n3161 = n3160 ^ n3074;
  assign n3165 = n3164 ^ n3161;
  assign n3038 = n2936 ^ n2925;
  assign n3039 = ~n2940 & n3038;
  assign n3040 = n3039 ^ n2925;
  assign n3033 = n2961 ^ n2954;
  assign n3034 = n2961 ^ n2957;
  assign n3035 = ~n3033 & ~n3034;
  assign n3036 = n3035 ^ n2954;
  assign n3029 = n2935 ^ n2928;
  assign n3030 = ~n2932 & n3029;
  assign n3031 = n3030 ^ n2935;
  assign n3019 = ~x11 & n1396;
  assign n3020 = ~x10 & n1400;
  assign n3021 = ~n3019 & ~n3020;
  assign n3022 = x11 & n1403;
  assign n3023 = x10 & n1405;
  assign n3024 = ~n3022 & ~n3023;
  assign n3025 = n3021 & n3024;
  assign n3012 = x13 & n1234;
  assign n3013 = x12 & n1238;
  assign n3014 = ~n3012 & ~n3013;
  assign n3015 = ~x13 & n1241;
  assign n3016 = ~x12 & n1243;
  assign n3017 = ~n3015 & ~n3016;
  assign n3018 = n3014 & n3017;
  assign n3026 = n3025 ^ n3018;
  assign n3005 = ~x27 & n146;
  assign n3006 = ~x26 & n150;
  assign n3007 = ~n3005 & ~n3006;
  assign n3008 = x27 & n153;
  assign n3009 = x26 & n155;
  assign n3010 = ~n3008 & ~n3009;
  assign n3011 = n3007 & n3010;
  assign n3027 = n3026 ^ n3011;
  assign n2996 = x21 & n430;
  assign n2997 = x20 & n434;
  assign n2998 = ~n2996 & ~n2997;
  assign n2999 = ~x21 & n437;
  assign n3000 = ~x20 & n439;
  assign n3001 = ~n2999 & ~n3000;
  assign n3002 = n2998 & n3001;
  assign n2989 = ~x9 & n1687;
  assign n2990 = ~x8 & n1691;
  assign n2991 = ~n2989 & ~n2990;
  assign n2992 = x9 & n1694;
  assign n2993 = x8 & n1696;
  assign n2994 = ~n2992 & ~n2993;
  assign n2995 = n2991 & n2994;
  assign n3003 = n3002 ^ n2995;
  assign n2982 = x7 & n1969;
  assign n2983 = x6 & n1971;
  assign n2984 = ~n2982 & ~n2983;
  assign n2985 = ~x7 & n1962;
  assign n2986 = ~x6 & n1966;
  assign n2987 = ~n2985 & ~n2986;
  assign n2988 = n2984 & n2987;
  assign n3004 = n3003 ^ n2988;
  assign n3028 = n3027 ^ n3004;
  assign n3032 = n3031 ^ n3028;
  assign n3037 = n3036 ^ n3032;
  assign n3041 = n3040 ^ n3037;
  assign n3166 = n3165 ^ n3041;
  assign n3170 = n3169 ^ n3166;
  assign n3175 = n3174 ^ n3170;
  assign n3179 = n3178 ^ n3175;
  assign n3363 = n3178 ^ n3170;
  assign n3364 = ~n3175 & n3363;
  assign n3365 = n3364 ^ n3178;
  assign n3359 = n3169 ^ n3165;
  assign n3360 = ~n3166 & ~n3359;
  assign n3361 = n3360 ^ n3041;
  assign n3354 = n3164 ^ n3160;
  assign n3355 = n3161 & ~n3354;
  assign n3356 = n3355 ^ n3074;
  assign n3351 = n3040 ^ n3036;
  assign n3352 = ~n3037 & n3351;
  assign n3353 = n3352 ^ n3032;
  assign n3357 = n3356 ^ n3353;
  assign n3346 = n3155 ^ n3151;
  assign n3347 = ~n3159 & n3346;
  assign n3348 = n3347 ^ n3151;
  assign n3342 = n3069 ^ n3058;
  assign n3343 = ~n3073 & n3342;
  assign n3344 = n3343 ^ n3058;
  assign n3338 = n3068 ^ n3064;
  assign n3339 = n3065 & ~n3338;
  assign n3340 = n3339 ^ n3061;
  assign n3328 = ~x26 & n210;
  assign n3329 = ~x25 & n214;
  assign n3330 = ~n3328 & ~n3329;
  assign n3331 = x26 & n217;
  assign n3332 = x25 & n219;
  assign n3333 = ~n3331 & ~n3332;
  assign n3334 = n3330 & n3333;
  assign n3321 = x2 & n3105;
  assign n3322 = x1 & n3107;
  assign n3323 = ~n3321 & ~n3322;
  assign n3324 = ~x2 & n3098;
  assign n3325 = ~x1 & n3102;
  assign n3326 = ~n3324 & ~n3325;
  assign n3327 = n3323 & n3326;
  assign n3335 = n3334 ^ n3327;
  assign n3314 = x18 & n780;
  assign n3315 = x17 & n784;
  assign n3316 = ~n3314 & ~n3315;
  assign n3317 = ~x18 & n787;
  assign n3318 = ~x17 & n789;
  assign n3319 = ~n3317 & ~n3318;
  assign n3320 = n3316 & n3319;
  assign n3336 = n3335 ^ n3320;
  assign n3305 = ~x4 & n2681;
  assign n3306 = ~x3 & n2685;
  assign n3307 = ~n3305 & ~n3306;
  assign n3308 = x4 & n2688;
  assign n3309 = x3 & n2690;
  assign n3310 = ~n3308 & ~n3309;
  assign n3311 = n3307 & n3310;
  assign n3298 = ~x6 & n2406;
  assign n3299 = ~x5 & n2408;
  assign n3300 = ~n3298 & ~n3299;
  assign n3301 = x6 & n2399;
  assign n3302 = x5 & n2403;
  assign n3303 = ~n3301 & ~n3302;
  assign n3304 = n3300 & n3303;
  assign n3312 = n3311 ^ n3304;
  assign n3297 = n3045 & n3049;
  assign n3313 = n3312 ^ n3297;
  assign n3337 = n3336 ^ n3313;
  assign n3341 = n3340 ^ n3337;
  assign n3345 = n3344 ^ n3341;
  assign n3349 = n3348 ^ n3345;
  assign n3292 = n3031 ^ n3027;
  assign n3293 = n3028 & ~n3292;
  assign n3294 = n3293 ^ n3004;
  assign n3286 = n3018 ^ n3011;
  assign n3287 = n3025 ^ n3011;
  assign n3288 = n3286 & ~n3287;
  assign n3289 = n3288 ^ n3018;
  assign n3282 = n3124 ^ n3110;
  assign n3283 = n3125 & ~n3282;
  assign n3284 = n3283 ^ n3117;
  assign n3279 = n3088 ^ n3081;
  assign n3280 = ~n3096 & n3279;
  assign n3281 = n3280 ^ n3081;
  assign n3285 = n3284 ^ n3281;
  assign n3290 = n3289 ^ n3285;
  assign n3268 = x12 & n1403;
  assign n3269 = x11 & n1405;
  assign n3270 = ~n3268 & ~n3269;
  assign n3271 = ~x12 & n1396;
  assign n3272 = ~x11 & n1400;
  assign n3273 = ~n3271 & ~n3272;
  assign n3274 = n3270 & n3273;
  assign n3261 = x28 & n153;
  assign n3262 = x27 & n155;
  assign n3263 = ~n3261 & ~n3262;
  assign n3264 = ~x28 & n146;
  assign n3265 = ~x27 & n150;
  assign n3266 = ~n3264 & ~n3265;
  assign n3267 = n3263 & n3266;
  assign n3275 = n3274 ^ n3267;
  assign n3254 = x22 & n430;
  assign n3255 = x21 & n434;
  assign n3256 = ~n3254 & ~n3255;
  assign n3257 = ~x22 & n437;
  assign n3258 = ~x21 & n439;
  assign n3259 = ~n3257 & ~n3258;
  assign n3260 = n3256 & n3259;
  assign n3276 = n3275 ^ n3260;
  assign n3245 = ~x16 & n1000;
  assign n3246 = ~x15 & n1004;
  assign n3247 = ~n3245 & ~n3246;
  assign n3248 = x16 & n1007;
  assign n3249 = x15 & n1009;
  assign n3250 = ~n3248 & ~n3249;
  assign n3251 = n3247 & n3250;
  assign n3238 = ~x24 & n329;
  assign n3239 = ~x23 & n333;
  assign n3240 = ~n3238 & ~n3239;
  assign n3241 = x24 & n336;
  assign n3242 = x23 & n338;
  assign n3243 = ~n3241 & ~n3242;
  assign n3244 = n3240 & n3243;
  assign n3252 = n3251 ^ n3244;
  assign n3231 = ~x14 & n1241;
  assign n3232 = ~x13 & n1243;
  assign n3233 = ~n3231 & ~n3232;
  assign n3234 = x14 & n1234;
  assign n3235 = x13 & n1238;
  assign n3236 = ~n3234 & ~n3235;
  assign n3237 = n3233 & n3236;
  assign n3253 = n3252 ^ n3237;
  assign n3277 = n3276 ^ n3253;
  assign n3222 = x8 & n1969;
  assign n3223 = x7 & n1971;
  assign n3224 = ~n3222 & ~n3223;
  assign n3225 = ~x8 & n1962;
  assign n3226 = ~x7 & n1966;
  assign n3227 = ~n3225 & ~n3226;
  assign n3228 = n3224 & n3227;
  assign n3215 = ~x10 & n1687;
  assign n3216 = ~x9 & n1691;
  assign n3217 = ~n3215 & ~n3216;
  assign n3218 = x10 & n1694;
  assign n3219 = x9 & n1696;
  assign n3220 = ~n3218 & ~n3219;
  assign n3221 = n3217 & n3220;
  assign n3229 = n3228 ^ n3221;
  assign n3208 = x20 & n598;
  assign n3209 = x19 & n600;
  assign n3210 = ~n3208 & ~n3209;
  assign n3211 = ~x20 & n591;
  assign n3212 = ~x19 & n595;
  assign n3213 = ~n3211 & ~n3212;
  assign n3214 = n3210 & n3213;
  assign n3230 = n3229 ^ n3214;
  assign n3278 = n3277 ^ n3230;
  assign n3291 = n3290 ^ n3278;
  assign n3295 = n3294 ^ n3291;
  assign n3203 = n3057 ^ n3053;
  assign n3204 = n3054 & n3203;
  assign n3205 = n3204 ^ n3050;
  assign n3200 = n3126 ^ n3097;
  assign n3201 = ~n3150 & n3200;
  assign n3202 = n3201 ^ n3097;
  assign n3206 = n3205 ^ n3202;
  assign n3195 = n3140 ^ n3133;
  assign n3196 = ~n3148 & n3195;
  assign n3197 = n3196 ^ n3133;
  assign n3192 = n2995 ^ n2988;
  assign n3193 = ~n3003 & n3192;
  assign n3194 = n3193 ^ n2988;
  assign n3198 = n3197 ^ n3194;
  assign n3184 = ~x30 & n82;
  assign n3185 = ~x29 & n86;
  assign n3186 = ~n3184 & ~n3185;
  assign n3187 = x30 & n89;
  assign n3188 = x29 & n91;
  assign n3189 = ~n3187 & ~n3188;
  assign n3190 = n3186 & n3189;
  assign n3181 = x31 & n68;
  assign n3182 = n3181 ^ x33;
  assign n3180 = x0 & x63;
  assign n3183 = n3182 ^ n3180;
  assign n3191 = n3190 ^ n3183;
  assign n3199 = n3198 ^ n3191;
  assign n3207 = n3206 ^ n3199;
  assign n3296 = n3295 ^ n3207;
  assign n3350 = n3349 ^ n3296;
  assign n3358 = n3357 ^ n3350;
  assign n3362 = n3361 ^ n3358;
  assign n3366 = n3365 ^ n3362;
  assign n3553 = n3365 ^ n3358;
  assign n3554 = n3362 & ~n3553;
  assign n3555 = n3554 ^ n3365;
  assign n3549 = n3353 ^ n3350;
  assign n3550 = ~n3357 & n3549;
  assign n3551 = n3550 ^ n3350;
  assign n3545 = n3349 ^ n3295;
  assign n3546 = ~n3296 & n3545;
  assign n3547 = n3546 ^ n3207;
  assign n3540 = n3348 ^ n3344;
  assign n3541 = ~n3345 & ~n3540;
  assign n3542 = n3541 ^ n3341;
  assign n3536 = n3294 ^ n3290;
  assign n3537 = n3291 & ~n3536;
  assign n3538 = n3537 ^ n3278;
  assign n3532 = n3340 ^ n3336;
  assign n3533 = ~n3337 & ~n3532;
  assign n3534 = n3533 ^ n3313;
  assign n3525 = n3267 ^ n3260;
  assign n3526 = n3274 ^ n3260;
  assign n3527 = n3525 & ~n3526;
  assign n3528 = n3527 ^ n3267;
  assign n3516 = ~x3 & n3098;
  assign n3517 = ~x2 & n3102;
  assign n3518 = ~n3516 & ~n3517;
  assign n3519 = x3 & n3105;
  assign n3520 = x2 & n3107;
  assign n3521 = ~n3519 & ~n3520;
  assign n3522 = n3518 & n3521;
  assign n3509 = ~x19 & n787;
  assign n3510 = ~x18 & n789;
  assign n3511 = ~n3509 & ~n3510;
  assign n3512 = x19 & n780;
  assign n3513 = x18 & n784;
  assign n3514 = ~n3512 & ~n3513;
  assign n3515 = n3511 & n3514;
  assign n3523 = n3522 ^ n3515;
  assign n3508 = x1 & x63;
  assign n3524 = n3523 ^ n3508;
  assign n3529 = n3528 ^ n3524;
  assign n3499 = ~x9 & n1962;
  assign n3500 = ~x8 & n1966;
  assign n3501 = ~n3499 & ~n3500;
  assign n3502 = x9 & n1969;
  assign n3503 = x8 & n1971;
  assign n3504 = ~n3502 & ~n3503;
  assign n3505 = n3501 & n3504;
  assign n3492 = ~x21 & n591;
  assign n3493 = ~x20 & n595;
  assign n3494 = ~n3492 & ~n3493;
  assign n3495 = x21 & n598;
  assign n3496 = x20 & n600;
  assign n3497 = ~n3495 & ~n3496;
  assign n3498 = n3494 & n3497;
  assign n3506 = n3505 ^ n3498;
  assign n3485 = x7 & n2399;
  assign n3486 = x6 & n2403;
  assign n3487 = ~n3485 & ~n3486;
  assign n3488 = ~x7 & n2406;
  assign n3489 = ~x6 & n2408;
  assign n3490 = ~n3488 & ~n3489;
  assign n3491 = n3487 & n3490;
  assign n3507 = n3506 ^ n3491;
  assign n3530 = n3529 ^ n3507;
  assign n3474 = ~x17 & n1000;
  assign n3475 = ~x16 & n1004;
  assign n3476 = ~n3474 & ~n3475;
  assign n3477 = x17 & n1007;
  assign n3478 = x16 & n1009;
  assign n3479 = ~n3477 & ~n3478;
  assign n3480 = n3476 & n3479;
  assign n3467 = ~x31 & n82;
  assign n3468 = ~x30 & n86;
  assign n3469 = ~n3467 & ~n3468;
  assign n3470 = x31 & n89;
  assign n3471 = x30 & n91;
  assign n3472 = ~n3470 & ~n3471;
  assign n3473 = n3469 & n3472;
  assign n3481 = n3480 ^ n3473;
  assign n3460 = x27 & n217;
  assign n3461 = x26 & n219;
  assign n3462 = ~n3460 & ~n3461;
  assign n3463 = ~x27 & n210;
  assign n3464 = ~x26 & n214;
  assign n3465 = ~n3463 & ~n3464;
  assign n3466 = n3462 & n3465;
  assign n3482 = n3481 ^ n3466;
  assign n3451 = x23 & n430;
  assign n3452 = x22 & n434;
  assign n3453 = ~n3451 & ~n3452;
  assign n3454 = ~x23 & n437;
  assign n3455 = ~x22 & n439;
  assign n3456 = ~n3454 & ~n3455;
  assign n3457 = n3453 & n3456;
  assign n3444 = ~x29 & n146;
  assign n3445 = ~x28 & n150;
  assign n3446 = ~n3444 & ~n3445;
  assign n3447 = x29 & n153;
  assign n3448 = x28 & n155;
  assign n3449 = ~n3447 & ~n3448;
  assign n3450 = n3446 & n3449;
  assign n3458 = n3457 ^ n3450;
  assign n3437 = ~x11 & n1687;
  assign n3438 = ~x10 & n1691;
  assign n3439 = ~n3437 & ~n3438;
  assign n3440 = x11 & n1694;
  assign n3441 = x10 & n1696;
  assign n3442 = ~n3440 & ~n3441;
  assign n3443 = n3439 & n3442;
  assign n3459 = n3458 ^ n3443;
  assign n3483 = n3482 ^ n3459;
  assign n3428 = ~x25 & n329;
  assign n3429 = ~x24 & n333;
  assign n3430 = ~n3428 & ~n3429;
  assign n3431 = x25 & n336;
  assign n3432 = x24 & n338;
  assign n3433 = ~n3431 & ~n3432;
  assign n3434 = n3430 & n3433;
  assign n3421 = x15 & n1234;
  assign n3422 = x14 & n1238;
  assign n3423 = ~n3421 & ~n3422;
  assign n3424 = ~x15 & n1241;
  assign n3425 = ~x14 & n1243;
  assign n3426 = ~n3424 & ~n3425;
  assign n3427 = n3423 & n3426;
  assign n3435 = n3434 ^ n3427;
  assign n3414 = ~x13 & n1396;
  assign n3415 = ~x12 & n1400;
  assign n3416 = ~n3414 & ~n3415;
  assign n3417 = x13 & n1403;
  assign n3418 = x12 & n1405;
  assign n3419 = ~n3417 & ~n3418;
  assign n3420 = n3416 & n3419;
  assign n3436 = n3435 ^ n3420;
  assign n3484 = n3483 ^ n3436;
  assign n3531 = n3530 ^ n3484;
  assign n3535 = n3534 ^ n3531;
  assign n3539 = n3538 ^ n3535;
  assign n3543 = n3542 ^ n3539;
  assign n3408 = n3202 ^ n3199;
  assign n3409 = n3205 ^ n3199;
  assign n3410 = n3408 & n3409;
  assign n3411 = n3410 ^ n3202;
  assign n3404 = n3194 ^ n3191;
  assign n3405 = ~n3198 & n3404;
  assign n3406 = n3405 ^ n3191;
  assign n3400 = n3289 ^ n3284;
  assign n3401 = n3285 & ~n3400;
  assign n3402 = n3401 ^ n3281;
  assign n3397 = n3311 ^ n3297;
  assign n3398 = n3312 & n3397;
  assign n3399 = n3398 ^ n3304;
  assign n3403 = n3402 ^ n3399;
  assign n3407 = n3406 ^ n3403;
  assign n3412 = n3411 ^ n3407;
  assign n3393 = n3276 ^ n3230;
  assign n3394 = n3277 & ~n3393;
  assign n3395 = n3394 ^ n3253;
  assign n3387 = n3221 ^ n3214;
  assign n3388 = n3228 ^ n3214;
  assign n3389 = n3387 & ~n3388;
  assign n3390 = n3389 ^ n3221;
  assign n3383 = n3251 ^ n3237;
  assign n3384 = n3252 & ~n3383;
  assign n3385 = n3384 ^ n3244;
  assign n3379 = n3327 ^ n3320;
  assign n3380 = n3334 ^ n3320;
  assign n3381 = n3379 & ~n3380;
  assign n3382 = n3381 ^ n3327;
  assign n3386 = n3385 ^ n3382;
  assign n3391 = n3390 ^ n3386;
  assign n3375 = n3190 ^ n3182;
  assign n3376 = n3183 & n3375;
  assign n3377 = n3376 ^ n3180;
  assign n3367 = ~x5 & n2681;
  assign n3368 = ~x4 & n2685;
  assign n3369 = ~n3367 & ~n3368;
  assign n3370 = x5 & n2688;
  assign n3371 = x4 & n2690;
  assign n3372 = ~n3370 & ~n3371;
  assign n3373 = n3369 & n3372;
  assign n3374 = n3373 ^ x33;
  assign n3378 = n3377 ^ n3374;
  assign n3392 = n3391 ^ n3378;
  assign n3396 = n3395 ^ n3392;
  assign n3413 = n3412 ^ n3396;
  assign n3544 = n3543 ^ n3413;
  assign n3548 = n3547 ^ n3544;
  assign n3552 = n3551 ^ n3548;
  assign n3556 = n3555 ^ n3552;
  assign n3739 = n3555 ^ n3548;
  assign n3740 = ~n3552 & ~n3739;
  assign n3741 = n3740 ^ n3555;
  assign n3735 = n3547 ^ n3543;
  assign n3736 = ~n3544 & ~n3735;
  assign n3737 = n3736 ^ n3413;
  assign n3731 = n3542 ^ n3538;
  assign n3732 = n3539 & n3731;
  assign n3733 = n3732 ^ n3535;
  assign n3726 = n3407 ^ n3396;
  assign n3727 = ~n3412 & n3726;
  assign n3728 = n3727 ^ n3396;
  assign n3722 = n3534 ^ n3530;
  assign n3723 = ~n3531 & ~n3722;
  assign n3724 = n3723 ^ n3484;
  assign n3717 = n3395 ^ n3378;
  assign n3718 = n3395 ^ n3391;
  assign n3719 = n3717 & ~n3718;
  assign n3720 = n3719 ^ n3378;
  assign n3710 = n3498 ^ n3491;
  assign n3711 = n3505 ^ n3491;
  assign n3712 = n3710 & ~n3711;
  assign n3713 = n3712 ^ n3498;
  assign n3701 = x20 & n780;
  assign n3702 = x19 & n784;
  assign n3703 = ~n3701 & ~n3702;
  assign n3704 = ~x20 & n787;
  assign n3705 = ~x19 & n789;
  assign n3706 = ~n3704 & ~n3705;
  assign n3707 = n3703 & n3706;
  assign n3694 = ~x6 & n2681;
  assign n3695 = ~x5 & n2685;
  assign n3696 = ~n3694 & ~n3695;
  assign n3697 = x6 & n2688;
  assign n3698 = x5 & n2690;
  assign n3699 = ~n3697 & ~n3698;
  assign n3700 = n3696 & n3699;
  assign n3708 = n3707 ^ n3700;
  assign n3687 = ~x4 & n3098;
  assign n3688 = ~x3 & n3102;
  assign n3689 = ~n3687 & ~n3688;
  assign n3690 = x4 & n3105;
  assign n3691 = x3 & n3107;
  assign n3692 = ~n3690 & ~n3691;
  assign n3693 = n3689 & n3692;
  assign n3709 = n3708 ^ n3693;
  assign n3714 = n3713 ^ n3709;
  assign n3678 = x16 & n1234;
  assign n3679 = x15 & n1238;
  assign n3680 = ~n3678 & ~n3679;
  assign n3681 = ~x16 & n1241;
  assign n3682 = ~x15 & n1243;
  assign n3683 = ~n3681 & ~n3682;
  assign n3684 = n3680 & n3683;
  assign n3671 = ~x18 & n1000;
  assign n3672 = ~x17 & n1004;
  assign n3673 = ~n3671 & ~n3672;
  assign n3674 = x18 & n1007;
  assign n3675 = x17 & n1009;
  assign n3676 = ~n3674 & ~n3675;
  assign n3677 = n3673 & n3676;
  assign n3685 = n3684 ^ n3677;
  assign n3664 = ~x24 & n437;
  assign n3665 = ~x23 & n439;
  assign n3666 = ~n3664 & ~n3665;
  assign n3667 = x24 & n430;
  assign n3668 = x23 & n434;
  assign n3669 = ~n3667 & ~n3668;
  assign n3670 = n3666 & n3669;
  assign n3686 = n3685 ^ n3670;
  assign n3715 = n3714 ^ n3686;
  assign n3653 = ~x14 & n1396;
  assign n3654 = ~x13 & n1400;
  assign n3655 = ~n3653 & ~n3654;
  assign n3656 = x14 & n1403;
  assign n3657 = x13 & n1405;
  assign n3658 = ~n3656 & ~n3657;
  assign n3659 = n3655 & n3658;
  assign n3646 = ~x12 & n1687;
  assign n3647 = ~x11 & n1691;
  assign n3648 = ~n3646 & ~n3647;
  assign n3649 = x12 & n1694;
  assign n3650 = x11 & n1696;
  assign n3651 = ~n3649 & ~n3650;
  assign n3652 = n3648 & n3651;
  assign n3660 = n3659 ^ n3652;
  assign n3639 = ~x28 & n210;
  assign n3640 = ~x27 & n214;
  assign n3641 = ~n3639 & ~n3640;
  assign n3642 = x28 & n217;
  assign n3643 = x27 & n219;
  assign n3644 = ~n3642 & ~n3643;
  assign n3645 = n3641 & n3644;
  assign n3661 = n3660 ^ n3645;
  assign n3630 = ~x30 & n146;
  assign n3631 = ~x29 & n150;
  assign n3632 = ~n3630 & ~n3631;
  assign n3633 = x30 & n153;
  assign n3634 = x29 & n155;
  assign n3635 = ~n3633 & ~n3634;
  assign n3636 = n3632 & n3635;
  assign n3623 = ~x26 & n329;
  assign n3624 = ~x25 & n333;
  assign n3625 = ~n3623 & ~n3624;
  assign n3626 = x26 & n336;
  assign n3627 = x25 & n338;
  assign n3628 = ~n3626 & ~n3627;
  assign n3629 = n3625 & n3628;
  assign n3637 = n3636 ^ n3629;
  assign n3622 = x2 & x63;
  assign n3638 = n3637 ^ n3622;
  assign n3662 = n3661 ^ n3638;
  assign n3613 = ~x10 & n1962;
  assign n3614 = ~x9 & n1966;
  assign n3615 = ~n3613 & ~n3614;
  assign n3616 = x10 & n1969;
  assign n3617 = x9 & n1971;
  assign n3618 = ~n3616 & ~n3617;
  assign n3619 = n3615 & n3618;
  assign n3606 = ~x22 & n591;
  assign n3607 = ~x21 & n595;
  assign n3608 = ~n3606 & ~n3607;
  assign n3609 = x22 & n598;
  assign n3610 = x21 & n600;
  assign n3611 = ~n3609 & ~n3610;
  assign n3612 = n3608 & n3611;
  assign n3620 = n3619 ^ n3612;
  assign n3599 = ~x8 & n2406;
  assign n3600 = ~x7 & n2408;
  assign n3601 = ~n3599 & ~n3600;
  assign n3602 = x8 & n2399;
  assign n3603 = x7 & n2403;
  assign n3604 = ~n3602 & ~n3603;
  assign n3605 = n3601 & n3604;
  assign n3621 = n3620 ^ n3605;
  assign n3663 = n3662 ^ n3621;
  assign n3716 = n3715 ^ n3663;
  assign n3721 = n3720 ^ n3716;
  assign n3725 = n3724 ^ n3721;
  assign n3729 = n3728 ^ n3725;
  assign n3593 = n3406 ^ n3399;
  assign n3594 = n3406 ^ n3402;
  assign n3595 = n3593 & ~n3594;
  assign n3596 = n3595 ^ n3399;
  assign n3588 = n3390 ^ n3382;
  assign n3589 = ~n3386 & n3588;
  assign n3590 = n3589 ^ n3390;
  assign n3585 = n3377 ^ n3373;
  assign n3586 = ~n3374 & n3585;
  assign n3587 = n3586 ^ x33;
  assign n3591 = n3590 ^ n3587;
  assign n3581 = n3450 ^ n3443;
  assign n3582 = ~n3458 & n3581;
  assign n3583 = n3582 ^ n3443;
  assign n3577 = n3473 ^ n3466;
  assign n3578 = ~n3481 & n3577;
  assign n3579 = n3578 ^ n3466;
  assign n3574 = n3434 ^ n3420;
  assign n3575 = n3435 & ~n3574;
  assign n3576 = n3575 ^ n3427;
  assign n3580 = n3579 ^ n3576;
  assign n3584 = n3583 ^ n3580;
  assign n3592 = n3591 ^ n3584;
  assign n3597 = n3596 ^ n3592;
  assign n3569 = n3459 ^ n3436;
  assign n3570 = n3482 ^ n3436;
  assign n3571 = n3569 & ~n3570;
  assign n3572 = n3571 ^ n3459;
  assign n3565 = n3524 ^ n3507;
  assign n3566 = n3529 & ~n3565;
  assign n3567 = n3566 ^ n3507;
  assign n3561 = n3515 ^ n3508;
  assign n3562 = ~n3523 & ~n3561;
  assign n3563 = n3562 ^ n3508;
  assign n3557 = x35 ^ x31;
  assign n3558 = n85 & n3557;
  assign n3559 = ~n82 & ~n3558;
  assign n3560 = n3559 ^ x33;
  assign n3564 = n3563 ^ n3560;
  assign n3568 = n3567 ^ n3564;
  assign n3573 = n3572 ^ n3568;
  assign n3598 = n3597 ^ n3573;
  assign n3730 = n3729 ^ n3598;
  assign n3734 = n3733 ^ n3730;
  assign n3738 = n3737 ^ n3734;
  assign n3742 = n3741 ^ n3738;
  assign n3923 = n3741 ^ n3734;
  assign n3924 = ~n3738 & ~n3923;
  assign n3925 = n3924 ^ n3741;
  assign n3919 = n3733 ^ n3729;
  assign n3920 = n3730 & n3919;
  assign n3921 = n3920 ^ n3598;
  assign n3914 = n3728 ^ n3721;
  assign n3915 = n3728 ^ n3724;
  assign n3916 = ~n3914 & ~n3915;
  assign n3917 = n3916 ^ n3721;
  assign n3909 = n3592 ^ n3573;
  assign n3910 = n3597 & ~n3909;
  assign n3911 = n3910 ^ n3573;
  assign n3905 = n3720 ^ n3715;
  assign n3906 = ~n3716 & ~n3905;
  assign n3907 = n3906 ^ n3663;
  assign n3900 = n3563 ^ n3559;
  assign n3901 = ~n3560 & ~n3900;
  assign n3902 = n3901 ^ x33;
  assign n3896 = n3583 ^ n3579;
  assign n3897 = n3580 & ~n3896;
  assign n3898 = n3897 ^ n3576;
  assign n3892 = n3629 ^ n3622;
  assign n3893 = ~n3637 & ~n3892;
  assign n3894 = n3893 ^ n3622;
  assign n3884 = x5 & n3105;
  assign n3885 = x4 & n3107;
  assign n3886 = ~n3884 & ~n3885;
  assign n3887 = ~x5 & n3098;
  assign n3888 = ~x4 & n3102;
  assign n3889 = ~n3887 & ~n3888;
  assign n3890 = n3886 & n3889;
  assign n3891 = n3890 ^ n3559;
  assign n3895 = n3894 ^ n3891;
  assign n3899 = n3898 ^ n3895;
  assign n3903 = n3902 ^ n3899;
  assign n3878 = n3700 ^ n3693;
  assign n3879 = ~n3708 & n3878;
  assign n3880 = n3879 ^ n3693;
  assign n3869 = ~x19 & n1000;
  assign n3870 = ~x18 & n1004;
  assign n3871 = ~n3869 & ~n3870;
  assign n3872 = x19 & n1007;
  assign n3873 = x18 & n1009;
  assign n3874 = ~n3872 & ~n3873;
  assign n3875 = n3871 & n3874;
  assign n3868 = x3 & x63;
  assign n3876 = n3875 ^ n3868;
  assign n3861 = ~x17 & n1241;
  assign n3862 = ~x16 & n1243;
  assign n3863 = ~n3861 & ~n3862;
  assign n3864 = x17 & n1234;
  assign n3865 = x16 & n1238;
  assign n3866 = ~n3864 & ~n3865;
  assign n3867 = n3863 & n3866;
  assign n3877 = n3876 ^ n3867;
  assign n3881 = n3880 ^ n3877;
  assign n3852 = x31 & n153;
  assign n3853 = x30 & n155;
  assign n3854 = ~n3852 & ~n3853;
  assign n3855 = ~x31 & n146;
  assign n3856 = ~x30 & n150;
  assign n3857 = ~n3855 & ~n3856;
  assign n3858 = n3854 & n3857;
  assign n3851 = ~n82 & ~n86;
  assign n3859 = n3858 ^ n3851;
  assign n3844 = x27 & n336;
  assign n3845 = x26 & n338;
  assign n3846 = ~n3844 & ~n3845;
  assign n3847 = ~x27 & n329;
  assign n3848 = ~x26 & n333;
  assign n3849 = ~n3847 & ~n3848;
  assign n3850 = n3846 & n3849;
  assign n3860 = n3859 ^ n3850;
  assign n3882 = n3881 ^ n3860;
  assign n3833 = ~x15 & n1396;
  assign n3834 = ~x14 & n1400;
  assign n3835 = ~n3833 & ~n3834;
  assign n3836 = x15 & n1403;
  assign n3837 = x14 & n1405;
  assign n3838 = ~n3836 & ~n3837;
  assign n3839 = n3835 & n3838;
  assign n3826 = ~x25 & n437;
  assign n3827 = ~x24 & n439;
  assign n3828 = ~n3826 & ~n3827;
  assign n3829 = x25 & n430;
  assign n3830 = x24 & n434;
  assign n3831 = ~n3829 & ~n3830;
  assign n3832 = n3828 & n3831;
  assign n3840 = n3839 ^ n3832;
  assign n3819 = ~x13 & n1687;
  assign n3820 = ~x12 & n1691;
  assign n3821 = ~n3819 & ~n3820;
  assign n3822 = x13 & n1694;
  assign n3823 = x12 & n1696;
  assign n3824 = ~n3822 & ~n3823;
  assign n3825 = n3821 & n3824;
  assign n3841 = n3840 ^ n3825;
  assign n3810 = x9 & n2399;
  assign n3811 = x8 & n2403;
  assign n3812 = ~n3810 & ~n3811;
  assign n3813 = ~x9 & n2406;
  assign n3814 = ~x8 & n2408;
  assign n3815 = ~n3813 & ~n3814;
  assign n3816 = n3812 & n3815;
  assign n3803 = ~x21 & n787;
  assign n3804 = ~x20 & n789;
  assign n3805 = ~n3803 & ~n3804;
  assign n3806 = x21 & n780;
  assign n3807 = x20 & n784;
  assign n3808 = ~n3806 & ~n3807;
  assign n3809 = n3805 & n3808;
  assign n3817 = n3816 ^ n3809;
  assign n3796 = ~x7 & n2681;
  assign n3797 = ~x6 & n2685;
  assign n3798 = ~n3796 & ~n3797;
  assign n3799 = x7 & n2688;
  assign n3800 = x6 & n2690;
  assign n3801 = ~n3799 & ~n3800;
  assign n3802 = n3798 & n3801;
  assign n3818 = n3817 ^ n3802;
  assign n3842 = n3841 ^ n3818;
  assign n3787 = x23 & n598;
  assign n3788 = x22 & n600;
  assign n3789 = ~n3787 & ~n3788;
  assign n3790 = ~x23 & n591;
  assign n3791 = ~x22 & n595;
  assign n3792 = ~n3790 & ~n3791;
  assign n3793 = n3789 & n3792;
  assign n3780 = ~x29 & n210;
  assign n3781 = ~x28 & n214;
  assign n3782 = ~n3780 & ~n3781;
  assign n3783 = x29 & n217;
  assign n3784 = x28 & n219;
  assign n3785 = ~n3783 & ~n3784;
  assign n3786 = n3782 & n3785;
  assign n3794 = n3793 ^ n3786;
  assign n3773 = x11 & n1969;
  assign n3774 = x10 & n1971;
  assign n3775 = ~n3773 & ~n3774;
  assign n3776 = ~x11 & n1962;
  assign n3777 = ~x10 & n1966;
  assign n3778 = ~n3776 & ~n3777;
  assign n3779 = n3775 & n3778;
  assign n3795 = n3794 ^ n3779;
  assign n3843 = n3842 ^ n3795;
  assign n3883 = n3882 ^ n3843;
  assign n3904 = n3903 ^ n3883;
  assign n3908 = n3907 ^ n3904;
  assign n3912 = n3911 ^ n3908;
  assign n3768 = n3587 ^ n3584;
  assign n3769 = n3591 & ~n3768;
  assign n3770 = n3769 ^ n3584;
  assign n3764 = n3572 ^ n3564;
  assign n3765 = n3572 ^ n3567;
  assign n3766 = n3764 & ~n3765;
  assign n3767 = n3766 ^ n3564;
  assign n3771 = n3770 ^ n3767;
  assign n3759 = n3709 ^ n3686;
  assign n3760 = n3713 ^ n3686;
  assign n3761 = n3759 & ~n3760;
  assign n3762 = n3761 ^ n3709;
  assign n3754 = n3638 ^ n3621;
  assign n3755 = n3661 ^ n3621;
  assign n3756 = ~n3754 & ~n3755;
  assign n3757 = n3756 ^ n3638;
  assign n3750 = n3619 ^ n3605;
  assign n3751 = n3620 & ~n3750;
  assign n3752 = n3751 ^ n3612;
  assign n3746 = n3684 ^ n3670;
  assign n3747 = n3685 & ~n3746;
  assign n3748 = n3747 ^ n3677;
  assign n3743 = n3652 ^ n3645;
  assign n3744 = ~n3660 & n3743;
  assign n3745 = n3744 ^ n3645;
  assign n3749 = n3748 ^ n3745;
  assign n3753 = n3752 ^ n3749;
  assign n3758 = n3757 ^ n3753;
  assign n3763 = n3762 ^ n3758;
  assign n3772 = n3771 ^ n3763;
  assign n3913 = n3912 ^ n3772;
  assign n3918 = n3917 ^ n3913;
  assign n3922 = n3921 ^ n3918;
  assign n3926 = n3925 ^ n3922;
  assign n4103 = n3925 ^ n3918;
  assign n4104 = n3922 & ~n4103;
  assign n4105 = n4104 ^ n3925;
  assign n4099 = n3917 ^ n3912;
  assign n4100 = ~n3913 & n4099;
  assign n4101 = n4100 ^ n3772;
  assign n4095 = n3911 ^ n3907;
  assign n4096 = n3908 & n4095;
  assign n4097 = n4096 ^ n3904;
  assign n4090 = n3767 ^ n3763;
  assign n4091 = ~n3771 & ~n4090;
  assign n4092 = n4091 ^ n3763;
  assign n4086 = n3903 ^ n3882;
  assign n4087 = n3883 & n4086;
  assign n4088 = n4087 ^ n3843;
  assign n4081 = n3902 ^ n3895;
  assign n4082 = n3902 ^ n3898;
  assign n4083 = ~n4081 & ~n4082;
  assign n4084 = n4083 ^ n3895;
  assign n4077 = n3818 ^ n3795;
  assign n4078 = ~n3842 & n4077;
  assign n4079 = n4078 ^ n3795;
  assign n4066 = ~x24 & n591;
  assign n4067 = ~x23 & n595;
  assign n4068 = ~n4066 & ~n4067;
  assign n4069 = x24 & n598;
  assign n4070 = x23 & n600;
  assign n4071 = ~n4069 & ~n4070;
  assign n4072 = n4068 & n4071;
  assign n4059 = ~x16 & n1396;
  assign n4060 = ~x15 & n1400;
  assign n4061 = ~n4059 & ~n4060;
  assign n4062 = x16 & n1403;
  assign n4063 = x15 & n1405;
  assign n4064 = ~n4062 & ~n4063;
  assign n4065 = n4061 & n4064;
  assign n4073 = n4072 ^ n4065;
  assign n4052 = x14 & n1694;
  assign n4053 = x13 & n1696;
  assign n4054 = ~n4052 & ~n4053;
  assign n4055 = ~x14 & n1687;
  assign n4056 = ~x13 & n1691;
  assign n4057 = ~n4055 & ~n4056;
  assign n4058 = n4054 & n4057;
  assign n4074 = n4073 ^ n4058;
  assign n4043 = x8 & n2688;
  assign n4044 = x7 & n2690;
  assign n4045 = ~n4043 & ~n4044;
  assign n4046 = ~x8 & n2681;
  assign n4047 = ~x7 & n2685;
  assign n4048 = ~n4046 & ~n4047;
  assign n4049 = n4045 & n4048;
  assign n4036 = x10 & n2399;
  assign n4037 = x9 & n2403;
  assign n4038 = ~n4036 & ~n4037;
  assign n4039 = ~x10 & n2406;
  assign n4040 = ~x9 & n2408;
  assign n4041 = ~n4039 & ~n4040;
  assign n4042 = n4038 & n4041;
  assign n4050 = n4049 ^ n4042;
  assign n4029 = ~x20 & n1000;
  assign n4030 = ~x19 & n1004;
  assign n4031 = ~n4029 & ~n4030;
  assign n4032 = x20 & n1007;
  assign n4033 = x19 & n1009;
  assign n4034 = ~n4032 & ~n4033;
  assign n4035 = n4031 & n4034;
  assign n4051 = n4050 ^ n4035;
  assign n4075 = n4074 ^ n4051;
  assign n4020 = ~x12 & n1962;
  assign n4021 = ~x11 & n1966;
  assign n4022 = ~n4020 & ~n4021;
  assign n4023 = x12 & n1969;
  assign n4024 = x11 & n1971;
  assign n4025 = ~n4023 & ~n4024;
  assign n4026 = n4022 & n4025;
  assign n4013 = ~x28 & n329;
  assign n4014 = ~x27 & n333;
  assign n4015 = ~n4013 & ~n4014;
  assign n4016 = x28 & n336;
  assign n4017 = x27 & n338;
  assign n4018 = ~n4016 & ~n4017;
  assign n4019 = n4015 & n4018;
  assign n4027 = n4026 ^ n4019;
  assign n4006 = x22 & n780;
  assign n4007 = x21 & n784;
  assign n4008 = ~n4006 & ~n4007;
  assign n4009 = ~x22 & n787;
  assign n4010 = ~x21 & n789;
  assign n4011 = ~n4009 & ~n4010;
  assign n4012 = n4008 & n4011;
  assign n4028 = n4027 ^ n4012;
  assign n4076 = n4075 ^ n4028;
  assign n4080 = n4079 ^ n4076;
  assign n4085 = n4084 ^ n4080;
  assign n4089 = n4088 ^ n4085;
  assign n4093 = n4092 ^ n4089;
  assign n4001 = n3762 ^ n3757;
  assign n4002 = ~n3758 & n4001;
  assign n4003 = n4002 ^ n3753;
  assign n3997 = n3894 ^ n3890;
  assign n3998 = n3891 & n3997;
  assign n3999 = n3998 ^ n3559;
  assign n3992 = n3752 ^ n3745;
  assign n3993 = n3752 ^ n3748;
  assign n3994 = n3992 & ~n3993;
  assign n3995 = n3994 ^ n3745;
  assign n3983 = x6 & n3105;
  assign n3984 = x5 & n3107;
  assign n3985 = ~n3983 & ~n3984;
  assign n3986 = ~x6 & n3098;
  assign n3987 = ~x5 & n3102;
  assign n3988 = ~n3986 & ~n3987;
  assign n3989 = n3985 & n3988;
  assign n3982 = x4 & x63;
  assign n3990 = n3989 ^ n3982;
  assign n3979 = x37 ^ x31;
  assign n3980 = n149 & n3979;
  assign n3981 = ~n146 & ~n3980;
  assign n3991 = n3990 ^ n3981;
  assign n3996 = n3995 ^ n3991;
  assign n4000 = n3999 ^ n3996;
  assign n4004 = n4003 ^ n4000;
  assign n3973 = n3877 ^ n3860;
  assign n3974 = n3880 ^ n3860;
  assign n3975 = n3973 & n3974;
  assign n3976 = n3975 ^ n3877;
  assign n3968 = n3832 ^ n3825;
  assign n3969 = n3839 ^ n3825;
  assign n3970 = n3968 & ~n3969;
  assign n3971 = n3970 ^ n3832;
  assign n3963 = n3868 ^ n3867;
  assign n3964 = n3875 ^ n3867;
  assign n3965 = ~n3963 & ~n3964;
  assign n3966 = n3965 ^ n3868;
  assign n3959 = n3851 ^ n3850;
  assign n3960 = n3858 ^ n3850;
  assign n3961 = ~n3959 & ~n3960;
  assign n3962 = n3961 ^ n3851;
  assign n3967 = n3966 ^ n3962;
  assign n3972 = n3971 ^ n3967;
  assign n3977 = n3976 ^ n3972;
  assign n3953 = n3809 ^ n3802;
  assign n3954 = n3816 ^ n3802;
  assign n3955 = n3953 & ~n3954;
  assign n3956 = n3955 ^ n3809;
  assign n3950 = n3793 ^ n3779;
  assign n3951 = n3794 & ~n3950;
  assign n3952 = n3951 ^ n3786;
  assign n3957 = n3956 ^ n3952;
  assign n3941 = ~x30 & n210;
  assign n3942 = ~x29 & n214;
  assign n3943 = ~n3941 & ~n3942;
  assign n3944 = x30 & n217;
  assign n3945 = x29 & n219;
  assign n3946 = ~n3944 & ~n3945;
  assign n3947 = n3943 & n3946;
  assign n3934 = ~x26 & n437;
  assign n3935 = ~x25 & n439;
  assign n3936 = ~n3934 & ~n3935;
  assign n3937 = x26 & n430;
  assign n3938 = x25 & n434;
  assign n3939 = ~n3937 & ~n3938;
  assign n3940 = n3936 & n3939;
  assign n3948 = n3947 ^ n3940;
  assign n3927 = x18 & n1234;
  assign n3928 = x17 & n1238;
  assign n3929 = ~n3927 & ~n3928;
  assign n3930 = ~x18 & n1241;
  assign n3931 = ~x17 & n1243;
  assign n3932 = ~n3930 & ~n3931;
  assign n3933 = n3929 & n3932;
  assign n3949 = n3948 ^ n3933;
  assign n3958 = n3957 ^ n3949;
  assign n3978 = n3977 ^ n3958;
  assign n4005 = n4004 ^ n3978;
  assign n4094 = n4093 ^ n4005;
  assign n4098 = n4097 ^ n4094;
  assign n4102 = n4101 ^ n4098;
  assign n4106 = n4105 ^ n4102;
  assign n4277 = n4105 ^ n4098;
  assign n4278 = n4102 & ~n4277;
  assign n4279 = n4278 ^ n4105;
  assign n4273 = n4097 ^ n4093;
  assign n4274 = ~n4094 & n4273;
  assign n4275 = n4274 ^ n4005;
  assign n4269 = n4092 ^ n4088;
  assign n4270 = ~n4089 & n4269;
  assign n4271 = n4270 ^ n4085;
  assign n4263 = n4000 ^ n3978;
  assign n4264 = n4003 ^ n3978;
  assign n4265 = ~n4263 & n4264;
  assign n4266 = n4265 ^ n4000;
  assign n4259 = n4084 ^ n4079;
  assign n4260 = n4080 & n4259;
  assign n4261 = n4260 ^ n4076;
  assign n4253 = n3971 ^ n3962;
  assign n4254 = n3971 ^ n3966;
  assign n4255 = ~n4253 & n4254;
  assign n4256 = n4255 ^ n3962;
  assign n4248 = n3982 ^ n3981;
  assign n4249 = n3989 ^ n3981;
  assign n4250 = n4248 & n4249;
  assign n4251 = n4250 ^ n3982;
  assign n4239 = x13 & n1969;
  assign n4240 = x12 & n1971;
  assign n4241 = ~n4239 & ~n4240;
  assign n4242 = ~x13 & n1962;
  assign n4243 = ~x12 & n1966;
  assign n4244 = ~n4242 & ~n4243;
  assign n4245 = n4241 & n4244;
  assign n4232 = ~x15 & n1687;
  assign n4233 = ~x14 & n1691;
  assign n4234 = ~n4232 & ~n4233;
  assign n4235 = x15 & n1694;
  assign n4236 = x14 & n1696;
  assign n4237 = ~n4235 & ~n4236;
  assign n4238 = n4234 & n4237;
  assign n4246 = n4245 ^ n4238;
  assign n4225 = ~x29 & n329;
  assign n4226 = ~x28 & n333;
  assign n4227 = ~n4225 & ~n4226;
  assign n4228 = x29 & n336;
  assign n4229 = x28 & n338;
  assign n4230 = ~n4228 & ~n4229;
  assign n4231 = n4227 & n4230;
  assign n4247 = n4246 ^ n4231;
  assign n4252 = n4251 ^ n4247;
  assign n4257 = n4256 ^ n4252;
  assign n4220 = n4051 ^ n4028;
  assign n4221 = n4074 ^ n4028;
  assign n4222 = n4220 & ~n4221;
  assign n4223 = n4222 ^ n4051;
  assign n4209 = ~x7 & n3098;
  assign n4210 = ~x6 & n3102;
  assign n4211 = ~n4209 & ~n4210;
  assign n4212 = x7 & n3105;
  assign n4213 = x6 & n3107;
  assign n4214 = ~n4212 & ~n4213;
  assign n4215 = n4211 & n4214;
  assign n4202 = ~x21 & n1000;
  assign n4203 = ~x20 & n1004;
  assign n4204 = ~n4202 & ~n4203;
  assign n4205 = x21 & n1007;
  assign n4206 = x20 & n1009;
  assign n4207 = ~n4205 & ~n4206;
  assign n4208 = n4204 & n4207;
  assign n4216 = n4215 ^ n4208;
  assign n4201 = x5 & x63;
  assign n4217 = n4216 ^ n4201;
  assign n4192 = ~x31 & n210;
  assign n4193 = ~x30 & n214;
  assign n4194 = ~n4192 & ~n4193;
  assign n4195 = x31 & n217;
  assign n4196 = x30 & n219;
  assign n4197 = ~n4195 & ~n4196;
  assign n4198 = n4194 & n4197;
  assign n4191 = ~n146 & ~n150;
  assign n4199 = n4198 ^ n4191;
  assign n4184 = ~x27 & n437;
  assign n4185 = ~x26 & n439;
  assign n4186 = ~n4184 & ~n4185;
  assign n4187 = x27 & n430;
  assign n4188 = x26 & n434;
  assign n4189 = ~n4187 & ~n4188;
  assign n4190 = n4186 & n4189;
  assign n4200 = n4199 ^ n4190;
  assign n4218 = n4217 ^ n4200;
  assign n4175 = ~x11 & n2406;
  assign n4176 = ~x10 & n2408;
  assign n4177 = ~n4175 & ~n4176;
  assign n4178 = x11 & n2399;
  assign n4179 = x10 & n2403;
  assign n4180 = ~n4178 & ~n4179;
  assign n4181 = n4177 & n4180;
  assign n4168 = ~x23 & n787;
  assign n4169 = ~x22 & n789;
  assign n4170 = ~n4168 & ~n4169;
  assign n4171 = x23 & n780;
  assign n4172 = x22 & n784;
  assign n4173 = ~n4171 & ~n4172;
  assign n4174 = n4170 & n4173;
  assign n4182 = n4181 ^ n4174;
  assign n4161 = ~x9 & n2681;
  assign n4162 = ~x8 & n2685;
  assign n4163 = ~n4161 & ~n4162;
  assign n4164 = x9 & n2688;
  assign n4165 = x8 & n2690;
  assign n4166 = ~n4164 & ~n4165;
  assign n4167 = n4163 & n4166;
  assign n4183 = n4182 ^ n4167;
  assign n4219 = n4218 ^ n4183;
  assign n4224 = n4223 ^ n4219;
  assign n4258 = n4257 ^ n4224;
  assign n4262 = n4261 ^ n4258;
  assign n4267 = n4266 ^ n4262;
  assign n4156 = n3972 ^ n3958;
  assign n4157 = n3977 & n4156;
  assign n4158 = n4157 ^ n3958;
  assign n4152 = n3999 ^ n3991;
  assign n4153 = n3999 ^ n3995;
  assign n4154 = n4152 & ~n4153;
  assign n4155 = n4154 ^ n3991;
  assign n4159 = n4158 ^ n4155;
  assign n4148 = n3952 ^ n3949;
  assign n4149 = ~n3957 & n4148;
  assign n4150 = n4149 ^ n3949;
  assign n4143 = n4072 ^ n4058;
  assign n4144 = n4073 & ~n4143;
  assign n4145 = n4144 ^ n4065;
  assign n4139 = n3947 ^ n3933;
  assign n4140 = n3948 & ~n4139;
  assign n4141 = n4140 ^ n3940;
  assign n4142 = n4141 ^ n3981;
  assign n4146 = n4145 ^ n4142;
  assign n4133 = n4019 ^ n4012;
  assign n4134 = n4026 ^ n4012;
  assign n4135 = n4133 & ~n4134;
  assign n4136 = n4135 ^ n4019;
  assign n4130 = n4042 ^ n4035;
  assign n4131 = ~n4050 & n4130;
  assign n4132 = n4131 ^ n4035;
  assign n4137 = n4136 ^ n4132;
  assign n4121 = x17 & n1403;
  assign n4122 = x16 & n1405;
  assign n4123 = ~n4121 & ~n4122;
  assign n4124 = ~x17 & n1396;
  assign n4125 = ~x16 & n1400;
  assign n4126 = ~n4124 & ~n4125;
  assign n4127 = n4123 & n4126;
  assign n4114 = ~x19 & n1241;
  assign n4115 = ~x18 & n1243;
  assign n4116 = ~n4114 & ~n4115;
  assign n4117 = x19 & n1234;
  assign n4118 = x18 & n1238;
  assign n4119 = ~n4117 & ~n4118;
  assign n4120 = n4116 & n4119;
  assign n4128 = n4127 ^ n4120;
  assign n4107 = ~x25 & n591;
  assign n4108 = ~x24 & n595;
  assign n4109 = ~n4107 & ~n4108;
  assign n4110 = x25 & n598;
  assign n4111 = x24 & n600;
  assign n4112 = ~n4110 & ~n4111;
  assign n4113 = n4109 & n4112;
  assign n4129 = n4128 ^ n4113;
  assign n4138 = n4137 ^ n4129;
  assign n4147 = n4146 ^ n4138;
  assign n4151 = n4150 ^ n4147;
  assign n4160 = n4159 ^ n4151;
  assign n4268 = n4267 ^ n4160;
  assign n4272 = n4271 ^ n4268;
  assign n4276 = n4275 ^ n4272;
  assign n4280 = n4279 ^ n4276;
  assign n4440 = n4279 ^ n4272;
  assign n4441 = ~n4276 & n4440;
  assign n4442 = n4441 ^ n4279;
  assign n4436 = n4271 ^ n4267;
  assign n4437 = n4268 & n4436;
  assign n4438 = n4437 ^ n4160;
  assign n4432 = n4266 ^ n4261;
  assign n4433 = n4262 & ~n4432;
  assign n4434 = n4433 ^ n4258;
  assign n4428 = n4155 ^ n4151;
  assign n4429 = ~n4159 & n4428;
  assign n4430 = n4429 ^ n4151;
  assign n4423 = n4257 ^ n4223;
  assign n4424 = n4224 & ~n4423;
  assign n4425 = n4424 ^ n4219;
  assign n4419 = n4256 ^ n4251;
  assign n4420 = ~n4252 & ~n4419;
  assign n4421 = n4420 ^ n4247;
  assign n4414 = n4200 ^ n4183;
  assign n4415 = n4217 ^ n4183;
  assign n4416 = ~n4414 & n4415;
  assign n4417 = n4416 ^ n4200;
  assign n4409 = n4208 ^ n4201;
  assign n4410 = ~n4216 & ~n4409;
  assign n4411 = n4410 ^ n4201;
  assign n4400 = ~x8 & n3098;
  assign n4401 = ~x7 & n3102;
  assign n4402 = ~n4400 & ~n4401;
  assign n4403 = x8 & n3105;
  assign n4404 = x7 & n3107;
  assign n4405 = ~n4403 & ~n4404;
  assign n4406 = n4402 & n4405;
  assign n4393 = ~x28 & n437;
  assign n4394 = ~x27 & n439;
  assign n4395 = ~n4393 & ~n4394;
  assign n4396 = x28 & n430;
  assign n4397 = x27 & n434;
  assign n4398 = ~n4396 & ~n4397;
  assign n4399 = n4395 & n4398;
  assign n4407 = n4406 ^ n4399;
  assign n4392 = x6 & x63;
  assign n4408 = n4407 ^ n4392;
  assign n4412 = n4411 ^ n4408;
  assign n4383 = ~x18 & n1396;
  assign n4384 = ~x17 & n1400;
  assign n4385 = ~n4383 & ~n4384;
  assign n4386 = x18 & n1403;
  assign n4387 = x17 & n1405;
  assign n4388 = ~n4386 & ~n4387;
  assign n4389 = n4385 & n4388;
  assign n4376 = ~x26 & n591;
  assign n4377 = ~x25 & n595;
  assign n4378 = ~n4376 & ~n4377;
  assign n4379 = x26 & n598;
  assign n4380 = x25 & n600;
  assign n4381 = ~n4379 & ~n4380;
  assign n4382 = n4378 & n4381;
  assign n4390 = n4389 ^ n4382;
  assign n4369 = ~x16 & n1687;
  assign n4370 = ~x15 & n1691;
  assign n4371 = ~n4369 & ~n4370;
  assign n4372 = x16 & n1694;
  assign n4373 = x15 & n1696;
  assign n4374 = ~n4372 & ~n4373;
  assign n4375 = n4371 & n4374;
  assign n4391 = n4390 ^ n4375;
  assign n4413 = n4412 ^ n4391;
  assign n4418 = n4417 ^ n4413;
  assign n4422 = n4421 ^ n4418;
  assign n4426 = n4425 ^ n4422;
  assign n4364 = n4150 ^ n4146;
  assign n4365 = n4147 & ~n4364;
  assign n4366 = n4365 ^ n4138;
  assign n4359 = n4174 ^ n4167;
  assign n4360 = ~n4182 & n4359;
  assign n4361 = n4360 ^ n4167;
  assign n4351 = ~x20 & n1241;
  assign n4352 = ~x19 & n1243;
  assign n4353 = ~n4351 & ~n4352;
  assign n4354 = x20 & n1234;
  assign n4355 = x19 & n1238;
  assign n4356 = ~n4354 & ~n4355;
  assign n4357 = n4353 & n4356;
  assign n4344 = ~x30 & n329;
  assign n4345 = ~x29 & n333;
  assign n4346 = ~n4344 & ~n4345;
  assign n4347 = x30 & n336;
  assign n4348 = x29 & n338;
  assign n4349 = ~n4347 & ~n4348;
  assign n4350 = n4346 & n4349;
  assign n4358 = n4357 ^ n4350;
  assign n4362 = n4361 ^ n4358;
  assign n4334 = ~x14 & n1962;
  assign n4335 = ~x13 & n1966;
  assign n4336 = ~n4334 & ~n4335;
  assign n4337 = x14 & n1969;
  assign n4338 = x13 & n1971;
  assign n4339 = ~n4337 & ~n4338;
  assign n4340 = n4336 & n4339;
  assign n4327 = ~x24 & n787;
  assign n4328 = ~x23 & n789;
  assign n4329 = ~n4327 & ~n4328;
  assign n4330 = x24 & n780;
  assign n4331 = x23 & n784;
  assign n4332 = ~n4330 & ~n4331;
  assign n4333 = n4329 & n4332;
  assign n4341 = n4340 ^ n4333;
  assign n4320 = x12 & n2399;
  assign n4321 = x11 & n2403;
  assign n4322 = ~n4320 & ~n4321;
  assign n4323 = ~x12 & n2406;
  assign n4324 = ~x11 & n2408;
  assign n4325 = ~n4323 & ~n4324;
  assign n4326 = n4322 & n4325;
  assign n4342 = n4341 ^ n4326;
  assign n4311 = ~x22 & n1000;
  assign n4312 = ~x21 & n1004;
  assign n4313 = ~n4311 & ~n4312;
  assign n4314 = x22 & n1007;
  assign n4315 = x21 & n1009;
  assign n4316 = ~n4314 & ~n4315;
  assign n4317 = n4313 & n4316;
  assign n4308 = x39 ^ x31;
  assign n4309 = n213 & n4308;
  assign n4310 = ~n210 & ~n4309;
  assign n4318 = n4317 ^ n4310;
  assign n4301 = ~x10 & n2681;
  assign n4302 = ~x9 & n2685;
  assign n4303 = ~n4301 & ~n4302;
  assign n4304 = x10 & n2688;
  assign n4305 = x9 & n2690;
  assign n4306 = ~n4304 & ~n4305;
  assign n4307 = n4303 & n4306;
  assign n4319 = n4318 ^ n4307;
  assign n4343 = n4342 ^ n4319;
  assign n4363 = n4362 ^ n4343;
  assign n4367 = n4366 ^ n4363;
  assign n4297 = n4132 ^ n4129;
  assign n4298 = ~n4137 & n4297;
  assign n4299 = n4298 ^ n4129;
  assign n4293 = n4145 ^ n4141;
  assign n4294 = n4142 & ~n4293;
  assign n4295 = n4294 ^ n3981;
  assign n4289 = n4245 ^ n4231;
  assign n4290 = n4246 & ~n4289;
  assign n4291 = n4290 ^ n4238;
  assign n4285 = n4120 ^ n4113;
  assign n4286 = ~n4128 & n4285;
  assign n4287 = n4286 ^ n4113;
  assign n4281 = n4191 ^ n4190;
  assign n4282 = n4198 ^ n4190;
  assign n4283 = ~n4281 & ~n4282;
  assign n4284 = n4283 ^ n4191;
  assign n4288 = n4287 ^ n4284;
  assign n4292 = n4291 ^ n4288;
  assign n4296 = n4295 ^ n4292;
  assign n4300 = n4299 ^ n4296;
  assign n4368 = n4367 ^ n4300;
  assign n4427 = n4426 ^ n4368;
  assign n4431 = n4430 ^ n4427;
  assign n4435 = n4434 ^ n4431;
  assign n4439 = n4438 ^ n4435;
  assign n4443 = n4442 ^ n4439;
  assign n4599 = n4442 ^ n4435;
  assign n4600 = n4439 & n4599;
  assign n4601 = n4600 ^ n4442;
  assign n4595 = n4434 ^ n4430;
  assign n4596 = ~n4431 & ~n4595;
  assign n4597 = n4596 ^ n4427;
  assign n4590 = n4422 ^ n4368;
  assign n4591 = n4425 ^ n4368;
  assign n4592 = ~n4590 & ~n4591;
  assign n4593 = n4592 ^ n4422;
  assign n4585 = n4363 ^ n4300;
  assign n4586 = n4366 ^ n4300;
  assign n4587 = n4585 & n4586;
  assign n4588 = n4587 ^ n4363;
  assign n4580 = n4421 ^ n4417;
  assign n4581 = ~n4418 & n4580;
  assign n4582 = n4581 ^ n4413;
  assign n4575 = n4408 ^ n4391;
  assign n4576 = ~n4412 & ~n4575;
  assign n4577 = n4576 ^ n4391;
  assign n4570 = n4399 ^ n4392;
  assign n4571 = ~n4407 & ~n4570;
  assign n4572 = n4571 ^ n4392;
  assign n4561 = ~x17 & n1687;
  assign n4562 = ~x16 & n1691;
  assign n4563 = ~n4561 & ~n4562;
  assign n4564 = x17 & n1694;
  assign n4565 = x16 & n1696;
  assign n4566 = ~n4564 & ~n4565;
  assign n4567 = n4563 & n4566;
  assign n4554 = ~x19 & n1396;
  assign n4555 = ~x18 & n1400;
  assign n4556 = ~n4554 & ~n4555;
  assign n4557 = x19 & n1403;
  assign n4558 = x18 & n1405;
  assign n4559 = ~n4557 & ~n4558;
  assign n4560 = n4556 & n4559;
  assign n4568 = n4567 ^ n4560;
  assign n4547 = ~x25 & n787;
  assign n4548 = ~x24 & n789;
  assign n4549 = ~n4547 & ~n4548;
  assign n4550 = x25 & n780;
  assign n4551 = x24 & n784;
  assign n4552 = ~n4550 & ~n4551;
  assign n4553 = n4549 & n4552;
  assign n4569 = n4568 ^ n4553;
  assign n4573 = n4572 ^ n4569;
  assign n4538 = ~x31 & n329;
  assign n4539 = ~x30 & n333;
  assign n4540 = ~n4538 & ~n4539;
  assign n4541 = x31 & n336;
  assign n4542 = x30 & n338;
  assign n4543 = ~n4541 & ~n4542;
  assign n4544 = n4540 & n4543;
  assign n4537 = ~n210 & ~n214;
  assign n4545 = n4544 ^ n4537;
  assign n4530 = x27 & n598;
  assign n4531 = x26 & n600;
  assign n4532 = ~n4530 & ~n4531;
  assign n4533 = ~x27 & n591;
  assign n4534 = ~x26 & n595;
  assign n4535 = ~n4533 & ~n4534;
  assign n4536 = n4532 & n4535;
  assign n4546 = n4545 ^ n4536;
  assign n4574 = n4573 ^ n4546;
  assign n4578 = n4577 ^ n4574;
  assign n4519 = ~x13 & n2406;
  assign n4520 = ~x12 & n2408;
  assign n4521 = ~n4519 & ~n4520;
  assign n4522 = x13 & n2399;
  assign n4523 = x12 & n2403;
  assign n4524 = ~n4522 & ~n4523;
  assign n4525 = n4521 & n4524;
  assign n4512 = x15 & n1969;
  assign n4513 = x14 & n1971;
  assign n4514 = ~n4512 & ~n4513;
  assign n4515 = ~x15 & n1962;
  assign n4516 = ~x14 & n1966;
  assign n4517 = ~n4515 & ~n4516;
  assign n4518 = n4514 & n4517;
  assign n4526 = n4525 ^ n4518;
  assign n4505 = ~x29 & n437;
  assign n4506 = ~x28 & n439;
  assign n4507 = ~n4505 & ~n4506;
  assign n4508 = x29 & n430;
  assign n4509 = x28 & n434;
  assign n4510 = ~n4508 & ~n4509;
  assign n4511 = n4507 & n4510;
  assign n4527 = n4526 ^ n4511;
  assign n4496 = ~x11 & n2681;
  assign n4497 = ~x10 & n2685;
  assign n4498 = ~n4496 & ~n4497;
  assign n4499 = x11 & n2688;
  assign n4500 = x10 & n2690;
  assign n4501 = ~n4499 & ~n4500;
  assign n4502 = n4498 & n4501;
  assign n4489 = x23 & n1007;
  assign n4490 = x22 & n1009;
  assign n4491 = ~n4489 & ~n4490;
  assign n4492 = ~x23 & n1000;
  assign n4493 = ~x22 & n1004;
  assign n4494 = ~n4492 & ~n4493;
  assign n4495 = n4491 & n4494;
  assign n4503 = n4502 ^ n4495;
  assign n4482 = x9 & n3105;
  assign n4483 = x8 & n3107;
  assign n4484 = ~n4482 & ~n4483;
  assign n4485 = ~x9 & n3098;
  assign n4486 = ~x8 & n3102;
  assign n4487 = ~n4485 & ~n4486;
  assign n4488 = n4484 & n4487;
  assign n4504 = n4503 ^ n4488;
  assign n4528 = n4527 ^ n4504;
  assign n4473 = ~x21 & n1241;
  assign n4474 = ~x20 & n1243;
  assign n4475 = ~n4473 & ~n4474;
  assign n4476 = x21 & n1234;
  assign n4477 = x20 & n1238;
  assign n4478 = ~n4476 & ~n4477;
  assign n4479 = n4475 & n4478;
  assign n4472 = x7 & x63;
  assign n4480 = n4479 ^ n4472;
  assign n4481 = n4480 ^ n4350;
  assign n4529 = n4528 ^ n4481;
  assign n4579 = n4578 ^ n4529;
  assign n4583 = n4582 ^ n4579;
  assign n4467 = n4299 ^ n4292;
  assign n4468 = n4299 ^ n4295;
  assign n4469 = ~n4467 & ~n4468;
  assign n4470 = n4469 ^ n4292;
  assign n4463 = n4362 ^ n4342;
  assign n4464 = n4343 & n4463;
  assign n4465 = n4464 ^ n4319;
  assign n4458 = n4291 ^ n4287;
  assign n4459 = ~n4288 & ~n4458;
  assign n4460 = n4459 ^ n4284;
  assign n4455 = n4361 ^ n4357;
  assign n4456 = ~n4358 & ~n4455;
  assign n4457 = n4456 ^ n4350;
  assign n4461 = n4460 ^ n4457;
  assign n4451 = n4317 ^ n4307;
  assign n4452 = n4318 & ~n4451;
  assign n4453 = n4452 ^ n4310;
  assign n4447 = n4382 ^ n4375;
  assign n4448 = ~n4390 & n4447;
  assign n4449 = n4448 ^ n4375;
  assign n4444 = n4333 ^ n4326;
  assign n4445 = ~n4341 & n4444;
  assign n4446 = n4445 ^ n4326;
  assign n4450 = n4449 ^ n4446;
  assign n4454 = n4453 ^ n4450;
  assign n4462 = n4461 ^ n4454;
  assign n4466 = n4465 ^ n4462;
  assign n4471 = n4470 ^ n4466;
  assign n4584 = n4583 ^ n4471;
  assign n4589 = n4588 ^ n4584;
  assign n4594 = n4593 ^ n4589;
  assign n4598 = n4597 ^ n4594;
  assign n4602 = n4601 ^ n4598;
  assign n4751 = n4601 ^ n4594;
  assign n4752 = n4598 & ~n4751;
  assign n4753 = n4752 ^ n4601;
  assign n4746 = n4593 ^ n4588;
  assign n4747 = n4593 ^ n4584;
  assign n4748 = n4746 & n4747;
  assign n4749 = n4748 ^ n4588;
  assign n4741 = n4579 ^ n4471;
  assign n4742 = n4582 ^ n4471;
  assign n4743 = n4741 & n4742;
  assign n4744 = n4743 ^ n4579;
  assign n4736 = n4470 ^ n4462;
  assign n4737 = n4466 & n4736;
  assign n4738 = n4737 ^ n4465;
  assign n4732 = n4574 ^ n4529;
  assign n4733 = ~n4578 & ~n4732;
  assign n4734 = n4733 ^ n4529;
  assign n4728 = n4504 ^ n4481;
  assign n4729 = ~n4528 & ~n4728;
  assign n4730 = n4729 ^ n4481;
  assign n4724 = n4569 ^ n4546;
  assign n4725 = n4573 & ~n4724;
  assign n4726 = n4725 ^ n4546;
  assign n4719 = n4502 ^ n4488;
  assign n4720 = n4503 & ~n4719;
  assign n4721 = n4720 ^ n4495;
  assign n4715 = n4537 ^ n4536;
  assign n4716 = n4544 ^ n4536;
  assign n4717 = ~n4715 & ~n4716;
  assign n4718 = n4717 ^ n4537;
  assign n4722 = n4721 ^ n4718;
  assign n4706 = x28 & n598;
  assign n4707 = x27 & n600;
  assign n4708 = ~n4706 & ~n4707;
  assign n4709 = ~x28 & n591;
  assign n4710 = ~x27 & n595;
  assign n4711 = ~n4709 & ~n4710;
  assign n4712 = n4708 & n4711;
  assign n4705 = x8 & x63;
  assign n4713 = n4712 ^ n4705;
  assign n4698 = ~x20 & n1396;
  assign n4699 = ~x19 & n1400;
  assign n4700 = ~n4698 & ~n4699;
  assign n4701 = x20 & n1403;
  assign n4702 = x19 & n1405;
  assign n4703 = ~n4701 & ~n4702;
  assign n4704 = n4700 & n4703;
  assign n4714 = n4713 ^ n4704;
  assign n4723 = n4722 ^ n4714;
  assign n4727 = n4726 ^ n4723;
  assign n4731 = n4730 ^ n4727;
  assign n4735 = n4734 ^ n4731;
  assign n4739 = n4738 ^ n4735;
  assign n4693 = n4457 ^ n4454;
  assign n4694 = ~n4461 & ~n4693;
  assign n4695 = n4694 ^ n4454;
  assign n4682 = x22 & n1234;
  assign n4683 = x21 & n1238;
  assign n4684 = ~n4682 & ~n4683;
  assign n4685 = ~x22 & n1241;
  assign n4686 = ~x21 & n1243;
  assign n4687 = ~n4685 & ~n4686;
  assign n4688 = n4684 & n4687;
  assign n4679 = x41 ^ x31;
  assign n4680 = n332 & n4679;
  assign n4681 = ~n329 & ~n4680;
  assign n4689 = n4688 ^ n4681;
  assign n4672 = ~x10 & n3098;
  assign n4673 = ~x9 & n3102;
  assign n4674 = ~n4672 & ~n4673;
  assign n4675 = x10 & n3105;
  assign n4676 = x9 & n3107;
  assign n4677 = ~n4675 & ~n4676;
  assign n4678 = n4674 & n4677;
  assign n4690 = n4689 ^ n4678;
  assign n4663 = x26 & n780;
  assign n4664 = x25 & n784;
  assign n4665 = ~n4663 & ~n4664;
  assign n4666 = ~x26 & n787;
  assign n4667 = ~x25 & n789;
  assign n4668 = ~n4666 & ~n4667;
  assign n4669 = n4665 & n4668;
  assign n4656 = ~x18 & n1687;
  assign n4657 = ~x17 & n1691;
  assign n4658 = ~n4656 & ~n4657;
  assign n4659 = x18 & n1694;
  assign n4660 = x17 & n1696;
  assign n4661 = ~n4659 & ~n4660;
  assign n4662 = n4658 & n4661;
  assign n4670 = n4669 ^ n4662;
  assign n4649 = ~x16 & n1962;
  assign n4650 = ~x15 & n1966;
  assign n4651 = ~n4649 & ~n4650;
  assign n4652 = x16 & n1969;
  assign n4653 = x15 & n1971;
  assign n4654 = ~n4652 & ~n4653;
  assign n4655 = n4651 & n4654;
  assign n4671 = n4670 ^ n4655;
  assign n4691 = n4690 ^ n4671;
  assign n4640 = ~x14 & n2406;
  assign n4641 = ~x13 & n2408;
  assign n4642 = ~n4640 & ~n4641;
  assign n4643 = x14 & n2399;
  assign n4644 = x13 & n2403;
  assign n4645 = ~n4643 & ~n4644;
  assign n4646 = n4642 & n4645;
  assign n4633 = ~x24 & n1000;
  assign n4634 = ~x23 & n1004;
  assign n4635 = ~n4633 & ~n4634;
  assign n4636 = x24 & n1007;
  assign n4637 = x23 & n1009;
  assign n4638 = ~n4636 & ~n4637;
  assign n4639 = n4635 & n4638;
  assign n4647 = n4646 ^ n4639;
  assign n4626 = ~x12 & n2681;
  assign n4627 = ~x11 & n2685;
  assign n4628 = ~n4626 & ~n4627;
  assign n4629 = x12 & n2688;
  assign n4630 = x11 & n2690;
  assign n4631 = ~n4629 & ~n4630;
  assign n4632 = n4628 & n4631;
  assign n4648 = n4647 ^ n4632;
  assign n4692 = n4691 ^ n4648;
  assign n4696 = n4695 ^ n4692;
  assign n4621 = n4453 ^ n4449;
  assign n4622 = n4450 & ~n4621;
  assign n4623 = n4622 ^ n4446;
  assign n4618 = n4479 ^ n4350;
  assign n4619 = ~n4480 & ~n4618;
  assign n4620 = n4619 ^ n4472;
  assign n4624 = n4623 ^ n4620;
  assign n4614 = n4518 ^ n4511;
  assign n4615 = ~n4526 & n4614;
  assign n4616 = n4615 ^ n4511;
  assign n4610 = n4560 ^ n4553;
  assign n4611 = ~n4568 & n4610;
  assign n4612 = n4611 ^ n4553;
  assign n4603 = ~x30 & n437;
  assign n4604 = ~x29 & n439;
  assign n4605 = ~n4603 & ~n4604;
  assign n4606 = x30 & n430;
  assign n4607 = x29 & n434;
  assign n4608 = ~n4606 & ~n4607;
  assign n4609 = n4605 & n4608;
  assign n4613 = n4612 ^ n4609;
  assign n4617 = n4616 ^ n4613;
  assign n4625 = n4624 ^ n4617;
  assign n4697 = n4696 ^ n4625;
  assign n4740 = n4739 ^ n4697;
  assign n4745 = n4744 ^ n4740;
  assign n4750 = n4749 ^ n4745;
  assign n4754 = n4753 ^ n4750;
  assign n4901 = n4753 ^ n4745;
  assign n4902 = n4750 & ~n4901;
  assign n4903 = n4902 ^ n4753;
  assign n4897 = n4744 ^ n4739;
  assign n4898 = ~n4740 & ~n4897;
  assign n4899 = n4898 ^ n4697;
  assign n4893 = n4738 ^ n4734;
  assign n4894 = ~n4735 & n4893;
  assign n4895 = n4894 ^ n4731;
  assign n4887 = n4692 ^ n4625;
  assign n4888 = n4695 ^ n4625;
  assign n4889 = n4887 & ~n4888;
  assign n4890 = n4889 ^ n4692;
  assign n4882 = n4730 ^ n4723;
  assign n4883 = n4730 ^ n4726;
  assign n4884 = ~n4882 & ~n4883;
  assign n4885 = n4884 ^ n4723;
  assign n4877 = n4671 ^ n4648;
  assign n4878 = n4690 ^ n4648;
  assign n4879 = n4877 & ~n4878;
  assign n4880 = n4879 ^ n4671;
  assign n4873 = n4718 ^ n4714;
  assign n4874 = n4722 & n4873;
  assign n4875 = n4874 ^ n4714;
  assign n4868 = n4662 ^ n4655;
  assign n4869 = n4669 ^ n4655;
  assign n4870 = n4868 & ~n4869;
  assign n4871 = n4870 ^ n4662;
  assign n4863 = n4681 ^ n4678;
  assign n4864 = n4688 ^ n4678;
  assign n4865 = n4863 & ~n4864;
  assign n4866 = n4865 ^ n4681;
  assign n4860 = n4712 ^ n4704;
  assign n4861 = ~n4713 & ~n4860;
  assign n4862 = n4861 ^ n4705;
  assign n4867 = n4866 ^ n4862;
  assign n4872 = n4871 ^ n4867;
  assign n4876 = n4875 ^ n4872;
  assign n4881 = n4880 ^ n4876;
  assign n4886 = n4885 ^ n4881;
  assign n4891 = n4890 ^ n4886;
  assign n4854 = n4620 ^ n4617;
  assign n4855 = n4623 ^ n4617;
  assign n4856 = n4854 & n4855;
  assign n4857 = n4856 ^ n4620;
  assign n4843 = ~x13 & n2681;
  assign n4844 = ~x12 & n2685;
  assign n4845 = ~n4843 & ~n4844;
  assign n4846 = x13 & n2688;
  assign n4847 = x12 & n2690;
  assign n4848 = ~n4846 & ~n4847;
  assign n4849 = n4845 & n4848;
  assign n4836 = ~x15 & n2406;
  assign n4837 = ~x14 & n2408;
  assign n4838 = ~n4836 & ~n4837;
  assign n4839 = x15 & n2399;
  assign n4840 = x14 & n2403;
  assign n4841 = ~n4839 & ~n4840;
  assign n4842 = n4838 & n4841;
  assign n4850 = n4849 ^ n4842;
  assign n4829 = ~x29 & n591;
  assign n4830 = ~x28 & n595;
  assign n4831 = ~n4829 & ~n4830;
  assign n4832 = x29 & n598;
  assign n4833 = x28 & n600;
  assign n4834 = ~n4832 & ~n4833;
  assign n4835 = n4831 & n4834;
  assign n4851 = n4850 ^ n4835;
  assign n4820 = ~x31 & n437;
  assign n4821 = ~x30 & n439;
  assign n4822 = ~n4820 & ~n4821;
  assign n4823 = x31 & n430;
  assign n4824 = x30 & n434;
  assign n4825 = ~n4823 & ~n4824;
  assign n4826 = n4822 & n4825;
  assign n4819 = ~n329 & ~n333;
  assign n4827 = n4826 ^ n4819;
  assign n4812 = x27 & n780;
  assign n4813 = x26 & n784;
  assign n4814 = ~n4812 & ~n4813;
  assign n4815 = ~x27 & n787;
  assign n4816 = ~x26 & n789;
  assign n4817 = ~n4815 & ~n4816;
  assign n4818 = n4814 & n4817;
  assign n4828 = n4827 ^ n4818;
  assign n4852 = n4851 ^ n4828;
  assign n4803 = ~x17 & n1962;
  assign n4804 = ~x16 & n1966;
  assign n4805 = ~n4803 & ~n4804;
  assign n4806 = x17 & n1969;
  assign n4807 = x16 & n1971;
  assign n4808 = ~n4806 & ~n4807;
  assign n4809 = n4805 & n4808;
  assign n4796 = x19 & n1694;
  assign n4797 = x18 & n1696;
  assign n4798 = ~n4796 & ~n4797;
  assign n4799 = ~x19 & n1687;
  assign n4800 = ~x18 & n1691;
  assign n4801 = ~n4799 & ~n4800;
  assign n4802 = n4798 & n4801;
  assign n4810 = n4809 ^ n4802;
  assign n4789 = x25 & n1007;
  assign n4790 = x24 & n1009;
  assign n4791 = ~n4789 & ~n4790;
  assign n4792 = ~x25 & n1000;
  assign n4793 = ~x24 & n1004;
  assign n4794 = ~n4792 & ~n4793;
  assign n4795 = n4791 & n4794;
  assign n4811 = n4810 ^ n4795;
  assign n4853 = n4852 ^ n4811;
  assign n4858 = n4857 ^ n4853;
  assign n4785 = n4616 ^ n4612;
  assign n4786 = ~n4613 & ~n4785;
  assign n4787 = n4786 ^ n4609;
  assign n4780 = n4639 ^ n4632;
  assign n4781 = ~n4647 & n4780;
  assign n4782 = n4781 ^ n4632;
  assign n4772 = ~x21 & n1396;
  assign n4773 = ~x20 & n1400;
  assign n4774 = ~n4772 & ~n4773;
  assign n4775 = x21 & n1403;
  assign n4776 = x20 & n1405;
  assign n4777 = ~n4775 & ~n4776;
  assign n4778 = n4774 & n4777;
  assign n4779 = n4778 ^ n4609;
  assign n4783 = n4782 ^ n4779;
  assign n4763 = ~x11 & n3098;
  assign n4764 = ~x10 & n3102;
  assign n4765 = ~n4763 & ~n4764;
  assign n4766 = x11 & n3105;
  assign n4767 = x10 & n3107;
  assign n4768 = ~n4766 & ~n4767;
  assign n4769 = n4765 & n4768;
  assign n4756 = ~x23 & n1241;
  assign n4757 = ~x22 & n1243;
  assign n4758 = ~n4756 & ~n4757;
  assign n4759 = x23 & n1234;
  assign n4760 = x22 & n1238;
  assign n4761 = ~n4759 & ~n4760;
  assign n4762 = n4758 & n4761;
  assign n4770 = n4769 ^ n4762;
  assign n4755 = x9 & x63;
  assign n4771 = n4770 ^ n4755;
  assign n4784 = n4783 ^ n4771;
  assign n4788 = n4787 ^ n4784;
  assign n4859 = n4858 ^ n4788;
  assign n4892 = n4891 ^ n4859;
  assign n4896 = n4895 ^ n4892;
  assign n4900 = n4899 ^ n4896;
  assign n4904 = n4903 ^ n4900;
  assign n5040 = n4903 ^ n4896;
  assign n5041 = ~n4900 & ~n5040;
  assign n5042 = n5041 ^ n4903;
  assign n5036 = n4895 ^ n4891;
  assign n5037 = n4892 & ~n5036;
  assign n5038 = n5037 ^ n4859;
  assign n5032 = n4890 ^ n4885;
  assign n5033 = n4886 & ~n5032;
  assign n5034 = n5033 ^ n4881;
  assign n5026 = n4853 ^ n4788;
  assign n5027 = n4857 ^ n4788;
  assign n5028 = ~n5026 & n5027;
  assign n5029 = n5028 ^ n4853;
  assign n5022 = n4880 ^ n4872;
  assign n5023 = ~n4876 & ~n5022;
  assign n5024 = n5023 ^ n4880;
  assign n5018 = n4851 ^ n4811;
  assign n5019 = ~n4852 & ~n5018;
  assign n5020 = n5019 ^ n4828;
  assign n5014 = n4782 ^ n4778;
  assign n5015 = n4779 & ~n5014;
  assign n5016 = n5015 ^ n4609;
  assign n5010 = n4826 ^ n4818;
  assign n5011 = ~n4827 & ~n5010;
  assign n5012 = n5011 ^ n4819;
  assign n5006 = n4762 ^ n4755;
  assign n5007 = ~n4770 & ~n5006;
  assign n5008 = n5007 ^ n4755;
  assign n5003 = n4842 ^ n4835;
  assign n5004 = ~n4850 & n5003;
  assign n5005 = n5004 ^ n4835;
  assign n5009 = n5008 ^ n5005;
  assign n5013 = n5012 ^ n5009;
  assign n5017 = n5016 ^ n5013;
  assign n5021 = n5020 ^ n5017;
  assign n5025 = n5024 ^ n5021;
  assign n5030 = n5029 ^ n5025;
  assign n4998 = n4787 ^ n4783;
  assign n4999 = ~n4784 & n4998;
  assign n5000 = n4999 ^ n4771;
  assign n4993 = n4809 ^ n4795;
  assign n4994 = n4810 & ~n4993;
  assign n4995 = n4994 ^ n4802;
  assign n4984 = ~x28 & n787;
  assign n4985 = ~x27 & n789;
  assign n4986 = ~n4984 & ~n4985;
  assign n4987 = x28 & n780;
  assign n4988 = x27 & n784;
  assign n4989 = ~n4987 & ~n4988;
  assign n4990 = n4986 & n4989;
  assign n4981 = x43 ^ x31;
  assign n4982 = n433 & n4981;
  assign n4983 = ~n437 & ~n4982;
  assign n4991 = n4990 ^ n4983;
  assign n4980 = x10 & x63;
  assign n4992 = n4991 ^ n4980;
  assign n4996 = n4995 ^ n4992;
  assign n4971 = ~x26 & n1000;
  assign n4972 = ~x25 & n1004;
  assign n4973 = ~n4971 & ~n4972;
  assign n4974 = x26 & n1007;
  assign n4975 = x25 & n1009;
  assign n4976 = ~n4974 & ~n4975;
  assign n4977 = n4973 & n4976;
  assign n4964 = ~x18 & n1962;
  assign n4965 = ~x17 & n1966;
  assign n4966 = ~n4964 & ~n4965;
  assign n4967 = x18 & n1969;
  assign n4968 = x17 & n1971;
  assign n4969 = ~n4967 & ~n4968;
  assign n4970 = n4966 & n4969;
  assign n4978 = n4977 ^ n4970;
  assign n4957 = ~x16 & n2406;
  assign n4958 = ~x15 & n2408;
  assign n4959 = ~n4957 & ~n4958;
  assign n4960 = x16 & n2399;
  assign n4961 = x15 & n2403;
  assign n4962 = ~n4960 & ~n4961;
  assign n4963 = n4959 & n4962;
  assign n4979 = n4978 ^ n4963;
  assign n4997 = n4996 ^ n4979;
  assign n5001 = n5000 ^ n4997;
  assign n4952 = n4871 ^ n4862;
  assign n4953 = n4871 ^ n4866;
  assign n4954 = ~n4952 & ~n4953;
  assign n4955 = n4954 ^ n4862;
  assign n4942 = x24 & n1234;
  assign n4943 = x23 & n1238;
  assign n4944 = ~n4942 & ~n4943;
  assign n4945 = ~x24 & n1241;
  assign n4946 = ~x23 & n1243;
  assign n4947 = ~n4945 & ~n4946;
  assign n4948 = n4944 & n4947;
  assign n4935 = x14 & n2688;
  assign n4936 = x13 & n2690;
  assign n4937 = ~n4935 & ~n4936;
  assign n4938 = ~x14 & n2681;
  assign n4939 = ~x13 & n2685;
  assign n4940 = ~n4938 & ~n4939;
  assign n4941 = n4937 & n4940;
  assign n4949 = n4948 ^ n4941;
  assign n4928 = ~x12 & n3098;
  assign n4929 = ~x11 & n3102;
  assign n4930 = ~n4928 & ~n4929;
  assign n4931 = x12 & n3105;
  assign n4932 = x11 & n3107;
  assign n4933 = ~n4931 & ~n4932;
  assign n4934 = n4930 & n4933;
  assign n4950 = n4949 ^ n4934;
  assign n4919 = x22 & n1403;
  assign n4920 = x21 & n1405;
  assign n4921 = ~n4919 & ~n4920;
  assign n4922 = ~x22 & n1396;
  assign n4923 = ~x21 & n1400;
  assign n4924 = ~n4922 & ~n4923;
  assign n4925 = n4921 & n4924;
  assign n4912 = ~x20 & n1687;
  assign n4913 = ~x19 & n1691;
  assign n4914 = ~n4912 & ~n4913;
  assign n4915 = x20 & n1694;
  assign n4916 = x19 & n1696;
  assign n4917 = ~n4915 & ~n4916;
  assign n4918 = n4914 & n4917;
  assign n4926 = n4925 ^ n4918;
  assign n4905 = ~x30 & n591;
  assign n4906 = ~x29 & n595;
  assign n4907 = ~n4905 & ~n4906;
  assign n4908 = x30 & n598;
  assign n4909 = x29 & n600;
  assign n4910 = ~n4908 & ~n4909;
  assign n4911 = n4907 & n4910;
  assign n4927 = n4926 ^ n4911;
  assign n4951 = n4950 ^ n4927;
  assign n4956 = n4955 ^ n4951;
  assign n5002 = n5001 ^ n4956;
  assign n5031 = n5030 ^ n5002;
  assign n5035 = n5034 ^ n5031;
  assign n5039 = n5038 ^ n5035;
  assign n5043 = n5042 ^ n5039;
  assign n5178 = n5042 ^ n5035;
  assign n5179 = ~n5039 & ~n5178;
  assign n5180 = n5179 ^ n5042;
  assign n5174 = n5034 ^ n5030;
  assign n5175 = n5031 & ~n5174;
  assign n5176 = n5175 ^ n5002;
  assign n5170 = n5029 ^ n5024;
  assign n5171 = ~n5025 & n5170;
  assign n5172 = n5171 ^ n5021;
  assign n5164 = n4997 ^ n4956;
  assign n5165 = n5000 ^ n4956;
  assign n5166 = ~n5164 & n5165;
  assign n5167 = n5166 ^ n4997;
  assign n5159 = n5020 ^ n5013;
  assign n5160 = n5020 ^ n5016;
  assign n5161 = ~n5159 & n5160;
  assign n5162 = n5161 ^ n5013;
  assign n5153 = n5012 ^ n5005;
  assign n5154 = n5012 ^ n5008;
  assign n5155 = ~n5153 & ~n5154;
  assign n5156 = n5155 ^ n5005;
  assign n5149 = n4992 ^ n4979;
  assign n5150 = n4995 ^ n4979;
  assign n5151 = ~n5149 & ~n5150;
  assign n5152 = n5151 ^ n4992;
  assign n5157 = n5156 ^ n5152;
  assign n5145 = n4977 ^ n4963;
  assign n5146 = n4978 & ~n5145;
  assign n5147 = n5146 ^ n4970;
  assign n5141 = n4983 ^ n4980;
  assign n5142 = ~n4991 & ~n5141;
  assign n5143 = n5142 ^ n4980;
  assign n5144 = n5143 ^ n4911;
  assign n5148 = n5147 ^ n5144;
  assign n5158 = n5157 ^ n5148;
  assign n5163 = n5162 ^ n5158;
  assign n5168 = n5167 ^ n5163;
  assign n5137 = n4955 ^ n4950;
  assign n5138 = ~n4951 & n5137;
  assign n5139 = n5138 ^ n4927;
  assign n5131 = n4918 ^ n4911;
  assign n5132 = n4925 ^ n4911;
  assign n5133 = ~n5131 & n5132;
  assign n5134 = n5133 ^ n4918;
  assign n5121 = ~x17 & n2406;
  assign n5122 = ~x16 & n2408;
  assign n5123 = ~n5121 & ~n5122;
  assign n5124 = x17 & n2399;
  assign n5125 = x16 & n2403;
  assign n5126 = ~n5124 & ~n5125;
  assign n5127 = n5123 & n5126;
  assign n5114 = x19 & n1969;
  assign n5115 = x18 & n1971;
  assign n5116 = ~n5114 & ~n5115;
  assign n5117 = ~x19 & n1962;
  assign n5118 = ~x18 & n1966;
  assign n5119 = ~n5117 & ~n5118;
  assign n5120 = n5116 & n5119;
  assign n5128 = n5127 ^ n5120;
  assign n5107 = ~x25 & n1241;
  assign n5108 = ~x24 & n1243;
  assign n5109 = ~n5107 & ~n5108;
  assign n5110 = x25 & n1234;
  assign n5111 = x24 & n1238;
  assign n5112 = ~n5110 & ~n5111;
  assign n5113 = n5109 & n5112;
  assign n5129 = n5128 ^ n5113;
  assign n5098 = ~x31 & n591;
  assign n5099 = ~x30 & n595;
  assign n5100 = ~n5098 & ~n5099;
  assign n5101 = x31 & n598;
  assign n5102 = x30 & n600;
  assign n5103 = ~n5101 & ~n5102;
  assign n5104 = n5100 & n5103;
  assign n5097 = ~n437 & ~n439;
  assign n5105 = n5104 ^ n5097;
  assign n5090 = ~x27 & n1000;
  assign n5091 = ~x26 & n1004;
  assign n5092 = ~n5090 & ~n5091;
  assign n5093 = x27 & n1007;
  assign n5094 = x26 & n1009;
  assign n5095 = ~n5093 & ~n5094;
  assign n5096 = n5092 & n5095;
  assign n5106 = n5105 ^ n5096;
  assign n5130 = n5129 ^ n5106;
  assign n5135 = n5134 ^ n5130;
  assign n5084 = n4941 ^ n4934;
  assign n5085 = n4948 ^ n4934;
  assign n5086 = n5084 & ~n5085;
  assign n5087 = n5086 ^ n4941;
  assign n5075 = ~x13 & n3098;
  assign n5076 = ~x12 & n3102;
  assign n5077 = ~n5075 & ~n5076;
  assign n5078 = x13 & n3105;
  assign n5079 = x12 & n3107;
  assign n5080 = ~n5078 & ~n5079;
  assign n5081 = n5077 & n5080;
  assign n5068 = ~x15 & n2681;
  assign n5069 = ~x14 & n2685;
  assign n5070 = ~n5068 & ~n5069;
  assign n5071 = x15 & n2688;
  assign n5072 = x14 & n2690;
  assign n5073 = ~n5071 & ~n5072;
  assign n5074 = n5070 & n5073;
  assign n5082 = n5081 ^ n5074;
  assign n5061 = ~x29 & n787;
  assign n5062 = ~x28 & n789;
  assign n5063 = ~n5061 & ~n5062;
  assign n5064 = x29 & n780;
  assign n5065 = x28 & n784;
  assign n5066 = ~n5064 & ~n5065;
  assign n5067 = n5063 & n5066;
  assign n5083 = n5082 ^ n5067;
  assign n5088 = n5087 ^ n5083;
  assign n5052 = x23 & n1403;
  assign n5053 = x22 & n1405;
  assign n5054 = ~n5052 & ~n5053;
  assign n5055 = ~x23 & n1396;
  assign n5056 = ~x22 & n1400;
  assign n5057 = ~n5055 & ~n5056;
  assign n5058 = n5054 & n5057;
  assign n5051 = x11 & x63;
  assign n5059 = n5058 ^ n5051;
  assign n5044 = ~x21 & n1687;
  assign n5045 = ~x20 & n1691;
  assign n5046 = ~n5044 & ~n5045;
  assign n5047 = x21 & n1694;
  assign n5048 = x20 & n1696;
  assign n5049 = ~n5047 & ~n5048;
  assign n5050 = n5046 & n5049;
  assign n5060 = n5059 ^ n5050;
  assign n5089 = n5088 ^ n5060;
  assign n5136 = n5135 ^ n5089;
  assign n5140 = n5139 ^ n5136;
  assign n5169 = n5168 ^ n5140;
  assign n5173 = n5172 ^ n5169;
  assign n5177 = n5176 ^ n5173;
  assign n5181 = n5180 ^ n5177;
  assign n5304 = n5180 ^ n5173;
  assign n5305 = n5177 & n5304;
  assign n5306 = n5305 ^ n5180;
  assign n5300 = n5172 ^ n5168;
  assign n5301 = n5169 & ~n5300;
  assign n5302 = n5301 ^ n5140;
  assign n5296 = n5167 ^ n5162;
  assign n5297 = n5163 & n5296;
  assign n5298 = n5297 ^ n5158;
  assign n5291 = n5139 ^ n5135;
  assign n5292 = n5136 & ~n5291;
  assign n5293 = n5292 ^ n5089;
  assign n5287 = n5152 ^ n5148;
  assign n5288 = n5157 & n5287;
  assign n5289 = n5288 ^ n5148;
  assign n5282 = n5147 ^ n5143;
  assign n5283 = ~n5144 & n5282;
  assign n5284 = n5283 ^ n4911;
  assign n5277 = n5074 ^ n5067;
  assign n5278 = n5081 ^ n5067;
  assign n5279 = n5277 & ~n5278;
  assign n5280 = n5279 ^ n5074;
  assign n5269 = ~x20 & n1962;
  assign n5270 = ~x19 & n1966;
  assign n5271 = ~n5269 & ~n5270;
  assign n5272 = x20 & n1969;
  assign n5273 = x19 & n1971;
  assign n5274 = ~n5272 & ~n5273;
  assign n5275 = n5271 & n5274;
  assign n5262 = ~x30 & n787;
  assign n5263 = ~x29 & n789;
  assign n5264 = ~n5262 & ~n5263;
  assign n5265 = x30 & n780;
  assign n5266 = x29 & n784;
  assign n5267 = ~n5265 & ~n5266;
  assign n5268 = n5264 & n5267;
  assign n5276 = n5275 ^ n5268;
  assign n5281 = n5280 ^ n5276;
  assign n5285 = n5284 ^ n5281;
  assign n5258 = n5127 ^ n5113;
  assign n5259 = n5128 & ~n5258;
  assign n5260 = n5259 ^ n5120;
  assign n5254 = n5104 ^ n5096;
  assign n5255 = ~n5105 & ~n5254;
  assign n5256 = n5255 ^ n5097;
  assign n5251 = n5058 ^ n5050;
  assign n5252 = ~n5059 & ~n5251;
  assign n5253 = n5252 ^ n5051;
  assign n5257 = n5256 ^ n5253;
  assign n5261 = n5260 ^ n5257;
  assign n5286 = n5285 ^ n5261;
  assign n5290 = n5289 ^ n5286;
  assign n5294 = n5293 ^ n5290;
  assign n5246 = n5134 ^ n5129;
  assign n5247 = ~n5130 & ~n5246;
  assign n5248 = n5247 ^ n5106;
  assign n5243 = n5083 ^ n5060;
  assign n5244 = ~n5088 & ~n5243;
  assign n5245 = n5244 ^ n5060;
  assign n5249 = n5248 ^ n5245;
  assign n5232 = x14 & n3105;
  assign n5233 = x13 & n3107;
  assign n5234 = ~n5232 & ~n5233;
  assign n5235 = ~x14 & n3098;
  assign n5236 = ~x13 & n3102;
  assign n5237 = ~n5235 & ~n5236;
  assign n5238 = n5234 & n5237;
  assign n5225 = x24 & n1403;
  assign n5226 = x23 & n1405;
  assign n5227 = ~n5225 & ~n5226;
  assign n5228 = ~x24 & n1396;
  assign n5229 = ~x23 & n1400;
  assign n5230 = ~n5228 & ~n5229;
  assign n5231 = n5227 & n5230;
  assign n5239 = n5238 ^ n5231;
  assign n5224 = x12 & x63;
  assign n5240 = n5239 ^ n5224;
  assign n5215 = ~x28 & n1000;
  assign n5216 = ~x27 & n1004;
  assign n5217 = ~n5215 & ~n5216;
  assign n5218 = x28 & n1007;
  assign n5219 = x27 & n1009;
  assign n5220 = ~n5218 & ~n5219;
  assign n5221 = n5217 & n5220;
  assign n5212 = x45 ^ x31;
  assign n5213 = n594 & n5212;
  assign n5214 = ~n591 & ~n5213;
  assign n5222 = n5221 ^ n5214;
  assign n5205 = ~x22 & n1687;
  assign n5206 = ~x21 & n1691;
  assign n5207 = ~n5205 & ~n5206;
  assign n5208 = x22 & n1694;
  assign n5209 = x21 & n1696;
  assign n5210 = ~n5208 & ~n5209;
  assign n5211 = n5207 & n5210;
  assign n5223 = n5222 ^ n5211;
  assign n5241 = n5240 ^ n5223;
  assign n5196 = x26 & n1234;
  assign n5197 = x25 & n1238;
  assign n5198 = ~n5196 & ~n5197;
  assign n5199 = ~x26 & n1241;
  assign n5200 = ~x25 & n1243;
  assign n5201 = ~n5199 & ~n5200;
  assign n5202 = n5198 & n5201;
  assign n5189 = x18 & n2399;
  assign n5190 = x17 & n2403;
  assign n5191 = ~n5189 & ~n5190;
  assign n5192 = ~x18 & n2406;
  assign n5193 = ~x17 & n2408;
  assign n5194 = ~n5192 & ~n5193;
  assign n5195 = n5191 & n5194;
  assign n5203 = n5202 ^ n5195;
  assign n5182 = ~x16 & n2681;
  assign n5183 = ~x15 & n2685;
  assign n5184 = ~n5182 & ~n5183;
  assign n5185 = x16 & n2688;
  assign n5186 = x15 & n2690;
  assign n5187 = ~n5185 & ~n5186;
  assign n5188 = n5184 & n5187;
  assign n5204 = n5203 ^ n5188;
  assign n5242 = n5241 ^ n5204;
  assign n5250 = n5249 ^ n5242;
  assign n5295 = n5294 ^ n5250;
  assign n5299 = n5298 ^ n5295;
  assign n5303 = n5302 ^ n5299;
  assign n5307 = n5306 ^ n5303;
  assign n5429 = n5306 ^ n5299;
  assign n5430 = n5303 & ~n5429;
  assign n5431 = n5430 ^ n5306;
  assign n5425 = n5298 ^ n5294;
  assign n5426 = n5295 & n5425;
  assign n5427 = n5426 ^ n5250;
  assign n5421 = n5293 ^ n5289;
  assign n5422 = n5290 & ~n5421;
  assign n5423 = n5422 ^ n5286;
  assign n5417 = n5245 ^ n5242;
  assign n5418 = ~n5249 & n5417;
  assign n5419 = n5418 ^ n5242;
  assign n5411 = n5281 ^ n5261;
  assign n5412 = n5284 ^ n5261;
  assign n5413 = ~n5411 & ~n5412;
  assign n5414 = n5413 ^ n5281;
  assign n5407 = n5280 ^ n5275;
  assign n5408 = ~n5276 & ~n5407;
  assign n5409 = n5408 ^ n5268;
  assign n5402 = n5260 ^ n5253;
  assign n5403 = n5260 ^ n5256;
  assign n5404 = ~n5402 & n5403;
  assign n5405 = n5404 ^ n5253;
  assign n5393 = x23 & n1694;
  assign n5394 = x22 & n1696;
  assign n5395 = ~n5393 & ~n5394;
  assign n5396 = ~x23 & n1687;
  assign n5397 = ~x22 & n1691;
  assign n5398 = ~n5396 & ~n5397;
  assign n5399 = n5395 & n5398;
  assign n5386 = ~x21 & n1962;
  assign n5387 = ~x20 & n1966;
  assign n5388 = ~n5386 & ~n5387;
  assign n5389 = x21 & n1969;
  assign n5390 = x20 & n1971;
  assign n5391 = ~n5389 & ~n5390;
  assign n5392 = n5388 & n5391;
  assign n5400 = n5399 ^ n5392;
  assign n5401 = n5400 ^ n5268;
  assign n5406 = n5405 ^ n5401;
  assign n5410 = n5409 ^ n5406;
  assign n5415 = n5414 ^ n5410;
  assign n5380 = n5223 ^ n5204;
  assign n5381 = n5240 ^ n5204;
  assign n5382 = n5380 & n5381;
  assign n5383 = n5382 ^ n5223;
  assign n5376 = n5231 ^ n5224;
  assign n5377 = ~n5239 & ~n5376;
  assign n5378 = n5377 ^ n5224;
  assign n5371 = n5195 ^ n5188;
  assign n5372 = n5202 ^ n5188;
  assign n5373 = n5371 & ~n5372;
  assign n5374 = n5373 ^ n5195;
  assign n5367 = n5214 ^ n5211;
  assign n5368 = n5221 ^ n5211;
  assign n5369 = n5367 & ~n5368;
  assign n5370 = n5369 ^ n5214;
  assign n5375 = n5374 ^ n5370;
  assign n5379 = n5378 ^ n5375;
  assign n5384 = n5383 ^ n5379;
  assign n5356 = x15 & n3105;
  assign n5357 = x14 & n3107;
  assign n5358 = ~n5356 & ~n5357;
  assign n5359 = ~x15 & n3098;
  assign n5360 = ~x14 & n3102;
  assign n5361 = ~n5359 & ~n5360;
  assign n5362 = n5358 & n5361;
  assign n5355 = x13 & x63;
  assign n5363 = n5362 ^ n5355;
  assign n5348 = ~x29 & n1000;
  assign n5349 = ~x28 & n1004;
  assign n5350 = ~n5348 & ~n5349;
  assign n5351 = x29 & n1007;
  assign n5352 = x28 & n1009;
  assign n5353 = ~n5351 & ~n5352;
  assign n5354 = n5350 & n5353;
  assign n5364 = n5363 ^ n5354;
  assign n5339 = ~x17 & n2681;
  assign n5340 = ~x16 & n2685;
  assign n5341 = ~n5339 & ~n5340;
  assign n5342 = x17 & n2688;
  assign n5343 = x16 & n2690;
  assign n5344 = ~n5342 & ~n5343;
  assign n5345 = n5341 & n5344;
  assign n5332 = x19 & n2399;
  assign n5333 = x18 & n2403;
  assign n5334 = ~n5332 & ~n5333;
  assign n5335 = ~x19 & n2406;
  assign n5336 = ~x18 & n2408;
  assign n5337 = ~n5335 & ~n5336;
  assign n5338 = n5334 & n5337;
  assign n5346 = n5345 ^ n5338;
  assign n5325 = ~x25 & n1396;
  assign n5326 = ~x24 & n1400;
  assign n5327 = ~n5325 & ~n5326;
  assign n5328 = x25 & n1403;
  assign n5329 = x24 & n1405;
  assign n5330 = ~n5328 & ~n5329;
  assign n5331 = n5327 & n5330;
  assign n5347 = n5346 ^ n5331;
  assign n5365 = n5364 ^ n5347;
  assign n5316 = ~x31 & n787;
  assign n5317 = ~x30 & n789;
  assign n5318 = ~n5316 & ~n5317;
  assign n5319 = x31 & n780;
  assign n5320 = x30 & n784;
  assign n5321 = ~n5319 & ~n5320;
  assign n5322 = n5318 & n5321;
  assign n5315 = ~n591 & ~n595;
  assign n5323 = n5322 ^ n5315;
  assign n5308 = x27 & n1234;
  assign n5309 = x26 & n1238;
  assign n5310 = ~n5308 & ~n5309;
  assign n5311 = ~x27 & n1241;
  assign n5312 = ~x26 & n1243;
  assign n5313 = ~n5311 & ~n5312;
  assign n5314 = n5310 & n5313;
  assign n5324 = n5323 ^ n5314;
  assign n5366 = n5365 ^ n5324;
  assign n5385 = n5384 ^ n5366;
  assign n5416 = n5415 ^ n5385;
  assign n5420 = n5419 ^ n5416;
  assign n5424 = n5423 ^ n5420;
  assign n5428 = n5427 ^ n5424;
  assign n5432 = n5431 ^ n5428;
  assign n5545 = n5431 ^ n5424;
  assign n5546 = n5428 & ~n5545;
  assign n5547 = n5546 ^ n5431;
  assign n5541 = n5423 ^ n5419;
  assign n5542 = ~n5420 & ~n5541;
  assign n5543 = n5542 ^ n5416;
  assign n5537 = n5410 ^ n5385;
  assign n5538 = n5415 & ~n5537;
  assign n5539 = n5538 ^ n5385;
  assign n5532 = n5383 ^ n5366;
  assign n5533 = n5384 & n5532;
  assign n5534 = n5533 ^ n5366;
  assign n5527 = n5409 ^ n5401;
  assign n5528 = n5409 ^ n5405;
  assign n5529 = ~n5527 & ~n5528;
  assign n5530 = n5529 ^ n5401;
  assign n5523 = n5378 ^ n5374;
  assign n5524 = n5375 & n5523;
  assign n5525 = n5524 ^ n5370;
  assign n5518 = n5392 ^ n5268;
  assign n5519 = n5399 ^ n5268;
  assign n5520 = n5518 & ~n5519;
  assign n5521 = n5520 ^ n5392;
  assign n5509 = ~x28 & n1241;
  assign n5510 = ~x27 & n1243;
  assign n5511 = ~n5509 & ~n5510;
  assign n5512 = x28 & n1234;
  assign n5513 = x27 & n1238;
  assign n5514 = ~n5512 & ~n5513;
  assign n5515 = n5511 & n5514;
  assign n5502 = ~x22 & n1962;
  assign n5503 = ~x21 & n1966;
  assign n5504 = ~n5502 & ~n5503;
  assign n5505 = x22 & n1969;
  assign n5506 = x21 & n1971;
  assign n5507 = ~n5505 & ~n5506;
  assign n5508 = n5504 & n5507;
  assign n5516 = n5515 ^ n5508;
  assign n5495 = x20 & n2399;
  assign n5496 = x19 & n2403;
  assign n5497 = ~n5495 & ~n5496;
  assign n5498 = ~x20 & n2406;
  assign n5499 = ~x19 & n2408;
  assign n5500 = ~n5498 & ~n5499;
  assign n5501 = n5497 & n5500;
  assign n5517 = n5516 ^ n5501;
  assign n5522 = n5521 ^ n5517;
  assign n5526 = n5525 ^ n5522;
  assign n5531 = n5530 ^ n5526;
  assign n5535 = n5534 ^ n5531;
  assign n5490 = n5347 ^ n5324;
  assign n5491 = n5365 & ~n5490;
  assign n5492 = n5491 ^ n5324;
  assign n5486 = n5338 ^ n5331;
  assign n5487 = ~n5346 & n5486;
  assign n5488 = n5487 ^ n5331;
  assign n5482 = n5322 ^ n5314;
  assign n5483 = ~n5323 & ~n5482;
  assign n5484 = n5483 ^ n5315;
  assign n5479 = x47 ^ x31;
  assign n5480 = n783 & n5479;
  assign n5481 = ~n787 & ~n5480;
  assign n5485 = n5484 ^ n5481;
  assign n5489 = n5488 ^ n5485;
  assign n5493 = n5492 ^ n5489;
  assign n5473 = n5355 ^ n5354;
  assign n5474 = n5362 ^ n5354;
  assign n5475 = ~n5473 & ~n5474;
  assign n5476 = n5475 ^ n5355;
  assign n5464 = ~x18 & n2681;
  assign n5465 = ~x17 & n2685;
  assign n5466 = ~n5464 & ~n5465;
  assign n5467 = x18 & n2688;
  assign n5468 = x17 & n2690;
  assign n5469 = ~n5467 & ~n5468;
  assign n5470 = n5466 & n5469;
  assign n5457 = ~x26 & n1396;
  assign n5458 = ~x25 & n1400;
  assign n5459 = ~n5457 & ~n5458;
  assign n5460 = x26 & n1403;
  assign n5461 = x25 & n1405;
  assign n5462 = ~n5460 & ~n5461;
  assign n5463 = n5459 & n5462;
  assign n5471 = n5470 ^ n5463;
  assign n5450 = ~x16 & n3098;
  assign n5451 = ~x15 & n3102;
  assign n5452 = ~n5450 & ~n5451;
  assign n5453 = x16 & n3105;
  assign n5454 = x15 & n3107;
  assign n5455 = ~n5453 & ~n5454;
  assign n5456 = n5452 & n5455;
  assign n5472 = n5471 ^ n5456;
  assign n5477 = n5476 ^ n5472;
  assign n5441 = ~x30 & n1000;
  assign n5442 = ~x29 & n1004;
  assign n5443 = ~n5441 & ~n5442;
  assign n5444 = x30 & n1007;
  assign n5445 = x29 & n1009;
  assign n5446 = ~n5444 & ~n5445;
  assign n5447 = n5443 & n5446;
  assign n5440 = x14 & x63;
  assign n5448 = n5447 ^ n5440;
  assign n5433 = ~x24 & n1687;
  assign n5434 = ~x23 & n1691;
  assign n5435 = ~n5433 & ~n5434;
  assign n5436 = x24 & n1694;
  assign n5437 = x23 & n1696;
  assign n5438 = ~n5436 & ~n5437;
  assign n5439 = n5435 & n5438;
  assign n5449 = n5448 ^ n5439;
  assign n5478 = n5477 ^ n5449;
  assign n5494 = n5493 ^ n5478;
  assign n5536 = n5535 ^ n5494;
  assign n5540 = n5539 ^ n5536;
  assign n5544 = n5543 ^ n5540;
  assign n5548 = n5547 ^ n5544;
  assign n5656 = n5547 ^ n5540;
  assign n5657 = ~n5544 & ~n5656;
  assign n5658 = n5657 ^ n5547;
  assign n5652 = n5539 ^ n5535;
  assign n5653 = ~n5536 & n5652;
  assign n5654 = n5653 ^ n5494;
  assign n5647 = n5534 ^ n5526;
  assign n5648 = n5534 ^ n5530;
  assign n5649 = n5647 & ~n5648;
  assign n5650 = n5649 ^ n5526;
  assign n5642 = n5489 ^ n5478;
  assign n5643 = n5493 & n5642;
  assign n5644 = n5643 ^ n5478;
  assign n5638 = n5525 ^ n5521;
  assign n5639 = n5522 & ~n5638;
  assign n5640 = n5639 ^ n5517;
  assign n5633 = n5470 ^ n5456;
  assign n5634 = n5471 & ~n5633;
  assign n5635 = n5634 ^ n5463;
  assign n5625 = x21 & n2399;
  assign n5626 = x20 & n2403;
  assign n5627 = ~n5625 & ~n5626;
  assign n5628 = ~x21 & n2406;
  assign n5629 = ~x20 & n2408;
  assign n5630 = ~n5628 & ~n5629;
  assign n5631 = n5627 & n5630;
  assign n5632 = n5631 ^ n5481;
  assign n5636 = n5635 ^ n5632;
  assign n5615 = ~x17 & n3098;
  assign n5616 = ~x16 & n3102;
  assign n5617 = ~n5615 & ~n5616;
  assign n5618 = x17 & n3105;
  assign n5619 = x16 & n3107;
  assign n5620 = ~n5618 & ~n5619;
  assign n5621 = n5617 & n5620;
  assign n5608 = ~x19 & n2681;
  assign n5609 = ~x18 & n2685;
  assign n5610 = ~n5608 & ~n5609;
  assign n5611 = x19 & n2688;
  assign n5612 = x18 & n2690;
  assign n5613 = ~n5611 & ~n5612;
  assign n5614 = n5610 & n5613;
  assign n5622 = n5621 ^ n5614;
  assign n5601 = x25 & n1694;
  assign n5602 = x24 & n1696;
  assign n5603 = ~n5601 & ~n5602;
  assign n5604 = ~x25 & n1687;
  assign n5605 = ~x24 & n1691;
  assign n5606 = ~n5604 & ~n5605;
  assign n5607 = n5603 & n5606;
  assign n5623 = n5622 ^ n5607;
  assign n5592 = ~x31 & n1000;
  assign n5593 = ~x30 & n1004;
  assign n5594 = ~n5592 & ~n5593;
  assign n5595 = x31 & n1007;
  assign n5596 = x30 & n1009;
  assign n5597 = ~n5595 & ~n5596;
  assign n5598 = n5594 & n5597;
  assign n5591 = ~n787 & ~n789;
  assign n5599 = n5598 ^ n5591;
  assign n5584 = ~x27 & n1396;
  assign n5585 = ~x26 & n1400;
  assign n5586 = ~n5584 & ~n5585;
  assign n5587 = x27 & n1403;
  assign n5588 = x26 & n1405;
  assign n5589 = ~n5587 & ~n5588;
  assign n5590 = n5586 & n5589;
  assign n5600 = n5599 ^ n5590;
  assign n5624 = n5623 ^ n5600;
  assign n5637 = n5636 ^ n5624;
  assign n5641 = n5640 ^ n5637;
  assign n5645 = n5644 ^ n5641;
  assign n5578 = n5488 ^ n5481;
  assign n5579 = n5488 ^ n5484;
  assign n5580 = ~n5578 & n5579;
  assign n5581 = n5580 ^ n5481;
  assign n5575 = n5472 ^ n5449;
  assign n5576 = n5477 & ~n5575;
  assign n5577 = n5576 ^ n5449;
  assign n5582 = n5581 ^ n5577;
  assign n5569 = n5508 ^ n5501;
  assign n5570 = n5515 ^ n5501;
  assign n5571 = n5569 & ~n5570;
  assign n5572 = n5571 ^ n5508;
  assign n5566 = n5447 ^ n5439;
  assign n5567 = ~n5448 & ~n5566;
  assign n5568 = n5567 ^ n5440;
  assign n5573 = n5572 ^ n5568;
  assign n5557 = x29 & n1234;
  assign n5558 = x28 & n1238;
  assign n5559 = ~n5557 & ~n5558;
  assign n5560 = ~x29 & n1241;
  assign n5561 = ~x28 & n1243;
  assign n5562 = ~n5560 & ~n5561;
  assign n5563 = n5559 & n5562;
  assign n5556 = x15 & x63;
  assign n5564 = n5563 ^ n5556;
  assign n5549 = ~x23 & n1962;
  assign n5550 = ~x22 & n1966;
  assign n5551 = ~n5549 & ~n5550;
  assign n5552 = x23 & n1969;
  assign n5553 = x22 & n1971;
  assign n5554 = ~n5552 & ~n5553;
  assign n5555 = n5551 & n5554;
  assign n5565 = n5564 ^ n5555;
  assign n5574 = n5573 ^ n5565;
  assign n5583 = n5582 ^ n5574;
  assign n5646 = n5645 ^ n5583;
  assign n5651 = n5650 ^ n5646;
  assign n5655 = n5654 ^ n5651;
  assign n5659 = n5658 ^ n5655;
  assign n5758 = n5658 ^ n5651;
  assign n5759 = ~n5655 & n5758;
  assign n5760 = n5759 ^ n5658;
  assign n5754 = n5650 ^ n5645;
  assign n5755 = ~n5646 & n5754;
  assign n5756 = n5755 ^ n5583;
  assign n5749 = n5644 ^ n5637;
  assign n5750 = n5644 ^ n5640;
  assign n5751 = ~n5749 & ~n5750;
  assign n5752 = n5751 ^ n5637;
  assign n5744 = n5577 ^ n5574;
  assign n5745 = ~n5582 & ~n5744;
  assign n5746 = n5745 ^ n5574;
  assign n5740 = n5636 ^ n5623;
  assign n5741 = ~n5624 & ~n5740;
  assign n5742 = n5741 ^ n5600;
  assign n5729 = x26 & n1694;
  assign n5730 = x25 & n1696;
  assign n5731 = ~n5729 & ~n5730;
  assign n5732 = ~x26 & n1687;
  assign n5733 = ~x25 & n1691;
  assign n5734 = ~n5732 & ~n5733;
  assign n5735 = n5731 & n5734;
  assign n5722 = ~x18 & n3098;
  assign n5723 = ~x17 & n3102;
  assign n5724 = ~n5722 & ~n5723;
  assign n5725 = x18 & n3105;
  assign n5726 = x17 & n3107;
  assign n5727 = ~n5725 & ~n5726;
  assign n5728 = n5724 & n5727;
  assign n5736 = n5735 ^ n5728;
  assign n5721 = x16 & x63;
  assign n5737 = n5736 ^ n5721;
  assign n5712 = x30 & n1234;
  assign n5713 = x29 & n1238;
  assign n5714 = ~n5712 & ~n5713;
  assign n5715 = ~x30 & n1241;
  assign n5716 = ~x29 & n1243;
  assign n5717 = ~n5715 & ~n5716;
  assign n5718 = n5714 & n5717;
  assign n5705 = x24 & n1969;
  assign n5706 = x23 & n1971;
  assign n5707 = ~n5705 & ~n5706;
  assign n5708 = ~x24 & n1962;
  assign n5709 = ~x23 & n1966;
  assign n5710 = ~n5708 & ~n5709;
  assign n5711 = n5707 & n5710;
  assign n5719 = n5718 ^ n5711;
  assign n5698 = x28 & n1403;
  assign n5699 = x27 & n1405;
  assign n5700 = ~n5698 & ~n5699;
  assign n5701 = ~x28 & n1396;
  assign n5702 = ~x27 & n1400;
  assign n5703 = ~n5701 & ~n5702;
  assign n5704 = n5700 & n5703;
  assign n5720 = n5719 ^ n5704;
  assign n5738 = n5737 ^ n5720;
  assign n5689 = ~x22 & n2406;
  assign n5690 = ~x21 & n2408;
  assign n5691 = ~n5689 & ~n5690;
  assign n5692 = x22 & n2399;
  assign n5693 = x21 & n2403;
  assign n5694 = ~n5692 & ~n5693;
  assign n5695 = n5691 & n5694;
  assign n5682 = ~x20 & n2681;
  assign n5683 = ~x19 & n2685;
  assign n5684 = ~n5682 & ~n5683;
  assign n5685 = x20 & n2688;
  assign n5686 = x19 & n2690;
  assign n5687 = ~n5685 & ~n5686;
  assign n5688 = n5684 & n5687;
  assign n5696 = n5695 ^ n5688;
  assign n5679 = x49 ^ x31;
  assign n5680 = n1003 & n5679;
  assign n5681 = ~n1000 & ~n5680;
  assign n5697 = n5696 ^ n5681;
  assign n5739 = n5738 ^ n5697;
  assign n5743 = n5742 ^ n5739;
  assign n5747 = n5746 ^ n5743;
  assign n5674 = n5568 ^ n5565;
  assign n5675 = n5573 & n5674;
  assign n5676 = n5675 ^ n5565;
  assign n5671 = n5635 ^ n5631;
  assign n5672 = n5632 & ~n5671;
  assign n5673 = n5672 ^ n5481;
  assign n5677 = n5676 ^ n5673;
  assign n5667 = n5563 ^ n5555;
  assign n5668 = ~n5564 & ~n5667;
  assign n5669 = n5668 ^ n5556;
  assign n5663 = n5621 ^ n5607;
  assign n5664 = n5622 & ~n5663;
  assign n5665 = n5664 ^ n5614;
  assign n5660 = n5598 ^ n5590;
  assign n5661 = ~n5599 & ~n5660;
  assign n5662 = n5661 ^ n5591;
  assign n5666 = n5665 ^ n5662;
  assign n5670 = n5669 ^ n5666;
  assign n5678 = n5677 ^ n5670;
  assign n5748 = n5747 ^ n5678;
  assign n5753 = n5752 ^ n5748;
  assign n5757 = n5756 ^ n5753;
  assign n5761 = n5760 ^ n5757;
  assign n5854 = n5760 ^ n5753;
  assign n5855 = n5757 & n5854;
  assign n5856 = n5855 ^ n5760;
  assign n5850 = n5752 ^ n5747;
  assign n5851 = n5748 & ~n5850;
  assign n5852 = n5851 ^ n5678;
  assign n5846 = n5746 ^ n5742;
  assign n5847 = ~n5743 & n5846;
  assign n5848 = n5847 ^ n5739;
  assign n5841 = n5673 ^ n5670;
  assign n5842 = n5677 & n5841;
  assign n5843 = n5842 ^ n5670;
  assign n5837 = n5720 ^ n5697;
  assign n5838 = n5738 & ~n5837;
  assign n5839 = n5838 ^ n5697;
  assign n5826 = ~x31 & n1241;
  assign n5827 = ~x30 & n1243;
  assign n5828 = ~n5826 & ~n5827;
  assign n5829 = x31 & n1234;
  assign n5830 = x30 & n1238;
  assign n5831 = ~n5829 & ~n5830;
  assign n5832 = n5828 & n5831;
  assign n5825 = ~n1000 & ~n1004;
  assign n5833 = n5832 ^ n5825;
  assign n5818 = ~x27 & n1687;
  assign n5819 = ~x26 & n1691;
  assign n5820 = ~n5818 & ~n5819;
  assign n5821 = x27 & n1694;
  assign n5822 = x26 & n1696;
  assign n5823 = ~n5821 & ~n5822;
  assign n5824 = n5820 & n5823;
  assign n5834 = n5833 ^ n5824;
  assign n5809 = ~x23 & n2406;
  assign n5810 = ~x22 & n2408;
  assign n5811 = ~n5809 & ~n5810;
  assign n5812 = x23 & n2399;
  assign n5813 = x22 & n2403;
  assign n5814 = ~n5812 & ~n5813;
  assign n5815 = n5811 & n5814;
  assign n5802 = ~x29 & n1396;
  assign n5803 = ~x28 & n1400;
  assign n5804 = ~n5802 & ~n5803;
  assign n5805 = x29 & n1403;
  assign n5806 = x28 & n1405;
  assign n5807 = ~n5805 & ~n5806;
  assign n5808 = n5804 & n5807;
  assign n5816 = n5815 ^ n5808;
  assign n5795 = x21 & n2688;
  assign n5796 = x20 & n2690;
  assign n5797 = ~n5795 & ~n5796;
  assign n5798 = ~x21 & n2681;
  assign n5799 = ~x20 & n2685;
  assign n5800 = ~n5798 & ~n5799;
  assign n5801 = n5797 & n5800;
  assign n5817 = n5816 ^ n5801;
  assign n5835 = n5834 ^ n5817;
  assign n5786 = x19 & n3105;
  assign n5787 = x18 & n3107;
  assign n5788 = ~n5786 & ~n5787;
  assign n5789 = ~x19 & n3098;
  assign n5790 = ~x18 & n3102;
  assign n5791 = ~n5789 & ~n5790;
  assign n5792 = n5788 & n5791;
  assign n5785 = x17 & x63;
  assign n5793 = n5792 ^ n5785;
  assign n5778 = ~x25 & n1962;
  assign n5779 = ~x24 & n1966;
  assign n5780 = ~n5778 & ~n5779;
  assign n5781 = x25 & n1969;
  assign n5782 = x24 & n1971;
  assign n5783 = ~n5781 & ~n5782;
  assign n5784 = n5780 & n5783;
  assign n5794 = n5793 ^ n5784;
  assign n5836 = n5835 ^ n5794;
  assign n5840 = n5839 ^ n5836;
  assign n5844 = n5843 ^ n5840;
  assign n5773 = n5669 ^ n5662;
  assign n5774 = n5666 & n5773;
  assign n5775 = n5774 ^ n5669;
  assign n5770 = n5688 ^ n5681;
  assign n5771 = ~n5696 & ~n5770;
  assign n5772 = n5771 ^ n5681;
  assign n5776 = n5775 ^ n5772;
  assign n5766 = n5718 ^ n5704;
  assign n5767 = n5719 & ~n5766;
  assign n5768 = n5767 ^ n5711;
  assign n5762 = n5728 ^ n5721;
  assign n5763 = ~n5736 & ~n5762;
  assign n5764 = n5763 ^ n5721;
  assign n5765 = n5764 ^ n5681;
  assign n5769 = n5768 ^ n5765;
  assign n5777 = n5776 ^ n5769;
  assign n5845 = n5844 ^ n5777;
  assign n5849 = n5848 ^ n5845;
  assign n5853 = n5852 ^ n5849;
  assign n5857 = n5856 ^ n5853;
  assign n5946 = n5856 ^ n5849;
  assign n5947 = n5853 & ~n5946;
  assign n5948 = n5947 ^ n5856;
  assign n5942 = n5848 ^ n5844;
  assign n5943 = n5845 & n5942;
  assign n5944 = n5943 ^ n5777;
  assign n5938 = n5843 ^ n5839;
  assign n5939 = ~n5840 & n5938;
  assign n5940 = n5939 ^ n5836;
  assign n5933 = n5772 ^ n5769;
  assign n5934 = n5775 ^ n5769;
  assign n5935 = n5933 & ~n5934;
  assign n5936 = n5935 ^ n5772;
  assign n5928 = n5768 ^ n5764;
  assign n5929 = ~n5765 & n5928;
  assign n5930 = n5929 ^ n5681;
  assign n5922 = n5825 ^ n5824;
  assign n5923 = n5832 ^ n5824;
  assign n5924 = ~n5922 & ~n5923;
  assign n5925 = n5924 ^ n5825;
  assign n5914 = x20 & n3105;
  assign n5915 = x19 & n3107;
  assign n5916 = ~n5914 & ~n5915;
  assign n5917 = ~x20 & n3098;
  assign n5918 = ~x19 & n3102;
  assign n5919 = ~n5917 & ~n5918;
  assign n5920 = n5916 & n5919;
  assign n5911 = x51 ^ x31;
  assign n5912 = n1237 & n5911;
  assign n5913 = ~n1241 & ~n5912;
  assign n5921 = n5920 ^ n5913;
  assign n5926 = n5925 ^ n5921;
  assign n5902 = ~x30 & n1396;
  assign n5903 = ~x29 & n1400;
  assign n5904 = ~n5902 & ~n5903;
  assign n5905 = x30 & n1403;
  assign n5906 = x29 & n1405;
  assign n5907 = ~n5905 & ~n5906;
  assign n5908 = n5904 & n5907;
  assign n5901 = x18 & x63;
  assign n5909 = n5908 ^ n5901;
  assign n5894 = x26 & n1969;
  assign n5895 = x25 & n1971;
  assign n5896 = ~n5894 & ~n5895;
  assign n5897 = ~x26 & n1962;
  assign n5898 = ~x25 & n1966;
  assign n5899 = ~n5897 & ~n5898;
  assign n5900 = n5896 & n5899;
  assign n5910 = n5909 ^ n5900;
  assign n5927 = n5926 ^ n5910;
  assign n5931 = n5930 ^ n5927;
  assign n5890 = n5834 ^ n5794;
  assign n5891 = ~n5835 & ~n5890;
  assign n5892 = n5891 ^ n5817;
  assign n5885 = n5815 ^ n5801;
  assign n5886 = n5816 & ~n5885;
  assign n5887 = n5886 ^ n5808;
  assign n5881 = n5785 ^ n5784;
  assign n5882 = n5792 ^ n5784;
  assign n5883 = ~n5881 & ~n5882;
  assign n5884 = n5883 ^ n5785;
  assign n5888 = n5887 ^ n5884;
  assign n5872 = x28 & n1694;
  assign n5873 = x27 & n1696;
  assign n5874 = ~n5872 & ~n5873;
  assign n5875 = ~x28 & n1687;
  assign n5876 = ~x27 & n1691;
  assign n5877 = ~n5875 & ~n5876;
  assign n5878 = n5874 & n5877;
  assign n5865 = ~x24 & n2406;
  assign n5866 = ~x23 & n2408;
  assign n5867 = ~n5865 & ~n5866;
  assign n5868 = x24 & n2399;
  assign n5869 = x23 & n2403;
  assign n5870 = ~n5868 & ~n5869;
  assign n5871 = n5867 & n5870;
  assign n5879 = n5878 ^ n5871;
  assign n5858 = ~x22 & n2681;
  assign n5859 = ~x21 & n2685;
  assign n5860 = ~n5858 & ~n5859;
  assign n5861 = x22 & n2688;
  assign n5862 = x21 & n2690;
  assign n5863 = ~n5861 & ~n5862;
  assign n5864 = n5860 & n5863;
  assign n5880 = n5879 ^ n5864;
  assign n5889 = n5888 ^ n5880;
  assign n5893 = n5892 ^ n5889;
  assign n5932 = n5931 ^ n5893;
  assign n5937 = n5936 ^ n5932;
  assign n5941 = n5940 ^ n5937;
  assign n5945 = n5944 ^ n5941;
  assign n5949 = n5948 ^ n5945;
  assign n6030 = n5948 ^ n5941;
  assign n6031 = ~n5945 & n6030;
  assign n6032 = n6031 ^ n5948;
  assign n6026 = n5940 ^ n5936;
  assign n6027 = ~n5937 & n6026;
  assign n6028 = n6027 ^ n5932;
  assign n6022 = n5931 ^ n5892;
  assign n6023 = ~n5893 & n6022;
  assign n6024 = n6023 ^ n5889;
  assign n6017 = n5930 ^ n5926;
  assign n6018 = ~n5927 & ~n6017;
  assign n6019 = n6018 ^ n5910;
  assign n6013 = n5884 ^ n5880;
  assign n6014 = n5888 & ~n6013;
  assign n6015 = n6014 ^ n5880;
  assign n6008 = n5871 ^ n5864;
  assign n6009 = ~n5879 & n6008;
  assign n6010 = n6009 ^ n5864;
  assign n6005 = n5908 ^ n5900;
  assign n6006 = ~n5909 & ~n6005;
  assign n6007 = n6006 ^ n5901;
  assign n6011 = n6010 ^ n6007;
  assign n5996 = ~x31 & n1396;
  assign n5997 = ~x30 & n1400;
  assign n5998 = ~n5996 & ~n5997;
  assign n5999 = x31 & n1403;
  assign n6000 = x30 & n1405;
  assign n6001 = ~n5999 & ~n6000;
  assign n6002 = n5998 & n6001;
  assign n5995 = ~n1241 & ~n1243;
  assign n6003 = n6002 ^ n5995;
  assign n5988 = ~x27 & n1962;
  assign n5989 = ~x26 & n1966;
  assign n5990 = ~n5988 & ~n5989;
  assign n5991 = x27 & n1969;
  assign n5992 = x26 & n1971;
  assign n5993 = ~n5991 & ~n5992;
  assign n5994 = n5990 & n5993;
  assign n6004 = n6003 ^ n5994;
  assign n6012 = n6011 ^ n6004;
  assign n6016 = n6015 ^ n6012;
  assign n6020 = n6019 ^ n6016;
  assign n5984 = n5925 ^ n5920;
  assign n5985 = ~n5921 & n5984;
  assign n5986 = n5985 ^ n5913;
  assign n5974 = ~x25 & n2406;
  assign n5975 = ~x24 & n2408;
  assign n5976 = ~n5974 & ~n5975;
  assign n5977 = x25 & n2399;
  assign n5978 = x24 & n2403;
  assign n5979 = ~n5977 & ~n5978;
  assign n5980 = n5976 & n5979;
  assign n5973 = x19 & x63;
  assign n5981 = n5980 ^ n5973;
  assign n5966 = ~x29 & n1687;
  assign n5967 = ~x28 & n1691;
  assign n5968 = ~n5966 & ~n5967;
  assign n5969 = x29 & n1694;
  assign n5970 = x28 & n1696;
  assign n5971 = ~n5969 & ~n5970;
  assign n5972 = n5968 & n5971;
  assign n5982 = n5981 ^ n5972;
  assign n5957 = ~x21 & n3098;
  assign n5958 = ~x20 & n3102;
  assign n5959 = ~n5957 & ~n5958;
  assign n5960 = x21 & n3105;
  assign n5961 = x20 & n3107;
  assign n5962 = ~n5960 & ~n5961;
  assign n5963 = n5959 & n5962;
  assign n5950 = x23 & n2688;
  assign n5951 = x22 & n2690;
  assign n5952 = ~n5950 & ~n5951;
  assign n5953 = ~x23 & n2681;
  assign n5954 = ~x22 & n2685;
  assign n5955 = ~n5953 & ~n5954;
  assign n5956 = n5952 & n5955;
  assign n5964 = n5963 ^ n5956;
  assign n5965 = n5964 ^ n5913;
  assign n5983 = n5982 ^ n5965;
  assign n5987 = n5986 ^ n5983;
  assign n6021 = n6020 ^ n5987;
  assign n6025 = n6024 ^ n6021;
  assign n6029 = n6028 ^ n6025;
  assign n6033 = n6032 ^ n6029;
  assign n6108 = n6032 ^ n6025;
  assign n6109 = ~n6029 & ~n6108;
  assign n6110 = n6109 ^ n6032;
  assign n6103 = n6024 ^ n5987;
  assign n6104 = n6024 ^ n6020;
  assign n6105 = ~n6103 & ~n6104;
  assign n6106 = n6105 ^ n5987;
  assign n6099 = n6019 ^ n6015;
  assign n6100 = n6016 & n6099;
  assign n6101 = n6100 ^ n6012;
  assign n6095 = n5986 ^ n5982;
  assign n6096 = ~n5983 & ~n6095;
  assign n6097 = n6096 ^ n5965;
  assign n6090 = n6007 ^ n6004;
  assign n6091 = n6011 & n6090;
  assign n6092 = n6091 ^ n6004;
  assign n6086 = n5980 ^ n5972;
  assign n6087 = ~n5981 & ~n6086;
  assign n6088 = n6087 ^ n5973;
  assign n6082 = n6002 ^ n5994;
  assign n6083 = ~n6003 & ~n6082;
  assign n6084 = n6083 ^ n5995;
  assign n6079 = x53 ^ x31;
  assign n6080 = n1399 & n6079;
  assign n6081 = ~n1396 & ~n6080;
  assign n6085 = n6084 ^ n6081;
  assign n6089 = n6088 ^ n6085;
  assign n6093 = n6092 ^ n6089;
  assign n6075 = n5956 ^ n5913;
  assign n6076 = ~n5964 & n6075;
  assign n6077 = n6076 ^ n5913;
  assign n6065 = x26 & n2399;
  assign n6066 = x25 & n2403;
  assign n6067 = ~n6065 & ~n6066;
  assign n6068 = ~x26 & n2406;
  assign n6069 = ~x25 & n2408;
  assign n6070 = ~n6068 & ~n6069;
  assign n6071 = n6067 & n6070;
  assign n6058 = ~x30 & n1687;
  assign n6059 = ~x29 & n1691;
  assign n6060 = ~n6058 & ~n6059;
  assign n6061 = x30 & n1694;
  assign n6062 = x29 & n1696;
  assign n6063 = ~n6061 & ~n6062;
  assign n6064 = n6060 & n6063;
  assign n6072 = n6071 ^ n6064;
  assign n6051 = ~x24 & n2681;
  assign n6052 = ~x23 & n2685;
  assign n6053 = ~n6051 & ~n6052;
  assign n6054 = x24 & n2688;
  assign n6055 = x23 & n2690;
  assign n6056 = ~n6054 & ~n6055;
  assign n6057 = n6053 & n6056;
  assign n6073 = n6072 ^ n6057;
  assign n6042 = ~x22 & n3098;
  assign n6043 = ~x21 & n3102;
  assign n6044 = ~n6042 & ~n6043;
  assign n6045 = x22 & n3105;
  assign n6046 = x21 & n3107;
  assign n6047 = ~n6045 & ~n6046;
  assign n6048 = n6044 & n6047;
  assign n6035 = ~x28 & n1962;
  assign n6036 = ~x27 & n1966;
  assign n6037 = ~n6035 & ~n6036;
  assign n6038 = x28 & n1969;
  assign n6039 = x27 & n1971;
  assign n6040 = ~n6038 & ~n6039;
  assign n6041 = n6037 & n6040;
  assign n6049 = n6048 ^ n6041;
  assign n6034 = x20 & x63;
  assign n6050 = n6049 ^ n6034;
  assign n6074 = n6073 ^ n6050;
  assign n6078 = n6077 ^ n6074;
  assign n6094 = n6093 ^ n6078;
  assign n6098 = n6097 ^ n6094;
  assign n6102 = n6101 ^ n6098;
  assign n6107 = n6106 ^ n6102;
  assign n6111 = n6110 ^ n6107;
  assign n6181 = n6110 ^ n6102;
  assign n6182 = n6107 & n6181;
  assign n6183 = n6182 ^ n6110;
  assign n6177 = n6101 ^ n6097;
  assign n6178 = ~n6098 & ~n6177;
  assign n6179 = n6178 ^ n6094;
  assign n6173 = n6089 ^ n6078;
  assign n6174 = ~n6093 & n6173;
  assign n6175 = n6174 ^ n6078;
  assign n6168 = n6077 ^ n6073;
  assign n6169 = ~n6074 & ~n6168;
  assign n6170 = n6169 ^ n6050;
  assign n6163 = n6088 ^ n6081;
  assign n6164 = n6088 ^ n6084;
  assign n6165 = n6163 & ~n6164;
  assign n6166 = n6165 ^ n6081;
  assign n6159 = n6071 ^ n6057;
  assign n6160 = n6072 & ~n6159;
  assign n6161 = n6160 ^ n6064;
  assign n6157 = x21 & x63;
  assign n6158 = n6157 ^ n6081;
  assign n6162 = n6161 ^ n6158;
  assign n6167 = n6166 ^ n6162;
  assign n6171 = n6170 ^ n6167;
  assign n6152 = n6041 ^ n6034;
  assign n6153 = ~n6049 & ~n6152;
  assign n6154 = n6153 ^ n6034;
  assign n6143 = x29 & n1969;
  assign n6144 = x28 & n1971;
  assign n6145 = ~n6143 & ~n6144;
  assign n6146 = ~x29 & n1962;
  assign n6147 = ~x28 & n1966;
  assign n6148 = ~n6146 & ~n6147;
  assign n6149 = n6145 & n6148;
  assign n6136 = ~x25 & n2681;
  assign n6137 = ~x24 & n2685;
  assign n6138 = ~n6136 & ~n6137;
  assign n6139 = x25 & n2688;
  assign n6140 = x24 & n2690;
  assign n6141 = ~n6139 & ~n6140;
  assign n6142 = n6138 & n6141;
  assign n6150 = n6149 ^ n6142;
  assign n6129 = x23 & n3105;
  assign n6130 = x22 & n3107;
  assign n6131 = ~n6129 & ~n6130;
  assign n6132 = ~x23 & n3098;
  assign n6133 = ~x22 & n3102;
  assign n6134 = ~n6132 & ~n6133;
  assign n6135 = n6131 & n6134;
  assign n6151 = n6150 ^ n6135;
  assign n6155 = n6154 ^ n6151;
  assign n6120 = x31 & n1694;
  assign n6121 = x30 & n1696;
  assign n6122 = ~n6120 & ~n6121;
  assign n6123 = ~x31 & n1687;
  assign n6124 = ~x30 & n1691;
  assign n6125 = ~n6123 & ~n6124;
  assign n6126 = n6122 & n6125;
  assign n6119 = ~n1396 & ~n1400;
  assign n6127 = n6126 ^ n6119;
  assign n6112 = ~x27 & n2406;
  assign n6113 = ~x26 & n2408;
  assign n6114 = ~n6112 & ~n6113;
  assign n6115 = x27 & n2399;
  assign n6116 = x26 & n2403;
  assign n6117 = ~n6115 & ~n6116;
  assign n6118 = n6114 & n6117;
  assign n6128 = n6127 ^ n6118;
  assign n6156 = n6155 ^ n6128;
  assign n6172 = n6171 ^ n6156;
  assign n6176 = n6175 ^ n6172;
  assign n6180 = n6179 ^ n6176;
  assign n6184 = n6183 ^ n6180;
  assign n6249 = n6183 ^ n6176;
  assign n6250 = n6180 & ~n6249;
  assign n6251 = n6250 ^ n6183;
  assign n6245 = n6175 ^ n6171;
  assign n6246 = ~n6172 & ~n6245;
  assign n6247 = n6246 ^ n6156;
  assign n6240 = n6170 ^ n6162;
  assign n6241 = n6170 ^ n6166;
  assign n6242 = n6240 & ~n6241;
  assign n6243 = n6242 ^ n6162;
  assign n6234 = n6151 ^ n6128;
  assign n6235 = n6154 ^ n6128;
  assign n6236 = ~n6234 & ~n6235;
  assign n6237 = n6236 ^ n6151;
  assign n6230 = n6161 ^ n6081;
  assign n6231 = ~n6158 & ~n6230;
  assign n6232 = n6231 ^ n6157;
  assign n6221 = ~x28 & n2406;
  assign n6222 = ~x27 & n2408;
  assign n6223 = ~n6221 & ~n6222;
  assign n6224 = x28 & n2399;
  assign n6225 = x27 & n2403;
  assign n6226 = ~n6224 & ~n6225;
  assign n6227 = n6223 & n6226;
  assign n6220 = x22 & x63;
  assign n6228 = n6227 ^ n6220;
  assign n6213 = x30 & n1969;
  assign n6214 = x29 & n1971;
  assign n6215 = ~n6213 & ~n6214;
  assign n6216 = ~x30 & n1962;
  assign n6217 = ~x29 & n1966;
  assign n6218 = ~n6216 & ~n6217;
  assign n6219 = n6215 & n6218;
  assign n6229 = n6228 ^ n6219;
  assign n6233 = n6232 ^ n6229;
  assign n6238 = n6237 ^ n6233;
  assign n6207 = n6142 ^ n6135;
  assign n6208 = n6149 ^ n6135;
  assign n6209 = n6207 & ~n6208;
  assign n6210 = n6209 ^ n6142;
  assign n6204 = n6126 ^ n6118;
  assign n6205 = ~n6127 & ~n6204;
  assign n6206 = n6205 ^ n6119;
  assign n6211 = n6210 ^ n6206;
  assign n6195 = ~x26 & n2681;
  assign n6196 = ~x25 & n2685;
  assign n6197 = ~n6195 & ~n6196;
  assign n6198 = x26 & n2688;
  assign n6199 = x25 & n2690;
  assign n6200 = ~n6198 & ~n6199;
  assign n6201 = n6197 & n6200;
  assign n6188 = x24 & n3105;
  assign n6189 = x23 & n3107;
  assign n6190 = ~n6188 & ~n6189;
  assign n6191 = ~x24 & n3098;
  assign n6192 = ~x23 & n3102;
  assign n6193 = ~n6191 & ~n6192;
  assign n6194 = n6190 & n6193;
  assign n6202 = n6201 ^ n6194;
  assign n6185 = x55 ^ x31;
  assign n6186 = n1690 & n6185;
  assign n6187 = ~n1687 & ~n6186;
  assign n6203 = n6202 ^ n6187;
  assign n6212 = n6211 ^ n6203;
  assign n6239 = n6238 ^ n6212;
  assign n6244 = n6243 ^ n6239;
  assign n6248 = n6247 ^ n6244;
  assign n6252 = n6251 ^ n6248;
  assign n6310 = n6251 ^ n6244;
  assign n6311 = n6248 & n6310;
  assign n6312 = n6311 ^ n6251;
  assign n6306 = n6243 ^ n6238;
  assign n6307 = n6239 & ~n6306;
  assign n6308 = n6307 ^ n6212;
  assign n6302 = n6237 ^ n6232;
  assign n6303 = ~n6233 & n6302;
  assign n6304 = n6303 ^ n6229;
  assign n6298 = n6206 ^ n6203;
  assign n6299 = n6211 & ~n6298;
  assign n6300 = n6299 ^ n6203;
  assign n6292 = n6220 ^ n6219;
  assign n6293 = n6227 ^ n6219;
  assign n6294 = n6292 & n6293;
  assign n6295 = n6294 ^ n6220;
  assign n6283 = ~x31 & n1962;
  assign n6284 = ~x30 & n1966;
  assign n6285 = ~n6283 & ~n6284;
  assign n6286 = x31 & n1969;
  assign n6287 = x30 & n1971;
  assign n6288 = ~n6286 & ~n6287;
  assign n6289 = n6285 & n6288;
  assign n6282 = ~n1687 & ~n1691;
  assign n6290 = n6289 ^ n6282;
  assign n6275 = ~x27 & n2681;
  assign n6276 = ~x26 & n2685;
  assign n6277 = ~n6275 & ~n6276;
  assign n6278 = x27 & n2688;
  assign n6279 = x26 & n2690;
  assign n6280 = ~n6278 & ~n6279;
  assign n6281 = n6277 & n6280;
  assign n6291 = n6290 ^ n6281;
  assign n6296 = n6295 ^ n6291;
  assign n6270 = n6194 ^ n6187;
  assign n6271 = ~n6202 & n6270;
  assign n6272 = n6271 ^ n6187;
  assign n6273 = n6272 ^ n6219;
  assign n6261 = ~x25 & n3098;
  assign n6262 = ~x24 & n3102;
  assign n6263 = ~n6261 & ~n6262;
  assign n6264 = x25 & n3105;
  assign n6265 = x24 & n3107;
  assign n6266 = ~n6264 & ~n6265;
  assign n6267 = n6263 & n6266;
  assign n6254 = x29 & n2399;
  assign n6255 = x28 & n2403;
  assign n6256 = ~n6254 & ~n6255;
  assign n6257 = ~x29 & n2406;
  assign n6258 = ~x28 & n2408;
  assign n6259 = ~n6257 & ~n6258;
  assign n6260 = n6256 & n6259;
  assign n6268 = n6267 ^ n6260;
  assign n6253 = x23 & x63;
  assign n6269 = n6268 ^ n6253;
  assign n6274 = n6273 ^ n6269;
  assign n6297 = n6296 ^ n6274;
  assign n6301 = n6300 ^ n6297;
  assign n6305 = n6304 ^ n6301;
  assign n6309 = n6308 ^ n6305;
  assign n6313 = n6312 ^ n6309;
  assign n6364 = n6312 ^ n6305;
  assign n6365 = ~n6309 & n6364;
  assign n6366 = n6365 ^ n6312;
  assign n6360 = n6304 ^ n6300;
  assign n6361 = ~n6301 & ~n6360;
  assign n6362 = n6361 ^ n6297;
  assign n6356 = n6295 ^ n6274;
  assign n6357 = n6296 & ~n6356;
  assign n6358 = n6357 ^ n6291;
  assign n6351 = n6269 ^ n6219;
  assign n6352 = n6272 ^ n6269;
  assign n6353 = ~n6351 & n6352;
  assign n6354 = n6353 ^ n6219;
  assign n6346 = n6289 ^ n6281;
  assign n6347 = ~n6290 & ~n6346;
  assign n6348 = n6347 ^ n6282;
  assign n6337 = x26 & n3105;
  assign n6338 = x25 & n3107;
  assign n6339 = ~n6337 & ~n6338;
  assign n6340 = ~x26 & n3098;
  assign n6341 = ~x25 & n3102;
  assign n6342 = ~n6340 & ~n6341;
  assign n6343 = n6339 & n6342;
  assign n6336 = x24 & x63;
  assign n6344 = n6343 ^ n6336;
  assign n6333 = x57 ^ x31;
  assign n6334 = n1965 & n6333;
  assign n6335 = ~n1962 & ~n6334;
  assign n6345 = n6344 ^ n6335;
  assign n6349 = n6348 ^ n6345;
  assign n6329 = n6260 ^ n6253;
  assign n6330 = ~n6268 & ~n6329;
  assign n6331 = n6330 ^ n6253;
  assign n6321 = ~x28 & n2681;
  assign n6322 = ~x27 & n2685;
  assign n6323 = ~n6321 & ~n6322;
  assign n6324 = x28 & n2688;
  assign n6325 = x27 & n2690;
  assign n6326 = ~n6324 & ~n6325;
  assign n6327 = n6323 & n6326;
  assign n6314 = ~x30 & n2406;
  assign n6315 = ~x29 & n2408;
  assign n6316 = ~n6314 & ~n6315;
  assign n6317 = x30 & n2399;
  assign n6318 = x29 & n2403;
  assign n6319 = ~n6317 & ~n6318;
  assign n6320 = n6316 & n6319;
  assign n6328 = n6327 ^ n6320;
  assign n6332 = n6331 ^ n6328;
  assign n6350 = n6349 ^ n6332;
  assign n6355 = n6354 ^ n6350;
  assign n6359 = n6358 ^ n6355;
  assign n6363 = n6362 ^ n6359;
  assign n6367 = n6366 ^ n6363;
  assign n6413 = n6366 ^ n6359;
  assign n6414 = ~n6363 & n6413;
  assign n6415 = n6414 ^ n6366;
  assign n6409 = n6358 ^ n6354;
  assign n6410 = n6355 & n6409;
  assign n6411 = n6410 ^ n6350;
  assign n6405 = n6348 ^ n6332;
  assign n6406 = n6349 & n6405;
  assign n6407 = n6406 ^ n6345;
  assign n6401 = n6331 ^ n6327;
  assign n6402 = ~n6328 & n6401;
  assign n6403 = n6402 ^ n6320;
  assign n6395 = n6336 ^ n6335;
  assign n6396 = n6343 ^ n6335;
  assign n6397 = ~n6395 & ~n6396;
  assign n6398 = n6397 ^ n6336;
  assign n6386 = ~x31 & n2406;
  assign n6387 = ~x30 & n2408;
  assign n6388 = ~n6386 & ~n6387;
  assign n6389 = x31 & n2399;
  assign n6390 = x30 & n2403;
  assign n6391 = ~n6389 & ~n6390;
  assign n6392 = n6388 & n6391;
  assign n6385 = ~n1962 & ~n1966;
  assign n6393 = n6392 ^ n6385;
  assign n6378 = x27 & n3105;
  assign n6379 = x26 & n3107;
  assign n6380 = ~n6378 & ~n6379;
  assign n6381 = ~x27 & n3098;
  assign n6382 = ~x26 & n3102;
  assign n6383 = ~n6381 & ~n6382;
  assign n6384 = n6380 & n6383;
  assign n6394 = n6393 ^ n6384;
  assign n6399 = n6398 ^ n6394;
  assign n6369 = ~x29 & n2681;
  assign n6370 = ~x28 & n2685;
  assign n6371 = ~n6369 & ~n6370;
  assign n6372 = x29 & n2688;
  assign n6373 = x28 & n2690;
  assign n6374 = ~n6372 & ~n6373;
  assign n6375 = n6371 & n6374;
  assign n6368 = x25 & x63;
  assign n6376 = n6375 ^ n6368;
  assign n6377 = n6376 ^ n6320;
  assign n6400 = n6399 ^ n6377;
  assign n6404 = n6403 ^ n6400;
  assign n6408 = n6407 ^ n6404;
  assign n6412 = n6411 ^ n6408;
  assign n6416 = n6415 ^ n6412;
  assign n6456 = n6415 ^ n6408;
  assign n6457 = n6412 & n6456;
  assign n6458 = n6457 ^ n6415;
  assign n6452 = n6407 ^ n6403;
  assign n6453 = n6404 & ~n6452;
  assign n6454 = n6453 ^ n6400;
  assign n6448 = n6394 ^ n6377;
  assign n6449 = ~n6399 & n6448;
  assign n6450 = n6449 ^ n6377;
  assign n6443 = n6368 ^ n6320;
  assign n6444 = n6375 ^ n6320;
  assign n6445 = ~n6443 & ~n6444;
  assign n6446 = n6445 ^ n6368;
  assign n6437 = n6385 ^ n6384;
  assign n6438 = n6392 ^ n6384;
  assign n6439 = ~n6437 & ~n6438;
  assign n6440 = n6439 ^ n6385;
  assign n6434 = x59 ^ x31;
  assign n6435 = n2402 & n6434;
  assign n6436 = ~n2406 & ~n6435;
  assign n6441 = n6440 ^ n6436;
  assign n6425 = ~x30 & n2681;
  assign n6426 = ~x29 & n2685;
  assign n6427 = ~n6425 & ~n6426;
  assign n6428 = x30 & n2688;
  assign n6429 = x29 & n2690;
  assign n6430 = ~n6428 & ~n6429;
  assign n6431 = n6427 & n6430;
  assign n6424 = x26 & x63;
  assign n6432 = n6431 ^ n6424;
  assign n6417 = x28 & n3105;
  assign n6418 = x27 & n3107;
  assign n6419 = ~n6417 & ~n6418;
  assign n6420 = ~x28 & n3098;
  assign n6421 = ~x27 & n3102;
  assign n6422 = ~n6420 & ~n6421;
  assign n6423 = n6419 & n6422;
  assign n6433 = n6432 ^ n6423;
  assign n6442 = n6441 ^ n6433;
  assign n6447 = n6446 ^ n6442;
  assign n6451 = n6450 ^ n6447;
  assign n6455 = n6454 ^ n6451;
  assign n6459 = n6458 ^ n6455;
  assign n6493 = n6458 ^ n6451;
  assign n6494 = ~n6455 & n6493;
  assign n6495 = n6494 ^ n6458;
  assign n6489 = n6450 ^ n6442;
  assign n6490 = n6447 & ~n6489;
  assign n6491 = n6490 ^ n6446;
  assign n6484 = n6436 ^ n6433;
  assign n6485 = n6440 ^ n6433;
  assign n6486 = n6484 & ~n6485;
  assign n6487 = n6486 ^ n6436;
  assign n6479 = n6431 ^ n6423;
  assign n6480 = ~n6432 & ~n6479;
  assign n6481 = n6480 ^ n6424;
  assign n6471 = ~x29 & n3098;
  assign n6472 = ~x28 & n3102;
  assign n6473 = ~n6471 & ~n6472;
  assign n6474 = x29 & n3105;
  assign n6475 = x28 & n3107;
  assign n6476 = ~n6474 & ~n6475;
  assign n6477 = n6473 & n6476;
  assign n6478 = n6477 ^ n6436;
  assign n6482 = n6481 ^ n6478;
  assign n6462 = x31 & n2688;
  assign n6463 = x30 & n2690;
  assign n6464 = ~n6462 & ~n6463;
  assign n6465 = ~x31 & n2681;
  assign n6466 = ~x30 & n2685;
  assign n6467 = ~n6465 & ~n6466;
  assign n6468 = n6464 & n6467;
  assign n6461 = ~n2406 & ~n2408;
  assign n6469 = n6468 ^ n6461;
  assign n6460 = x27 & x63;
  assign n6470 = n6469 ^ n6460;
  assign n6483 = n6482 ^ n6470;
  assign n6488 = n6487 ^ n6483;
  assign n6492 = n6491 ^ n6488;
  assign n6496 = n6495 ^ n6492;
  assign n6522 = n6495 ^ n6488;
  assign n6523 = n6492 & ~n6522;
  assign n6524 = n6523 ^ n6495;
  assign n6518 = n6487 ^ n6482;
  assign n6519 = ~n6483 & ~n6518;
  assign n6520 = n6519 ^ n6470;
  assign n6514 = n6481 ^ n6477;
  assign n6515 = n6478 & n6514;
  assign n6516 = n6515 ^ n6436;
  assign n6510 = n6461 ^ n6460;
  assign n6511 = n6469 & n6510;
  assign n6512 = n6511 ^ n6460;
  assign n6501 = ~x30 & n3098;
  assign n6502 = ~x29 & n3102;
  assign n6503 = ~n6501 & ~n6502;
  assign n6504 = x30 & n3105;
  assign n6505 = x29 & n3107;
  assign n6506 = ~n6504 & ~n6505;
  assign n6507 = n6503 & n6506;
  assign n6500 = x28 & x63;
  assign n6508 = n6507 ^ n6500;
  assign n6497 = x61 ^ x31;
  assign n6498 = n2684 & n6497;
  assign n6499 = ~n2681 & ~n6498;
  assign n6509 = n6508 ^ n6499;
  assign n6513 = n6512 ^ n6509;
  assign n6517 = n6516 ^ n6513;
  assign n6521 = n6520 ^ n6517;
  assign n6525 = n6524 ^ n6521;
  assign n6547 = n6524 ^ n6517;
  assign n6548 = n6521 & n6547;
  assign n6549 = n6548 ^ n6524;
  assign n6543 = n6516 ^ n6512;
  assign n6544 = ~n6513 & n6543;
  assign n6545 = n6544 ^ n6509;
  assign n6538 = n6500 ^ n6499;
  assign n6539 = n6507 ^ n6499;
  assign n6540 = n6538 & n6539;
  assign n6541 = n6540 ^ n6500;
  assign n6528 = x31 & n3105;
  assign n6529 = x30 & n3107;
  assign n6530 = ~n6528 & ~n6529;
  assign n6531 = ~x31 & n3098;
  assign n6532 = ~x30 & n3102;
  assign n6533 = ~n6531 & ~n6532;
  assign n6534 = n6530 & n6533;
  assign n6527 = ~n2681 & ~n2685;
  assign n6535 = n6534 ^ n6527;
  assign n6526 = x29 & x63;
  assign n6536 = n6535 ^ n6526;
  assign n6537 = n6536 ^ n6499;
  assign n6542 = n6541 ^ n6537;
  assign n6546 = n6545 ^ n6542;
  assign n6550 = n6549 ^ n6546;
  assign n6564 = n6549 ^ n6542;
  assign n6565 = n6546 & n6564;
  assign n6566 = n6565 ^ n6549;
  assign n6560 = n6541 ^ n6536;
  assign n6561 = n6537 & n6560;
  assign n6562 = n6561 ^ n6499;
  assign n6556 = n6527 ^ n6526;
  assign n6557 = n6535 & n6556;
  assign n6558 = n6557 ^ n6526;
  assign n6552 = x63 ^ x31;
  assign n6553 = n3101 & n6552;
  assign n6554 = ~n3098 & ~n6553;
  assign n6551 = x30 & x63;
  assign n6555 = n6554 ^ n6551;
  assign n6559 = n6558 ^ n6555;
  assign n6563 = n6562 ^ n6559;
  assign n6567 = n6566 ^ n6563;
  assign n6576 = n6566 ^ n6559;
  assign n6577 = n6563 & n6576;
  assign n6578 = n6577 ^ n6566;
  assign n6572 = n6558 ^ n6554;
  assign n6573 = n6555 & n6572;
  assign n6574 = n6573 ^ n6551;
  assign n6568 = ~n2830 & ~n3101;
  assign n6569 = n6568 ^ x31;
  assign n6570 = x63 & ~n6569;
  assign n6571 = n6570 ^ n6551;
  assign n6575 = n6574 ^ n6571;
  assign n6579 = n6578 ^ n6575;
  assign y0 = n65;
  assign y1 = n72;
  assign y2 = n81;
  assign y3 = ~n108;
  assign y4 = ~n129;
  assign y5 = n169;
  assign y6 = ~n202;
  assign y7 = n253;
  assign y8 = n300;
  assign y9 = n364;
  assign y10 = ~n422;
  assign y11 = ~n498;
  assign y12 = ~n567;
  assign y13 = n655;
  assign y14 = ~n736;
  assign y15 = n836;
  assign y16 = ~n932;
  assign y17 = n1044;
  assign y18 = n1150;
  assign y19 = ~n1274;
  assign y20 = n1395;
  assign y21 = ~n1532;
  assign y22 = ~n1663;
  assign y23 = n1812;
  assign y24 = n1954;
  assign y25 = ~n2117;
  assign y26 = n2274;
  assign y27 = ~n2448;
  assign y28 = n2616;
  assign y29 = ~n2802;
  assign y30 = n2981;
  assign y31 = n3179;
  assign y32 = ~n3366;
  assign y33 = n3556;
  assign y34 = n3742;
  assign y35 = ~n3926;
  assign y36 = ~n4106;
  assign y37 = n4280;
  assign y38 = ~n4443;
  assign y39 = ~n4602;
  assign y40 = ~n4754;
  assign y41 = n4904;
  assign y42 = n5043;
  assign y43 = ~n5181;
  assign y44 = ~n5307;
  assign y45 = ~n5432;
  assign y46 = n5548;
  assign y47 = n5659;
  assign y48 = ~n5761;
  assign y49 = ~n5857;
  assign y50 = n5949;
  assign y51 = n6033;
  assign y52 = ~n6111;
  assign y53 = ~n6184;
  assign y54 = ~n6252;
  assign y55 = n6313;
  assign y56 = n6367;
  assign y57 = ~n6416;
  assign y58 = n6459;
  assign y59 = ~n6496;
  assign y60 = ~n6525;
  assign y61 = ~n6550;
  assign y62 = ~n6567;
  assign y63 = n6579;
endmodule
