module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127;
  wire n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958;
  assign n65 = ~x0 & x1;
  assign n66 = x2 ^ x1;
  assign n67 = x0 & n66;
  assign n69 = ~x1 & x2;
  assign n68 = x3 ^ x2;
  assign n70 = n69 ^ n68;
  assign n71 = x0 & n70;
  assign n72 = n71 ^ n69;
  assign n73 = x1 & n68;
  assign n74 = ~x3 & ~x4;
  assign n75 = ~n73 & ~n74;
  assign n76 = x4 ^ x2;
  assign n77 = x3 & ~n76;
  assign n78 = n75 & ~n77;
  assign n79 = x0 & n78;
  assign n80 = x0 & x1;
  assign n81 = x4 & n80;
  assign n82 = n73 & ~n81;
  assign n83 = ~n79 & ~n82;
  assign n85 = ~x2 & x3;
  assign n89 = x3 & x4;
  assign n90 = ~n85 & ~n89;
  assign n91 = x1 & n78;
  assign n92 = n90 & ~n91;
  assign n93 = n92 ^ x5;
  assign n84 = x4 ^ x3;
  assign n86 = n85 ^ n84;
  assign n87 = x1 & n86;
  assign n88 = n87 ^ n85;
  assign n94 = n93 ^ n88;
  assign n95 = ~x0 & ~n94;
  assign n96 = n95 ^ n93;
  assign n97 = ~x3 & ~x5;
  assign n105 = x2 & x4;
  assign n106 = n97 & n105;
  assign n107 = x3 & x5;
  assign n108 = ~n106 & ~n107;
  assign n109 = n80 & ~n108;
  assign n110 = x0 & x5;
  assign n111 = ~n90 & n110;
  assign n112 = n65 & n89;
  assign n113 = ~n111 & ~n112;
  assign n114 = ~n109 & n113;
  assign n102 = x2 & n84;
  assign n100 = x0 & x6;
  assign n99 = x1 & x5;
  assign n101 = n100 ^ n99;
  assign n103 = n102 ^ n101;
  assign n98 = n81 & ~n97;
  assign n104 = n103 ^ n98;
  assign n115 = n114 ^ n104;
  assign n142 = ~n98 & n114;
  assign n127 = x5 & x6;
  assign n143 = n89 & n127;
  assign n144 = ~n103 & ~n143;
  assign n145 = ~n142 & ~n144;
  assign n117 = x2 & x5;
  assign n131 = x4 & x6;
  assign n132 = x1 & n131;
  assign n133 = ~n117 & n132;
  assign n134 = x1 & x6;
  assign n135 = ~x4 & ~n134;
  assign n136 = ~n133 & ~n135;
  assign n137 = ~x6 & n105;
  assign n138 = n99 & n137;
  assign n139 = n136 & ~n138;
  assign n120 = x3 & x6;
  assign n121 = x0 & n120;
  assign n122 = n99 ^ x4;
  assign n123 = ~n121 & ~n122;
  assign n124 = ~x3 & ~n100;
  assign n125 = x2 & ~n124;
  assign n126 = ~n123 & n125;
  assign n128 = n80 & ~n105;
  assign n129 = n127 & n128;
  assign n130 = ~n126 & ~n129;
  assign n140 = n139 ^ n130;
  assign n118 = n117 ^ n89;
  assign n116 = x0 & x7;
  assign n119 = n118 ^ n116;
  assign n141 = n140 ^ n119;
  assign n146 = n145 ^ n141;
  assign n161 = ~n130 & n139;
  assign n162 = n161 ^ n138;
  assign n156 = n132 ^ x2;
  assign n157 = x6 & n156;
  assign n155 = x0 & x8;
  assign n158 = n157 ^ n155;
  assign n153 = x1 & x7;
  assign n154 = n153 ^ n107;
  assign n159 = n158 ^ n154;
  assign n150 = n117 ^ n116;
  assign n151 = n118 & ~n150;
  assign n152 = n151 ^ n89;
  assign n160 = n159 ^ n152;
  assign n163 = n162 ^ n160;
  assign n147 = n145 ^ n140;
  assign n148 = n141 & ~n147;
  assign n149 = n148 ^ n145;
  assign n164 = n163 ^ n149;
  assign n184 = x3 & x7;
  assign n185 = x5 & x8;
  assign n186 = ~n184 & n185;
  assign n187 = x1 & n186;
  assign n188 = x1 & x8;
  assign n189 = ~x5 & ~n188;
  assign n190 = ~n187 & ~n189;
  assign n191 = n99 & n184;
  assign n192 = ~x8 & n191;
  assign n193 = n190 & ~n192;
  assign n183 = x0 & x9;
  assign n194 = n193 ^ n183;
  assign n176 = x4 & x8;
  assign n177 = n80 & n176;
  assign n178 = ~x2 & ~n177;
  assign n179 = x6 & n155;
  assign n180 = ~n132 & ~n179;
  assign n181 = ~n178 & ~n180;
  assign n173 = x4 & x5;
  assign n174 = n173 ^ n120;
  assign n172 = x2 & x7;
  assign n175 = n174 ^ n172;
  assign n182 = n181 ^ n175;
  assign n195 = n194 ^ n182;
  assign n168 = n162 ^ n149;
  assign n169 = n162 ^ n152;
  assign n170 = n168 & ~n169;
  assign n171 = n170 ^ n149;
  assign n196 = n195 ^ n171;
  assign n165 = n164 ^ n154;
  assign n166 = n159 & n165;
  assign n167 = n166 ^ n158;
  assign n197 = n196 ^ n167;
  assign n214 = n183 & n193;
  assign n215 = n214 ^ n192;
  assign n211 = x2 & x8;
  assign n212 = n211 ^ n184;
  assign n210 = x0 & x10;
  assign n213 = n212 ^ n210;
  assign n216 = n215 ^ n213;
  assign n207 = n172 & n174;
  assign n208 = ~n143 & ~n207;
  assign n204 = n185 ^ x9;
  assign n205 = x1 & n204;
  assign n206 = n205 ^ n131;
  assign n209 = n208 ^ n206;
  assign n217 = n216 ^ n209;
  assign n201 = n194 ^ n181;
  assign n202 = ~n182 & n201;
  assign n203 = n202 ^ n194;
  assign n218 = n217 ^ n203;
  assign n198 = n195 ^ n167;
  assign n199 = n196 & ~n198;
  assign n200 = n199 ^ n171;
  assign n219 = n218 ^ n200;
  assign n244 = n131 ^ x9;
  assign n245 = n185 & n244;
  assign n246 = n208 & ~n245;
  assign n247 = ~n185 & ~n244;
  assign n248 = x1 & ~n247;
  assign n249 = ~n246 & n248;
  assign n250 = ~x1 & n131;
  assign n251 = ~n208 & n250;
  assign n252 = ~n249 & ~n251;
  assign n241 = x4 & x7;
  assign n242 = n241 ^ n127;
  assign n240 = x0 & x11;
  assign n243 = n242 ^ n240;
  assign n253 = n252 ^ n243;
  assign n236 = x9 & n156;
  assign n235 = x3 & x8;
  assign n237 = n236 ^ n235;
  assign n232 = n211 ^ n210;
  assign n233 = n212 & ~n232;
  assign n234 = n233 ^ n184;
  assign n238 = n237 ^ n234;
  assign n230 = x1 & x10;
  assign n231 = n230 ^ x6;
  assign n239 = n238 ^ n231;
  assign n254 = n253 ^ n239;
  assign n225 = n203 & ~n209;
  assign n224 = ~n203 & n209;
  assign n226 = n225 ^ n224;
  assign n227 = ~n200 & n226;
  assign n228 = n227 ^ n225;
  assign n220 = n213 ^ n209;
  assign n221 = n220 ^ n203;
  assign n222 = n221 ^ n200;
  assign n223 = ~n216 & ~n222;
  assign n229 = n228 ^ n223;
  assign n255 = n254 ^ n229;
  assign n287 = n213 & n215;
  assign n288 = ~n200 & ~n287;
  assign n289 = ~n213 & ~n215;
  assign n290 = ~n225 & n254;
  assign n291 = ~n289 & ~n290;
  assign n292 = ~n288 & n291;
  assign n293 = n225 & ~n254;
  assign n294 = ~n292 & ~n293;
  assign n295 = n254 & ~n287;
  assign n296 = ~n224 & ~n295;
  assign n297 = n219 & n296;
  assign n298 = n294 & ~n297;
  assign n278 = x2 & n235;
  assign n279 = ~n132 & ~n278;
  assign n280 = ~x2 & ~n235;
  assign n281 = x9 & ~n280;
  assign n282 = ~n279 & n281;
  assign n274 = x6 & x10;
  assign n275 = x1 & n274;
  assign n276 = n275 ^ n176;
  assign n272 = x1 & x11;
  assign n271 = x5 & x7;
  assign n273 = n272 ^ n271;
  assign n277 = n276 ^ n273;
  assign n283 = n282 ^ n277;
  assign n267 = x3 & x9;
  assign n266 = x2 & x10;
  assign n268 = n267 ^ n266;
  assign n265 = x0 & x12;
  assign n269 = n268 ^ n265;
  assign n262 = n241 ^ n240;
  assign n263 = n242 & ~n262;
  assign n264 = n263 ^ n127;
  assign n270 = n269 ^ n264;
  assign n284 = n283 ^ n270;
  assign n259 = n234 ^ n231;
  assign n260 = n238 & ~n259;
  assign n261 = n260 ^ n237;
  assign n285 = n284 ^ n261;
  assign n256 = n243 ^ n239;
  assign n257 = ~n253 & ~n256;
  assign n258 = n257 ^ n252;
  assign n286 = n285 ^ n258;
  assign n299 = n298 ^ n286;
  assign n328 = x5 & x11;
  assign n329 = x1 & n328;
  assign n330 = x7 & ~n329;
  assign n327 = x1 & x12;
  assign n331 = n330 ^ n327;
  assign n324 = n266 ^ n265;
  assign n325 = n268 & ~n324;
  assign n326 = n325 ^ n267;
  assign n332 = n331 ^ n326;
  assign n321 = n282 ^ n261;
  assign n322 = ~n283 & ~n321;
  assign n318 = n283 ^ n269;
  assign n319 = n318 ^ n261;
  assign n320 = ~n270 & n319;
  assign n323 = n322 ^ n320;
  assign n333 = n332 ^ n323;
  assign n313 = n273 & n276;
  assign n314 = x8 & x10;
  assign n315 = n132 & n314;
  assign n316 = ~n313 & ~n315;
  assign n309 = x4 & x9;
  assign n308 = x3 & x10;
  assign n310 = n309 ^ n308;
  assign n307 = x0 & x13;
  assign n311 = n310 ^ n307;
  assign n304 = x6 & x7;
  assign n305 = n304 ^ n185;
  assign n303 = x2 & x11;
  assign n306 = n305 ^ n303;
  assign n312 = n311 ^ n306;
  assign n317 = n316 ^ n312;
  assign n334 = n333 ^ n317;
  assign n300 = n298 ^ n258;
  assign n301 = n286 & n300;
  assign n302 = n301 ^ n298;
  assign n335 = n334 ^ n302;
  assign n371 = ~n277 & ~n282;
  assign n372 = n264 & n333;
  assign n373 = n277 & n282;
  assign n374 = ~n261 & ~n373;
  assign n375 = n332 & ~n374;
  assign n376 = ~n372 & ~n375;
  assign n377 = ~n371 & ~n376;
  assign n378 = ~n332 & ~n373;
  assign n379 = n333 & ~n378;
  assign n380 = ~n377 & ~n379;
  assign n364 = n326 & n331;
  assign n365 = ~x12 & n153;
  assign n366 = n328 & n365;
  assign n367 = ~n364 & ~n366;
  assign n360 = x7 & n327;
  assign n359 = x5 & x9;
  assign n361 = n360 ^ n359;
  assign n358 = x4 & x10;
  assign n362 = n361 ^ n358;
  assign n355 = x3 & x11;
  assign n354 = x2 & x12;
  assign n356 = n355 ^ n354;
  assign n353 = x0 & x14;
  assign n357 = n356 ^ n353;
  assign n363 = n362 ^ n357;
  assign n368 = n367 ^ n363;
  assign n348 = n308 ^ n307;
  assign n349 = n310 & ~n348;
  assign n350 = n349 ^ n309;
  assign n345 = n304 ^ n303;
  assign n346 = n305 & ~n345;
  assign n347 = n346 ^ n185;
  assign n351 = n350 ^ n347;
  assign n343 = x6 & x8;
  assign n342 = x1 & x13;
  assign n344 = n343 ^ n342;
  assign n352 = n351 ^ n344;
  assign n369 = n368 ^ n352;
  assign n339 = n316 ^ n311;
  assign n340 = ~n312 & ~n339;
  assign n341 = n340 ^ n316;
  assign n370 = n369 ^ n341;
  assign n381 = n380 ^ n370;
  assign n336 = n333 ^ n302;
  assign n337 = ~n334 & n336;
  assign n338 = n337 ^ n302;
  assign n382 = n381 ^ n338;
  assign n417 = n380 ^ n341;
  assign n422 = n341 ^ n338;
  assign n423 = ~n417 & ~n422;
  assign n418 = n380 ^ n338;
  assign n419 = ~n417 & n418;
  assign n420 = n419 ^ n338;
  assign n421 = n420 ^ n352;
  assign n424 = n423 ^ n421;
  assign n425 = ~n369 & n424;
  assign n426 = n425 ^ n421;
  assign n410 = x5 & x10;
  assign n409 = x3 & x12;
  assign n411 = n410 ^ n409;
  assign n408 = x0 & x15;
  assign n412 = n411 ^ n408;
  assign n405 = n354 ^ n353;
  assign n406 = n356 & ~n405;
  assign n407 = n406 ^ n355;
  assign n413 = n412 ^ n407;
  assign n402 = n359 ^ n358;
  assign n403 = n361 & ~n402;
  assign n404 = n403 ^ n360;
  assign n414 = n413 ^ n404;
  assign n399 = n367 ^ n362;
  assign n400 = ~n363 & ~n399;
  assign n401 = n400 ^ n367;
  assign n415 = n414 ^ n401;
  assign n393 = n342 & n343;
  assign n394 = x8 & ~n393;
  assign n392 = x1 & x14;
  assign n395 = n394 ^ n392;
  assign n391 = x4 & x11;
  assign n396 = n395 ^ n391;
  assign n388 = x7 & x8;
  assign n387 = x6 & x9;
  assign n389 = n388 ^ n387;
  assign n386 = x2 & x13;
  assign n390 = n389 ^ n386;
  assign n397 = n396 ^ n390;
  assign n383 = n347 ^ n344;
  assign n384 = n351 & ~n383;
  assign n385 = n384 ^ n350;
  assign n398 = n397 ^ n385;
  assign n416 = n415 ^ n398;
  assign n427 = n426 ^ n416;
  assign n467 = ~n352 & n368;
  assign n468 = n467 ^ n420;
  assign n469 = n467 ^ n416;
  assign n470 = n468 & ~n469;
  assign n471 = n470 ^ n420;
  assign n475 = ~n341 & ~n380;
  assign n476 = ~n338 & n475;
  assign n477 = ~n369 & ~n476;
  assign n472 = ~n369 & n423;
  assign n473 = n472 ^ n369;
  assign n474 = ~n416 & ~n473;
  assign n478 = n477 ^ n474;
  assign n479 = ~n471 & ~n478;
  assign n461 = n391 & n395;
  assign n462 = ~x14 & n393;
  assign n463 = ~n461 & ~n462;
  assign n458 = n328 ^ n274;
  assign n457 = x0 & x16;
  assign n459 = n458 ^ n457;
  assign n454 = n409 ^ n408;
  assign n455 = n411 & ~n454;
  assign n456 = n455 ^ n410;
  assign n460 = n459 ^ n456;
  assign n464 = n463 ^ n460;
  assign n451 = n414 ^ n398;
  assign n452 = ~n415 & ~n451;
  assign n453 = n452 ^ n401;
  assign n465 = n464 ^ n453;
  assign n443 = x8 & x14;
  assign n444 = n443 ^ x15;
  assign n445 = x1 & n444;
  assign n442 = x7 & x9;
  assign n446 = n445 ^ n442;
  assign n439 = n387 ^ n386;
  assign n440 = n389 & ~n439;
  assign n441 = n440 ^ n388;
  assign n447 = n446 ^ n441;
  assign n436 = x4 & x12;
  assign n435 = x3 & x13;
  assign n437 = n436 ^ n435;
  assign n434 = x2 & x14;
  assign n438 = n437 ^ n434;
  assign n448 = n447 ^ n438;
  assign n431 = n407 ^ n404;
  assign n432 = ~n413 & n431;
  assign n433 = n432 ^ n404;
  assign n449 = n448 ^ n433;
  assign n428 = n396 ^ n385;
  assign n429 = ~n397 & n428;
  assign n430 = n429 ^ n385;
  assign n450 = n449 ^ n430;
  assign n466 = n465 ^ n450;
  assign n480 = n479 ^ n466;
  assign n525 = n442 ^ x15;
  assign n526 = n443 & n525;
  assign n527 = ~n441 & ~n526;
  assign n528 = ~n443 & ~n525;
  assign n529 = x1 & ~n528;
  assign n530 = ~n527 & n529;
  assign n531 = ~x1 & n442;
  assign n532 = n441 & n531;
  assign n533 = ~n530 & ~n532;
  assign n520 = n435 ^ n434;
  assign n521 = n437 & ~n520;
  assign n522 = n521 ^ n436;
  assign n517 = n457 ^ n328;
  assign n518 = n458 & ~n517;
  assign n519 = n518 ^ n274;
  assign n523 = n522 ^ n519;
  assign n515 = x1 & x16;
  assign n516 = n515 ^ x9;
  assign n524 = n523 ^ n516;
  assign n534 = n533 ^ n524;
  assign n512 = n463 ^ n456;
  assign n513 = ~n460 & ~n512;
  assign n514 = n513 ^ n463;
  assign n535 = n534 ^ n514;
  assign n509 = n447 ^ n433;
  assign n510 = ~n448 & n509;
  assign n511 = n510 ^ n433;
  assign n536 = n535 ^ n511;
  assign n504 = x9 & x15;
  assign n505 = n153 & n504;
  assign n502 = x0 & x17;
  assign n501 = x5 & x12;
  assign n503 = n502 ^ n501;
  assign n506 = n505 ^ n503;
  assign n498 = x6 & x11;
  assign n497 = x4 & x13;
  assign n499 = n498 ^ n497;
  assign n496 = x2 & x15;
  assign n500 = n499 ^ n496;
  assign n507 = n506 ^ n500;
  assign n493 = x8 & x9;
  assign n492 = x7 & x10;
  assign n494 = n493 ^ n492;
  assign n491 = x3 & x14;
  assign n495 = n494 ^ n491;
  assign n508 = n507 ^ n495;
  assign n537 = n536 ^ n508;
  assign n486 = n479 ^ n464;
  assign n487 = ~n465 & n486;
  assign n488 = n450 & n487;
  assign n489 = n488 ^ n450;
  assign n482 = n479 ^ n453;
  assign n483 = ~n465 & ~n482;
  assign n481 = n479 ^ n430;
  assign n484 = n483 ^ n481;
  assign n485 = ~n450 & n484;
  assign n490 = n489 ^ n485;
  assign n538 = n537 ^ n490;
  assign n587 = n483 ^ n479;
  assign n586 = ~n430 & ~n449;
  assign n588 = n587 ^ n586;
  assign n589 = n586 ^ n537;
  assign n590 = ~n588 & n589;
  assign n591 = n590 ^ n587;
  assign n595 = n489 & n537;
  assign n592 = ~n453 & ~n464;
  assign n593 = n479 & n592;
  assign n594 = n450 & ~n593;
  assign n596 = n595 ^ n594;
  assign n597 = n591 & ~n596;
  assign n578 = n519 ^ n516;
  assign n579 = n523 & ~n578;
  assign n580 = n579 ^ n522;
  assign n575 = n500 ^ n495;
  assign n576 = n507 & ~n575;
  assign n577 = n576 ^ n506;
  assign n581 = n580 ^ n577;
  assign n570 = n492 ^ n491;
  assign n571 = n494 & ~n570;
  assign n572 = n571 ^ n493;
  assign n567 = n497 ^ n496;
  assign n568 = n499 & ~n567;
  assign n569 = n568 ^ n498;
  assign n573 = n572 ^ n569;
  assign n563 = n503 & n505;
  assign n564 = x5 & x17;
  assign n565 = n265 & n564;
  assign n566 = ~n563 & ~n565;
  assign n574 = n573 ^ n566;
  assign n582 = n581 ^ n574;
  assign n559 = x9 & n515;
  assign n558 = x6 & x12;
  assign n560 = n559 ^ n558;
  assign n556 = x1 & x17;
  assign n557 = n556 ^ n314;
  assign n561 = n560 ^ n557;
  assign n552 = x7 & x11;
  assign n551 = x5 & x13;
  assign n553 = n552 ^ n551;
  assign n550 = x0 & x18;
  assign n554 = n553 ^ n550;
  assign n547 = x4 & x14;
  assign n546 = x3 & x15;
  assign n548 = n547 ^ n546;
  assign n545 = x2 & x16;
  assign n549 = n548 ^ n545;
  assign n555 = n554 ^ n549;
  assign n562 = n561 ^ n555;
  assign n583 = n582 ^ n562;
  assign n542 = n533 ^ n514;
  assign n543 = n534 & n542;
  assign n544 = n543 ^ n514;
  assign n584 = n583 ^ n544;
  assign n539 = n511 ^ n508;
  assign n540 = n536 & ~n539;
  assign n541 = n540 ^ n535;
  assign n585 = n584 ^ n541;
  assign n598 = n597 ^ n585;
  assign n646 = n582 ^ n544;
  assign n647 = n583 & n646;
  assign n648 = n647 ^ n544;
  assign n649 = n541 & ~n648;
  assign n650 = n562 & ~n582;
  assign n651 = ~n544 & n650;
  assign n652 = ~n649 & ~n651;
  assign n653 = n597 & ~n652;
  assign n654 = n541 & n651;
  assign n655 = ~n562 & n582;
  assign n656 = n544 & n655;
  assign n657 = ~n541 & n656;
  assign n658 = ~n654 & ~n657;
  assign n659 = ~n653 & n658;
  assign n660 = n541 & ~n656;
  assign n661 = n648 & ~n660;
  assign n662 = ~n597 & n661;
  assign n663 = n659 & ~n662;
  assign n637 = x8 & x17;
  assign n638 = n230 & n637;
  assign n639 = x10 & ~n638;
  assign n636 = x1 & x18;
  assign n640 = n639 ^ n636;
  assign n633 = n546 ^ n545;
  assign n634 = n548 & ~n633;
  assign n635 = n634 ^ n547;
  assign n641 = n640 ^ n635;
  assign n630 = n561 ^ n554;
  assign n631 = ~n555 & n630;
  assign n632 = n631 ^ n561;
  assign n642 = n641 ^ n632;
  assign n625 = x9 & x10;
  assign n624 = x8 & x11;
  assign n626 = n625 ^ n624;
  assign n623 = x3 & x16;
  assign n627 = n626 ^ n623;
  assign n620 = n551 ^ n550;
  assign n621 = n553 & ~n620;
  assign n622 = n621 ^ n552;
  assign n628 = n627 ^ n622;
  assign n617 = n558 ^ n557;
  assign n618 = n560 & ~n617;
  assign n619 = n618 ^ n559;
  assign n629 = n628 ^ n619;
  assign n643 = n642 ^ n629;
  assign n612 = x6 & x13;
  assign n611 = x7 & x12;
  assign n613 = n612 ^ n611;
  assign n610 = x5 & x14;
  assign n614 = n613 ^ n610;
  assign n607 = x4 & x15;
  assign n606 = x2 & x17;
  assign n608 = n607 ^ n606;
  assign n605 = x0 & x19;
  assign n609 = n608 ^ n605;
  assign n615 = n614 ^ n609;
  assign n602 = n569 ^ n566;
  assign n603 = n573 & n602;
  assign n604 = n603 ^ n572;
  assign n616 = n615 ^ n604;
  assign n644 = n643 ^ n616;
  assign n599 = n577 ^ n574;
  assign n600 = n581 & n599;
  assign n601 = n600 ^ n580;
  assign n645 = n644 ^ n601;
  assign n664 = n663 ^ n645;
  assign n718 = ~n645 & n652;
  assign n719 = ~n657 & ~n718;
  assign n720 = n597 & n719;
  assign n721 = ~n645 & ~n654;
  assign n722 = ~n661 & ~n721;
  assign n723 = ~n720 & ~n722;
  assign n709 = n606 ^ n605;
  assign n710 = n608 & ~n709;
  assign n711 = n710 ^ n607;
  assign n706 = n624 ^ n623;
  assign n707 = n626 & ~n706;
  assign n708 = n707 ^ n625;
  assign n712 = n711 ^ n708;
  assign n704 = x1 & x19;
  assign n703 = x9 & x11;
  assign n705 = n704 ^ n703;
  assign n713 = n712 ^ n705;
  assign n700 = n614 ^ n604;
  assign n701 = ~n615 & n700;
  assign n702 = n701 ^ n604;
  assign n714 = n713 ^ n702;
  assign n695 = x10 & n636;
  assign n694 = x0 & x20;
  assign n696 = n695 ^ n694;
  assign n693 = x7 & x13;
  assign n697 = n696 ^ n693;
  assign n690 = x8 & x12;
  assign n689 = x6 & x14;
  assign n691 = n690 ^ n689;
  assign n688 = x5 & x15;
  assign n692 = n691 ^ n688;
  assign n698 = n697 ^ n692;
  assign n685 = n611 ^ n610;
  assign n686 = n613 & ~n685;
  assign n687 = n686 ^ n612;
  assign n699 = n698 ^ n687;
  assign n715 = n714 ^ n699;
  assign n679 = n635 & n640;
  assign n680 = ~x18 & n638;
  assign n681 = ~n679 & ~n680;
  assign n676 = x4 & x16;
  assign n675 = x3 & x17;
  assign n677 = n676 ^ n675;
  assign n674 = x2 & x18;
  assign n678 = n677 ^ n674;
  assign n682 = n681 ^ n678;
  assign n671 = n622 ^ n619;
  assign n672 = ~n628 & n671;
  assign n673 = n672 ^ n619;
  assign n683 = n682 ^ n673;
  assign n668 = n641 ^ n629;
  assign n669 = n642 & ~n668;
  assign n670 = n669 ^ n632;
  assign n684 = n683 ^ n670;
  assign n716 = n715 ^ n684;
  assign n665 = n643 ^ n601;
  assign n666 = ~n644 & n665;
  assign n667 = n666 ^ n601;
  assign n717 = n716 ^ n667;
  assign n724 = n723 ^ n717;
  assign n777 = n670 & ~n683;
  assign n778 = n715 & n777;
  assign n779 = ~n667 & ~n778;
  assign n780 = n715 ^ n670;
  assign n781 = n684 & n780;
  assign n782 = n781 ^ n715;
  assign n783 = ~n779 & n782;
  assign n784 = ~n723 & n783;
  assign n785 = ~n670 & n683;
  assign n786 = ~n715 & n785;
  assign n787 = n786 ^ n778;
  assign n788 = ~n667 & n787;
  assign n789 = n788 ^ n778;
  assign n790 = ~n784 & ~n789;
  assign n791 = n667 & ~n786;
  assign n792 = ~n782 & ~n791;
  assign n793 = n723 & n792;
  assign n794 = n790 & ~n793;
  assign n768 = x10 & x11;
  assign n767 = x9 & x12;
  assign n769 = n768 ^ n767;
  assign n766 = x4 & x17;
  assign n770 = n769 ^ n766;
  assign n763 = x8 & x13;
  assign n762 = x7 & x14;
  assign n764 = n763 ^ n762;
  assign n761 = x6 & x15;
  assign n765 = n764 ^ n761;
  assign n771 = n770 ^ n765;
  assign n758 = x5 & x16;
  assign n757 = x3 & x18;
  assign n759 = n758 ^ n757;
  assign n756 = x2 & x19;
  assign n760 = n759 ^ n756;
  assign n772 = n771 ^ n760;
  assign n753 = n681 ^ n673;
  assign n754 = n682 & ~n753;
  assign n755 = n754 ^ n673;
  assign n773 = n772 ^ n755;
  assign n748 = n675 ^ n674;
  assign n749 = n677 & ~n748;
  assign n750 = n749 ^ n676;
  assign n745 = n689 ^ n688;
  assign n746 = n691 & ~n745;
  assign n747 = n746 ^ n690;
  assign n751 = n750 ^ n747;
  assign n742 = n694 ^ n693;
  assign n743 = n696 & ~n742;
  assign n744 = n743 ^ n695;
  assign n752 = n751 ^ n744;
  assign n774 = n773 ^ n752;
  assign n739 = n713 ^ n699;
  assign n740 = n714 & ~n739;
  assign n741 = n740 ^ n702;
  assign n775 = n774 ^ n741;
  assign n734 = n703 & n704;
  assign n735 = x11 & ~n734;
  assign n732 = x0 & x21;
  assign n731 = x1 & x20;
  assign n733 = n732 ^ n731;
  assign n736 = n735 ^ n733;
  assign n728 = n708 ^ n705;
  assign n729 = n712 & ~n728;
  assign n730 = n729 ^ n711;
  assign n737 = n736 ^ n730;
  assign n725 = n692 ^ n687;
  assign n726 = n698 & ~n725;
  assign n727 = n726 ^ n697;
  assign n738 = n737 ^ n727;
  assign n776 = n775 ^ n738;
  assign n795 = n794 ^ n776;
  assign n853 = ~n667 & ~n715;
  assign n854 = ~n723 & ~n853;
  assign n855 = n776 & ~n785;
  assign n856 = n667 & n715;
  assign n857 = ~n855 & ~n856;
  assign n858 = ~n854 & n857;
  assign n859 = ~n776 & n785;
  assign n860 = ~n858 & ~n859;
  assign n861 = n776 & ~n853;
  assign n862 = ~n777 & ~n861;
  assign n863 = n724 & n862;
  assign n864 = n860 & ~n863;
  assign n843 = x11 & x20;
  assign n844 = n843 ^ x21;
  assign n845 = x1 & n844;
  assign n842 = x10 & x12;
  assign n846 = n845 ^ n842;
  assign n839 = n767 ^ n766;
  assign n840 = n769 & ~n839;
  assign n841 = n840 ^ n768;
  assign n847 = n846 ^ n841;
  assign n836 = n750 ^ n744;
  assign n837 = ~n751 & n836;
  assign n838 = n837 ^ n744;
  assign n848 = n847 ^ n838;
  assign n833 = n765 ^ n760;
  assign n834 = n771 & ~n833;
  assign n835 = n834 ^ n770;
  assign n849 = n848 ^ n835;
  assign n830 = n772 ^ n752;
  assign n831 = n773 & ~n830;
  assign n832 = n831 ^ n755;
  assign n850 = n849 ^ n832;
  assign n823 = x7 & x15;
  assign n824 = n823 ^ n443;
  assign n822 = x0 & x22;
  assign n825 = n824 ^ n822;
  assign n819 = x9 & x13;
  assign n818 = x6 & x16;
  assign n820 = n819 ^ n818;
  assign n817 = x2 & x20;
  assign n821 = n820 ^ n817;
  assign n826 = n825 ^ n821;
  assign n814 = x4 & x18;
  assign n815 = n814 ^ n564;
  assign n813 = x3 & x19;
  assign n816 = n815 ^ n813;
  assign n827 = n826 ^ n816;
  assign n810 = n736 ^ n727;
  assign n811 = n737 & ~n810;
  assign n812 = n811 ^ n730;
  assign n828 = n827 ^ n812;
  assign n806 = n732 & ~n736;
  assign n807 = ~x20 & n734;
  assign n808 = ~n806 & ~n807;
  assign n802 = n762 ^ n761;
  assign n803 = n764 & ~n802;
  assign n804 = n803 ^ n763;
  assign n799 = n757 ^ n756;
  assign n800 = n759 & ~n799;
  assign n801 = n800 ^ n758;
  assign n805 = n804 ^ n801;
  assign n809 = n808 ^ n805;
  assign n829 = n828 ^ n809;
  assign n851 = n850 ^ n829;
  assign n796 = n774 ^ n738;
  assign n797 = n775 & ~n796;
  assign n798 = n797 ^ n741;
  assign n852 = n851 ^ n798;
  assign n865 = n864 ^ n852;
  assign n921 = n842 ^ x21;
  assign n922 = n843 & n921;
  assign n923 = ~n841 & ~n922;
  assign n924 = ~n843 & ~n921;
  assign n925 = x1 & ~n924;
  assign n926 = ~n923 & n925;
  assign n927 = ~x1 & n842;
  assign n928 = n841 & n927;
  assign n929 = ~n926 & ~n928;
  assign n918 = x6 & x17;
  assign n917 = x5 & x18;
  assign n919 = n918 ^ n917;
  assign n916 = x3 & x20;
  assign n920 = n919 ^ n916;
  assign n930 = n929 ^ n920;
  assign n913 = x11 & x12;
  assign n912 = x10 & x13;
  assign n914 = n913 ^ n912;
  assign n911 = x4 & x19;
  assign n915 = n914 ^ n911;
  assign n931 = n930 ^ n915;
  assign n908 = n847 ^ n835;
  assign n909 = n848 & ~n908;
  assign n910 = n909 ^ n838;
  assign n932 = n931 ^ n910;
  assign n903 = x9 & x14;
  assign n902 = x8 & x15;
  assign n904 = n903 ^ n902;
  assign n901 = x7 & x16;
  assign n905 = n904 ^ n901;
  assign n898 = n823 ^ n822;
  assign n899 = n824 & ~n898;
  assign n900 = n899 ^ n443;
  assign n906 = n905 ^ n900;
  assign n894 = x10 & n327;
  assign n895 = n894 ^ x2;
  assign n896 = x21 & n895;
  assign n893 = x0 & x23;
  assign n897 = n896 ^ n893;
  assign n907 = n906 ^ n897;
  assign n933 = n932 ^ n907;
  assign n886 = n814 ^ n813;
  assign n887 = n815 & ~n886;
  assign n888 = n887 ^ n564;
  assign n883 = n818 ^ n817;
  assign n884 = n820 & ~n883;
  assign n885 = n884 ^ n819;
  assign n889 = n888 ^ n885;
  assign n881 = x1 & x22;
  assign n882 = n881 ^ x12;
  assign n890 = n889 ^ n882;
  assign n878 = n821 ^ n816;
  assign n879 = n826 & ~n878;
  assign n880 = n879 ^ n825;
  assign n891 = n890 ^ n880;
  assign n875 = n808 ^ n804;
  assign n876 = ~n805 & ~n875;
  assign n877 = n876 ^ n808;
  assign n892 = n891 ^ n877;
  assign n934 = n933 ^ n892;
  assign n872 = n827 ^ n809;
  assign n873 = n828 & n872;
  assign n874 = n873 ^ n812;
  assign n935 = n934 ^ n874;
  assign n869 = n849 ^ n829;
  assign n870 = n850 & n869;
  assign n871 = n870 ^ n832;
  assign n936 = n935 ^ n871;
  assign n866 = n864 ^ n798;
  assign n867 = n852 & n866;
  assign n868 = n867 ^ n864;
  assign n937 = n936 ^ n868;
  assign n1005 = x22 & n327;
  assign n1003 = x1 & x23;
  assign n1002 = x11 & x13;
  assign n1004 = n1003 ^ n1002;
  assign n1006 = n1005 ^ n1004;
  assign n1001 = x0 & x24;
  assign n1007 = n1006 ^ n1001;
  assign n998 = x7 & x17;
  assign n997 = x6 & x18;
  assign n999 = n998 ^ n997;
  assign n996 = x2 & x22;
  assign n1000 = n999 ^ n996;
  assign n1008 = n1007 ^ n1000;
  assign n993 = n885 ^ n882;
  assign n994 = n889 & ~n993;
  assign n995 = n994 ^ n888;
  assign n1009 = n1008 ^ n995;
  assign n990 = n880 ^ n877;
  assign n991 = ~n891 & ~n990;
  assign n992 = n991 ^ n877;
  assign n1010 = n1009 ^ n992;
  assign n985 = n893 & n895;
  assign n986 = n266 & n327;
  assign n987 = ~n985 & ~n986;
  assign n988 = x21 & ~n987;
  assign n981 = x5 & x19;
  assign n980 = x4 & x20;
  assign n982 = n981 ^ n980;
  assign n979 = x3 & x21;
  assign n983 = n982 ^ n979;
  assign n976 = x10 & x14;
  assign n977 = n976 ^ n504;
  assign n975 = x8 & x16;
  assign n978 = n977 ^ n975;
  assign n984 = n983 ^ n978;
  assign n989 = n988 ^ n984;
  assign n1011 = n1010 ^ n989;
  assign n968 = n902 ^ n901;
  assign n969 = n904 & ~n968;
  assign n970 = n969 ^ n903;
  assign n965 = n917 ^ n916;
  assign n966 = n919 & ~n965;
  assign n967 = n966 ^ n918;
  assign n971 = n970 ^ n967;
  assign n962 = n912 ^ n911;
  assign n963 = n914 & ~n962;
  assign n964 = n963 ^ n913;
  assign n972 = n971 ^ n964;
  assign n959 = n920 ^ n915;
  assign n960 = ~n930 & ~n959;
  assign n961 = n960 ^ n929;
  assign n973 = n972 ^ n961;
  assign n956 = n905 ^ n897;
  assign n957 = n906 & ~n956;
  assign n958 = n957 ^ n900;
  assign n974 = n973 ^ n958;
  assign n1012 = n1011 ^ n974;
  assign n953 = n931 ^ n907;
  assign n954 = ~n932 & n953;
  assign n955 = n954 ^ n910;
  assign n1013 = n1012 ^ n955;
  assign n938 = n933 ^ n871;
  assign n939 = n892 ^ n874;
  assign n940 = ~n934 & n939;
  assign n941 = n938 & n940;
  assign n942 = ~n871 & ~n874;
  assign n943 = n892 & n933;
  assign n944 = ~n942 & ~n943;
  assign n945 = n944 ^ n868;
  assign n946 = n871 & n874;
  assign n947 = ~n892 & ~n933;
  assign n948 = ~n946 & ~n947;
  assign n949 = n948 ^ n944;
  assign n950 = ~n945 & n949;
  assign n951 = ~n941 & n950;
  assign n952 = n951 ^ n941;
  assign n1014 = n1013 ^ n952;
  assign n1084 = ~n868 & ~n946;
  assign n1085 = ~n947 & ~n1013;
  assign n1086 = ~n942 & ~n1085;
  assign n1087 = ~n1084 & n1086;
  assign n1088 = n947 & n1013;
  assign n1089 = ~n1087 & ~n1088;
  assign n1090 = ~n946 & ~n1013;
  assign n1091 = ~n943 & ~n1090;
  assign n1092 = ~n937 & n1091;
  assign n1093 = n1089 & ~n1092;
  assign n1075 = x10 & x15;
  assign n1074 = x2 & x23;
  assign n1076 = n1075 ^ n1074;
  assign n1073 = x0 & x25;
  assign n1077 = n1076 ^ n1073;
  assign n1070 = x6 & x19;
  assign n1069 = x4 & x21;
  assign n1071 = n1070 ^ n1069;
  assign n1068 = x3 & x22;
  assign n1072 = n1071 ^ n1068;
  assign n1078 = n1077 ^ n1072;
  assign n1065 = x9 & x16;
  assign n1066 = n1065 ^ n637;
  assign n1064 = x7 & x18;
  assign n1067 = n1066 ^ n1064;
  assign n1079 = n1078 ^ n1067;
  assign n1061 = n972 ^ n958;
  assign n1062 = ~n973 & ~n1061;
  assign n1063 = n1062 ^ n961;
  assign n1080 = n1079 ^ n1063;
  assign n1056 = x1 & x24;
  assign n1052 = x11 & x23;
  assign n1053 = x13 & n1052;
  assign n1054 = x1 & n1053;
  assign n1055 = n1054 ^ x13;
  assign n1057 = n1056 ^ n1055;
  assign n1049 = n980 ^ n979;
  assign n1050 = n982 & ~n1049;
  assign n1051 = n1050 ^ n981;
  assign n1058 = n1057 ^ n1051;
  assign n1046 = x12 & x13;
  assign n1045 = x11 & x14;
  assign n1047 = n1046 ^ n1045;
  assign n1044 = x5 & x20;
  assign n1048 = n1047 ^ n1044;
  assign n1059 = n1058 ^ n1048;
  assign n1041 = n967 ^ n964;
  assign n1042 = n971 & ~n1041;
  assign n1043 = n1042 ^ n970;
  assign n1060 = n1059 ^ n1043;
  assign n1081 = n1080 ^ n1060;
  assign n1038 = n1009 ^ n989;
  assign n1039 = ~n1010 & ~n1038;
  assign n1040 = n1039 ^ n992;
  assign n1082 = n1081 ^ n1040;
  assign n1032 = n1007 ^ n995;
  assign n1033 = ~n1008 & n1032;
  assign n1034 = n1033 ^ n995;
  assign n1029 = n988 ^ n983;
  assign n1030 = ~n984 & n1029;
  assign n1031 = n1030 ^ n988;
  assign n1035 = n1034 ^ n1031;
  assign n1024 = n976 ^ n975;
  assign n1025 = n977 & ~n1024;
  assign n1026 = n1025 ^ n504;
  assign n1021 = n997 ^ n996;
  assign n1022 = n999 & ~n1021;
  assign n1023 = n1022 ^ n998;
  assign n1027 = n1026 ^ n1023;
  assign n1018 = n1004 ^ n1001;
  assign n1019 = n1006 & ~n1018;
  assign n1020 = n1019 ^ n1005;
  assign n1028 = n1027 ^ n1020;
  assign n1036 = n1035 ^ n1028;
  assign n1015 = n1011 ^ n955;
  assign n1016 = ~n1012 & ~n1015;
  assign n1017 = n1016 ^ n955;
  assign n1037 = n1036 ^ n1017;
  assign n1083 = n1082 ^ n1037;
  assign n1094 = n1093 ^ n1083;
  assign n1168 = n1017 & n1036;
  assign n1169 = n1093 ^ n1081;
  assign n1170 = ~n1082 & n1169;
  assign n1171 = n1170 ^ n1093;
  assign n1172 = n1168 & ~n1171;
  assign n1173 = ~n1040 & ~n1081;
  assign n1174 = ~n1017 & ~n1036;
  assign n1175 = n1173 & ~n1174;
  assign n1176 = ~n1093 & n1175;
  assign n1177 = n1040 & n1081;
  assign n1178 = n1174 & n1177;
  assign n1179 = ~n1176 & ~n1178;
  assign n1180 = ~n1173 & n1174;
  assign n1181 = ~n1168 & n1177;
  assign n1182 = ~n1180 & ~n1181;
  assign n1183 = n1093 & ~n1182;
  assign n1184 = n1179 & ~n1183;
  assign n1185 = ~n1172 & n1184;
  assign n1153 = x24 & n1051;
  assign n1154 = ~n1053 & ~n1153;
  assign n1155 = x13 & x24;
  assign n1156 = x1 & ~n1155;
  assign n1157 = ~n1154 & n1156;
  assign n1158 = ~n1052 & n1056;
  assign n1159 = x13 & ~n1158;
  assign n1160 = n1051 & n1159;
  assign n1161 = ~n1157 & ~n1160;
  assign n1148 = n1065 ^ n1064;
  assign n1149 = n1066 & ~n1148;
  assign n1150 = n1149 ^ n637;
  assign n1145 = n1074 ^ n1073;
  assign n1146 = n1076 & ~n1145;
  assign n1147 = n1146 ^ n1075;
  assign n1151 = n1150 ^ n1147;
  assign n1143 = x24 & n342;
  assign n1141 = x0 & x26;
  assign n1140 = x8 & x18;
  assign n1142 = n1141 ^ n1140;
  assign n1144 = n1143 ^ n1142;
  assign n1152 = n1151 ^ n1144;
  assign n1162 = n1161 ^ n1152;
  assign n1137 = n1026 ^ n1020;
  assign n1138 = ~n1027 & n1137;
  assign n1139 = n1138 ^ n1020;
  assign n1163 = n1162 ^ n1139;
  assign n1134 = n1031 ^ n1028;
  assign n1135 = n1035 & ~n1134;
  assign n1136 = n1135 ^ n1034;
  assign n1164 = n1163 ^ n1136;
  assign n1129 = x7 & x19;
  assign n1128 = x3 & x23;
  assign n1130 = n1129 ^ n1128;
  assign n1127 = x2 & x24;
  assign n1131 = n1130 ^ n1127;
  assign n1124 = x6 & x20;
  assign n1123 = x5 & x21;
  assign n1125 = n1124 ^ n1123;
  assign n1122 = x4 & x22;
  assign n1126 = n1125 ^ n1122;
  assign n1132 = n1131 ^ n1126;
  assign n1119 = x11 & x15;
  assign n1118 = x10 & x16;
  assign n1120 = n1119 ^ n1118;
  assign n1117 = x9 & x17;
  assign n1121 = n1120 ^ n1117;
  assign n1133 = n1132 ^ n1121;
  assign n1165 = n1164 ^ n1133;
  assign n1114 = n1079 ^ n1060;
  assign n1115 = ~n1080 & ~n1114;
  assign n1116 = n1115 ^ n1063;
  assign n1166 = n1165 ^ n1116;
  assign n1107 = n1045 ^ n1044;
  assign n1108 = n1047 & ~n1107;
  assign n1109 = n1108 ^ n1046;
  assign n1104 = n1069 ^ n1068;
  assign n1105 = n1071 & ~n1104;
  assign n1106 = n1105 ^ n1070;
  assign n1110 = n1109 ^ n1106;
  assign n1102 = x1 & x25;
  assign n1101 = x12 & x14;
  assign n1103 = n1102 ^ n1101;
  assign n1111 = n1110 ^ n1103;
  assign n1098 = n1058 ^ n1043;
  assign n1099 = ~n1059 & n1098;
  assign n1100 = n1099 ^ n1043;
  assign n1112 = n1111 ^ n1100;
  assign n1095 = n1072 ^ n1067;
  assign n1096 = n1078 & ~n1095;
  assign n1097 = n1096 ^ n1077;
  assign n1113 = n1112 ^ n1097;
  assign n1167 = n1166 ^ n1113;
  assign n1186 = n1185 ^ n1167;
  assign n1263 = n1167 & ~n1174;
  assign n1264 = n1171 & ~n1263;
  assign n1265 = n1167 & ~n1177;
  assign n1266 = ~n1168 & ~n1265;
  assign n1267 = ~n1094 & n1266;
  assign n1268 = ~n1167 & n1174;
  assign n1269 = ~n1267 & ~n1268;
  assign n1270 = ~n1264 & n1269;
  assign n1253 = n1128 ^ n1127;
  assign n1254 = n1130 & ~n1253;
  assign n1255 = n1254 ^ n1129;
  assign n1250 = n1118 ^ n1117;
  assign n1251 = n1120 & ~n1250;
  assign n1252 = n1251 ^ n1119;
  assign n1256 = n1255 ^ n1252;
  assign n1247 = n1123 ^ n1122;
  assign n1248 = n1125 & ~n1247;
  assign n1249 = n1248 ^ n1124;
  assign n1257 = n1256 ^ n1249;
  assign n1244 = n1152 ^ n1139;
  assign n1245 = ~n1162 & ~n1244;
  assign n1246 = n1245 ^ n1161;
  assign n1258 = n1257 ^ n1246;
  assign n1239 = x13 & x14;
  assign n1238 = x12 & x15;
  assign n1240 = n1239 ^ n1238;
  assign n1237 = x5 & x22;
  assign n1241 = n1240 ^ n1237;
  assign n1234 = x6 & x21;
  assign n1233 = x4 & x23;
  assign n1235 = n1234 ^ n1233;
  assign n1232 = x3 & x24;
  assign n1236 = n1235 ^ n1232;
  assign n1242 = n1241 ^ n1236;
  assign n1228 = x14 & x25;
  assign n1229 = n327 & n1228;
  assign n1230 = x14 & ~n1229;
  assign n1226 = x0 & x27;
  assign n1225 = x1 & x26;
  assign n1227 = n1226 ^ n1225;
  assign n1231 = n1230 ^ n1227;
  assign n1243 = n1242 ^ n1231;
  assign n1259 = n1258 ^ n1243;
  assign n1218 = n1106 ^ n1103;
  assign n1219 = n1110 & ~n1218;
  assign n1220 = n1219 ^ n1109;
  assign n1215 = n1147 ^ n1144;
  assign n1216 = n1151 & ~n1215;
  assign n1217 = n1216 ^ n1150;
  assign n1221 = n1220 ^ n1217;
  assign n1212 = n1126 ^ n1121;
  assign n1213 = n1132 & ~n1212;
  assign n1214 = n1213 ^ n1131;
  assign n1222 = n1221 ^ n1214;
  assign n1207 = n1142 & n1143;
  assign n1208 = x18 & x26;
  assign n1209 = n155 & n1208;
  assign n1210 = ~n1207 & ~n1209;
  assign n1203 = x10 & x17;
  assign n1202 = x9 & x18;
  assign n1204 = n1203 ^ n1202;
  assign n1201 = x8 & x19;
  assign n1205 = n1204 ^ n1201;
  assign n1198 = x11 & x16;
  assign n1197 = x7 & x20;
  assign n1199 = n1198 ^ n1197;
  assign n1196 = x2 & x25;
  assign n1200 = n1199 ^ n1196;
  assign n1206 = n1205 ^ n1200;
  assign n1211 = n1210 ^ n1206;
  assign n1223 = n1222 ^ n1211;
  assign n1193 = n1111 ^ n1097;
  assign n1194 = n1112 & ~n1193;
  assign n1195 = n1194 ^ n1100;
  assign n1224 = n1223 ^ n1195;
  assign n1260 = n1259 ^ n1224;
  assign n1190 = n1163 ^ n1133;
  assign n1191 = ~n1164 & n1190;
  assign n1192 = n1191 ^ n1136;
  assign n1261 = n1260 ^ n1192;
  assign n1187 = n1165 ^ n1113;
  assign n1188 = n1166 & n1187;
  assign n1189 = n1188 ^ n1116;
  assign n1262 = n1261 ^ n1189;
  assign n1271 = n1270 ^ n1262;
  assign n1346 = x9 & x19;
  assign n1345 = x10 & x18;
  assign n1347 = n1346 ^ n1345;
  assign n1344 = x2 & x26;
  assign n1348 = n1347 ^ n1344;
  assign n1341 = x12 & x16;
  assign n1340 = x11 & x17;
  assign n1342 = n1341 ^ n1340;
  assign n1339 = x0 & x28;
  assign n1343 = n1342 ^ n1339;
  assign n1349 = n1348 ^ n1343;
  assign n1336 = n1252 ^ n1249;
  assign n1337 = n1256 & ~n1336;
  assign n1338 = n1337 ^ n1255;
  assign n1350 = n1349 ^ n1338;
  assign n1333 = n1217 ^ n1214;
  assign n1334 = n1221 & ~n1333;
  assign n1335 = n1334 ^ n1220;
  assign n1351 = n1350 ^ n1335;
  assign n1328 = n1233 ^ n1232;
  assign n1329 = n1235 & ~n1328;
  assign n1330 = n1329 ^ n1234;
  assign n1325 = n1197 ^ n1196;
  assign n1326 = n1199 & ~n1325;
  assign n1327 = n1326 ^ n1198;
  assign n1331 = n1330 ^ n1327;
  assign n1322 = n1202 ^ n1201;
  assign n1323 = n1204 & ~n1322;
  assign n1324 = n1323 ^ n1203;
  assign n1332 = n1331 ^ n1324;
  assign n1352 = n1351 ^ n1332;
  assign n1312 = n1259 ^ n1195;
  assign n1315 = n1259 ^ n1192;
  assign n1316 = n1312 & ~n1315;
  assign n1317 = n1316 ^ n1192;
  assign n1318 = n1317 ^ n1211;
  assign n1313 = n1195 ^ n1192;
  assign n1314 = n1312 & ~n1313;
  assign n1319 = n1318 ^ n1314;
  assign n1320 = n1223 & n1319;
  assign n1321 = n1320 ^ n1314;
  assign n1353 = n1352 ^ n1321;
  assign n1303 = x14 & x26;
  assign n1304 = n1303 ^ x27;
  assign n1305 = x1 & n1304;
  assign n1302 = x13 & x15;
  assign n1306 = n1305 ^ n1302;
  assign n1299 = n1238 ^ n1237;
  assign n1300 = n1240 & ~n1299;
  assign n1301 = n1300 ^ n1239;
  assign n1307 = n1306 ^ n1301;
  assign n1296 = n1210 ^ n1205;
  assign n1297 = ~n1206 & ~n1296;
  assign n1298 = n1297 ^ n1210;
  assign n1308 = n1307 ^ n1298;
  assign n1293 = n1236 ^ n1231;
  assign n1294 = n1242 & ~n1293;
  assign n1295 = n1294 ^ n1241;
  assign n1309 = n1308 ^ n1295;
  assign n1289 = n1226 & ~n1231;
  assign n1290 = ~x26 & n1229;
  assign n1291 = ~n1289 & ~n1290;
  assign n1285 = x8 & x20;
  assign n1284 = x4 & x24;
  assign n1286 = n1285 ^ n1284;
  assign n1283 = x3 & x25;
  assign n1287 = n1286 ^ n1283;
  assign n1280 = x7 & x21;
  assign n1279 = x6 & x22;
  assign n1281 = n1280 ^ n1279;
  assign n1278 = x5 & x23;
  assign n1282 = n1281 ^ n1278;
  assign n1288 = n1287 ^ n1282;
  assign n1292 = n1291 ^ n1288;
  assign n1310 = n1309 ^ n1292;
  assign n1275 = n1257 ^ n1243;
  assign n1276 = ~n1258 & ~n1275;
  assign n1277 = n1276 ^ n1246;
  assign n1311 = n1310 ^ n1277;
  assign n1354 = n1353 ^ n1311;
  assign n1272 = n1270 ^ n1189;
  assign n1273 = n1262 & ~n1272;
  assign n1274 = n1273 ^ n1270;
  assign n1355 = n1354 ^ n1274;
  assign n1441 = n1192 & n1353;
  assign n1442 = ~n1195 & n1259;
  assign n1443 = n1352 & ~n1442;
  assign n1444 = ~n1441 & ~n1443;
  assign n1445 = ~n1223 & ~n1444;
  assign n1446 = n1317 & n1353;
  assign n1447 = ~n1211 & n1222;
  assign n1448 = n1352 & n1447;
  assign n1449 = ~n1446 & ~n1448;
  assign n1450 = ~n1445 & n1449;
  assign n1430 = n1345 ^ n1344;
  assign n1431 = n1347 & ~n1430;
  assign n1432 = n1431 ^ n1346;
  assign n1427 = n1340 ^ n1339;
  assign n1428 = n1342 & ~n1427;
  assign n1429 = n1428 ^ n1341;
  assign n1433 = n1432 ^ n1429;
  assign n1423 = x1 & n1302;
  assign n1424 = n1423 ^ x2;
  assign n1425 = x27 & n1424;
  assign n1422 = x0 & x29;
  assign n1426 = n1425 ^ n1422;
  assign n1434 = n1433 ^ n1426;
  assign n1419 = n1291 ^ n1287;
  assign n1420 = ~n1288 & ~n1419;
  assign n1421 = n1420 ^ n1291;
  assign n1435 = n1434 ^ n1421;
  assign n1416 = n1348 ^ n1338;
  assign n1417 = ~n1349 & n1416;
  assign n1418 = n1417 ^ n1338;
  assign n1436 = n1435 ^ n1418;
  assign n1413 = n1350 ^ n1332;
  assign n1414 = n1351 & ~n1413;
  assign n1415 = n1414 ^ n1335;
  assign n1437 = n1436 ^ n1415;
  assign n1410 = n1307 ^ n1295;
  assign n1411 = ~n1308 & ~n1410;
  assign n1412 = n1411 ^ n1298;
  assign n1438 = n1437 ^ n1412;
  assign n1397 = n1302 ^ x27;
  assign n1398 = n1303 & n1397;
  assign n1399 = ~n1301 & ~n1398;
  assign n1400 = ~n1303 & ~n1397;
  assign n1401 = x1 & ~n1400;
  assign n1402 = ~n1399 & n1401;
  assign n1403 = ~x1 & n1302;
  assign n1404 = n1301 & n1403;
  assign n1405 = ~n1402 & ~n1404;
  assign n1394 = n1327 ^ n1324;
  assign n1395 = n1331 & ~n1394;
  assign n1396 = n1395 ^ n1330;
  assign n1406 = n1405 ^ n1396;
  assign n1391 = x14 & x15;
  assign n1390 = x13 & x16;
  assign n1392 = n1391 ^ n1390;
  assign n1389 = x6 & x23;
  assign n1393 = n1392 ^ n1389;
  assign n1407 = n1406 ^ n1393;
  assign n1384 = n1284 ^ n1283;
  assign n1385 = n1286 & ~n1384;
  assign n1386 = n1385 ^ n1285;
  assign n1381 = n1279 ^ n1278;
  assign n1382 = n1281 & ~n1381;
  assign n1383 = n1382 ^ n1280;
  assign n1387 = n1386 ^ n1383;
  assign n1379 = x1 & x28;
  assign n1380 = n1379 ^ x15;
  assign n1388 = n1387 ^ n1380;
  assign n1408 = n1407 ^ n1388;
  assign n1374 = x12 & x17;
  assign n1373 = x8 & x21;
  assign n1375 = n1374 ^ n1373;
  assign n1372 = x3 & x26;
  assign n1376 = n1375 ^ n1372;
  assign n1369 = x11 & x18;
  assign n1368 = x10 & x19;
  assign n1370 = n1369 ^ n1368;
  assign n1367 = x9 & x20;
  assign n1371 = n1370 ^ n1367;
  assign n1377 = n1376 ^ n1371;
  assign n1364 = x7 & x22;
  assign n1363 = x5 & x24;
  assign n1365 = n1364 ^ n1363;
  assign n1362 = x4 & x25;
  assign n1366 = n1365 ^ n1362;
  assign n1378 = n1377 ^ n1366;
  assign n1409 = n1408 ^ n1378;
  assign n1439 = n1438 ^ n1409;
  assign n1359 = n1309 ^ n1277;
  assign n1360 = ~n1310 & n1359;
  assign n1361 = n1360 ^ n1277;
  assign n1440 = n1439 ^ n1361;
  assign n1451 = n1450 ^ n1440;
  assign n1356 = n1353 ^ n1274;
  assign n1357 = ~n1354 & ~n1356;
  assign n1358 = n1357 ^ n1274;
  assign n1452 = n1451 ^ n1358;
  assign n1533 = n1450 ^ n1409;
  assign n1534 = n1409 ^ n1361;
  assign n1535 = n1533 & ~n1534;
  assign n1536 = n1535 ^ n1450;
  assign n1537 = ~n1438 & n1536;
  assign n1538 = n1361 & n1450;
  assign n1539 = n1409 & n1538;
  assign n1540 = ~n1537 & ~n1539;
  assign n1541 = ~n1358 & ~n1540;
  assign n1542 = ~n1361 & ~n1450;
  assign n1543 = ~n1409 & n1542;
  assign n1544 = ~n1539 & ~n1543;
  assign n1545 = n1439 & ~n1544;
  assign n1546 = ~n1541 & ~n1545;
  assign n1547 = ~n1438 & ~n1543;
  assign n1548 = ~n1536 & ~n1547;
  assign n1549 = n1358 & n1548;
  assign n1550 = n1546 & ~n1549;
  assign n1524 = x8 & x22;
  assign n1523 = x4 & x26;
  assign n1525 = n1524 ^ n1523;
  assign n1522 = x3 & x27;
  assign n1526 = n1525 ^ n1522;
  assign n1519 = x12 & x18;
  assign n1518 = x11 & x19;
  assign n1520 = n1519 ^ n1518;
  assign n1517 = x10 & x20;
  assign n1521 = n1520 ^ n1517;
  assign n1527 = n1526 ^ n1521;
  assign n1514 = x7 & x23;
  assign n1513 = x6 & x24;
  assign n1515 = n1514 ^ n1513;
  assign n1512 = x5 & x25;
  assign n1516 = n1515 ^ n1512;
  assign n1528 = n1527 ^ n1516;
  assign n1509 = n1396 ^ n1393;
  assign n1510 = ~n1406 & ~n1509;
  assign n1511 = n1510 ^ n1405;
  assign n1529 = n1528 ^ n1511;
  assign n1506 = n1421 ^ n1418;
  assign n1507 = n1435 & ~n1506;
  assign n1508 = n1507 ^ n1418;
  assign n1530 = n1529 ^ n1508;
  assign n1503 = n1436 ^ n1412;
  assign n1504 = ~n1437 & ~n1503;
  assign n1505 = n1504 ^ n1415;
  assign n1531 = n1530 ^ n1505;
  assign n1496 = x15 & n1379;
  assign n1495 = x0 & x30;
  assign n1497 = n1496 ^ n1495;
  assign n1493 = x1 & x29;
  assign n1492 = x14 & x16;
  assign n1494 = n1493 ^ n1492;
  assign n1498 = n1497 ^ n1494;
  assign n1489 = n1383 ^ n1380;
  assign n1490 = n1387 & ~n1489;
  assign n1491 = n1490 ^ n1386;
  assign n1499 = n1498 ^ n1491;
  assign n1486 = n1429 ^ n1426;
  assign n1487 = n1433 & ~n1486;
  assign n1488 = n1487 ^ n1432;
  assign n1500 = n1499 ^ n1488;
  assign n1483 = n1388 ^ n1378;
  assign n1484 = ~n1408 & ~n1483;
  assign n1485 = n1484 ^ n1407;
  assign n1501 = n1500 ^ n1485;
  assign n1476 = x13 & x17;
  assign n1475 = x9 & x21;
  assign n1477 = n1476 ^ n1475;
  assign n1474 = x2 & x28;
  assign n1478 = n1477 ^ n1474;
  assign n1471 = n1363 ^ n1362;
  assign n1472 = n1365 & ~n1471;
  assign n1473 = n1472 ^ n1364;
  assign n1479 = n1478 ^ n1473;
  assign n1468 = n1390 ^ n1389;
  assign n1469 = n1392 & ~n1468;
  assign n1470 = n1469 ^ n1391;
  assign n1480 = n1479 ^ n1470;
  assign n1463 = n1423 ^ n1422;
  assign n1464 = n1424 & ~n1463;
  assign n1465 = n1464 ^ x2;
  assign n1466 = x27 & n1465;
  assign n1459 = n1373 ^ n1372;
  assign n1460 = n1375 & ~n1459;
  assign n1461 = n1460 ^ n1374;
  assign n1456 = n1368 ^ n1367;
  assign n1457 = n1370 & ~n1456;
  assign n1458 = n1457 ^ n1369;
  assign n1462 = n1461 ^ n1458;
  assign n1467 = n1466 ^ n1462;
  assign n1481 = n1480 ^ n1467;
  assign n1453 = n1371 ^ n1366;
  assign n1454 = n1377 & ~n1453;
  assign n1455 = n1454 ^ n1376;
  assign n1482 = n1481 ^ n1455;
  assign n1502 = n1501 ^ n1482;
  assign n1532 = n1531 ^ n1502;
  assign n1551 = n1550 ^ n1532;
  assign n1639 = ~n1532 & n1544;
  assign n1640 = n1639 ^ n1539;
  assign n1641 = n1438 & ~n1640;
  assign n1642 = n1532 & ~n1536;
  assign n1643 = ~n1641 & ~n1642;
  assign n1644 = ~n1358 & n1643;
  assign n1645 = ~n1438 & n1640;
  assign n1646 = ~n1532 & n1536;
  assign n1647 = ~n1645 & ~n1646;
  assign n1648 = ~n1644 & n1647;
  assign n1629 = x12 & x19;
  assign n1628 = x13 & x18;
  assign n1630 = n1629 ^ n1628;
  assign n1631 = n1630 ^ n843;
  assign n1625 = x10 & x21;
  assign n1624 = x9 & x22;
  assign n1626 = n1625 ^ n1624;
  assign n1623 = x0 & x31;
  assign n1627 = n1626 ^ n1623;
  assign n1632 = n1631 ^ n1627;
  assign n1620 = n1495 ^ n1494;
  assign n1621 = n1497 & ~n1620;
  assign n1622 = n1621 ^ n1496;
  assign n1633 = n1632 ^ n1622;
  assign n1615 = x8 & x23;
  assign n1614 = x7 & x24;
  assign n1616 = n1615 ^ n1614;
  assign n1613 = x5 & x26;
  assign n1617 = n1616 ^ n1613;
  assign n1610 = x4 & x27;
  assign n1609 = x3 & x28;
  assign n1611 = n1610 ^ n1609;
  assign n1608 = x2 & x29;
  assign n1612 = n1611 ^ n1608;
  assign n1618 = n1617 ^ n1612;
  assign n1605 = x15 & x16;
  assign n1604 = x14 & x17;
  assign n1606 = n1605 ^ n1604;
  assign n1603 = x6 & x25;
  assign n1607 = n1606 ^ n1603;
  assign n1619 = n1618 ^ n1607;
  assign n1634 = n1633 ^ n1619;
  assign n1600 = n1467 ^ n1455;
  assign n1601 = n1481 & ~n1600;
  assign n1602 = n1601 ^ n1480;
  assign n1635 = n1634 ^ n1602;
  assign n1597 = n1500 ^ n1482;
  assign n1598 = ~n1501 & ~n1597;
  assign n1599 = n1598 ^ n1485;
  assign n1636 = n1635 ^ n1599;
  assign n1590 = n1498 ^ n1488;
  assign n1591 = n1499 & ~n1590;
  assign n1592 = n1591 ^ n1491;
  assign n1587 = n1521 ^ n1516;
  assign n1588 = n1527 & ~n1587;
  assign n1589 = n1588 ^ n1526;
  assign n1593 = n1592 ^ n1589;
  assign n1582 = n1523 ^ n1522;
  assign n1583 = n1525 & ~n1582;
  assign n1584 = n1583 ^ n1524;
  assign n1579 = n1475 ^ n1474;
  assign n1580 = n1477 & ~n1579;
  assign n1581 = n1580 ^ n1476;
  assign n1585 = n1584 ^ n1581;
  assign n1576 = n1518 ^ n1517;
  assign n1577 = n1520 & ~n1576;
  assign n1578 = n1577 ^ n1519;
  assign n1586 = n1585 ^ n1578;
  assign n1594 = n1593 ^ n1586;
  assign n1571 = x1 & x30;
  assign n1567 = x14 & x29;
  assign n1568 = x16 & n1567;
  assign n1569 = x1 & n1568;
  assign n1570 = n1569 ^ x16;
  assign n1572 = n1571 ^ n1570;
  assign n1564 = n1513 ^ n1512;
  assign n1565 = n1515 & ~n1564;
  assign n1566 = n1565 ^ n1514;
  assign n1573 = n1572 ^ n1566;
  assign n1561 = n1478 ^ n1470;
  assign n1562 = n1479 & ~n1561;
  assign n1563 = n1562 ^ n1473;
  assign n1574 = n1573 ^ n1563;
  assign n1558 = n1466 ^ n1461;
  assign n1559 = ~n1462 & n1558;
  assign n1560 = n1559 ^ n1466;
  assign n1575 = n1574 ^ n1560;
  assign n1595 = n1594 ^ n1575;
  assign n1555 = n1511 ^ n1508;
  assign n1556 = n1529 & ~n1555;
  assign n1557 = n1556 ^ n1508;
  assign n1596 = n1595 ^ n1557;
  assign n1637 = n1636 ^ n1596;
  assign n1552 = n1530 ^ n1502;
  assign n1553 = ~n1531 & ~n1552;
  assign n1554 = n1553 ^ n1505;
  assign n1638 = n1637 ^ n1554;
  assign n1649 = n1648 ^ n1638;
  assign n1739 = x0 & x32;
  assign n1737 = n515 ^ x2;
  assign n1738 = x30 & n1737;
  assign n1740 = n1739 ^ n1738;
  assign n1733 = x13 & x19;
  assign n1732 = x12 & x20;
  assign n1734 = n1733 ^ n1732;
  assign n1731 = x11 & x21;
  assign n1735 = n1734 ^ n1731;
  assign n1728 = x14 & x18;
  assign n1727 = x10 & x22;
  assign n1729 = n1728 ^ n1727;
  assign n1726 = x3 & x29;
  assign n1730 = n1729 ^ n1726;
  assign n1736 = n1735 ^ n1730;
  assign n1741 = n1740 ^ n1736;
  assign n1723 = n1589 ^ n1586;
  assign n1724 = n1593 & ~n1723;
  assign n1725 = n1724 ^ n1592;
  assign n1742 = n1741 ^ n1725;
  assign n1713 = x30 & n1566;
  assign n1714 = ~n1568 & ~n1713;
  assign n1715 = x16 & x30;
  assign n1716 = x1 & ~n1715;
  assign n1717 = ~n1714 & n1716;
  assign n1718 = ~n1567 & n1571;
  assign n1719 = x16 & ~n1718;
  assign n1720 = n1566 & n1719;
  assign n1721 = ~n1717 & ~n1720;
  assign n1709 = x9 & x23;
  assign n1708 = x5 & x27;
  assign n1710 = n1709 ^ n1708;
  assign n1707 = x4 & x28;
  assign n1711 = n1710 ^ n1707;
  assign n1704 = x8 & x24;
  assign n1703 = x7 & x25;
  assign n1705 = n1704 ^ n1703;
  assign n1702 = x6 & x26;
  assign n1706 = n1705 ^ n1702;
  assign n1712 = n1711 ^ n1706;
  assign n1722 = n1721 ^ n1712;
  assign n1743 = n1742 ^ n1722;
  assign n1693 = n1604 ^ n1603;
  assign n1694 = n1606 & ~n1693;
  assign n1695 = n1694 ^ n1605;
  assign n1690 = n1614 ^ n1613;
  assign n1691 = n1616 & ~n1690;
  assign n1692 = n1691 ^ n1615;
  assign n1696 = n1695 ^ n1692;
  assign n1688 = x1 & x31;
  assign n1687 = x15 & x17;
  assign n1689 = n1688 ^ n1687;
  assign n1697 = n1696 ^ n1689;
  assign n1684 = n1573 ^ n1560;
  assign n1685 = n1574 & ~n1684;
  assign n1686 = n1685 ^ n1563;
  assign n1698 = n1697 ^ n1686;
  assign n1679 = n1609 ^ n1608;
  assign n1680 = n1611 & ~n1679;
  assign n1681 = n1680 ^ n1610;
  assign n1676 = n1629 ^ n843;
  assign n1677 = ~n1630 & n1676;
  assign n1678 = n1677 ^ n843;
  assign n1682 = n1681 ^ n1678;
  assign n1673 = n1624 ^ n1623;
  assign n1674 = n1626 & ~n1673;
  assign n1675 = n1674 ^ n1625;
  assign n1683 = n1682 ^ n1675;
  assign n1699 = n1698 ^ n1683;
  assign n1668 = n1631 ^ n1622;
  assign n1669 = ~n1632 & n1668;
  assign n1670 = n1669 ^ n1622;
  assign n1665 = n1612 ^ n1607;
  assign n1666 = n1618 & ~n1665;
  assign n1667 = n1666 ^ n1617;
  assign n1671 = n1670 ^ n1667;
  assign n1662 = n1581 ^ n1578;
  assign n1663 = n1585 & ~n1662;
  assign n1664 = n1663 ^ n1584;
  assign n1672 = n1671 ^ n1664;
  assign n1700 = n1699 ^ n1672;
  assign n1659 = n1633 ^ n1602;
  assign n1660 = ~n1634 & n1659;
  assign n1661 = n1660 ^ n1602;
  assign n1701 = n1700 ^ n1661;
  assign n1744 = n1743 ^ n1701;
  assign n1656 = n1594 ^ n1557;
  assign n1657 = ~n1595 & n1656;
  assign n1658 = n1657 ^ n1557;
  assign n1745 = n1744 ^ n1658;
  assign n1653 = n1635 ^ n1596;
  assign n1654 = ~n1636 & ~n1653;
  assign n1655 = n1654 ^ n1599;
  assign n1746 = n1745 ^ n1655;
  assign n1650 = n1648 ^ n1554;
  assign n1651 = n1638 & n1650;
  assign n1652 = n1651 ^ n1648;
  assign n1747 = n1746 ^ n1652;
  assign n1834 = ~x2 & ~n515;
  assign n1835 = x30 & ~n1834;
  assign n1833 = n1738 & ~n1739;
  assign n1836 = n1835 ^ n1833;
  assign n1830 = n1732 ^ n1731;
  assign n1831 = n1734 & ~n1830;
  assign n1832 = n1831 ^ n1733;
  assign n1837 = n1836 ^ n1832;
  assign n1827 = n1727 ^ n1726;
  assign n1828 = n1729 & ~n1827;
  assign n1829 = n1828 ^ n1728;
  assign n1838 = n1837 ^ n1829;
  assign n1822 = x9 & x24;
  assign n1821 = x4 & x29;
  assign n1823 = n1822 ^ n1821;
  assign n1820 = x3 & x30;
  assign n1824 = n1823 ^ n1820;
  assign n1817 = x8 & x25;
  assign n1816 = x6 & x27;
  assign n1818 = n1817 ^ n1816;
  assign n1815 = x5 & x28;
  assign n1819 = n1818 ^ n1815;
  assign n1825 = n1824 ^ n1819;
  assign n1812 = x16 & x17;
  assign n1811 = x15 & x18;
  assign n1813 = n1812 ^ n1811;
  assign n1810 = x7 & x26;
  assign n1814 = n1813 ^ n1810;
  assign n1826 = n1825 ^ n1814;
  assign n1839 = n1838 ^ n1826;
  assign n1805 = x11 & x22;
  assign n1804 = x2 & x31;
  assign n1806 = n1805 ^ n1804;
  assign n1803 = x0 & x33;
  assign n1807 = n1806 ^ n1803;
  assign n1800 = n1703 ^ n1702;
  assign n1801 = n1705 & ~n1800;
  assign n1802 = n1801 ^ n1704;
  assign n1808 = n1807 ^ n1802;
  assign n1797 = n1708 ^ n1707;
  assign n1798 = n1710 & ~n1797;
  assign n1799 = n1798 ^ n1709;
  assign n1809 = n1808 ^ n1799;
  assign n1840 = n1839 ^ n1809;
  assign n1794 = n1741 ^ n1722;
  assign n1795 = n1742 & n1794;
  assign n1796 = n1795 ^ n1725;
  assign n1841 = n1840 ^ n1796;
  assign n1789 = n1721 ^ n1711;
  assign n1790 = ~n1712 & ~n1789;
  assign n1791 = n1790 ^ n1721;
  assign n1786 = n1740 ^ n1735;
  assign n1787 = ~n1736 & n1786;
  assign n1788 = n1787 ^ n1740;
  assign n1792 = n1791 ^ n1788;
  assign n1783 = n1678 ^ n1675;
  assign n1784 = n1682 & ~n1783;
  assign n1785 = n1784 ^ n1681;
  assign n1793 = n1792 ^ n1785;
  assign n1842 = n1841 ^ n1793;
  assign n1780 = n1672 ^ n1661;
  assign n1781 = n1700 & ~n1780;
  assign n1782 = n1781 ^ n1699;
  assign n1843 = n1842 ^ n1782;
  assign n1773 = x14 & x19;
  assign n1772 = x13 & x20;
  assign n1774 = n1773 ^ n1772;
  assign n1771 = x12 & x21;
  assign n1775 = n1774 ^ n1771;
  assign n1768 = n1692 ^ n1689;
  assign n1769 = n1696 & ~n1768;
  assign n1770 = n1769 ^ n1695;
  assign n1776 = n1775 ^ n1770;
  assign n1764 = x15 & x31;
  assign n1765 = x1 & n1764;
  assign n1766 = x17 & ~n1765;
  assign n1762 = x10 & x23;
  assign n1761 = x1 & x32;
  assign n1763 = n1762 ^ n1761;
  assign n1767 = n1766 ^ n1763;
  assign n1777 = n1776 ^ n1767;
  assign n1758 = n1667 ^ n1664;
  assign n1759 = n1671 & ~n1758;
  assign n1760 = n1759 ^ n1670;
  assign n1778 = n1777 ^ n1760;
  assign n1755 = n1697 ^ n1683;
  assign n1756 = n1698 & ~n1755;
  assign n1757 = n1756 ^ n1686;
  assign n1779 = n1778 ^ n1757;
  assign n1844 = n1843 ^ n1779;
  assign n1749 = n1701 ^ n1658;
  assign n1752 = n1744 & ~n1749;
  assign n1750 = n1749 ^ n1743;
  assign n1751 = n1655 & ~n1750;
  assign n1753 = n1752 ^ n1751;
  assign n1748 = n1652 & n1746;
  assign n1754 = n1753 ^ n1748;
  assign n1845 = n1844 ^ n1754;
  assign n1952 = ~n1744 & ~n1749;
  assign n1953 = n1952 ^ n1743;
  assign n1954 = n1701 & ~n1743;
  assign n1955 = n1658 & n1954;
  assign n1956 = n1655 & ~n1955;
  assign n1957 = ~n1953 & ~n1956;
  assign n1949 = ~n1655 & n1750;
  assign n1950 = n1949 ^ n1752;
  assign n1951 = ~n1844 & ~n1950;
  assign n1958 = n1957 ^ n1951;
  assign n1959 = n1652 & n1958;
  assign n1961 = ~n1753 & ~n1844;
  assign n1960 = ~n1655 & n1955;
  assign n1962 = n1961 ^ n1960;
  assign n1963 = ~n1959 & ~n1962;
  assign n1929 = x10 & x32;
  assign n1930 = x23 & n1929;
  assign n1931 = x17 & x31;
  assign n1932 = x15 & n1931;
  assign n1933 = ~n1930 & ~n1932;
  assign n1883 = x17 & x32;
  assign n1934 = x1 & ~n1883;
  assign n1935 = ~n1933 & n1934;
  assign n1936 = n1761 & ~n1764;
  assign n1937 = x17 & x23;
  assign n1938 = x10 & n1937;
  assign n1939 = ~n1936 & n1938;
  assign n1940 = ~n1935 & ~n1939;
  assign n1925 = x12 & x22;
  assign n1926 = n1925 ^ n1052;
  assign n1924 = x2 & x32;
  assign n1927 = n1926 ^ n1924;
  assign n1921 = n1772 ^ n1771;
  assign n1922 = n1774 & ~n1921;
  assign n1923 = n1922 ^ n1773;
  assign n1928 = n1927 ^ n1923;
  assign n1941 = n1940 ^ n1928;
  assign n1916 = x10 & x24;
  assign n1915 = x9 & x25;
  assign n1917 = n1916 ^ n1915;
  assign n1914 = x5 & x29;
  assign n1918 = n1917 ^ n1914;
  assign n1911 = x15 & x19;
  assign n1910 = x14 & x20;
  assign n1912 = n1911 ^ n1910;
  assign n1909 = x13 & x21;
  assign n1913 = n1912 ^ n1909;
  assign n1919 = n1918 ^ n1913;
  assign n1906 = x8 & x26;
  assign n1905 = x7 & x27;
  assign n1907 = n1906 ^ n1905;
  assign n1904 = x6 & x28;
  assign n1908 = n1907 ^ n1904;
  assign n1920 = n1919 ^ n1908;
  assign n1942 = n1941 ^ n1920;
  assign n1901 = n1775 ^ n1767;
  assign n1902 = n1776 & ~n1901;
  assign n1903 = n1902 ^ n1770;
  assign n1943 = n1942 ^ n1903;
  assign n1894 = n1804 ^ n1803;
  assign n1895 = n1806 & ~n1894;
  assign n1896 = n1895 ^ n1805;
  assign n1891 = n1816 ^ n1815;
  assign n1892 = n1818 & ~n1891;
  assign n1893 = n1892 ^ n1817;
  assign n1897 = n1896 ^ n1893;
  assign n1888 = n1821 ^ n1820;
  assign n1889 = n1823 & ~n1888;
  assign n1890 = n1889 ^ n1822;
  assign n1898 = n1897 ^ n1890;
  assign n1884 = n1883 ^ x33;
  assign n1885 = x1 & n1884;
  assign n1882 = x16 & x18;
  assign n1886 = n1885 ^ n1882;
  assign n1879 = n1811 ^ n1810;
  assign n1880 = n1813 & ~n1879;
  assign n1881 = n1880 ^ n1812;
  assign n1887 = n1886 ^ n1881;
  assign n1899 = n1898 ^ n1887;
  assign n1876 = n1819 ^ n1814;
  assign n1877 = n1825 & ~n1876;
  assign n1878 = n1877 ^ n1824;
  assign n1900 = n1899 ^ n1878;
  assign n1944 = n1943 ^ n1900;
  assign n1873 = n1760 ^ n1757;
  assign n1874 = ~n1778 & n1873;
  assign n1875 = n1874 ^ n1757;
  assign n1945 = n1944 ^ n1875;
  assign n1866 = x4 & x30;
  assign n1865 = x3 & x31;
  assign n1867 = n1866 ^ n1865;
  assign n1864 = x0 & x34;
  assign n1868 = n1867 ^ n1864;
  assign n1861 = n1832 ^ n1829;
  assign n1862 = n1837 & ~n1861;
  assign n1863 = n1862 ^ n1836;
  assign n1869 = n1868 ^ n1863;
  assign n1858 = n1807 ^ n1799;
  assign n1859 = n1808 & ~n1858;
  assign n1860 = n1859 ^ n1802;
  assign n1870 = n1869 ^ n1860;
  assign n1855 = n1826 ^ n1809;
  assign n1856 = n1839 & ~n1855;
  assign n1857 = n1856 ^ n1838;
  assign n1871 = n1870 ^ n1857;
  assign n1852 = n1788 ^ n1785;
  assign n1853 = ~n1792 & ~n1852;
  assign n1854 = n1853 ^ n1791;
  assign n1872 = n1871 ^ n1854;
  assign n1946 = n1945 ^ n1872;
  assign n1849 = n1840 ^ n1793;
  assign n1850 = n1841 & n1849;
  assign n1851 = n1850 ^ n1796;
  assign n1947 = n1946 ^ n1851;
  assign n1846 = n1782 ^ n1779;
  assign n1847 = ~n1843 & ~n1846;
  assign n1848 = n1847 ^ n1842;
  assign n1948 = n1947 ^ n1848;
  assign n1964 = n1963 ^ n1948;
  assign n2065 = n1872 & n1945;
  assign n2066 = ~n1851 & n2065;
  assign n2067 = ~n1848 & ~n2066;
  assign n2068 = n1945 ^ n1851;
  assign n2069 = ~n1946 & ~n2068;
  assign n2070 = n2069 ^ n1851;
  assign n2071 = ~n2067 & ~n2070;
  assign n2072 = n1963 & n2071;
  assign n2073 = n1848 & n2066;
  assign n2074 = ~n2072 & ~n2073;
  assign n2075 = ~n1872 & ~n1945;
  assign n2076 = n1851 & n2075;
  assign n2077 = n1848 & ~n2076;
  assign n2078 = n2070 & ~n2077;
  assign n2079 = ~n1963 & n2078;
  assign n2080 = ~n1848 & n2076;
  assign n2081 = ~n2079 & ~n2080;
  assign n2082 = n2074 & n2081;
  assign n2054 = x16 & n636;
  assign n2055 = n2054 ^ x2;
  assign n2056 = x33 & n2055;
  assign n2053 = x0 & x35;
  assign n2057 = n2056 ^ n2053;
  assign n2049 = x12 & x23;
  assign n2048 = x11 & x24;
  assign n2050 = n2049 ^ n2048;
  assign n2047 = x3 & x32;
  assign n2051 = n2050 ^ n2047;
  assign n2044 = x15 & x20;
  assign n2043 = x14 & x21;
  assign n2045 = n2044 ^ n2043;
  assign n2042 = x13 & x22;
  assign n2046 = n2045 ^ n2042;
  assign n2052 = n2051 ^ n2046;
  assign n2058 = n2057 ^ n2052;
  assign n2037 = x17 & x18;
  assign n2036 = x16 & x19;
  assign n2038 = n2037 ^ n2036;
  assign n2035 = x7 & x28;
  assign n2039 = n2038 ^ n2035;
  assign n2032 = x8 & x27;
  assign n2031 = x6 & x29;
  assign n2033 = n2032 ^ n2031;
  assign n2030 = x5 & x30;
  assign n2034 = n2033 ^ n2030;
  assign n2040 = n2039 ^ n2034;
  assign n2027 = x10 & x25;
  assign n2026 = x9 & x26;
  assign n2028 = n2027 ^ n2026;
  assign n2025 = x4 & x31;
  assign n2029 = n2028 ^ n2025;
  assign n2041 = n2040 ^ n2029;
  assign n2059 = n2058 ^ n2041;
  assign n2022 = n1868 ^ n1860;
  assign n2023 = n1869 & ~n2022;
  assign n2024 = n2023 ^ n1863;
  assign n2060 = n2059 ^ n2024;
  assign n2015 = n1905 ^ n1904;
  assign n2016 = n1907 & ~n2015;
  assign n2017 = n2016 ^ n1906;
  assign n2012 = n1915 ^ n1914;
  assign n2013 = n1917 & ~n2012;
  assign n2014 = n2013 ^ n1916;
  assign n2018 = n2017 ^ n2014;
  assign n2010 = x1 & x34;
  assign n2011 = n2010 ^ x18;
  assign n2019 = n2018 ^ n2011;
  assign n2007 = n1913 ^ n1908;
  assign n2008 = n1919 & ~n2007;
  assign n2009 = n2008 ^ n1918;
  assign n2020 = n2019 ^ n2009;
  assign n2002 = n1925 ^ n1924;
  assign n2003 = n1926 & ~n2002;
  assign n2004 = n2003 ^ n1052;
  assign n1999 = n1865 ^ n1864;
  assign n2000 = n1867 & ~n1999;
  assign n2001 = n2000 ^ n1866;
  assign n2005 = n2004 ^ n2001;
  assign n1996 = n1910 ^ n1909;
  assign n1997 = n1912 & ~n1996;
  assign n1998 = n1997 ^ n1911;
  assign n2006 = n2005 ^ n1998;
  assign n2021 = n2020 ^ n2006;
  assign n2061 = n2060 ^ n2021;
  assign n1993 = n1857 ^ n1854;
  assign n1994 = ~n1871 & ~n1993;
  assign n1995 = n1994 ^ n1854;
  assign n2062 = n2061 ^ n1995;
  assign n1980 = n1882 ^ x33;
  assign n1981 = n1883 & n1980;
  assign n1982 = ~n1881 & ~n1981;
  assign n1983 = ~n1883 & ~n1980;
  assign n1984 = x1 & ~n1983;
  assign n1985 = ~n1982 & n1984;
  assign n1986 = ~x1 & n1882;
  assign n1987 = n1881 & n1986;
  assign n1988 = ~n1985 & ~n1987;
  assign n1977 = n1893 ^ n1890;
  assign n1978 = n1897 & ~n1977;
  assign n1979 = n1978 ^ n1896;
  assign n1989 = n1988 ^ n1979;
  assign n1974 = n1940 ^ n1923;
  assign n1975 = ~n1928 & ~n1974;
  assign n1976 = n1975 ^ n1940;
  assign n1990 = n1989 ^ n1976;
  assign n1971 = n1887 ^ n1878;
  assign n1972 = n1899 & ~n1971;
  assign n1973 = n1972 ^ n1898;
  assign n1991 = n1990 ^ n1973;
  assign n1968 = n1941 ^ n1903;
  assign n1969 = n1942 & ~n1968;
  assign n1970 = n1969 ^ n1903;
  assign n1992 = n1991 ^ n1970;
  assign n2063 = n2062 ^ n1992;
  assign n1965 = n1943 ^ n1875;
  assign n1966 = n1944 & ~n1965;
  assign n1967 = n1966 ^ n1875;
  assign n2064 = n2063 ^ n1967;
  assign n2083 = n2082 ^ n2064;
  assign n2187 = ~n2064 & ~n2073;
  assign n2188 = ~n2078 & ~n2187;
  assign n2189 = ~n1963 & ~n2188;
  assign n2190 = ~n2064 & ~n2071;
  assign n2191 = ~n2080 & ~n2190;
  assign n2192 = ~n2189 & n2191;
  assign n2175 = x16 & x20;
  assign n2174 = x15 & x21;
  assign n2176 = n2175 ^ n2174;
  assign n2173 = x14 & x22;
  assign n2177 = n2176 ^ n2173;
  assign n2170 = x11 & x25;
  assign n2169 = x4 & x32;
  assign n2171 = n2170 ^ n2169;
  assign n2168 = x3 & x33;
  assign n2172 = n2171 ^ n2168;
  assign n2178 = n2177 ^ n2172;
  assign n2165 = x34 & n636;
  assign n2163 = x1 & x35;
  assign n2162 = x17 & x19;
  assign n2164 = n2163 ^ n2162;
  assign n2166 = n2165 ^ n2164;
  assign n2161 = x0 & x36;
  assign n2167 = n2166 ^ n2161;
  assign n2179 = n2178 ^ n2167;
  assign n2158 = n1979 ^ n1976;
  assign n2159 = ~n1989 & n2158;
  assign n2160 = n2159 ^ n1988;
  assign n2180 = n2179 ^ n2160;
  assign n2153 = x13 & x23;
  assign n2152 = x12 & x24;
  assign n2154 = n2153 ^ n2152;
  assign n2151 = x2 & x34;
  assign n2155 = n2154 ^ n2151;
  assign n2148 = x10 & x26;
  assign n2147 = x9 & x27;
  assign n2149 = n2148 ^ n2147;
  assign n2146 = x5 & x31;
  assign n2150 = n2149 ^ n2146;
  assign n2156 = n2155 ^ n2150;
  assign n2143 = x8 & x28;
  assign n2142 = x7 & x29;
  assign n2144 = n2143 ^ n2142;
  assign n2141 = x6 & x30;
  assign n2145 = n2144 ^ n2141;
  assign n2157 = n2156 ^ n2145;
  assign n2181 = n2180 ^ n2157;
  assign n2134 = ~x2 & ~n2054;
  assign n2135 = n2053 & ~n2134;
  assign n2136 = n545 & n636;
  assign n2137 = ~n2135 & ~n2136;
  assign n2138 = x33 & ~n2137;
  assign n2130 = n2048 ^ n2047;
  assign n2131 = n2050 & ~n2130;
  assign n2132 = n2131 ^ n2049;
  assign n2127 = n2043 ^ n2042;
  assign n2128 = n2045 & ~n2127;
  assign n2129 = n2128 ^ n2044;
  assign n2133 = n2132 ^ n2129;
  assign n2139 = n2138 ^ n2133;
  assign n2121 = n2031 ^ n2030;
  assign n2122 = n2033 & ~n2121;
  assign n2123 = n2122 ^ n2032;
  assign n2118 = n2026 ^ n2025;
  assign n2119 = n2028 & ~n2118;
  assign n2120 = n2119 ^ n2027;
  assign n2124 = n2123 ^ n2120;
  assign n2115 = n2036 ^ n2035;
  assign n2116 = n2038 & ~n2115;
  assign n2117 = n2116 ^ n2037;
  assign n2125 = n2124 ^ n2117;
  assign n2112 = n2034 ^ n2029;
  assign n2113 = n2040 & ~n2112;
  assign n2114 = n2113 ^ n2039;
  assign n2126 = n2125 ^ n2114;
  assign n2140 = n2139 ^ n2126;
  assign n2182 = n2181 ^ n2140;
  assign n2109 = n1973 ^ n1970;
  assign n2110 = ~n1991 & n2109;
  assign n2111 = n2110 ^ n1970;
  assign n2183 = n2182 ^ n2111;
  assign n2102 = n2014 ^ n2011;
  assign n2103 = n2018 & ~n2102;
  assign n2104 = n2103 ^ n2017;
  assign n2099 = n2001 ^ n1998;
  assign n2100 = n2005 & ~n2099;
  assign n2101 = n2100 ^ n2004;
  assign n2105 = n2104 ^ n2101;
  assign n2096 = n2057 ^ n2051;
  assign n2097 = ~n2052 & n2096;
  assign n2098 = n2097 ^ n2057;
  assign n2106 = n2105 ^ n2098;
  assign n2093 = n2019 ^ n2006;
  assign n2094 = n2020 & ~n2093;
  assign n2095 = n2094 ^ n2009;
  assign n2107 = n2106 ^ n2095;
  assign n2090 = n2058 ^ n2024;
  assign n2091 = ~n2059 & n2090;
  assign n2092 = n2091 ^ n2024;
  assign n2108 = n2107 ^ n2092;
  assign n2184 = n2183 ^ n2108;
  assign n2087 = n2060 ^ n1995;
  assign n2088 = ~n2061 & ~n2087;
  assign n2089 = n2088 ^ n1995;
  assign n2185 = n2184 ^ n2089;
  assign n2084 = n2062 ^ n1967;
  assign n2085 = n2063 & ~n2084;
  assign n2086 = n2085 ^ n1967;
  assign n2186 = n2185 ^ n2086;
  assign n2193 = n2192 ^ n2186;
  assign n2295 = n2183 ^ n2089;
  assign n2296 = n2184 & n2295;
  assign n2297 = n2296 ^ n2089;
  assign n2298 = ~n2086 & n2297;
  assign n2299 = ~n2108 & n2183;
  assign n2300 = n2089 & n2299;
  assign n2301 = ~n2298 & ~n2300;
  assign n2302 = n2192 & ~n2301;
  assign n2303 = n2108 & ~n2183;
  assign n2304 = ~n2089 & n2303;
  assign n2305 = n2086 & n2304;
  assign n2306 = ~n2302 & ~n2305;
  assign n2307 = ~n2086 & ~n2304;
  assign n2308 = ~n2297 & ~n2307;
  assign n2309 = ~n2192 & n2308;
  assign n2310 = ~n2086 & n2300;
  assign n2311 = ~n2309 & ~n2310;
  assign n2312 = n2306 & n2311;
  assign n2285 = x15 & x22;
  assign n2284 = x14 & x23;
  assign n2286 = n2285 ^ n2284;
  assign n2287 = n2286 ^ n1155;
  assign n2281 = n2147 ^ n2146;
  assign n2282 = n2149 & ~n2281;
  assign n2283 = n2282 ^ n2148;
  assign n2288 = n2287 ^ n2283;
  assign n2278 = n2164 ^ n2161;
  assign n2279 = n2166 & ~n2278;
  assign n2280 = n2279 ^ n2165;
  assign n2289 = n2288 ^ n2280;
  assign n2272 = n2169 ^ n2168;
  assign n2273 = n2171 & ~n2272;
  assign n2274 = n2273 ^ n2170;
  assign n2269 = n2174 ^ n2173;
  assign n2270 = n2176 & ~n2269;
  assign n2271 = n2270 ^ n2175;
  assign n2275 = n2274 ^ n2271;
  assign n2266 = n2152 ^ n2151;
  assign n2267 = n2154 & ~n2266;
  assign n2268 = n2267 ^ n2153;
  assign n2276 = n2275 ^ n2268;
  assign n2263 = n2172 ^ n2167;
  assign n2264 = n2178 & ~n2263;
  assign n2265 = n2264 ^ n2177;
  assign n2277 = n2276 ^ n2265;
  assign n2290 = n2289 ^ n2277;
  assign n2260 = n2095 ^ n2092;
  assign n2261 = ~n2107 & n2260;
  assign n2262 = n2261 ^ n2092;
  assign n2291 = n2290 ^ n2262;
  assign n2253 = x18 & x19;
  assign n2252 = x17 & x20;
  assign n2254 = n2253 ^ n2252;
  assign n2251 = x8 & x29;
  assign n2255 = n2254 ^ n2251;
  assign n2248 = x11 & x26;
  assign n2247 = x10 & x27;
  assign n2249 = n2248 ^ n2247;
  assign n2246 = x5 & x32;
  assign n2250 = n2249 ^ n2246;
  assign n2256 = n2255 ^ n2250;
  assign n2243 = n2138 ^ n2132;
  assign n2244 = ~n2133 & n2243;
  assign n2245 = n2244 ^ n2138;
  assign n2257 = n2256 ^ n2245;
  assign n2238 = x9 & x28;
  assign n2237 = x7 & x30;
  assign n2239 = n2238 ^ n2237;
  assign n2236 = x6 & x31;
  assign n2240 = n2239 ^ n2236;
  assign n2233 = x16 & x21;
  assign n2232 = x3 & x34;
  assign n2234 = n2233 ^ n2232;
  assign n2231 = x2 & x35;
  assign n2235 = n2234 ^ n2231;
  assign n2241 = n2240 ^ n2235;
  assign n2228 = x12 & x25;
  assign n2227 = x4 & x33;
  assign n2229 = n2228 ^ n2227;
  assign n2226 = x0 & x37;
  assign n2230 = n2229 ^ n2226;
  assign n2242 = n2241 ^ n2230;
  assign n2258 = n2257 ^ n2242;
  assign n2223 = n2101 ^ n2098;
  assign n2224 = n2105 & ~n2223;
  assign n2225 = n2224 ^ n2104;
  assign n2259 = n2258 ^ n2225;
  assign n2292 = n2291 ^ n2259;
  assign n2220 = n2181 ^ n2111;
  assign n2221 = n2182 & ~n2220;
  assign n2222 = n2221 ^ n2111;
  assign n2293 = n2292 ^ n2222;
  assign n2213 = x1 & x36;
  assign n2209 = x17 & x35;
  assign n2210 = x19 & n2209;
  assign n2211 = x1 & n2210;
  assign n2212 = n2211 ^ x19;
  assign n2214 = n2213 ^ n2212;
  assign n2206 = n2142 ^ n2141;
  assign n2207 = n2144 & ~n2206;
  assign n2208 = n2207 ^ n2143;
  assign n2215 = n2214 ^ n2208;
  assign n2203 = n2150 ^ n2145;
  assign n2204 = n2156 & ~n2203;
  assign n2205 = n2204 ^ n2155;
  assign n2216 = n2215 ^ n2205;
  assign n2200 = n2120 ^ n2117;
  assign n2201 = n2124 & ~n2200;
  assign n2202 = n2201 ^ n2123;
  assign n2217 = n2216 ^ n2202;
  assign n2197 = n2139 ^ n2114;
  assign n2198 = ~n2126 & n2197;
  assign n2199 = n2198 ^ n2139;
  assign n2218 = n2217 ^ n2199;
  assign n2194 = n2179 ^ n2157;
  assign n2195 = ~n2180 & ~n2194;
  assign n2196 = n2195 ^ n2160;
  assign n2219 = n2218 ^ n2196;
  assign n2294 = n2293 ^ n2219;
  assign n2313 = n2312 ^ n2294;
  assign n2426 = n2294 & ~n2305;
  assign n2427 = n2301 & ~n2426;
  assign n2428 = n2192 & ~n2427;
  assign n2429 = n2294 & ~n2308;
  assign n2430 = ~n2310 & ~n2429;
  assign n2431 = ~n2428 & n2430;
  assign n2414 = x17 & x21;
  assign n2413 = x16 & x22;
  assign n2415 = n2414 ^ n2413;
  assign n2412 = x15 & x23;
  assign n2416 = n2415 ^ n2412;
  assign n2409 = x10 & x28;
  assign n2408 = x6 & x32;
  assign n2410 = n2409 ^ n2408;
  assign n2407 = x5 & x33;
  assign n2411 = n2410 ^ n2407;
  assign n2417 = n2416 ^ n2411;
  assign n2404 = x9 & x29;
  assign n2403 = x8 & x30;
  assign n2405 = n2404 ^ n2403;
  assign n2402 = x7 & x31;
  assign n2406 = n2405 ^ n2402;
  assign n2418 = n2417 ^ n2406;
  assign n2399 = n2255 ^ n2245;
  assign n2400 = ~n2256 & n2399;
  assign n2401 = n2400 ^ n2245;
  assign n2419 = n2418 ^ n2401;
  assign n2394 = n2285 ^ n1155;
  assign n2395 = ~n2286 & n2394;
  assign n2396 = n2395 ^ n1155;
  assign n2391 = n2232 ^ n2231;
  assign n2392 = n2234 & ~n2391;
  assign n2393 = n2392 ^ n2233;
  assign n2397 = n2396 ^ n2393;
  assign n2388 = n2227 ^ n2226;
  assign n2389 = n2229 & ~n2388;
  assign n2390 = n2389 ^ n2228;
  assign n2398 = n2397 ^ n2390;
  assign n2420 = n2419 ^ n2398;
  assign n2385 = n2289 ^ n2265;
  assign n2386 = ~n2277 & n2385;
  assign n2387 = n2386 ^ n2289;
  assign n2421 = n2420 ^ n2387;
  assign n2382 = n2257 ^ n2225;
  assign n2383 = ~n2258 & n2382;
  assign n2384 = n2383 ^ n2225;
  assign n2422 = n2421 ^ n2384;
  assign n2379 = n2290 ^ n2259;
  assign n2380 = n2291 & ~n2379;
  assign n2381 = n2380 ^ n2262;
  assign n2423 = n2422 ^ n2381;
  assign n2365 = x36 & n2208;
  assign n2366 = ~n2210 & ~n2365;
  assign n2367 = x19 & x36;
  assign n2368 = x1 & ~n2367;
  assign n2369 = ~n2366 & n2368;
  assign n2370 = ~n2209 & n2213;
  assign n2371 = x19 & ~n2370;
  assign n2372 = n2208 & n2371;
  assign n2373 = ~n2369 & ~n2372;
  assign n2362 = x12 & x26;
  assign n2361 = x11 & x27;
  assign n2363 = n2362 ^ n2361;
  assign n2360 = x4 & x34;
  assign n2364 = n2363 ^ n2360;
  assign n2374 = n2373 ^ n2364;
  assign n2357 = n2271 ^ n2268;
  assign n2358 = n2275 & ~n2357;
  assign n2359 = n2358 ^ n2274;
  assign n2375 = n2374 ^ n2359;
  assign n2352 = x0 & x38;
  assign n2350 = n704 ^ x2;
  assign n2351 = x36 & n2350;
  assign n2353 = n2352 ^ n2351;
  assign n2347 = x14 & x24;
  assign n2346 = x13 & x25;
  assign n2348 = n2347 ^ n2346;
  assign n2345 = x3 & x35;
  assign n2349 = n2348 ^ n2345;
  assign n2354 = n2353 ^ n2349;
  assign n2342 = n2247 ^ n2246;
  assign n2343 = n2249 & ~n2342;
  assign n2344 = n2343 ^ n2248;
  assign n2355 = n2354 ^ n2344;
  assign n2339 = n2205 ^ n2202;
  assign n2340 = ~n2216 & n2339;
  assign n2341 = n2340 ^ n2202;
  assign n2356 = n2355 ^ n2341;
  assign n2376 = n2375 ^ n2356;
  assign n2332 = n2237 ^ n2236;
  assign n2333 = n2239 & ~n2332;
  assign n2334 = n2333 ^ n2238;
  assign n2329 = n2252 ^ n2251;
  assign n2330 = n2254 & ~n2329;
  assign n2331 = n2330 ^ n2253;
  assign n2335 = n2334 ^ n2331;
  assign n2327 = x1 & x37;
  assign n2326 = x18 & x20;
  assign n2328 = n2327 ^ n2326;
  assign n2336 = n2335 ^ n2328;
  assign n2323 = n2235 ^ n2230;
  assign n2324 = n2241 & ~n2323;
  assign n2325 = n2324 ^ n2240;
  assign n2337 = n2336 ^ n2325;
  assign n2320 = n2283 ^ n2280;
  assign n2321 = ~n2288 & n2320;
  assign n2322 = n2321 ^ n2280;
  assign n2338 = n2337 ^ n2322;
  assign n2377 = n2376 ^ n2338;
  assign n2317 = n2199 ^ n2196;
  assign n2318 = ~n2218 & ~n2317;
  assign n2319 = n2318 ^ n2196;
  assign n2378 = n2377 ^ n2319;
  assign n2424 = n2423 ^ n2378;
  assign n2314 = n2292 ^ n2219;
  assign n2315 = n2293 & n2314;
  assign n2316 = n2315 ^ n2222;
  assign n2425 = n2424 ^ n2316;
  assign n2432 = n2431 ^ n2425;
  assign n2540 = n2378 & n2422;
  assign n2541 = ~n2431 & ~n2540;
  assign n2542 = ~n2316 & ~n2381;
  assign n2543 = ~n2378 & ~n2422;
  assign n2544 = ~n2542 & ~n2543;
  assign n2545 = n2316 & n2381;
  assign n2546 = ~n2544 & ~n2545;
  assign n2547 = n2541 & n2546;
  assign n2548 = ~n2540 & ~n2545;
  assign n2549 = n2544 & ~n2548;
  assign n2550 = n2431 & n2549;
  assign n2551 = n2381 ^ n2316;
  assign n2552 = n2422 ^ n2378;
  assign n2553 = ~n2423 & ~n2552;
  assign n2554 = ~n2551 & n2553;
  assign n2555 = ~n2550 & ~n2554;
  assign n2556 = ~n2547 & n2555;
  assign n2529 = x19 & x20;
  assign n2528 = x18 & x21;
  assign n2530 = n2529 ^ n2528;
  assign n2527 = x8 & x31;
  assign n2531 = n2530 ^ n2527;
  assign n2524 = x17 & x22;
  assign n2523 = x12 & x27;
  assign n2525 = n2524 ^ n2523;
  assign n2522 = x4 & x35;
  assign n2526 = n2525 ^ n2522;
  assign n2532 = n2531 ^ n2526;
  assign n2519 = x11 & x28;
  assign n2518 = x10 & x29;
  assign n2520 = n2519 ^ n2518;
  assign n2517 = x5 & x34;
  assign n2521 = n2520 ^ n2517;
  assign n2533 = n2532 ^ n2521;
  assign n2514 = n2364 ^ n2359;
  assign n2515 = ~n2374 & ~n2514;
  assign n2516 = n2515 ^ n2373;
  assign n2534 = n2533 ^ n2516;
  assign n2509 = n2408 ^ n2407;
  assign n2510 = n2410 & ~n2509;
  assign n2511 = n2510 ^ n2409;
  assign n2506 = n2403 ^ n2402;
  assign n2507 = n2405 & ~n2506;
  assign n2508 = n2507 ^ n2404;
  assign n2512 = n2511 ^ n2508;
  assign n2503 = n2361 ^ n2360;
  assign n2504 = n2363 & ~n2503;
  assign n2505 = n2504 ^ n2362;
  assign n2513 = n2512 ^ n2505;
  assign n2535 = n2534 ^ n2513;
  assign n2500 = n2387 ^ n2384;
  assign n2501 = n2421 & ~n2500;
  assign n2502 = n2501 ^ n2420;
  assign n2536 = n2535 ^ n2502;
  assign n2493 = x13 & x26;
  assign n2492 = x3 & x36;
  assign n2494 = n2493 ^ n2492;
  assign n2491 = x2 & x37;
  assign n2495 = n2494 ^ n2491;
  assign n2488 = x16 & x23;
  assign n2487 = x15 & x24;
  assign n2489 = n2488 ^ n2487;
  assign n2490 = n2489 ^ n1228;
  assign n2496 = n2495 ^ n2490;
  assign n2484 = x9 & x30;
  assign n2483 = x7 & x32;
  assign n2485 = n2484 ^ n2483;
  assign n2482 = x6 & x33;
  assign n2486 = n2485 ^ n2482;
  assign n2497 = n2496 ^ n2486;
  assign n2479 = n2325 ^ n2322;
  assign n2480 = ~n2337 & n2479;
  assign n2481 = n2480 ^ n2322;
  assign n2498 = n2497 ^ n2481;
  assign n2476 = n2418 ^ n2398;
  assign n2477 = n2419 & ~n2476;
  assign n2478 = n2477 ^ n2401;
  assign n2499 = n2498 ^ n2478;
  assign n2537 = n2536 ^ n2499;
  assign n2473 = n2376 ^ n2319;
  assign n2474 = n2377 & n2473;
  assign n2475 = n2474 ^ n2319;
  assign n2538 = n2537 ^ n2475;
  assign n2464 = ~x2 & ~n704;
  assign n2465 = x36 & ~n2464;
  assign n2463 = n2351 & ~n2352;
  assign n2466 = n2465 ^ n2463;
  assign n2460 = n2413 ^ n2412;
  assign n2461 = n2415 & ~n2460;
  assign n2462 = n2461 ^ n2414;
  assign n2467 = n2466 ^ n2462;
  assign n2457 = n2346 ^ n2345;
  assign n2458 = n2348 & ~n2457;
  assign n2459 = n2458 ^ n2347;
  assign n2468 = n2467 ^ n2459;
  assign n2454 = n2349 ^ n2344;
  assign n2455 = n2354 & ~n2454;
  assign n2456 = n2455 ^ n2353;
  assign n2469 = n2468 ^ n2456;
  assign n2451 = n2411 ^ n2406;
  assign n2452 = n2417 & ~n2451;
  assign n2453 = n2452 ^ n2416;
  assign n2470 = n2469 ^ n2453;
  assign n2445 = x20 & x37;
  assign n2446 = n636 & n2445;
  assign n2447 = x20 & ~n2446;
  assign n2443 = x0 & x39;
  assign n2442 = x1 & x38;
  assign n2444 = n2443 ^ n2442;
  assign n2448 = n2447 ^ n2444;
  assign n2439 = n2331 ^ n2328;
  assign n2440 = n2335 & ~n2439;
  assign n2441 = n2440 ^ n2334;
  assign n2449 = n2448 ^ n2441;
  assign n2436 = n2393 ^ n2390;
  assign n2437 = n2397 & ~n2436;
  assign n2438 = n2437 ^ n2396;
  assign n2450 = n2449 ^ n2438;
  assign n2471 = n2470 ^ n2450;
  assign n2433 = n2375 ^ n2341;
  assign n2434 = ~n2356 & ~n2433;
  assign n2435 = n2434 ^ n2375;
  assign n2472 = n2471 ^ n2435;
  assign n2539 = n2538 ^ n2472;
  assign n2557 = n2556 ^ n2539;
  assign n2669 = n2539 & ~n2545;
  assign n2670 = ~n2543 & ~n2669;
  assign n2671 = ~n2541 & n2670;
  assign n2672 = n2539 & ~n2540;
  assign n2673 = ~n2542 & ~n2672;
  assign n2674 = n2431 & n2673;
  assign n2675 = ~n2539 & ~n2546;
  assign n2676 = ~n2674 & ~n2675;
  assign n2677 = ~n2671 & n2676;
  assign n2659 = n2490 ^ n2486;
  assign n2660 = n2496 & ~n2659;
  assign n2661 = n2660 ^ n2495;
  assign n2656 = n2526 ^ n2521;
  assign n2657 = n2532 & ~n2656;
  assign n2658 = n2657 ^ n2531;
  assign n2662 = n2661 ^ n2658;
  assign n2651 = n2492 ^ n2491;
  assign n2652 = n2494 & ~n2651;
  assign n2653 = n2652 ^ n2493;
  assign n2648 = n2518 ^ n2517;
  assign n2649 = n2520 & ~n2648;
  assign n2650 = n2649 ^ n2519;
  assign n2654 = n2653 ^ n2650;
  assign n2645 = n2523 ^ n2522;
  assign n2646 = n2525 & ~n2645;
  assign n2647 = n2646 ^ n2524;
  assign n2655 = n2654 ^ n2647;
  assign n2663 = n2662 ^ n2655;
  assign n2642 = n2533 ^ n2513;
  assign n2643 = ~n2534 & ~n2642;
  assign n2644 = n2643 ^ n2516;
  assign n2664 = n2663 ^ n2644;
  assign n2639 = n2481 ^ n2478;
  assign n2640 = ~n2498 & n2639;
  assign n2641 = n2640 ^ n2478;
  assign n2665 = n2664 ^ n2641;
  assign n2628 = x20 & x38;
  assign n2629 = n2628 ^ x39;
  assign n2630 = x1 & n2629;
  assign n2627 = x19 & x21;
  assign n2631 = n2630 ^ n2627;
  assign n2624 = n2528 ^ n2527;
  assign n2625 = n2530 & ~n2624;
  assign n2626 = n2625 ^ n2529;
  assign n2632 = n2631 ^ n2626;
  assign n2621 = n2508 ^ n2505;
  assign n2622 = n2512 & ~n2621;
  assign n2623 = n2622 ^ n2511;
  assign n2633 = n2632 ^ n2623;
  assign n2618 = n2462 ^ n2459;
  assign n2619 = n2467 & ~n2618;
  assign n2620 = n2619 ^ n2466;
  assign n2634 = n2633 ^ n2620;
  assign n2615 = n2468 ^ n2453;
  assign n2616 = n2469 & ~n2615;
  assign n2617 = n2616 ^ n2456;
  assign n2635 = n2634 ^ n2617;
  assign n2610 = x11 & x29;
  assign n2609 = x10 & x30;
  assign n2611 = n2610 ^ n2609;
  assign n2608 = x6 & x34;
  assign n2612 = n2611 ^ n2608;
  assign n2605 = x13 & x27;
  assign n2606 = n2605 ^ n1303;
  assign n2604 = x3 & x37;
  assign n2607 = n2606 ^ n2604;
  assign n2613 = n2612 ^ n2607;
  assign n2601 = x16 & x24;
  assign n2602 = n2601 ^ n1937;
  assign n2600 = x15 & x25;
  assign n2603 = n2602 ^ n2600;
  assign n2614 = n2613 ^ n2603;
  assign n2636 = n2635 ^ n2614;
  assign n2593 = x9 & x31;
  assign n2592 = x8 & x32;
  assign n2594 = n2593 ^ n2592;
  assign n2591 = x7 & x33;
  assign n2595 = n2594 ^ n2591;
  assign n2588 = x12 & x28;
  assign n2587 = x5 & x35;
  assign n2589 = n2588 ^ n2587;
  assign n2586 = x4 & x36;
  assign n2590 = n2589 ^ n2586;
  assign n2596 = n2595 ^ n2590;
  assign n2583 = x18 & x22;
  assign n2582 = x2 & x38;
  assign n2584 = n2583 ^ n2582;
  assign n2581 = x0 & x40;
  assign n2585 = n2584 ^ n2581;
  assign n2597 = n2596 ^ n2585;
  assign n2578 = n2448 ^ n2438;
  assign n2579 = n2449 & ~n2578;
  assign n2580 = n2579 ^ n2441;
  assign n2598 = n2597 ^ n2580;
  assign n2574 = n2443 & ~n2448;
  assign n2575 = ~x38 & n2446;
  assign n2576 = ~n2574 & ~n2575;
  assign n2570 = n2483 ^ n2482;
  assign n2571 = n2485 & ~n2570;
  assign n2572 = n2571 ^ n2484;
  assign n2567 = n2488 ^ n1228;
  assign n2568 = ~n2489 & n2567;
  assign n2569 = n2568 ^ n1228;
  assign n2573 = n2572 ^ n2569;
  assign n2577 = n2576 ^ n2573;
  assign n2599 = n2598 ^ n2577;
  assign n2637 = n2636 ^ n2599;
  assign n2564 = n2470 ^ n2435;
  assign n2565 = ~n2471 & ~n2564;
  assign n2566 = n2565 ^ n2435;
  assign n2638 = n2637 ^ n2566;
  assign n2666 = n2665 ^ n2638;
  assign n2561 = n2535 ^ n2499;
  assign n2562 = ~n2536 & n2561;
  assign n2563 = n2562 ^ n2502;
  assign n2667 = n2666 ^ n2563;
  assign n2558 = n2537 ^ n2472;
  assign n2559 = n2538 & ~n2558;
  assign n2560 = n2559 ^ n2475;
  assign n2668 = n2667 ^ n2560;
  assign n2678 = n2677 ^ n2668;
  assign n2797 = ~n2560 & ~n2677;
  assign n2798 = n2638 & ~n2665;
  assign n2799 = n2797 & n2798;
  assign n2800 = ~n2638 & n2665;
  assign n2801 = n2560 & n2800;
  assign n2802 = ~n2799 & ~n2801;
  assign n2803 = ~n2563 & ~n2802;
  assign n2804 = ~n2797 & ~n2798;
  assign n2805 = n2560 & n2677;
  assign n2806 = n2563 & ~n2800;
  assign n2807 = ~n2805 & n2806;
  assign n2808 = ~n2804 & n2807;
  assign n2809 = ~n2798 & ~n2806;
  assign n2810 = n2560 & n2809;
  assign n2811 = ~n2563 & n2800;
  assign n2812 = ~n2810 & ~n2811;
  assign n2813 = n2677 & ~n2812;
  assign n2814 = ~n2808 & ~n2813;
  assign n2815 = ~n2803 & n2814;
  assign n2786 = n2576 ^ n2572;
  assign n2787 = ~n2573 & ~n2786;
  assign n2788 = n2787 ^ n2576;
  assign n2783 = n2650 ^ n2647;
  assign n2784 = n2654 & ~n2783;
  assign n2785 = n2784 ^ n2653;
  assign n2789 = n2788 ^ n2785;
  assign n2780 = n2607 ^ n2603;
  assign n2781 = n2613 & ~n2780;
  assign n2782 = n2781 ^ n2612;
  assign n2790 = n2789 ^ n2782;
  assign n2777 = n2658 ^ n2655;
  assign n2778 = n2662 & ~n2777;
  assign n2779 = n2778 ^ n2661;
  assign n2791 = n2790 ^ n2779;
  assign n2772 = x15 & x26;
  assign n2771 = x13 & x28;
  assign n2773 = n2772 ^ n2771;
  assign n2770 = x3 & x38;
  assign n2774 = n2773 ^ n2770;
  assign n2767 = n2587 ^ n2586;
  assign n2768 = n2589 & ~n2767;
  assign n2769 = n2768 ^ n2588;
  assign n2775 = n2774 ^ n2769;
  assign n2763 = x1 & n2627;
  assign n2764 = n2763 ^ x2;
  assign n2765 = x39 & n2764;
  assign n2762 = x0 & x41;
  assign n2766 = n2765 ^ n2762;
  assign n2776 = n2775 ^ n2766;
  assign n2792 = n2791 ^ n2776;
  assign n2759 = n2644 ^ n2641;
  assign n2760 = n2664 & ~n2759;
  assign n2761 = n2760 ^ n2641;
  assign n2793 = n2792 ^ n2761;
  assign n2746 = n2627 ^ x39;
  assign n2747 = n2628 & n2746;
  assign n2748 = ~n2626 & ~n2747;
  assign n2749 = ~n2628 & ~n2746;
  assign n2750 = x1 & ~n2749;
  assign n2751 = ~n2748 & n2750;
  assign n2752 = ~x1 & n2627;
  assign n2753 = n2626 & n2752;
  assign n2754 = ~n2751 & ~n2753;
  assign n2743 = x11 & x30;
  assign n2742 = x6 & x35;
  assign n2744 = n2743 ^ n2742;
  assign n2741 = x5 & x36;
  assign n2745 = n2744 ^ n2741;
  assign n2755 = n2754 ^ n2745;
  assign n2738 = x20 & x21;
  assign n2737 = x19 & x22;
  assign n2739 = n2738 ^ n2737;
  assign n2736 = x8 & x33;
  assign n2740 = n2739 ^ n2736;
  assign n2756 = n2755 ^ n2740;
  assign n2731 = x18 & x23;
  assign n2730 = x17 & x24;
  assign n2732 = n2731 ^ n2730;
  assign n2729 = x16 & x25;
  assign n2733 = n2732 ^ n2729;
  assign n2726 = x10 & x31;
  assign n2725 = x9 & x32;
  assign n2727 = n2726 ^ n2725;
  assign n2724 = x7 & x34;
  assign n2728 = n2727 ^ n2724;
  assign n2734 = n2733 ^ n2728;
  assign n2721 = x14 & x27;
  assign n2720 = x12 & x29;
  assign n2722 = n2721 ^ n2720;
  assign n2719 = x4 & x37;
  assign n2723 = n2722 ^ n2719;
  assign n2735 = n2734 ^ n2723;
  assign n2757 = n2756 ^ n2735;
  assign n2716 = n2632 ^ n2620;
  assign n2717 = n2633 & ~n2716;
  assign n2718 = n2717 ^ n2623;
  assign n2758 = n2757 ^ n2718;
  assign n2794 = n2793 ^ n2758;
  assign n2713 = n2636 ^ n2566;
  assign n2714 = n2637 & ~n2713;
  assign n2715 = n2714 ^ n2566;
  assign n2795 = n2794 ^ n2715;
  assign n2704 = n2609 ^ n2608;
  assign n2705 = n2611 & ~n2704;
  assign n2706 = n2705 ^ n2610;
  assign n2701 = n2592 ^ n2591;
  assign n2702 = n2594 & ~n2701;
  assign n2703 = n2702 ^ n2593;
  assign n2707 = n2706 ^ n2703;
  assign n2699 = x1 & x40;
  assign n2700 = n2699 ^ x21;
  assign n2708 = n2707 ^ n2700;
  assign n2696 = n2590 ^ n2585;
  assign n2697 = n2596 & ~n2696;
  assign n2698 = n2697 ^ n2595;
  assign n2709 = n2708 ^ n2698;
  assign n2691 = n2582 ^ n2581;
  assign n2692 = n2584 & ~n2691;
  assign n2693 = n2692 ^ n2583;
  assign n2688 = n2605 ^ n2604;
  assign n2689 = n2606 & ~n2688;
  assign n2690 = n2689 ^ n1303;
  assign n2694 = n2693 ^ n2690;
  assign n2685 = n2601 ^ n2600;
  assign n2686 = n2602 & ~n2685;
  assign n2687 = n2686 ^ n1937;
  assign n2695 = n2694 ^ n2687;
  assign n2710 = n2709 ^ n2695;
  assign n2682 = n2597 ^ n2577;
  assign n2683 = n2598 & n2682;
  assign n2684 = n2683 ^ n2580;
  assign n2711 = n2710 ^ n2684;
  assign n2679 = n2634 ^ n2614;
  assign n2680 = n2635 & ~n2679;
  assign n2681 = n2680 ^ n2617;
  assign n2712 = n2711 ^ n2681;
  assign n2796 = n2795 ^ n2712;
  assign n2816 = n2815 ^ n2796;
  assign n2936 = n2665 ^ n2563;
  assign n2937 = n2796 ^ n2638;
  assign n2938 = n2666 & ~n2937;
  assign n2939 = n2936 & n2938;
  assign n2940 = n2939 ^ n2796;
  assign n2941 = ~n2797 & n2940;
  assign n2942 = ~n2796 & ~n2809;
  assign n2943 = n2805 & ~n2942;
  assign n2944 = ~n2941 & ~n2943;
  assign n2945 = n2796 & n2809;
  assign n2946 = n2944 & ~n2945;
  assign n2924 = x9 & x33;
  assign n2925 = n2924 ^ n1929;
  assign n2923 = x8 & x34;
  assign n2926 = n2925 ^ n2923;
  assign n2920 = n2725 ^ n2724;
  assign n2921 = n2727 & ~n2920;
  assign n2922 = n2921 ^ n2726;
  assign n2927 = n2926 ^ n2922;
  assign n2917 = x11 & x31;
  assign n2916 = x7 & x35;
  assign n2918 = n2917 ^ n2916;
  assign n2915 = x6 & x36;
  assign n2919 = n2918 ^ n2915;
  assign n2928 = n2927 ^ n2919;
  assign n2910 = x19 & x23;
  assign n2909 = x18 & x24;
  assign n2911 = n2910 ^ n2909;
  assign n2908 = x17 & x25;
  assign n2912 = n2911 ^ n2908;
  assign n2905 = x15 & x27;
  assign n2904 = x14 & x28;
  assign n2906 = n2905 ^ n2904;
  assign n2903 = x4 & x38;
  assign n2907 = n2906 ^ n2903;
  assign n2913 = n2912 ^ n2907;
  assign n2900 = x16 & x26;
  assign n2899 = x3 & x39;
  assign n2901 = n2900 ^ n2899;
  assign n2898 = x2 & x40;
  assign n2902 = n2901 ^ n2898;
  assign n2914 = n2913 ^ n2902;
  assign n2929 = n2928 ^ n2914;
  assign n2895 = n2785 ^ n2782;
  assign n2896 = ~n2789 & ~n2895;
  assign n2897 = n2896 ^ n2788;
  assign n2930 = n2929 ^ n2897;
  assign n2892 = n2684 ^ n2681;
  assign n2893 = ~n2711 & n2892;
  assign n2894 = n2893 ^ n2681;
  assign n2931 = n2930 ^ n2894;
  assign n2884 = n2720 ^ n2719;
  assign n2885 = n2722 & ~n2884;
  assign n2886 = n2885 ^ n2721;
  assign n2881 = n2742 ^ n2741;
  assign n2882 = n2744 & ~n2881;
  assign n2883 = n2882 ^ n2743;
  assign n2887 = n2886 ^ n2883;
  assign n2878 = n2737 ^ n2736;
  assign n2879 = n2739 & ~n2878;
  assign n2880 = n2879 ^ n2738;
  assign n2888 = n2887 ^ n2880;
  assign n2875 = n2745 ^ n2740;
  assign n2876 = ~n2755 & ~n2875;
  assign n2877 = n2876 ^ n2754;
  assign n2889 = n2888 ^ n2877;
  assign n2870 = n2763 ^ n2762;
  assign n2871 = n2764 & ~n2870;
  assign n2872 = n2871 ^ x2;
  assign n2873 = x39 & n2872;
  assign n2866 = n2771 ^ n2770;
  assign n2867 = n2773 & ~n2866;
  assign n2868 = n2867 ^ n2772;
  assign n2863 = n2730 ^ n2729;
  assign n2864 = n2732 & ~n2863;
  assign n2865 = n2864 ^ n2731;
  assign n2869 = n2868 ^ n2865;
  assign n2874 = n2873 ^ n2869;
  assign n2890 = n2889 ^ n2874;
  assign n2856 = x21 & x40;
  assign n2857 = n2856 ^ x41;
  assign n2858 = x1 & n2857;
  assign n2854 = x0 & x42;
  assign n2853 = x20 & x22;
  assign n2855 = n2854 ^ n2853;
  assign n2859 = n2858 ^ n2855;
  assign n2850 = x13 & x29;
  assign n2849 = x12 & x30;
  assign n2851 = n2850 ^ n2849;
  assign n2848 = x5 & x37;
  assign n2852 = n2851 ^ n2848;
  assign n2860 = n2859 ^ n2852;
  assign n2845 = n2703 ^ n2700;
  assign n2846 = n2707 & ~n2845;
  assign n2847 = n2846 ^ n2706;
  assign n2861 = n2860 ^ n2847;
  assign n2842 = n2708 ^ n2695;
  assign n2843 = n2709 & ~n2842;
  assign n2844 = n2843 ^ n2698;
  assign n2862 = n2861 ^ n2844;
  assign n2891 = n2890 ^ n2862;
  assign n2932 = n2931 ^ n2891;
  assign n2835 = n2690 ^ n2687;
  assign n2836 = n2694 & ~n2835;
  assign n2837 = n2836 ^ n2693;
  assign n2832 = n2728 ^ n2723;
  assign n2833 = n2734 & ~n2832;
  assign n2834 = n2833 ^ n2733;
  assign n2838 = n2837 ^ n2834;
  assign n2829 = n2774 ^ n2766;
  assign n2830 = n2775 & ~n2829;
  assign n2831 = n2830 ^ n2769;
  assign n2839 = n2838 ^ n2831;
  assign n2826 = n2756 ^ n2718;
  assign n2827 = n2757 & ~n2826;
  assign n2828 = n2827 ^ n2718;
  assign n2840 = n2839 ^ n2828;
  assign n2823 = n2779 ^ n2776;
  assign n2824 = ~n2791 & ~n2823;
  assign n2825 = n2824 ^ n2790;
  assign n2841 = n2840 ^ n2825;
  assign n2933 = n2932 ^ n2841;
  assign n2820 = n2792 ^ n2758;
  assign n2821 = ~n2793 & ~n2820;
  assign n2822 = n2821 ^ n2761;
  assign n2934 = n2933 ^ n2822;
  assign n2817 = n2715 ^ n2712;
  assign n2818 = ~n2795 & n2817;
  assign n2819 = n2818 ^ n2794;
  assign n2935 = n2934 ^ n2819;
  assign n2947 = n2946 ^ n2935;
  assign n3072 = ~n2819 & ~n2822;
  assign n3073 = n2841 & ~n2932;
  assign n3074 = ~n3072 & ~n3073;
  assign n3075 = n2819 & n2822;
  assign n3076 = ~n2841 & n2932;
  assign n3077 = ~n3075 & ~n3076;
  assign n3078 = ~n3074 & n3077;
  assign n3079 = ~n2946 & n3078;
  assign n3080 = n3075 & n3076;
  assign n3081 = ~n3079 & ~n3080;
  assign n3082 = n3074 & ~n3077;
  assign n3083 = n2946 & n3082;
  assign n3084 = n3072 & n3073;
  assign n3085 = ~n3083 & ~n3084;
  assign n3086 = n3081 & n3085;
  assign n3059 = n2916 ^ n2915;
  assign n3060 = n2918 & ~n3059;
  assign n3061 = n3060 ^ n2917;
  assign n3056 = n2909 ^ n2908;
  assign n3057 = n2911 & ~n3056;
  assign n3058 = n3057 ^ n2910;
  assign n3062 = n3061 ^ n3058;
  assign n3053 = n2904 ^ n2903;
  assign n3054 = n2906 & ~n3053;
  assign n3055 = n3054 ^ n2905;
  assign n3063 = n3062 ^ n3055;
  assign n3048 = n2899 ^ n2898;
  assign n3049 = n2901 & ~n3048;
  assign n3050 = n3049 ^ n2900;
  assign n3045 = n2849 ^ n2848;
  assign n3046 = n2851 & ~n3045;
  assign n3047 = n3046 ^ n2850;
  assign n3051 = n3050 ^ n3047;
  assign n3036 = ~n2854 & ~n2856;
  assign n3037 = n2853 ^ x41;
  assign n3038 = ~n3036 & n3037;
  assign n3039 = n2854 & n2856;
  assign n3040 = x1 & ~n3039;
  assign n3041 = ~n3038 & n3040;
  assign n3042 = n2853 & n2854;
  assign n3043 = ~x1 & ~n3042;
  assign n3044 = ~n3041 & ~n3043;
  assign n3052 = n3051 ^ n3044;
  assign n3064 = n3063 ^ n3052;
  assign n3033 = n2859 ^ n2847;
  assign n3034 = ~n2860 & n3033;
  assign n3035 = n3034 ^ n2847;
  assign n3065 = n3064 ^ n3035;
  assign n3028 = x12 & x31;
  assign n3027 = x11 & x32;
  assign n3029 = n3028 ^ n3027;
  assign n3026 = x6 & x37;
  assign n3030 = n3029 ^ n3026;
  assign n3023 = n2883 ^ n2880;
  assign n3024 = n2887 & ~n3023;
  assign n3025 = n3024 ^ n2886;
  assign n3031 = n3030 ^ n3025;
  assign n3020 = n2873 ^ n2868;
  assign n3021 = ~n2869 & n3020;
  assign n3022 = n3021 ^ n2873;
  assign n3032 = n3031 ^ n3022;
  assign n3066 = n3065 ^ n3032;
  assign n3017 = n2888 ^ n2874;
  assign n3018 = ~n2889 & ~n3017;
  assign n3019 = n3018 ^ n2877;
  assign n3067 = n3066 ^ n3019;
  assign n3010 = x21 & x22;
  assign n3009 = x20 & x23;
  assign n3011 = n3010 ^ n3009;
  assign n3008 = x9 & x34;
  assign n3012 = n3011 ^ n3008;
  assign n3005 = x13 & x30;
  assign n3004 = x5 & x38;
  assign n3006 = n3005 ^ n3004;
  assign n3003 = x2 & x41;
  assign n3007 = n3006 ^ n3003;
  assign n3013 = n3012 ^ n3007;
  assign n3000 = x10 & x33;
  assign n2999 = x8 & x35;
  assign n3001 = n3000 ^ n2999;
  assign n2998 = x7 & x36;
  assign n3002 = n3001 ^ n2998;
  assign n3014 = n3013 ^ n3002;
  assign n2995 = n2834 ^ n2831;
  assign n2996 = n2838 & ~n2995;
  assign n2997 = n2996 ^ n2837;
  assign n3015 = n3014 ^ n2997;
  assign n2990 = x15 & x28;
  assign n2989 = x16 & x27;
  assign n2991 = n2990 ^ n2989;
  assign n2992 = n2991 ^ n1567;
  assign n2986 = x19 & x24;
  assign n2985 = x18 & x25;
  assign n2987 = n2986 ^ n2985;
  assign n2984 = x17 & x26;
  assign n2988 = n2987 ^ n2984;
  assign n2993 = n2992 ^ n2988;
  assign n2981 = x4 & x39;
  assign n2980 = x3 & x40;
  assign n2982 = n2981 ^ n2980;
  assign n2979 = x0 & x43;
  assign n2983 = n2982 ^ n2979;
  assign n2994 = n2993 ^ n2983;
  assign n3016 = n3015 ^ n2994;
  assign n3068 = n3067 ^ n3016;
  assign n2976 = n2828 ^ n2825;
  assign n2977 = ~n2840 & ~n2976;
  assign n2978 = n2977 ^ n2825;
  assign n3069 = n3068 ^ n2978;
  assign n2969 = x1 & x42;
  assign n2966 = n2924 ^ n2923;
  assign n2967 = n2925 & ~n2966;
  assign n2968 = n2967 ^ n1929;
  assign n2970 = n2969 ^ n2968;
  assign n2963 = x20 & x41;
  assign n2964 = x1 & n2963;
  assign n2965 = x22 & ~n2964;
  assign n2971 = n2970 ^ n2965;
  assign n2960 = n2907 ^ n2902;
  assign n2961 = n2913 & ~n2960;
  assign n2962 = n2961 ^ n2912;
  assign n2972 = n2971 ^ n2962;
  assign n2957 = n2926 ^ n2919;
  assign n2958 = n2927 & ~n2957;
  assign n2959 = n2958 ^ n2922;
  assign n2973 = n2972 ^ n2959;
  assign n2954 = n2928 ^ n2897;
  assign n2955 = ~n2929 & ~n2954;
  assign n2956 = n2955 ^ n2897;
  assign n2974 = n2973 ^ n2956;
  assign n2951 = n2890 ^ n2844;
  assign n2952 = ~n2862 & ~n2951;
  assign n2953 = n2952 ^ n2890;
  assign n2975 = n2974 ^ n2953;
  assign n3070 = n3069 ^ n2975;
  assign n2948 = n2930 ^ n2891;
  assign n2949 = ~n2931 & ~n2948;
  assign n2950 = n2949 ^ n2894;
  assign n3071 = n3070 ^ n2950;
  assign n3087 = n3086 ^ n3071;
  assign n3216 = n3071 & ~n3072;
  assign n3217 = ~n3076 & ~n3216;
  assign n3218 = n3071 & ~n3073;
  assign n3219 = ~n3075 & ~n3218;
  assign n3220 = ~n3217 & ~n3219;
  assign n3221 = ~n2946 & ~n3220;
  assign n3222 = n3071 & ~n3084;
  assign n3223 = ~n3082 & ~n3222;
  assign n3224 = ~n3221 & ~n3223;
  assign n3200 = x22 & x42;
  assign n3201 = ~n2965 & ~n3200;
  assign n3202 = n2968 & n2969;
  assign n3203 = ~n2963 & n3202;
  assign n3204 = n3203 ^ n2968;
  assign n3205 = ~n3201 & ~n3204;
  assign n3206 = ~x22 & ~n3202;
  assign n3207 = ~n3205 & ~n3206;
  assign n3196 = n3047 ^ n3044;
  assign n3197 = n3051 & ~n3196;
  assign n3198 = n3197 ^ n3050;
  assign n3193 = n3058 ^ n3055;
  assign n3194 = n3062 & ~n3193;
  assign n3195 = n3194 ^ n3061;
  assign n3199 = n3198 ^ n3195;
  assign n3208 = n3207 ^ n3199;
  assign n3190 = n3063 ^ n3035;
  assign n3191 = ~n3064 & n3190;
  assign n3192 = n3191 ^ n3035;
  assign n3209 = n3208 ^ n3192;
  assign n3184 = x0 & x44;
  assign n3182 = n881 ^ x2;
  assign n3183 = x42 & n3182;
  assign n3185 = n3184 ^ n3183;
  assign n3179 = n2990 ^ n1567;
  assign n3180 = ~n2991 & n3179;
  assign n3181 = n3180 ^ n1567;
  assign n3186 = n3185 ^ n3181;
  assign n3176 = n3027 ^ n3026;
  assign n3177 = n3029 & ~n3176;
  assign n3178 = n3177 ^ n3028;
  assign n3187 = n3186 ^ n3178;
  assign n3171 = n3009 ^ n3008;
  assign n3172 = n3011 & ~n3171;
  assign n3173 = n3172 ^ n3010;
  assign n3168 = n2999 ^ n2998;
  assign n3169 = n3001 & ~n3168;
  assign n3170 = n3169 ^ n3000;
  assign n3174 = n3173 ^ n3170;
  assign n3166 = x1 & x43;
  assign n3165 = x21 & x23;
  assign n3167 = n3166 ^ n3165;
  assign n3175 = n3174 ^ n3167;
  assign n3188 = n3187 ^ n3175;
  assign n3162 = n3025 ^ n3022;
  assign n3163 = ~n3031 & n3162;
  assign n3164 = n3163 ^ n3022;
  assign n3189 = n3188 ^ n3164;
  assign n3210 = n3209 ^ n3189;
  assign n3155 = x11 & x33;
  assign n3154 = x7 & x37;
  assign n3156 = n3155 ^ n3154;
  assign n3153 = x6 & x38;
  assign n3157 = n3156 ^ n3153;
  assign n3150 = x17 & x27;
  assign n3149 = x15 & x29;
  assign n3151 = n3150 ^ n3149;
  assign n3148 = x3 & x41;
  assign n3152 = n3151 ^ n3148;
  assign n3158 = n3157 ^ n3152;
  assign n3145 = x20 & x24;
  assign n3144 = x19 & x25;
  assign n3146 = n3145 ^ n3144;
  assign n3147 = n3146 ^ n1208;
  assign n3159 = n3158 ^ n3147;
  assign n3141 = n2971 ^ n2959;
  assign n3142 = n2972 & ~n3141;
  assign n3143 = n3142 ^ n2962;
  assign n3160 = n3159 ^ n3143;
  assign n3136 = x10 & x34;
  assign n3135 = x9 & x35;
  assign n3137 = n3136 ^ n3135;
  assign n3134 = x8 & x36;
  assign n3138 = n3137 ^ n3134;
  assign n3131 = x16 & x28;
  assign n3130 = x14 & x30;
  assign n3132 = n3131 ^ n3130;
  assign n3129 = x4 & x40;
  assign n3133 = n3132 ^ n3129;
  assign n3139 = n3138 ^ n3133;
  assign n3126 = x13 & x31;
  assign n3125 = x12 & x32;
  assign n3127 = n3126 ^ n3125;
  assign n3124 = x5 & x39;
  assign n3128 = n3127 ^ n3124;
  assign n3140 = n3139 ^ n3128;
  assign n3161 = n3160 ^ n3140;
  assign n3211 = n3210 ^ n3161;
  assign n3121 = n2956 ^ n2953;
  assign n3122 = n2974 & n3121;
  assign n3123 = n3122 ^ n2953;
  assign n3212 = n3211 ^ n3123;
  assign n3114 = n3007 ^ n3002;
  assign n3115 = n3013 & ~n3114;
  assign n3116 = n3115 ^ n3012;
  assign n3111 = n2988 ^ n2983;
  assign n3112 = n2993 & ~n3111;
  assign n3113 = n3112 ^ n2992;
  assign n3117 = n3116 ^ n3113;
  assign n3106 = n2985 ^ n2984;
  assign n3107 = n2987 & ~n3106;
  assign n3108 = n3107 ^ n2986;
  assign n3103 = n2980 ^ n2979;
  assign n3104 = n2982 & ~n3103;
  assign n3105 = n3104 ^ n2981;
  assign n3109 = n3108 ^ n3105;
  assign n3100 = n3004 ^ n3003;
  assign n3101 = n3006 & ~n3100;
  assign n3102 = n3101 ^ n3005;
  assign n3110 = n3109 ^ n3102;
  assign n3118 = n3117 ^ n3110;
  assign n3097 = n3014 ^ n2994;
  assign n3098 = n3015 & ~n3097;
  assign n3099 = n3098 ^ n2997;
  assign n3119 = n3118 ^ n3099;
  assign n3094 = n3065 ^ n3019;
  assign n3095 = ~n3066 & ~n3094;
  assign n3096 = n3095 ^ n3019;
  assign n3120 = n3119 ^ n3096;
  assign n3213 = n3212 ^ n3120;
  assign n3091 = n3067 ^ n2978;
  assign n3092 = n3068 & n3091;
  assign n3093 = n3092 ^ n2978;
  assign n3214 = n3213 ^ n3093;
  assign n3088 = n3069 ^ n2950;
  assign n3089 = ~n3070 & n3088;
  assign n3090 = n3089 ^ n2950;
  assign n3215 = n3214 ^ n3090;
  assign n3225 = n3224 ^ n3215;
  assign n3353 = n3120 ^ n3093;
  assign n3354 = n3213 & ~n3353;
  assign n3355 = n3354 ^ n3212;
  assign n3356 = ~n3090 & n3355;
  assign n3357 = n3093 & n3120;
  assign n3358 = n3212 & n3357;
  assign n3359 = ~n3356 & ~n3358;
  assign n3360 = ~n3224 & ~n3359;
  assign n3361 = ~n3093 & ~n3120;
  assign n3362 = ~n3212 & n3361;
  assign n3363 = n3090 & n3362;
  assign n3364 = ~n3360 & ~n3363;
  assign n3365 = ~n3090 & ~n3362;
  assign n3366 = ~n3355 & ~n3365;
  assign n3367 = n3224 & n3366;
  assign n3368 = ~n3090 & n3358;
  assign n3369 = ~n3367 & ~n3368;
  assign n3370 = n3364 & n3369;
  assign n3342 = n3181 ^ n3178;
  assign n3343 = n3186 & ~n3342;
  assign n3344 = n3343 ^ n3185;
  assign n3339 = n3170 ^ n3167;
  assign n3340 = n3174 & ~n3339;
  assign n3341 = n3340 ^ n3173;
  assign n3345 = n3344 ^ n3341;
  assign n3336 = n3105 ^ n3102;
  assign n3337 = n3109 & ~n3336;
  assign n3338 = n3337 ^ n3108;
  assign n3346 = n3345 ^ n3338;
  assign n3331 = n3152 ^ n3147;
  assign n3332 = n3158 & ~n3331;
  assign n3333 = n3332 ^ n3157;
  assign n3328 = n3133 ^ n3128;
  assign n3329 = n3139 & ~n3328;
  assign n3330 = n3329 ^ n3138;
  assign n3334 = n3333 ^ n3330;
  assign n3323 = n3125 ^ n3124;
  assign n3324 = n3127 & ~n3323;
  assign n3325 = n3324 ^ n3126;
  assign n3320 = n3130 ^ n3129;
  assign n3321 = n3132 & ~n3320;
  assign n3322 = n3321 ^ n3131;
  assign n3326 = n3325 ^ n3322;
  assign n3317 = n3154 ^ n3153;
  assign n3318 = n3156 & ~n3317;
  assign n3319 = n3318 ^ n3155;
  assign n3327 = n3326 ^ n3319;
  assign n3335 = n3334 ^ n3327;
  assign n3347 = n3346 ^ n3335;
  assign n3314 = n3187 ^ n3164;
  assign n3315 = ~n3188 & n3314;
  assign n3316 = n3315 ^ n3164;
  assign n3348 = n3347 ^ n3316;
  assign n3307 = x22 & x23;
  assign n3306 = x21 & x24;
  assign n3308 = n3307 ^ n3306;
  assign n3305 = x10 & x35;
  assign n3309 = n3308 ^ n3305;
  assign n3302 = x9 & x36;
  assign n3301 = x8 & x37;
  assign n3303 = n3302 ^ n3301;
  assign n3300 = x7 & x38;
  assign n3304 = n3303 ^ n3300;
  assign n3310 = n3309 ^ n3304;
  assign n3297 = x4 & x41;
  assign n3296 = x2 & x43;
  assign n3298 = n3297 ^ n3296;
  assign n3295 = x0 & x45;
  assign n3299 = n3298 ^ n3295;
  assign n3311 = n3310 ^ n3299;
  assign n3292 = n3113 ^ n3110;
  assign n3293 = n3117 & ~n3292;
  assign n3294 = n3293 ^ n3116;
  assign n3312 = n3311 ^ n3294;
  assign n3287 = x20 & x25;
  assign n3286 = x19 & x26;
  assign n3288 = n3287 ^ n3286;
  assign n3285 = x18 & x27;
  assign n3289 = n3288 ^ n3285;
  assign n3282 = n3135 ^ n3134;
  assign n3283 = n3137 & ~n3282;
  assign n3284 = n3283 ^ n3136;
  assign n3290 = n3289 ^ n3284;
  assign n3279 = x14 & x31;
  assign n3278 = x13 & x32;
  assign n3280 = n3279 ^ n3278;
  assign n3277 = x5 & x40;
  assign n3281 = n3280 ^ n3277;
  assign n3291 = n3290 ^ n3281;
  assign n3313 = n3312 ^ n3291;
  assign n3349 = n3348 ^ n3313;
  assign n3274 = n3099 ^ n3096;
  assign n3275 = ~n3119 & ~n3274;
  assign n3276 = n3275 ^ n3096;
  assign n3350 = n3349 ^ n3276;
  assign n3265 = ~x2 & ~n881;
  assign n3266 = x42 & ~n3265;
  assign n3264 = n3183 & ~n3184;
  assign n3267 = n3266 ^ n3264;
  assign n3261 = n3145 ^ n1208;
  assign n3262 = ~n3146 & n3261;
  assign n3263 = n3262 ^ n1208;
  assign n3268 = n3267 ^ n3263;
  assign n3258 = n3149 ^ n3148;
  assign n3259 = n3151 & ~n3258;
  assign n3260 = n3259 ^ n3150;
  assign n3269 = n3268 ^ n3260;
  assign n3253 = x12 & x33;
  assign n3252 = x11 & x34;
  assign n3254 = n3253 ^ n3252;
  assign n3251 = x6 & x39;
  assign n3255 = n3254 ^ n3251;
  assign n3248 = x16 & x29;
  assign n3247 = x17 & x28;
  assign n3249 = n3248 ^ n3247;
  assign n3246 = x15 & x30;
  assign n3250 = n3249 ^ n3246;
  assign n3256 = n3255 ^ n3250;
  assign n3243 = x3 & x42;
  assign n3242 = x1 & x44;
  assign n3244 = n3243 ^ n3242;
  assign n3238 = x21 & x43;
  assign n3239 = x23 & n3238;
  assign n3240 = x1 & n3239;
  assign n3241 = n3240 ^ x23;
  assign n3245 = n3244 ^ n3241;
  assign n3257 = n3256 ^ n3245;
  assign n3270 = n3269 ^ n3257;
  assign n3235 = n3207 ^ n3198;
  assign n3236 = ~n3199 & n3235;
  assign n3237 = n3236 ^ n3207;
  assign n3271 = n3270 ^ n3237;
  assign n3232 = n3159 ^ n3140;
  assign n3233 = n3160 & ~n3232;
  assign n3234 = n3233 ^ n3143;
  assign n3272 = n3271 ^ n3234;
  assign n3229 = n3208 ^ n3189;
  assign n3230 = n3209 & ~n3229;
  assign n3231 = n3230 ^ n3192;
  assign n3273 = n3272 ^ n3231;
  assign n3351 = n3350 ^ n3273;
  assign n3226 = n3210 ^ n3123;
  assign n3227 = ~n3211 & ~n3226;
  assign n3228 = n3227 ^ n3123;
  assign n3352 = n3351 ^ n3228;
  assign n3371 = n3370 ^ n3352;
  assign n3508 = ~n3352 & ~n3363;
  assign n3509 = n3359 & ~n3508;
  assign n3510 = ~n3224 & ~n3509;
  assign n3511 = ~n3352 & ~n3366;
  assign n3512 = ~n3368 & ~n3511;
  assign n3513 = ~n3510 & n3512;
  assign n3496 = n3289 ^ n3281;
  assign n3497 = n3290 & ~n3496;
  assign n3498 = n3497 ^ n3284;
  assign n3493 = n3304 ^ n3299;
  assign n3494 = n3310 & ~n3493;
  assign n3495 = n3494 ^ n3309;
  assign n3499 = n3498 ^ n3495;
  assign n3490 = n3250 ^ n3245;
  assign n3491 = n3256 & ~n3490;
  assign n3492 = n3491 ^ n3255;
  assign n3500 = n3499 ^ n3492;
  assign n3483 = n3296 ^ n3295;
  assign n3484 = n3298 & ~n3483;
  assign n3485 = n3484 ^ n3297;
  assign n3480 = n3301 ^ n3300;
  assign n3481 = n3303 & ~n3480;
  assign n3482 = n3481 ^ n3302;
  assign n3486 = n3485 ^ n3482;
  assign n3477 = n3278 ^ n3277;
  assign n3478 = n3280 & ~n3477;
  assign n3479 = n3478 ^ n3279;
  assign n3487 = n3486 ^ n3479;
  assign n3432 = x23 & x44;
  assign n3473 = n3432 ^ x45;
  assign n3474 = x1 & n3473;
  assign n3472 = x22 & x24;
  assign n3475 = n3474 ^ n3472;
  assign n3469 = n3306 ^ n3305;
  assign n3470 = n3308 & ~n3469;
  assign n3471 = n3470 ^ n3307;
  assign n3476 = n3475 ^ n3471;
  assign n3488 = n3487 ^ n3476;
  assign n3466 = n3263 ^ n3260;
  assign n3467 = n3268 & ~n3466;
  assign n3468 = n3467 ^ n3267;
  assign n3489 = n3488 ^ n3468;
  assign n3501 = n3500 ^ n3489;
  assign n3463 = n3269 ^ n3237;
  assign n3464 = ~n3270 & n3463;
  assign n3465 = n3464 ^ n3237;
  assign n3502 = n3501 ^ n3465;
  assign n3456 = x4 & x42;
  assign n3455 = x3 & x43;
  assign n3457 = n3456 ^ n3455;
  assign n3454 = x0 & x46;
  assign n3458 = n3457 ^ n3454;
  assign n3451 = x11 & x35;
  assign n3450 = x10 & x36;
  assign n3452 = n3451 ^ n3450;
  assign n3449 = x9 & x37;
  assign n3453 = n3452 ^ n3449;
  assign n3459 = n3458 ^ n3453;
  assign n3446 = x21 & x25;
  assign n3445 = x20 & x26;
  assign n3447 = n3446 ^ n3445;
  assign n3444 = x19 & x27;
  assign n3448 = n3447 ^ n3444;
  assign n3460 = n3459 ^ n3448;
  assign n3441 = n3330 ^ n3327;
  assign n3442 = n3334 & ~n3441;
  assign n3443 = n3442 ^ n3333;
  assign n3461 = n3460 ^ n3443;
  assign n3429 = x3 & x44;
  assign n3430 = x42 & n3429;
  assign n3431 = ~n3239 & ~n3430;
  assign n3433 = x1 & ~n3432;
  assign n3434 = ~n3431 & n3433;
  assign n3435 = ~n3238 & n3242;
  assign n3436 = x23 & x42;
  assign n3437 = x3 & n3436;
  assign n3438 = ~n3435 & n3437;
  assign n3439 = ~n3434 & ~n3438;
  assign n3425 = x18 & x28;
  assign n3424 = x17 & x29;
  assign n3426 = n3425 ^ n3424;
  assign n3427 = n3426 ^ n1715;
  assign n3421 = x12 & x34;
  assign n3420 = x8 & x38;
  assign n3422 = n3421 ^ n3420;
  assign n3419 = x7 & x39;
  assign n3423 = n3422 ^ n3419;
  assign n3428 = n3427 ^ n3423;
  assign n3440 = n3439 ^ n3428;
  assign n3462 = n3461 ^ n3440;
  assign n3503 = n3502 ^ n3462;
  assign n3416 = n3234 ^ n3231;
  assign n3417 = ~n3272 & n3416;
  assign n3418 = n3417 ^ n3231;
  assign n3504 = n3503 ^ n3418;
  assign n3407 = x14 & x32;
  assign n3406 = x13 & x33;
  assign n3408 = n3407 ^ n3406;
  assign n3405 = x6 & x40;
  assign n3409 = n3408 ^ n3405;
  assign n3402 = x5 & x41;
  assign n3403 = n3402 ^ n1764;
  assign n3401 = x2 & x44;
  assign n3404 = n3403 ^ n3401;
  assign n3410 = n3409 ^ n3404;
  assign n3398 = n3322 ^ n3319;
  assign n3399 = n3326 & ~n3398;
  assign n3400 = n3399 ^ n3325;
  assign n3411 = n3410 ^ n3400;
  assign n3393 = n3252 ^ n3251;
  assign n3394 = n3254 & ~n3393;
  assign n3395 = n3394 ^ n3253;
  assign n3390 = n3247 ^ n3246;
  assign n3391 = n3249 & ~n3390;
  assign n3392 = n3391 ^ n3248;
  assign n3396 = n3395 ^ n3392;
  assign n3387 = n3286 ^ n3285;
  assign n3388 = n3288 & ~n3387;
  assign n3389 = n3388 ^ n3287;
  assign n3397 = n3396 ^ n3389;
  assign n3412 = n3411 ^ n3397;
  assign n3384 = n3341 ^ n3338;
  assign n3385 = n3345 & ~n3384;
  assign n3386 = n3385 ^ n3344;
  assign n3413 = n3412 ^ n3386;
  assign n3381 = n3311 ^ n3291;
  assign n3382 = n3312 & ~n3381;
  assign n3383 = n3382 ^ n3294;
  assign n3414 = n3413 ^ n3383;
  assign n3378 = n3346 ^ n3316;
  assign n3379 = ~n3347 & n3378;
  assign n3380 = n3379 ^ n3316;
  assign n3415 = n3414 ^ n3380;
  assign n3505 = n3504 ^ n3415;
  assign n3375 = n3348 ^ n3276;
  assign n3376 = ~n3349 & ~n3375;
  assign n3377 = n3376 ^ n3276;
  assign n3506 = n3505 ^ n3377;
  assign n3372 = n3350 ^ n3228;
  assign n3373 = n3351 & n3372;
  assign n3374 = n3373 ^ n3228;
  assign n3507 = n3506 ^ n3374;
  assign n3514 = n3513 ^ n3507;
  assign n3650 = n3504 ^ n3377;
  assign n3651 = n3505 & n3650;
  assign n3652 = n3651 ^ n3377;
  assign n3653 = ~n3374 & ~n3652;
  assign n3654 = n3415 & ~n3504;
  assign n3655 = ~n3377 & n3654;
  assign n3656 = ~n3653 & ~n3655;
  assign n3657 = n3513 & ~n3656;
  assign n3658 = ~n3374 & n3655;
  assign n3659 = ~n3657 & ~n3658;
  assign n3660 = ~n3415 & n3504;
  assign n3661 = n3377 & n3660;
  assign n3662 = ~n3374 & ~n3661;
  assign n3663 = n3652 & ~n3662;
  assign n3664 = ~n3513 & n3663;
  assign n3665 = n3374 & n3661;
  assign n3666 = ~n3664 & ~n3665;
  assign n3667 = n3659 & n3666;
  assign n3637 = n3445 ^ n3444;
  assign n3638 = n3447 & ~n3637;
  assign n3639 = n3638 ^ n3446;
  assign n3634 = n3455 ^ n3454;
  assign n3635 = n3457 & ~n3634;
  assign n3636 = n3635 ^ n3456;
  assign n3640 = n3639 ^ n3636;
  assign n3631 = n3402 ^ n3401;
  assign n3632 = n3403 & ~n3631;
  assign n3633 = n3632 ^ n1764;
  assign n3641 = n3640 ^ n3633;
  assign n3628 = n3409 ^ n3400;
  assign n3629 = ~n3410 & n3628;
  assign n3630 = n3629 ^ n3400;
  assign n3642 = n3641 ^ n3630;
  assign n3625 = n3453 ^ n3448;
  assign n3626 = n3459 & ~n3625;
  assign n3627 = n3626 ^ n3458;
  assign n3643 = n3642 ^ n3627;
  assign n3622 = n3460 ^ n3440;
  assign n3623 = n3461 & n3622;
  assign n3624 = n3623 ^ n3443;
  assign n3644 = n3643 ^ n3624;
  assign n3619 = n3411 ^ n3386;
  assign n3620 = ~n3412 & n3619;
  assign n3621 = n3620 ^ n3386;
  assign n3645 = n3644 ^ n3621;
  assign n3616 = n3500 ^ n3465;
  assign n3617 = ~n3501 & n3616;
  assign n3618 = n3617 ^ n3465;
  assign n3646 = n3645 ^ n3618;
  assign n3613 = n3383 ^ n3380;
  assign n3614 = ~n3414 & n3613;
  assign n3615 = n3614 ^ n3380;
  assign n3647 = n3646 ^ n3615;
  assign n3599 = n3472 ^ x45;
  assign n3600 = n3432 & n3599;
  assign n3601 = ~n3471 & ~n3600;
  assign n3602 = ~n3432 & ~n3599;
  assign n3603 = x1 & ~n3602;
  assign n3604 = ~n3601 & n3603;
  assign n3605 = ~x1 & n3472;
  assign n3606 = n3471 & n3605;
  assign n3607 = ~n3604 & ~n3606;
  assign n3596 = x13 & x34;
  assign n3595 = x12 & x35;
  assign n3597 = n3596 ^ n3595;
  assign n3594 = x7 & x40;
  assign n3598 = n3597 ^ n3594;
  assign n3608 = n3607 ^ n3598;
  assign n3591 = n3392 ^ n3389;
  assign n3592 = n3396 & ~n3591;
  assign n3593 = n3592 ^ n3395;
  assign n3609 = n3608 ^ n3593;
  assign n3588 = n3487 ^ n3468;
  assign n3589 = ~n3488 & n3588;
  assign n3590 = n3589 ^ n3468;
  assign n3610 = n3609 ^ n3590;
  assign n3585 = n3495 ^ n3492;
  assign n3586 = n3499 & ~n3585;
  assign n3587 = n3586 ^ n3498;
  assign n3611 = n3610 ^ n3587;
  assign n3577 = n3420 ^ n3419;
  assign n3578 = n3422 & ~n3577;
  assign n3579 = n3578 ^ n3421;
  assign n3574 = n3450 ^ n3449;
  assign n3575 = n3452 & ~n3574;
  assign n3576 = n3575 ^ n3451;
  assign n3580 = n3579 ^ n3576;
  assign n3572 = x1 & x46;
  assign n3573 = n3572 ^ x24;
  assign n3581 = n3580 ^ n3573;
  assign n3569 = n3439 ^ n3427;
  assign n3570 = ~n3428 & ~n3569;
  assign n3571 = n3570 ^ n3439;
  assign n3582 = n3581 ^ n3571;
  assign n3566 = n3482 ^ n3479;
  assign n3567 = n3486 & ~n3566;
  assign n3568 = n3567 ^ n3485;
  assign n3583 = n3582 ^ n3568;
  assign n3559 = n3425 ^ n1715;
  assign n3560 = ~n3426 & n3559;
  assign n3561 = n3560 ^ n1715;
  assign n3556 = n3406 ^ n3405;
  assign n3557 = n3408 & ~n3556;
  assign n3558 = n3557 ^ n3407;
  assign n3562 = n3561 ^ n3558;
  assign n3553 = x15 & x32;
  assign n3552 = x4 & x43;
  assign n3554 = n3553 ^ n3552;
  assign n3555 = n3554 ^ n3429;
  assign n3563 = n3562 ^ n3555;
  assign n3547 = x24 & n881;
  assign n3548 = n3547 ^ x2;
  assign n3549 = x45 & n3548;
  assign n3546 = x0 & x47;
  assign n3550 = n3549 ^ n3546;
  assign n3542 = x21 & x26;
  assign n3541 = x20 & x27;
  assign n3543 = n3542 ^ n3541;
  assign n3540 = x19 & x28;
  assign n3544 = n3543 ^ n3540;
  assign n3537 = x18 & x29;
  assign n3536 = x17 & x30;
  assign n3538 = n3537 ^ n3536;
  assign n3535 = x16 & x31;
  assign n3539 = n3538 ^ n3535;
  assign n3545 = n3544 ^ n3539;
  assign n3551 = n3550 ^ n3545;
  assign n3564 = n3563 ^ n3551;
  assign n3530 = x14 & x33;
  assign n3529 = x6 & x41;
  assign n3531 = n3530 ^ n3529;
  assign n3528 = x5 & x42;
  assign n3532 = n3531 ^ n3528;
  assign n3525 = x11 & x36;
  assign n3524 = x9 & x38;
  assign n3526 = n3525 ^ n3524;
  assign n3523 = x8 & x39;
  assign n3527 = n3526 ^ n3523;
  assign n3533 = n3532 ^ n3527;
  assign n3520 = x23 & x24;
  assign n3519 = x22 & x25;
  assign n3521 = n3520 ^ n3519;
  assign n3518 = x10 & x37;
  assign n3522 = n3521 ^ n3518;
  assign n3534 = n3533 ^ n3522;
  assign n3565 = n3564 ^ n3534;
  assign n3584 = n3583 ^ n3565;
  assign n3612 = n3611 ^ n3584;
  assign n3648 = n3647 ^ n3612;
  assign n3515 = n3502 ^ n3418;
  assign n3516 = n3503 & n3515;
  assign n3517 = n3516 ^ n3418;
  assign n3649 = n3648 ^ n3517;
  assign n3668 = n3667 ^ n3649;
  assign n3806 = ~n3649 & ~n3658;
  assign n3807 = ~n3663 & ~n3806;
  assign n3808 = ~n3513 & ~n3807;
  assign n3809 = n3649 & ~n3665;
  assign n3810 = n3656 & ~n3809;
  assign n3811 = ~n3808 & ~n3810;
  assign n3794 = x14 & x34;
  assign n3793 = x13 & x35;
  assign n3795 = n3794 ^ n3793;
  assign n3792 = x6 & x42;
  assign n3796 = n3795 ^ n3792;
  assign n3789 = x12 & x36;
  assign n3788 = x8 & x40;
  assign n3790 = n3789 ^ n3788;
  assign n3787 = x7 & x41;
  assign n3791 = n3790 ^ n3787;
  assign n3797 = n3796 ^ n3791;
  assign n3784 = x11 & x37;
  assign n3783 = x10 & x38;
  assign n3785 = n3784 ^ n3783;
  assign n3782 = x9 & x39;
  assign n3786 = n3785 ^ n3782;
  assign n3798 = n3797 ^ n3786;
  assign n3779 = n3598 ^ n3593;
  assign n3780 = ~n3608 & ~n3779;
  assign n3781 = n3780 ^ n3607;
  assign n3799 = n3798 ^ n3781;
  assign n3774 = x19 & x29;
  assign n3773 = x18 & x30;
  assign n3775 = n3774 ^ n3773;
  assign n3776 = n3775 ^ n1931;
  assign n3770 = x15 & x33;
  assign n3769 = x5 & x43;
  assign n3771 = n3770 ^ n3769;
  assign n3768 = x4 & x44;
  assign n3772 = n3771 ^ n3768;
  assign n3777 = n3776 ^ n3772;
  assign n3765 = x22 & x26;
  assign n3764 = x21 & x27;
  assign n3766 = n3765 ^ n3764;
  assign n3763 = x20 & x28;
  assign n3767 = n3766 ^ n3763;
  assign n3778 = n3777 ^ n3767;
  assign n3800 = n3799 ^ n3778;
  assign n3760 = n3590 ^ n3587;
  assign n3761 = n3610 & n3760;
  assign n3762 = n3761 ^ n3587;
  assign n3801 = n3800 ^ n3762;
  assign n3757 = n3624 ^ n3621;
  assign n3758 = ~n3644 & n3757;
  assign n3759 = n3758 ^ n3621;
  assign n3802 = n3801 ^ n3759;
  assign n3746 = n3547 ^ n3546;
  assign n3747 = n3548 & ~n3746;
  assign n3748 = n3747 ^ x2;
  assign n3749 = x45 & n3748;
  assign n3742 = n3536 ^ n3535;
  assign n3743 = n3538 & ~n3742;
  assign n3744 = n3743 ^ n3537;
  assign n3739 = n3553 ^ n3429;
  assign n3740 = ~n3554 & n3739;
  assign n3741 = n3740 ^ n3429;
  assign n3745 = n3744 ^ n3741;
  assign n3750 = n3749 ^ n3745;
  assign n3736 = n3576 ^ n3573;
  assign n3737 = n3580 & ~n3736;
  assign n3738 = n3737 ^ n3579;
  assign n3751 = n3750 ^ n3738;
  assign n3733 = n3550 ^ n3544;
  assign n3734 = ~n3545 & n3733;
  assign n3735 = n3734 ^ n3550;
  assign n3752 = n3751 ^ n3735;
  assign n3726 = x16 & x32;
  assign n3725 = x3 & x45;
  assign n3727 = n3726 ^ n3725;
  assign n3724 = x2 & x46;
  assign n3728 = n3727 ^ n3724;
  assign n3721 = n3595 ^ n3594;
  assign n3722 = n3597 & ~n3721;
  assign n3723 = n3722 ^ n3596;
  assign n3729 = n3728 ^ n3723;
  assign n3718 = n3519 ^ n3518;
  assign n3719 = n3521 & ~n3718;
  assign n3720 = n3719 ^ n3520;
  assign n3730 = n3729 ^ n3720;
  assign n3715 = n3527 ^ n3522;
  assign n3716 = n3533 & ~n3715;
  assign n3717 = n3716 ^ n3532;
  assign n3731 = n3730 ^ n3717;
  assign n3710 = n3529 ^ n3528;
  assign n3711 = n3531 & ~n3710;
  assign n3712 = n3711 ^ n3530;
  assign n3707 = n3541 ^ n3540;
  assign n3708 = n3543 & ~n3707;
  assign n3709 = n3708 ^ n3542;
  assign n3713 = n3712 ^ n3709;
  assign n3704 = n3524 ^ n3523;
  assign n3705 = n3526 & ~n3704;
  assign n3706 = n3705 ^ n3525;
  assign n3714 = n3713 ^ n3706;
  assign n3732 = n3731 ^ n3714;
  assign n3753 = n3752 ^ n3732;
  assign n3701 = n3551 ^ n3534;
  assign n3702 = n3564 & ~n3701;
  assign n3703 = n3702 ^ n3563;
  assign n3754 = n3753 ^ n3703;
  assign n3698 = n3611 ^ n3583;
  assign n3699 = n3584 & n3698;
  assign n3700 = n3699 ^ n3611;
  assign n3755 = n3754 ^ n3700;
  assign n3691 = x46 & n1056;
  assign n3689 = x1 & x47;
  assign n3688 = x23 & x25;
  assign n3690 = n3689 ^ n3688;
  assign n3692 = n3691 ^ n3690;
  assign n3687 = x0 & x48;
  assign n3693 = n3692 ^ n3687;
  assign n3684 = n3636 ^ n3633;
  assign n3685 = n3640 & ~n3684;
  assign n3686 = n3685 ^ n3639;
  assign n3694 = n3693 ^ n3686;
  assign n3681 = n3558 ^ n3555;
  assign n3682 = n3562 & ~n3681;
  assign n3683 = n3682 ^ n3561;
  assign n3695 = n3694 ^ n3683;
  assign n3678 = n3581 ^ n3568;
  assign n3679 = ~n3582 & ~n3678;
  assign n3680 = n3679 ^ n3571;
  assign n3696 = n3695 ^ n3680;
  assign n3675 = n3641 ^ n3627;
  assign n3676 = n3642 & ~n3675;
  assign n3677 = n3676 ^ n3630;
  assign n3697 = n3696 ^ n3677;
  assign n3756 = n3755 ^ n3697;
  assign n3803 = n3802 ^ n3756;
  assign n3672 = n3618 ^ n3615;
  assign n3673 = ~n3646 & n3672;
  assign n3674 = n3673 ^ n3615;
  assign n3804 = n3803 ^ n3674;
  assign n3669 = n3612 ^ n3517;
  assign n3670 = n3648 & ~n3669;
  assign n3671 = n3670 ^ n3647;
  assign n3805 = n3804 ^ n3671;
  assign n3812 = n3811 ^ n3805;
  assign n3945 = n3693 ^ n3683;
  assign n3946 = n3694 & ~n3945;
  assign n3947 = n3946 ^ n3686;
  assign n3942 = n3772 ^ n3767;
  assign n3943 = n3777 & ~n3942;
  assign n3944 = n3943 ^ n3776;
  assign n3948 = n3947 ^ n3944;
  assign n3937 = n3774 ^ n1931;
  assign n3938 = ~n3775 & n3937;
  assign n3939 = n3938 ^ n1931;
  assign n3934 = n3788 ^ n3787;
  assign n3935 = n3790 & ~n3934;
  assign n3936 = n3935 ^ n3789;
  assign n3940 = n3939 ^ n3936;
  assign n3931 = n3793 ^ n3792;
  assign n3932 = n3795 & ~n3931;
  assign n3933 = n3932 ^ n3794;
  assign n3941 = n3940 ^ n3933;
  assign n3949 = n3948 ^ n3941;
  assign n3924 = x23 & x47;
  assign n3925 = x1 & n3924;
  assign n3926 = x25 & ~n3925;
  assign n3923 = x1 & x48;
  assign n3927 = n3926 ^ n3923;
  assign n3920 = n3783 ^ n3782;
  assign n3921 = n3785 & ~n3920;
  assign n3922 = n3921 ^ n3784;
  assign n3928 = n3927 ^ n3922;
  assign n3917 = n3791 ^ n3786;
  assign n3918 = n3797 & ~n3917;
  assign n3919 = n3918 ^ n3796;
  assign n3929 = n3928 ^ n3919;
  assign n3912 = n3769 ^ n3768;
  assign n3913 = n3771 & ~n3912;
  assign n3914 = n3913 ^ n3770;
  assign n3909 = n3725 ^ n3724;
  assign n3910 = n3727 & ~n3909;
  assign n3911 = n3910 ^ n3726;
  assign n3915 = n3914 ^ n3911;
  assign n3906 = n3764 ^ n3763;
  assign n3907 = n3766 & ~n3906;
  assign n3908 = n3907 ^ n3765;
  assign n3916 = n3915 ^ n3908;
  assign n3930 = n3929 ^ n3916;
  assign n3950 = n3949 ^ n3930;
  assign n3903 = n3798 ^ n3778;
  assign n3904 = ~n3799 & ~n3903;
  assign n3905 = n3904 ^ n3781;
  assign n3951 = n3950 ^ n3905;
  assign n3896 = n3709 ^ n3706;
  assign n3897 = n3713 & ~n3896;
  assign n3898 = n3897 ^ n3712;
  assign n3893 = n3728 ^ n3720;
  assign n3894 = n3729 & ~n3893;
  assign n3895 = n3894 ^ n3723;
  assign n3899 = n3898 ^ n3895;
  assign n3890 = n3749 ^ n3744;
  assign n3891 = ~n3745 & n3890;
  assign n3892 = n3891 ^ n3749;
  assign n3900 = n3899 ^ n3892;
  assign n3887 = n3730 ^ n3714;
  assign n3888 = n3731 & ~n3887;
  assign n3889 = n3888 ^ n3717;
  assign n3901 = n3900 ^ n3889;
  assign n3884 = n3750 ^ n3735;
  assign n3885 = n3751 & ~n3884;
  assign n3886 = n3885 ^ n3738;
  assign n3902 = n3901 ^ n3886;
  assign n3952 = n3951 ^ n3902;
  assign n3881 = n3800 ^ n3759;
  assign n3882 = n3801 & ~n3881;
  assign n3883 = n3882 ^ n3759;
  assign n3953 = n3952 ^ n3883;
  assign n3871 = x18 & x31;
  assign n3872 = n3871 ^ n1883;
  assign n3870 = x16 & x33;
  assign n3873 = n3872 ^ n3870;
  assign n3867 = x5 & x44;
  assign n3866 = x4 & x45;
  assign n3868 = n3867 ^ n3866;
  assign n3865 = x0 & x49;
  assign n3869 = n3868 ^ n3865;
  assign n3874 = n3873 ^ n3869;
  assign n3862 = n3690 ^ n3687;
  assign n3863 = n3692 & ~n3862;
  assign n3864 = n3863 ^ n3691;
  assign n3875 = n3874 ^ n3864;
  assign n3857 = x24 & x25;
  assign n3856 = x23 & x26;
  assign n3858 = n3857 ^ n3856;
  assign n3855 = x11 & x38;
  assign n3859 = n3858 ^ n3855;
  assign n3852 = x15 & x34;
  assign n3851 = x14 & x35;
  assign n3853 = n3852 ^ n3851;
  assign n3850 = x6 & x43;
  assign n3854 = n3853 ^ n3850;
  assign n3860 = n3859 ^ n3854;
  assign n3847 = x13 & x36;
  assign n3846 = x8 & x41;
  assign n3848 = n3847 ^ n3846;
  assign n3845 = x7 & x42;
  assign n3849 = n3848 ^ n3845;
  assign n3861 = n3860 ^ n3849;
  assign n3876 = n3875 ^ n3861;
  assign n3840 = x21 & x28;
  assign n3839 = x20 & x29;
  assign n3841 = n3840 ^ n3839;
  assign n3838 = x19 & x30;
  assign n3842 = n3841 ^ n3838;
  assign n3835 = x22 & x27;
  assign n3834 = x3 & x46;
  assign n3836 = n3835 ^ n3834;
  assign n3833 = x2 & x47;
  assign n3837 = n3836 ^ n3833;
  assign n3843 = n3842 ^ n3837;
  assign n3830 = x12 & x37;
  assign n3829 = x10 & x39;
  assign n3831 = n3830 ^ n3829;
  assign n3828 = x9 & x40;
  assign n3832 = n3831 ^ n3828;
  assign n3844 = n3843 ^ n3832;
  assign n3877 = n3876 ^ n3844;
  assign n3825 = n3732 ^ n3703;
  assign n3826 = n3753 & ~n3825;
  assign n3827 = n3826 ^ n3752;
  assign n3878 = n3877 ^ n3827;
  assign n3822 = n3680 ^ n3677;
  assign n3823 = n3696 & ~n3822;
  assign n3824 = n3823 ^ n3677;
  assign n3879 = n3878 ^ n3824;
  assign n3819 = n3754 ^ n3697;
  assign n3820 = ~n3755 & n3819;
  assign n3821 = n3820 ^ n3700;
  assign n3880 = n3879 ^ n3821;
  assign n3954 = n3953 ^ n3880;
  assign n3816 = n3802 ^ n3674;
  assign n3817 = n3803 & ~n3816;
  assign n3818 = n3817 ^ n3674;
  assign n3955 = n3954 ^ n3818;
  assign n3813 = n3811 ^ n3671;
  assign n3814 = n3805 & n3813;
  assign n3815 = n3814 ^ n3811;
  assign n3956 = n3955 ^ n3815;
  assign n4103 = n3821 & ~n3879;
  assign n4104 = n3953 & n4103;
  assign n4105 = n3818 & ~n4104;
  assign n4106 = n3953 ^ n3821;
  assign n4107 = n3880 & n4106;
  assign n4108 = n4107 ^ n3953;
  assign n4109 = ~n4105 & n4108;
  assign n4110 = ~n3815 & n4109;
  assign n4111 = ~n3818 & n4104;
  assign n4112 = ~n4110 & ~n4111;
  assign n4113 = n3818 & ~n4108;
  assign n4114 = ~n3821 & n3879;
  assign n4115 = ~n3953 & n4114;
  assign n4116 = ~n4113 & ~n4115;
  assign n4117 = n3815 & ~n4116;
  assign n4118 = n3818 & n4115;
  assign n4119 = ~n4117 & ~n4118;
  assign n4120 = n4112 & n4119;
  assign n4092 = n3936 ^ n3933;
  assign n4093 = n3940 & ~n4092;
  assign n4094 = n4093 ^ n3939;
  assign n4089 = n3911 ^ n3908;
  assign n4090 = n3915 & ~n4089;
  assign n4091 = n4090 ^ n3914;
  assign n4095 = n4094 ^ n4091;
  assign n4084 = n3851 ^ n3850;
  assign n4085 = n3853 & ~n4084;
  assign n4086 = n4085 ^ n3852;
  assign n4081 = n3834 ^ n3833;
  assign n4082 = n3836 & ~n4081;
  assign n4083 = n4082 ^ n3835;
  assign n4087 = n4086 ^ n4083;
  assign n4078 = n3866 ^ n3865;
  assign n4079 = n3868 & ~n4078;
  assign n4080 = n4079 ^ n3867;
  assign n4088 = n4087 ^ n4080;
  assign n4096 = n4095 ^ n4088;
  assign n4075 = n3928 ^ n3916;
  assign n4076 = n3929 & ~n4075;
  assign n4077 = n4076 ^ n3919;
  assign n4097 = n4096 ^ n4077;
  assign n4072 = n3944 ^ n3941;
  assign n4073 = n3948 & ~n4072;
  assign n4074 = n4073 ^ n3947;
  assign n4098 = n4097 ^ n4074;
  assign n4063 = n3829 ^ n3828;
  assign n4064 = n3831 & ~n4063;
  assign n4065 = n4064 ^ n3830;
  assign n4060 = n3856 ^ n3855;
  assign n4061 = n3858 & ~n4060;
  assign n4062 = n4061 ^ n3857;
  assign n4066 = n4065 ^ n4062;
  assign n4058 = x1 & x49;
  assign n4057 = x24 & x26;
  assign n4059 = n4058 ^ n4057;
  assign n4067 = n4066 ^ n4059;
  assign n4054 = n3837 ^ n3832;
  assign n4055 = n3843 & ~n4054;
  assign n4056 = n4055 ^ n3842;
  assign n4068 = n4067 ^ n4056;
  assign n4051 = n3873 ^ n3864;
  assign n4052 = ~n3874 & n4051;
  assign n4053 = n4052 ^ n3864;
  assign n4069 = n4068 ^ n4053;
  assign n4048 = n3861 ^ n3844;
  assign n4049 = n3876 & ~n4048;
  assign n4050 = n4049 ^ n3875;
  assign n4070 = n4069 ^ n4050;
  assign n4041 = n3839 ^ n3838;
  assign n4042 = n3841 & ~n4041;
  assign n4043 = n4042 ^ n3840;
  assign n4038 = n3846 ^ n3845;
  assign n4039 = n3848 & ~n4038;
  assign n4040 = n4039 ^ n3847;
  assign n4044 = n4043 ^ n4040;
  assign n4035 = n3871 ^ n3870;
  assign n4036 = n3872 & ~n4035;
  assign n4037 = n4036 ^ n1883;
  assign n4045 = n4044 ^ n4037;
  assign n4032 = n3854 ^ n3849;
  assign n4033 = n3860 & ~n4032;
  assign n4034 = n4033 ^ n3859;
  assign n4046 = n4045 ^ n4034;
  assign n4029 = n3895 ^ n3892;
  assign n4030 = n3899 & ~n4029;
  assign n4031 = n4030 ^ n3898;
  assign n4047 = n4046 ^ n4031;
  assign n4071 = n4070 ^ n4047;
  assign n4099 = n4098 ^ n4071;
  assign n4026 = n3827 ^ n3824;
  assign n4027 = ~n3878 & n4026;
  assign n4028 = n4027 ^ n3824;
  assign n4100 = n4099 ^ n4028;
  assign n4011 = x48 & n3922;
  assign n4012 = x25 & x47;
  assign n4013 = x23 & n4012;
  assign n4014 = ~n4011 & ~n4013;
  assign n4015 = x25 & x48;
  assign n4016 = x1 & ~n4015;
  assign n4017 = ~n4014 & n4016;
  assign n4018 = n3923 & ~n3924;
  assign n4019 = x25 & ~n4018;
  assign n4020 = n3922 & n4019;
  assign n4021 = ~n4017 & ~n4020;
  assign n4007 = x23 & x27;
  assign n4006 = x22 & x28;
  assign n4008 = n4007 ^ n4006;
  assign n4005 = x18 & x32;
  assign n4009 = n4008 ^ n4005;
  assign n4002 = x16 & x34;
  assign n4001 = x15 & x35;
  assign n4003 = n4002 ^ n4001;
  assign n4000 = x5 & x45;
  assign n4004 = n4003 ^ n4000;
  assign n4010 = n4009 ^ n4004;
  assign n4022 = n4021 ^ n4010;
  assign n3996 = x0 & x50;
  assign n3994 = n1102 ^ x2;
  assign n3995 = x48 & n3994;
  assign n3997 = n3996 ^ n3995;
  assign n3990 = x17 & x33;
  assign n3989 = x4 & x46;
  assign n3991 = n3990 ^ n3989;
  assign n3988 = x3 & x47;
  assign n3992 = n3991 ^ n3988;
  assign n3985 = x21 & x29;
  assign n3984 = x20 & x30;
  assign n3986 = n3985 ^ n3984;
  assign n3983 = x19 & x31;
  assign n3987 = n3986 ^ n3983;
  assign n3993 = n3992 ^ n3987;
  assign n3998 = n3997 ^ n3993;
  assign n3978 = x14 & x36;
  assign n3977 = x7 & x43;
  assign n3979 = n3978 ^ n3977;
  assign n3976 = x6 & x44;
  assign n3980 = n3979 ^ n3976;
  assign n3973 = x12 & x38;
  assign n3972 = x11 & x39;
  assign n3974 = n3973 ^ n3972;
  assign n3971 = x10 & x40;
  assign n3975 = n3974 ^ n3971;
  assign n3981 = n3980 ^ n3975;
  assign n3968 = x13 & x37;
  assign n3967 = x9 & x41;
  assign n3969 = n3968 ^ n3967;
  assign n3966 = x8 & x42;
  assign n3970 = n3969 ^ n3966;
  assign n3982 = n3981 ^ n3970;
  assign n3999 = n3998 ^ n3982;
  assign n4023 = n4022 ^ n3999;
  assign n3963 = n3889 ^ n3886;
  assign n3964 = ~n3901 & n3963;
  assign n3965 = n3964 ^ n3886;
  assign n4024 = n4023 ^ n3965;
  assign n3960 = n3949 ^ n3905;
  assign n3961 = ~n3950 & ~n3960;
  assign n3962 = n3961 ^ n3905;
  assign n4025 = n4024 ^ n3962;
  assign n4101 = n4100 ^ n4025;
  assign n3957 = n3951 ^ n3883;
  assign n3958 = n3952 & ~n3957;
  assign n3959 = n3958 ^ n3883;
  assign n4102 = n4101 ^ n3959;
  assign n4121 = n4120 ^ n4102;
  assign n4271 = n4102 & ~n4109;
  assign n4272 = ~n4118 & ~n4271;
  assign n4273 = ~n3815 & n4272;
  assign n4274 = n4102 & ~n4111;
  assign n4275 = n4116 & ~n4274;
  assign n4276 = ~n4273 & ~n4275;
  assign n4260 = x0 & x51;
  assign n4259 = x1 & x50;
  assign n4261 = n4260 ^ n4259;
  assign n4255 = x24 & x49;
  assign n4256 = x26 & n4255;
  assign n4257 = x1 & n4256;
  assign n4258 = n4257 ^ x26;
  assign n4262 = n4261 ^ n4258;
  assign n4252 = n4040 ^ n4037;
  assign n4253 = n4044 & ~n4252;
  assign n4254 = n4253 ^ n4043;
  assign n4263 = n4262 ^ n4254;
  assign n4249 = x20 & x31;
  assign n4248 = x19 & x32;
  assign n4250 = n4249 ^ n4248;
  assign n4247 = x17 & x34;
  assign n4251 = n4250 ^ n4247;
  assign n4264 = n4263 ^ n4251;
  assign n4241 = x25 & x26;
  assign n4240 = x24 & x27;
  assign n4242 = n4241 ^ n4240;
  assign n4239 = x11 & x40;
  assign n4243 = n4242 ^ n4239;
  assign n4236 = x13 & x38;
  assign n4235 = x8 & x43;
  assign n4237 = n4236 ^ n4235;
  assign n4234 = x7 & x44;
  assign n4238 = n4237 ^ n4234;
  assign n4244 = n4243 ^ n4238;
  assign n4231 = x12 & x39;
  assign n4230 = x10 & x41;
  assign n4232 = n4231 ^ n4230;
  assign n4229 = x9 & x42;
  assign n4233 = n4232 ^ n4229;
  assign n4245 = n4244 ^ n4233;
  assign n4224 = x15 & x36;
  assign n4223 = x14 & x37;
  assign n4225 = n4224 ^ n4223;
  assign n4222 = x6 & x45;
  assign n4226 = n4225 ^ n4222;
  assign n4219 = x23 & x28;
  assign n4218 = x22 & x29;
  assign n4220 = n4219 ^ n4218;
  assign n4217 = x21 & x30;
  assign n4221 = n4220 ^ n4217;
  assign n4227 = n4226 ^ n4221;
  assign n4214 = x18 & x33;
  assign n4213 = x16 & x35;
  assign n4215 = n4214 ^ n4213;
  assign n4212 = x5 & x46;
  assign n4216 = n4215 ^ n4212;
  assign n4228 = n4227 ^ n4216;
  assign n4246 = n4245 ^ n4228;
  assign n4265 = n4264 ^ n4246;
  assign n4209 = n4069 ^ n4047;
  assign n4210 = n4070 & ~n4209;
  assign n4211 = n4210 ^ n4050;
  assign n4266 = n4265 ^ n4211;
  assign n4206 = n4077 ^ n4074;
  assign n4207 = ~n4097 & n4206;
  assign n4208 = n4207 ^ n4074;
  assign n4267 = n4266 ^ n4208;
  assign n4203 = n4098 ^ n4028;
  assign n4204 = ~n4099 & n4203;
  assign n4205 = n4204 ^ n4028;
  assign n4268 = n4267 ^ n4205;
  assign n4192 = n4006 ^ n4005;
  assign n4193 = n4008 & ~n4192;
  assign n4194 = n4193 ^ n4007;
  assign n4189 = n3977 ^ n3976;
  assign n4190 = n3979 & ~n4189;
  assign n4191 = n4190 ^ n3978;
  assign n4195 = n4194 ^ n4191;
  assign n4186 = n3967 ^ n3966;
  assign n4187 = n3969 & ~n4186;
  assign n4188 = n4187 ^ n3968;
  assign n4196 = n4195 ^ n4188;
  assign n4183 = n3975 ^ n3970;
  assign n4184 = n3981 & ~n4183;
  assign n4185 = n4184 ^ n3980;
  assign n4197 = n4196 ^ n4185;
  assign n4178 = ~x2 & ~n1102;
  assign n4179 = x48 & ~n4178;
  assign n4177 = n3995 & ~n3996;
  assign n4180 = n4179 ^ n4177;
  assign n4174 = n3989 ^ n3988;
  assign n4175 = n3991 & ~n4174;
  assign n4176 = n4175 ^ n3990;
  assign n4181 = n4180 ^ n4176;
  assign n4171 = n3984 ^ n3983;
  assign n4172 = n3986 & ~n4171;
  assign n4173 = n4172 ^ n3985;
  assign n4182 = n4181 ^ n4173;
  assign n4198 = n4197 ^ n4182;
  assign n4168 = n4022 ^ n3998;
  assign n4169 = ~n3999 & ~n4168;
  assign n4170 = n4169 ^ n4022;
  assign n4199 = n4198 ^ n4170;
  assign n4161 = x4 & x47;
  assign n4160 = x3 & x48;
  assign n4162 = n4161 ^ n4160;
  assign n4159 = x2 & x49;
  assign n4163 = n4162 ^ n4159;
  assign n4156 = n3972 ^ n3971;
  assign n4157 = n3974 & ~n4156;
  assign n4158 = n4157 ^ n3973;
  assign n4164 = n4163 ^ n4158;
  assign n4153 = n4001 ^ n4000;
  assign n4154 = n4003 & ~n4153;
  assign n4155 = n4154 ^ n4002;
  assign n4165 = n4164 ^ n4155;
  assign n4150 = n4021 ^ n4009;
  assign n4151 = ~n4010 & ~n4150;
  assign n4152 = n4151 ^ n4021;
  assign n4166 = n4165 ^ n4152;
  assign n4147 = n4091 ^ n4088;
  assign n4148 = n4095 & ~n4147;
  assign n4149 = n4148 ^ n4094;
  assign n4167 = n4166 ^ n4149;
  assign n4200 = n4199 ^ n4167;
  assign n4140 = n4062 ^ n4059;
  assign n4141 = n4066 & ~n4140;
  assign n4142 = n4141 ^ n4065;
  assign n4137 = n4083 ^ n4080;
  assign n4138 = n4087 & ~n4137;
  assign n4139 = n4138 ^ n4086;
  assign n4143 = n4142 ^ n4139;
  assign n4134 = n3997 ^ n3992;
  assign n4135 = ~n3993 & n4134;
  assign n4136 = n4135 ^ n3997;
  assign n4144 = n4143 ^ n4136;
  assign n4131 = n4056 ^ n4053;
  assign n4132 = ~n4068 & n4131;
  assign n4133 = n4132 ^ n4053;
  assign n4145 = n4144 ^ n4133;
  assign n4128 = n4034 ^ n4031;
  assign n4129 = ~n4046 & n4128;
  assign n4130 = n4129 ^ n4031;
  assign n4146 = n4145 ^ n4130;
  assign n4201 = n4200 ^ n4146;
  assign n4125 = n3965 ^ n3962;
  assign n4126 = n4024 & ~n4125;
  assign n4127 = n4126 ^ n3962;
  assign n4202 = n4201 ^ n4127;
  assign n4269 = n4268 ^ n4202;
  assign n4122 = n4100 ^ n3959;
  assign n4123 = ~n4101 & n4122;
  assign n4124 = n4123 ^ n3959;
  assign n4270 = n4269 ^ n4124;
  assign n4277 = n4276 ^ n4270;
  assign n4423 = x19 & x33;
  assign n4422 = x3 & x49;
  assign n4424 = n4423 ^ n4422;
  assign n4421 = x2 & x50;
  assign n4425 = n4424 ^ n4421;
  assign n4418 = n4191 ^ n4188;
  assign n4419 = n4195 & ~n4418;
  assign n4420 = n4419 ^ n4194;
  assign n4426 = n4425 ^ n4420;
  assign n4415 = n4176 ^ n4173;
  assign n4416 = n4181 & ~n4415;
  assign n4417 = n4416 ^ n4180;
  assign n4427 = n4426 ^ n4417;
  assign n4353 = x26 & x50;
  assign n4409 = n4353 ^ x51;
  assign n4410 = x1 & n4409;
  assign n4408 = x25 & x27;
  assign n4411 = n4410 ^ n4408;
  assign n4405 = n4240 ^ n4239;
  assign n4406 = n4242 & ~n4405;
  assign n4407 = n4406 ^ n4241;
  assign n4412 = n4411 ^ n4407;
  assign n4402 = n4238 ^ n4233;
  assign n4403 = n4244 & ~n4402;
  assign n4404 = n4403 ^ n4243;
  assign n4413 = n4412 ^ n4404;
  assign n4399 = n4163 ^ n4155;
  assign n4400 = n4164 & ~n4399;
  assign n4401 = n4400 ^ n4158;
  assign n4414 = n4413 ^ n4401;
  assign n4428 = n4427 ^ n4414;
  assign n4396 = n4165 ^ n4149;
  assign n4397 = ~n4166 & ~n4396;
  assign n4398 = n4397 ^ n4152;
  assign n4429 = n4428 ^ n4398;
  assign n4387 = n4223 ^ n4222;
  assign n4388 = n4225 & ~n4387;
  assign n4389 = n4388 ^ n4224;
  assign n4384 = n4248 ^ n4247;
  assign n4385 = n4250 & ~n4384;
  assign n4386 = n4385 ^ n4249;
  assign n4390 = n4389 ^ n4386;
  assign n4381 = n4160 ^ n4159;
  assign n4382 = n4162 & ~n4381;
  assign n4383 = n4382 ^ n4161;
  assign n4391 = n4390 ^ n4383;
  assign n4378 = n4221 ^ n4216;
  assign n4379 = n4227 & ~n4378;
  assign n4380 = n4379 ^ n4226;
  assign n4392 = n4391 ^ n4380;
  assign n4373 = n4218 ^ n4217;
  assign n4374 = n4220 & ~n4373;
  assign n4375 = n4374 ^ n4219;
  assign n4370 = n4235 ^ n4234;
  assign n4371 = n4237 & ~n4370;
  assign n4372 = n4371 ^ n4236;
  assign n4376 = n4375 ^ n4372;
  assign n4367 = n4213 ^ n4212;
  assign n4368 = n4215 & ~n4367;
  assign n4369 = n4368 ^ n4214;
  assign n4377 = n4376 ^ n4369;
  assign n4393 = n4392 ^ n4377;
  assign n4364 = n4264 ^ n4245;
  assign n4365 = ~n4246 & n4364;
  assign n4366 = n4365 ^ n4264;
  assign n4394 = n4393 ^ n4366;
  assign n4351 = x51 & n3996;
  assign n4352 = ~n4256 & ~n4351;
  assign n4354 = x1 & ~n4353;
  assign n4355 = ~n4352 & n4354;
  assign n4356 = ~n4255 & n4259;
  assign n4357 = x26 & x51;
  assign n4358 = x0 & n4357;
  assign n4359 = ~n4356 & n4358;
  assign n4360 = ~n4355 & ~n4359;
  assign n4347 = x4 & x48;
  assign n4348 = n4347 ^ n2209;
  assign n4346 = x0 & x52;
  assign n4349 = n4348 ^ n4346;
  assign n4343 = n4230 ^ n4229;
  assign n4344 = n4232 & ~n4343;
  assign n4345 = n4344 ^ n4231;
  assign n4350 = n4349 ^ n4345;
  assign n4361 = n4360 ^ n4350;
  assign n4340 = n4262 ^ n4251;
  assign n4341 = n4263 & ~n4340;
  assign n4342 = n4341 ^ n4254;
  assign n4362 = n4361 ^ n4342;
  assign n4337 = n4139 ^ n4136;
  assign n4338 = n4143 & ~n4337;
  assign n4339 = n4338 ^ n4142;
  assign n4363 = n4362 ^ n4339;
  assign n4395 = n4394 ^ n4363;
  assign n4430 = n4429 ^ n4395;
  assign n4334 = n4211 ^ n4208;
  assign n4335 = ~n4266 & n4334;
  assign n4336 = n4335 ^ n4208;
  assign n4431 = n4430 ^ n4336;
  assign n4325 = x12 & x40;
  assign n4324 = x11 & x41;
  assign n4326 = n4325 ^ n4324;
  assign n4323 = x10 & x42;
  assign n4327 = n4326 ^ n4323;
  assign n4320 = x15 & x37;
  assign n4319 = x8 & x44;
  assign n4321 = n4320 ^ n4319;
  assign n4318 = x7 & x45;
  assign n4322 = n4321 ^ n4318;
  assign n4328 = n4327 ^ n4322;
  assign n4315 = x16 & x36;
  assign n4314 = x6 & x46;
  assign n4316 = n4315 ^ n4314;
  assign n4313 = x5 & x47;
  assign n4317 = n4316 ^ n4313;
  assign n4329 = n4328 ^ n4317;
  assign n4308 = x24 & x28;
  assign n4307 = x23 & x29;
  assign n4309 = n4308 ^ n4307;
  assign n4306 = x22 & x30;
  assign n4310 = n4309 ^ n4306;
  assign n4303 = x14 & x38;
  assign n4302 = x13 & x39;
  assign n4304 = n4303 ^ n4302;
  assign n4301 = x9 & x43;
  assign n4305 = n4304 ^ n4301;
  assign n4311 = n4310 ^ n4305;
  assign n4298 = x21 & x31;
  assign n4297 = x20 & x32;
  assign n4299 = n4298 ^ n4297;
  assign n4296 = x18 & x34;
  assign n4300 = n4299 ^ n4296;
  assign n4312 = n4311 ^ n4300;
  assign n4330 = n4329 ^ n4312;
  assign n4293 = n4196 ^ n4182;
  assign n4294 = n4197 & ~n4293;
  assign n4295 = n4294 ^ n4185;
  assign n4331 = n4330 ^ n4295;
  assign n4290 = n4133 ^ n4130;
  assign n4291 = ~n4145 & n4290;
  assign n4292 = n4291 ^ n4130;
  assign n4332 = n4331 ^ n4292;
  assign n4287 = n4198 ^ n4167;
  assign n4288 = ~n4199 & n4287;
  assign n4289 = n4288 ^ n4170;
  assign n4333 = n4332 ^ n4289;
  assign n4432 = n4431 ^ n4333;
  assign n4284 = n4200 ^ n4127;
  assign n4285 = ~n4201 & ~n4284;
  assign n4286 = n4285 ^ n4127;
  assign n4433 = n4432 ^ n4286;
  assign n4281 = n4267 ^ n4202;
  assign n4282 = n4268 & n4281;
  assign n4283 = n4282 ^ n4205;
  assign n4434 = n4433 ^ n4283;
  assign n4278 = n4276 ^ n4124;
  assign n4279 = n4270 & n4278;
  assign n4280 = n4279 ^ n4276;
  assign n4435 = n4434 ^ n4280;
  assign n4590 = ~n4283 & ~n4431;
  assign n4591 = ~n4286 & ~n4333;
  assign n4592 = n4590 & ~n4591;
  assign n4593 = n4283 & n4431;
  assign n4594 = n4286 & n4333;
  assign n4595 = ~n4593 & n4594;
  assign n4596 = ~n4592 & ~n4595;
  assign n4597 = ~n4280 & ~n4596;
  assign n4598 = n4286 ^ n4283;
  assign n4599 = n4431 ^ n4286;
  assign n4600 = n4432 & n4599;
  assign n4601 = n4598 & n4600;
  assign n4602 = ~n4597 & ~n4601;
  assign n4603 = ~n4590 & n4591;
  assign n4604 = n4593 & ~n4594;
  assign n4605 = ~n4603 & ~n4604;
  assign n4606 = n4280 & ~n4605;
  assign n4607 = n4602 & ~n4606;
  assign n4579 = n4360 ^ n4345;
  assign n4580 = ~n4350 & ~n4579;
  assign n4581 = n4580 ^ n4360;
  assign n4576 = n4305 ^ n4300;
  assign n4577 = n4311 & ~n4576;
  assign n4578 = n4577 ^ n4310;
  assign n4582 = n4581 ^ n4578;
  assign n4571 = n4307 ^ n4306;
  assign n4572 = n4309 & ~n4571;
  assign n4573 = n4572 ^ n4308;
  assign n4568 = n4347 ^ n4346;
  assign n4569 = n4348 & ~n4568;
  assign n4570 = n4569 ^ n2209;
  assign n4574 = n4573 ^ n4570;
  assign n4565 = n4422 ^ n4421;
  assign n4566 = n4424 & ~n4565;
  assign n4567 = n4566 ^ n4423;
  assign n4575 = n4574 ^ n4567;
  assign n4583 = n4582 ^ n4575;
  assign n4558 = n4314 ^ n4313;
  assign n4559 = n4316 & ~n4558;
  assign n4560 = n4559 ^ n4315;
  assign n4555 = n4319 ^ n4318;
  assign n4556 = n4321 & ~n4555;
  assign n4557 = n4556 ^ n4320;
  assign n4561 = n4560 ^ n4557;
  assign n4552 = n4297 ^ n4296;
  assign n4553 = n4299 & ~n4552;
  assign n4554 = n4553 ^ n4298;
  assign n4562 = n4561 ^ n4554;
  assign n4547 = n4302 ^ n4301;
  assign n4548 = n4304 & ~n4547;
  assign n4549 = n4548 ^ n4303;
  assign n4544 = n4324 ^ n4323;
  assign n4545 = n4326 & ~n4544;
  assign n4546 = n4545 ^ n4325;
  assign n4550 = n4549 ^ n4546;
  assign n4542 = x1 & x52;
  assign n4543 = n4542 ^ x27;
  assign n4551 = n4550 ^ n4543;
  assign n4563 = n4562 ^ n4551;
  assign n4539 = n4322 ^ n4317;
  assign n4540 = n4328 & ~n4539;
  assign n4541 = n4540 ^ n4327;
  assign n4564 = n4563 ^ n4541;
  assign n4584 = n4583 ^ n4564;
  assign n4536 = n4427 ^ n4398;
  assign n4537 = ~n4428 & ~n4536;
  assign n4538 = n4537 ^ n4398;
  assign n4585 = n4584 ^ n4538;
  assign n4523 = n4408 ^ x51;
  assign n4524 = n4353 & n4523;
  assign n4525 = ~n4407 & ~n4524;
  assign n4526 = ~n4353 & ~n4523;
  assign n4527 = x1 & ~n4526;
  assign n4528 = ~n4525 & n4527;
  assign n4529 = ~x1 & n4408;
  assign n4530 = n4407 & n4529;
  assign n4531 = ~n4528 & ~n4530;
  assign n4520 = n4386 ^ n4383;
  assign n4521 = n4390 & ~n4520;
  assign n4522 = n4521 ^ n4389;
  assign n4532 = n4531 ^ n4522;
  assign n4517 = n4372 ^ n4369;
  assign n4518 = n4376 & ~n4517;
  assign n4519 = n4518 ^ n4375;
  assign n4533 = n4532 ^ n4519;
  assign n4514 = n4329 ^ n4295;
  assign n4515 = ~n4330 & n4514;
  assign n4516 = n4515 ^ n4295;
  assign n4534 = n4533 ^ n4516;
  assign n4511 = n4361 ^ n4339;
  assign n4512 = ~n4362 & n4511;
  assign n4513 = n4512 ^ n4342;
  assign n4535 = n4534 ^ n4513;
  assign n4586 = n4585 ^ n4535;
  assign n4508 = n4331 ^ n4289;
  assign n4509 = n4332 & n4508;
  assign n4510 = n4509 ^ n4292;
  assign n4587 = n4586 ^ n4510;
  assign n4499 = x1 & n4408;
  assign n4500 = n4499 ^ x2;
  assign n4501 = x51 & n4500;
  assign n4498 = x3 & x50;
  assign n4502 = n4501 ^ n4498;
  assign n4494 = x18 & x35;
  assign n4493 = x17 & x36;
  assign n4495 = n4494 ^ n4493;
  assign n4492 = x4 & x49;
  assign n4496 = n4495 ^ n4492;
  assign n4489 = x21 & x32;
  assign n4488 = x20 & x33;
  assign n4490 = n4489 ^ n4488;
  assign n4487 = x19 & x34;
  assign n4491 = n4490 ^ n4487;
  assign n4497 = n4496 ^ n4491;
  assign n4503 = n4502 ^ n4497;
  assign n4484 = n4425 ^ n4417;
  assign n4485 = n4426 & ~n4484;
  assign n4486 = n4485 ^ n4420;
  assign n4504 = n4503 ^ n4486;
  assign n4479 = x15 & x38;
  assign n4478 = x7 & x46;
  assign n4480 = n4479 ^ n4478;
  assign n4477 = x6 & x47;
  assign n4481 = n4480 ^ n4477;
  assign n4474 = x16 & x37;
  assign n4473 = x5 & x48;
  assign n4475 = n4474 ^ n4473;
  assign n4472 = x0 & x53;
  assign n4476 = n4475 ^ n4472;
  assign n4482 = n4481 ^ n4476;
  assign n4469 = x14 & x39;
  assign n4468 = x9 & x44;
  assign n4470 = n4469 ^ n4468;
  assign n4467 = x8 & x45;
  assign n4471 = n4470 ^ n4467;
  assign n4483 = n4482 ^ n4471;
  assign n4505 = n4504 ^ n4483;
  assign n4460 = x13 & x40;
  assign n4459 = x12 & x41;
  assign n4461 = n4460 ^ n4459;
  assign n4458 = x10 & x43;
  assign n4462 = n4461 ^ n4458;
  assign n4455 = x24 & x29;
  assign n4454 = x23 & x30;
  assign n4456 = n4455 ^ n4454;
  assign n4453 = x22 & x31;
  assign n4457 = n4456 ^ n4453;
  assign n4463 = n4462 ^ n4457;
  assign n4450 = x26 & x27;
  assign n4449 = x25 & x28;
  assign n4451 = n4450 ^ n4449;
  assign n4448 = x11 & x42;
  assign n4452 = n4451 ^ n4448;
  assign n4464 = n4463 ^ n4452;
  assign n4445 = n4404 ^ n4401;
  assign n4446 = ~n4413 & n4445;
  assign n4447 = n4446 ^ n4401;
  assign n4465 = n4464 ^ n4447;
  assign n4442 = n4380 ^ n4377;
  assign n4443 = n4392 & ~n4442;
  assign n4444 = n4443 ^ n4391;
  assign n4466 = n4465 ^ n4444;
  assign n4506 = n4505 ^ n4466;
  assign n4439 = n4393 ^ n4363;
  assign n4440 = n4394 & n4439;
  assign n4441 = n4440 ^ n4366;
  assign n4507 = n4506 ^ n4441;
  assign n4588 = n4587 ^ n4507;
  assign n4436 = n4429 ^ n4336;
  assign n4437 = ~n4430 & ~n4436;
  assign n4438 = n4437 ^ n4336;
  assign n4589 = n4588 ^ n4438;
  assign n4608 = n4607 ^ n4589;
  assign n4767 = ~n4280 & ~n4593;
  assign n4768 = n4589 & ~n4591;
  assign n4769 = ~n4590 & ~n4768;
  assign n4770 = ~n4767 & n4769;
  assign n4771 = ~n4589 & ~n4592;
  assign n4772 = ~n4280 & ~n4771;
  assign n4773 = n4589 & ~n4593;
  assign n4774 = ~n4594 & ~n4773;
  assign n4775 = ~n4772 & n4774;
  assign n4776 = ~n4770 & ~n4775;
  assign n4755 = x27 & x52;
  assign n4756 = x1 & n4755;
  assign n4753 = x1 & x53;
  assign n4752 = x26 & x28;
  assign n4754 = n4753 ^ n4752;
  assign n4757 = n4756 ^ n4754;
  assign n4751 = x0 & x54;
  assign n4758 = n4757 ^ n4751;
  assign n4747 = x22 & x32;
  assign n4746 = x21 & x33;
  assign n4748 = n4747 ^ n4746;
  assign n4745 = x19 & x35;
  assign n4749 = n4748 ^ n4745;
  assign n4742 = x25 & x29;
  assign n4741 = x24 & x30;
  assign n4743 = n4742 ^ n4741;
  assign n4740 = x23 & x31;
  assign n4744 = n4743 ^ n4740;
  assign n4750 = n4749 ^ n4744;
  assign n4759 = n4758 ^ n4750;
  assign n4737 = n4551 ^ n4541;
  assign n4738 = n4563 & ~n4737;
  assign n4739 = n4738 ^ n4562;
  assign n4760 = n4759 ^ n4739;
  assign n4734 = n4578 ^ n4575;
  assign n4735 = ~n4582 & ~n4734;
  assign n4736 = n4735 ^ n4581;
  assign n4761 = n4760 ^ n4736;
  assign n4731 = n4516 ^ n4513;
  assign n4732 = n4534 & n4731;
  assign n4733 = n4732 ^ n4513;
  assign n4762 = n4761 ^ n4733;
  assign n4728 = n4583 ^ n4538;
  assign n4729 = n4584 & n4728;
  assign n4730 = n4729 ^ n4538;
  assign n4763 = n4762 ^ n4730;
  assign n4719 = n4557 ^ n4554;
  assign n4720 = n4561 & ~n4719;
  assign n4721 = n4720 ^ n4560;
  assign n4716 = n4546 ^ n4543;
  assign n4717 = n4550 & ~n4716;
  assign n4718 = n4717 ^ n4549;
  assign n4722 = n4721 ^ n4718;
  assign n4713 = n4570 ^ n4567;
  assign n4714 = n4574 & ~n4713;
  assign n4715 = n4714 ^ n4573;
  assign n4723 = n4722 ^ n4715;
  assign n4706 = n4493 ^ n4492;
  assign n4707 = n4495 & ~n4706;
  assign n4708 = n4707 ^ n4494;
  assign n4703 = n4454 ^ n4453;
  assign n4704 = n4456 & ~n4703;
  assign n4705 = n4704 ^ n4455;
  assign n4709 = n4708 ^ n4705;
  assign n4700 = n4488 ^ n4487;
  assign n4701 = n4490 & ~n4700;
  assign n4702 = n4701 ^ n4489;
  assign n4710 = n4709 ^ n4702;
  assign n4697 = n4476 ^ n4471;
  assign n4698 = n4482 & ~n4697;
  assign n4699 = n4698 ^ n4481;
  assign n4711 = n4710 ^ n4699;
  assign n4692 = n4449 ^ n4448;
  assign n4693 = n4451 & ~n4692;
  assign n4694 = n4693 ^ n4450;
  assign n4689 = n4478 ^ n4477;
  assign n4690 = n4480 & ~n4689;
  assign n4691 = n4690 ^ n4479;
  assign n4695 = n4694 ^ n4691;
  assign n4686 = n4473 ^ n4472;
  assign n4687 = n4475 & ~n4686;
  assign n4688 = n4687 ^ n4474;
  assign n4696 = n4695 ^ n4688;
  assign n4712 = n4711 ^ n4696;
  assign n4724 = n4723 ^ n4712;
  assign n4683 = n4503 ^ n4483;
  assign n4684 = n4504 & ~n4683;
  assign n4685 = n4684 ^ n4486;
  assign n4725 = n4724 ^ n4685;
  assign n4674 = x14 & x40;
  assign n4673 = x10 & x44;
  assign n4675 = n4674 ^ n4673;
  assign n4672 = x9 & x45;
  assign n4676 = n4675 ^ n4672;
  assign n4669 = x15 & x39;
  assign n4668 = x8 & x46;
  assign n4670 = n4669 ^ n4668;
  assign n4667 = x7 & x47;
  assign n4671 = n4670 ^ n4667;
  assign n4677 = n4676 ^ n4671;
  assign n4664 = x4 & x50;
  assign n4663 = x3 & x51;
  assign n4665 = n4664 ^ n4663;
  assign n4662 = x2 & x52;
  assign n4666 = n4665 ^ n4662;
  assign n4678 = n4677 ^ n4666;
  assign n4657 = x17 & x37;
  assign n4656 = x16 & x38;
  assign n4658 = n4657 ^ n4656;
  assign n4655 = x6 & x48;
  assign n4659 = n4658 ^ n4655;
  assign n4652 = x13 & x41;
  assign n4651 = x12 & x42;
  assign n4653 = n4652 ^ n4651;
  assign n4650 = x11 & x43;
  assign n4654 = n4653 ^ n4650;
  assign n4660 = n4659 ^ n4654;
  assign n4647 = x20 & x34;
  assign n4646 = x18 & x36;
  assign n4648 = n4647 ^ n4646;
  assign n4645 = x5 & x49;
  assign n4649 = n4648 ^ n4645;
  assign n4661 = n4660 ^ n4649;
  assign n4679 = n4678 ^ n4661;
  assign n4642 = n4522 ^ n4519;
  assign n4643 = ~n4532 & ~n4642;
  assign n4644 = n4643 ^ n4531;
  assign n4680 = n4679 ^ n4644;
  assign n4635 = n4459 ^ n4458;
  assign n4636 = n4461 & ~n4635;
  assign n4637 = n4636 ^ n4460;
  assign n4632 = n4468 ^ n4467;
  assign n4633 = n4470 & ~n4632;
  assign n4634 = n4633 ^ n4469;
  assign n4638 = n4637 ^ n4634;
  assign n4627 = x2 & n4498;
  assign n4628 = ~n4499 & ~n4627;
  assign n4629 = ~x2 & ~n4498;
  assign n4630 = x51 & ~n4629;
  assign n4631 = ~n4628 & n4630;
  assign n4639 = n4638 ^ n4631;
  assign n4624 = n4457 ^ n4452;
  assign n4625 = n4463 & ~n4624;
  assign n4626 = n4625 ^ n4462;
  assign n4640 = n4639 ^ n4626;
  assign n4621 = n4502 ^ n4496;
  assign n4622 = ~n4497 & n4621;
  assign n4623 = n4622 ^ n4502;
  assign n4641 = n4640 ^ n4623;
  assign n4681 = n4680 ^ n4641;
  assign n4618 = n4464 ^ n4444;
  assign n4619 = n4465 & ~n4618;
  assign n4620 = n4619 ^ n4447;
  assign n4682 = n4681 ^ n4620;
  assign n4726 = n4725 ^ n4682;
  assign n4615 = n4505 ^ n4441;
  assign n4616 = ~n4506 & n4615;
  assign n4617 = n4616 ^ n4441;
  assign n4727 = n4726 ^ n4617;
  assign n4764 = n4763 ^ n4727;
  assign n4612 = n4535 ^ n4510;
  assign n4613 = ~n4586 & n4612;
  assign n4614 = n4613 ^ n4585;
  assign n4765 = n4764 ^ n4614;
  assign n4609 = n4587 ^ n4438;
  assign n4610 = n4588 & ~n4609;
  assign n4611 = n4610 ^ n4438;
  assign n4766 = n4765 ^ n4611;
  assign n4777 = n4776 ^ n4766;
  assign n4926 = x26 & x53;
  assign n4927 = x1 & n4926;
  assign n4928 = x28 & ~n4927;
  assign n4925 = x1 & x54;
  assign n4929 = n4928 ^ n4925;
  assign n4922 = n4651 ^ n4650;
  assign n4923 = n4653 & ~n4922;
  assign n4924 = n4923 ^ n4652;
  assign n4930 = n4929 ^ n4924;
  assign n4919 = n4691 ^ n4688;
  assign n4920 = n4695 & ~n4919;
  assign n4921 = n4920 ^ n4694;
  assign n4931 = n4930 ^ n4921;
  assign n4916 = n4634 ^ n4631;
  assign n4917 = n4638 & ~n4916;
  assign n4918 = n4917 ^ n4637;
  assign n4932 = n4931 ^ n4918;
  assign n4909 = x18 & x37;
  assign n4910 = n4909 ^ n2367;
  assign n4908 = x5 & x50;
  assign n4911 = n4910 ^ n4908;
  assign n4905 = n4668 ^ n4667;
  assign n4906 = n4670 & ~n4905;
  assign n4907 = n4906 ^ n4669;
  assign n4912 = n4911 ^ n4907;
  assign n4902 = n4754 ^ n4751;
  assign n4903 = n4757 & ~n4902;
  assign n4904 = n4903 ^ n4756;
  assign n4913 = n4912 ^ n4904;
  assign n4897 = n4663 ^ n4662;
  assign n4898 = n4665 & ~n4897;
  assign n4899 = n4898 ^ n4664;
  assign n4894 = n4646 ^ n4645;
  assign n4895 = n4648 & ~n4894;
  assign n4896 = n4895 ^ n4647;
  assign n4900 = n4899 ^ n4896;
  assign n4891 = n4673 ^ n4672;
  assign n4892 = n4675 & ~n4891;
  assign n4893 = n4892 ^ n4674;
  assign n4901 = n4900 ^ n4893;
  assign n4914 = n4913 ^ n4901;
  assign n4888 = n4758 ^ n4749;
  assign n4889 = ~n4750 & n4888;
  assign n4890 = n4889 ^ n4758;
  assign n4915 = n4914 ^ n4890;
  assign n4933 = n4932 ^ n4915;
  assign n4885 = n4678 ^ n4644;
  assign n4886 = ~n4679 & ~n4885;
  assign n4887 = n4886 ^ n4644;
  assign n4934 = n4933 ^ n4887;
  assign n4876 = x22 & x33;
  assign n4875 = x21 & x34;
  assign n4877 = n4876 ^ n4875;
  assign n4874 = x20 & x35;
  assign n4878 = n4877 ^ n4874;
  assign n4871 = x25 & x30;
  assign n4870 = x24 & x31;
  assign n4872 = n4871 ^ n4870;
  assign n4869 = x23 & x32;
  assign n4873 = n4872 ^ n4869;
  assign n4879 = n4878 ^ n4873;
  assign n4866 = x4 & x51;
  assign n4865 = x2 & x53;
  assign n4867 = n4866 ^ n4865;
  assign n4864 = x0 & x55;
  assign n4868 = n4867 ^ n4864;
  assign n4880 = n4879 ^ n4868;
  assign n4859 = x27 & x28;
  assign n4858 = x26 & x29;
  assign n4860 = n4859 ^ n4858;
  assign n4857 = x12 & x43;
  assign n4861 = n4860 ^ n4857;
  assign n4854 = x13 & x42;
  assign n4853 = x11 & x44;
  assign n4855 = n4854 ^ n4853;
  assign n4852 = x10 & x45;
  assign n4856 = n4855 ^ n4852;
  assign n4862 = n4861 ^ n4856;
  assign n4849 = x16 & x39;
  assign n4848 = x8 & x47;
  assign n4850 = n4849 ^ n4848;
  assign n4847 = x7 & x48;
  assign n4851 = n4850 ^ n4847;
  assign n4863 = n4862 ^ n4851;
  assign n4881 = n4880 ^ n4863;
  assign n4844 = n4718 ^ n4715;
  assign n4845 = n4722 & ~n4844;
  assign n4846 = n4845 ^ n4721;
  assign n4882 = n4881 ^ n4846;
  assign n4837 = n4746 ^ n4745;
  assign n4838 = n4748 & ~n4837;
  assign n4839 = n4838 ^ n4747;
  assign n4834 = n4656 ^ n4655;
  assign n4835 = n4658 & ~n4834;
  assign n4836 = n4835 ^ n4657;
  assign n4840 = n4839 ^ n4836;
  assign n4831 = n4741 ^ n4740;
  assign n4832 = n4743 & ~n4831;
  assign n4833 = n4832 ^ n4742;
  assign n4841 = n4840 ^ n4833;
  assign n4828 = n4654 ^ n4649;
  assign n4829 = n4660 & ~n4828;
  assign n4830 = n4829 ^ n4659;
  assign n4842 = n4841 ^ n4830;
  assign n4825 = n4671 ^ n4666;
  assign n4826 = n4677 & ~n4825;
  assign n4827 = n4826 ^ n4676;
  assign n4843 = n4842 ^ n4827;
  assign n4883 = n4882 ^ n4843;
  assign n4822 = n4739 ^ n4736;
  assign n4823 = ~n4760 & ~n4822;
  assign n4824 = n4823 ^ n4736;
  assign n4884 = n4883 ^ n4824;
  assign n4935 = n4934 ^ n4884;
  assign n4819 = n4733 ^ n4730;
  assign n4820 = n4762 & ~n4819;
  assign n4821 = n4820 ^ n4730;
  assign n4936 = n4935 ^ n4821;
  assign n4809 = x17 & x38;
  assign n4808 = x6 & x49;
  assign n4810 = n4809 ^ n4808;
  assign n4807 = x3 & x52;
  assign n4811 = n4810 ^ n4807;
  assign n4804 = x15 & x40;
  assign n4803 = x14 & x41;
  assign n4805 = n4804 ^ n4803;
  assign n4802 = x9 & x46;
  assign n4806 = n4805 ^ n4802;
  assign n4812 = n4811 ^ n4806;
  assign n4799 = n4705 ^ n4702;
  assign n4800 = n4709 & ~n4799;
  assign n4801 = n4800 ^ n4708;
  assign n4813 = n4812 ^ n4801;
  assign n4796 = n4710 ^ n4696;
  assign n4797 = n4711 & ~n4796;
  assign n4798 = n4797 ^ n4699;
  assign n4814 = n4813 ^ n4798;
  assign n4793 = n4626 ^ n4623;
  assign n4794 = ~n4640 & n4793;
  assign n4795 = n4794 ^ n4623;
  assign n4815 = n4814 ^ n4795;
  assign n4790 = n4680 ^ n4620;
  assign n4791 = n4681 & ~n4790;
  assign n4792 = n4791 ^ n4620;
  assign n4816 = n4815 ^ n4792;
  assign n4787 = n4723 ^ n4685;
  assign n4788 = ~n4724 & n4787;
  assign n4789 = n4788 ^ n4685;
  assign n4817 = n4816 ^ n4789;
  assign n4784 = n4725 ^ n4617;
  assign n4785 = n4726 & n4784;
  assign n4786 = n4785 ^ n4617;
  assign n4818 = n4817 ^ n4786;
  assign n4937 = n4936 ^ n4818;
  assign n4781 = n4763 ^ n4614;
  assign n4782 = n4764 & n4781;
  assign n4783 = n4782 ^ n4614;
  assign n4938 = n4937 ^ n4783;
  assign n4778 = n4776 ^ n4611;
  assign n4779 = n4766 & ~n4778;
  assign n4780 = n4779 ^ n4776;
  assign n4939 = n4938 ^ n4780;
  assign n5097 = n4808 ^ n4807;
  assign n5098 = n4810 & ~n5097;
  assign n5099 = n5098 ^ n4809;
  assign n5094 = n4875 ^ n4874;
  assign n5095 = n4877 & ~n5094;
  assign n5096 = n5095 ^ n4876;
  assign n5100 = n5099 ^ n5096;
  assign n5091 = n4870 ^ n4869;
  assign n5092 = n4872 & ~n5091;
  assign n5093 = n5092 ^ n4871;
  assign n5101 = n5100 ^ n5093;
  assign n5086 = n4853 ^ n4852;
  assign n5087 = n4855 & ~n5086;
  assign n5088 = n5087 ^ n4854;
  assign n5083 = n4858 ^ n4857;
  assign n5084 = n4860 & ~n5083;
  assign n5085 = n5084 ^ n4859;
  assign n5089 = n5088 ^ n5085;
  assign n5081 = x1 & x55;
  assign n5080 = x27 & x29;
  assign n5082 = n5081 ^ n5080;
  assign n5090 = n5089 ^ n5082;
  assign n5102 = n5101 ^ n5090;
  assign n5077 = n4856 ^ n4851;
  assign n5078 = n4862 & ~n5077;
  assign n5079 = n5078 ^ n4861;
  assign n5103 = n5102 ^ n5079;
  assign n5072 = x0 & x56;
  assign n5070 = n1379 ^ x2;
  assign n5071 = x54 & n5070;
  assign n5073 = n5072 ^ n5071;
  assign n5067 = x19 & x37;
  assign n5066 = x4 & x52;
  assign n5068 = n5067 ^ n5066;
  assign n5065 = x3 & x53;
  assign n5069 = n5068 ^ n5065;
  assign n5074 = n5073 ^ n5069;
  assign n5062 = n4848 ^ n4847;
  assign n5063 = n4850 & ~n5062;
  assign n5064 = n5063 ^ n4849;
  assign n5075 = n5074 ^ n5064;
  assign n5056 = x14 & x42;
  assign n5055 = x10 & x46;
  assign n5057 = n5056 ^ n5055;
  assign n5054 = x9 & x47;
  assign n5058 = n5057 ^ n5054;
  assign n5051 = x26 & x30;
  assign n5050 = x25 & x31;
  assign n5052 = n5051 ^ n5050;
  assign n5049 = x24 & x32;
  assign n5053 = n5052 ^ n5049;
  assign n5059 = n5058 ^ n5053;
  assign n5046 = x23 & x33;
  assign n5045 = x22 & x34;
  assign n5047 = n5046 ^ n5045;
  assign n5044 = x20 & x36;
  assign n5048 = n5047 ^ n5044;
  assign n5060 = n5059 ^ n5048;
  assign n5039 = x13 & x43;
  assign n5038 = x12 & x44;
  assign n5040 = n5039 ^ n5038;
  assign n5037 = x11 & x45;
  assign n5041 = n5040 ^ n5037;
  assign n5034 = x16 & x40;
  assign n5033 = x15 & x41;
  assign n5035 = n5034 ^ n5033;
  assign n5032 = x8 & x48;
  assign n5036 = n5035 ^ n5032;
  assign n5042 = n5041 ^ n5036;
  assign n5029 = x17 & x39;
  assign n5028 = x7 & x49;
  assign n5030 = n5029 ^ n5028;
  assign n5027 = x6 & x50;
  assign n5031 = n5030 ^ n5027;
  assign n5043 = n5042 ^ n5031;
  assign n5061 = n5060 ^ n5043;
  assign n5076 = n5075 ^ n5061;
  assign n5104 = n5103 ^ n5076;
  assign n5024 = n4813 ^ n4795;
  assign n5025 = n4814 & ~n5024;
  assign n5026 = n5025 ^ n4798;
  assign n5105 = n5104 ^ n5026;
  assign n5015 = n4909 ^ n4908;
  assign n5016 = n4910 & ~n5015;
  assign n5017 = n5016 ^ n2367;
  assign n5012 = n4865 ^ n4864;
  assign n5013 = n4867 & ~n5012;
  assign n5014 = n5013 ^ n4866;
  assign n5018 = n5017 ^ n5014;
  assign n5009 = n4803 ^ n4802;
  assign n5010 = n4805 & ~n5009;
  assign n5011 = n5010 ^ n4804;
  assign n5019 = n5018 ^ n5011;
  assign n5006 = n4811 ^ n4801;
  assign n5007 = ~n4812 & n5006;
  assign n5008 = n5007 ^ n4801;
  assign n5020 = n5019 ^ n5008;
  assign n5003 = n4930 ^ n4918;
  assign n5004 = n4931 & ~n5003;
  assign n5005 = n5004 ^ n4921;
  assign n5021 = n5020 ^ n5005;
  assign n4998 = n4907 ^ n4904;
  assign n4999 = ~n4912 & n4998;
  assign n5000 = n4999 ^ n4904;
  assign n4995 = n4836 ^ n4833;
  assign n4996 = n4840 & ~n4995;
  assign n4997 = n4996 ^ n4839;
  assign n5001 = n5000 ^ n4997;
  assign n4992 = n4873 ^ n4868;
  assign n4993 = n4879 & ~n4992;
  assign n4994 = n4993 ^ n4878;
  assign n5002 = n5001 ^ n4994;
  assign n5022 = n5021 ^ n5002;
  assign n4989 = n4880 ^ n4846;
  assign n4990 = ~n4881 & n4989;
  assign n4991 = n4990 ^ n4846;
  assign n5023 = n5022 ^ n4991;
  assign n5106 = n5105 ^ n5023;
  assign n4986 = n4815 ^ n4789;
  assign n4987 = n4816 & ~n4986;
  assign n4988 = n4987 ^ n4792;
  assign n5107 = n5106 ^ n4988;
  assign n4970 = x54 & n4924;
  assign n4971 = x28 & x53;
  assign n4972 = x26 & n4971;
  assign n4973 = ~n4970 & ~n4972;
  assign n4974 = x28 & x54;
  assign n4975 = x1 & ~n4974;
  assign n4976 = ~n4973 & n4975;
  assign n4977 = n4925 & ~n4926;
  assign n4978 = x28 & ~n4977;
  assign n4979 = n4924 & n4978;
  assign n4980 = ~n4976 & ~n4979;
  assign n4967 = x21 & x35;
  assign n4966 = x18 & x38;
  assign n4968 = n4967 ^ n4966;
  assign n4965 = x5 & x51;
  assign n4969 = n4968 ^ n4965;
  assign n4981 = n4980 ^ n4969;
  assign n4962 = n4896 ^ n4893;
  assign n4963 = n4900 & ~n4962;
  assign n4964 = n4963 ^ n4899;
  assign n4982 = n4981 ^ n4964;
  assign n4958 = n4830 ^ n4827;
  assign n4959 = n4842 & ~n4958;
  assign n4960 = n4959 ^ n4841;
  assign n4955 = n4901 ^ n4890;
  assign n4956 = n4914 & ~n4955;
  assign n4957 = n4956 ^ n4913;
  assign n4961 = n4960 ^ n4957;
  assign n4983 = n4982 ^ n4961;
  assign n4952 = n4932 ^ n4887;
  assign n4953 = ~n4933 & ~n4952;
  assign n4954 = n4953 ^ n4887;
  assign n4984 = n4983 ^ n4954;
  assign n4949 = n4843 ^ n4824;
  assign n4950 = n4883 & n4949;
  assign n4951 = n4950 ^ n4882;
  assign n4985 = n4984 ^ n4951;
  assign n5108 = n5107 ^ n4985;
  assign n4946 = n4934 ^ n4821;
  assign n4947 = ~n4935 & n4946;
  assign n4948 = n4947 ^ n4821;
  assign n5109 = n5108 ^ n4948;
  assign n4943 = n4936 ^ n4786;
  assign n4944 = ~n4818 & ~n4943;
  assign n4945 = n4944 ^ n4936;
  assign n5110 = n5109 ^ n4945;
  assign n4940 = n4783 ^ n4780;
  assign n4941 = n4938 & ~n4940;
  assign n4942 = n4941 ^ n4780;
  assign n5111 = n5110 ^ n4942;
  assign n5266 = x4 & x53;
  assign n5265 = x3 & x54;
  assign n5267 = n5266 ^ n5265;
  assign n5264 = x2 & x55;
  assign n5268 = n5267 ^ n5264;
  assign n5261 = x19 & x38;
  assign n5262 = n5261 ^ n2445;
  assign n5260 = x5 & x52;
  assign n5263 = n5262 ^ n5260;
  assign n5269 = n5268 ^ n5263;
  assign n5257 = x15 & x42;
  assign n5256 = x10 & x47;
  assign n5258 = n5257 ^ n5256;
  assign n5255 = x9 & x48;
  assign n5259 = n5258 ^ n5255;
  assign n5270 = n5269 ^ n5259;
  assign n5250 = x14 & x43;
  assign n5249 = x13 & x44;
  assign n5251 = n5250 ^ n5249;
  assign n5248 = x11 & x46;
  assign n5252 = n5251 ^ n5248;
  assign n5245 = x18 & x39;
  assign n5244 = x17 & x40;
  assign n5246 = n5245 ^ n5244;
  assign n5243 = x6 & x51;
  assign n5247 = n5246 ^ n5243;
  assign n5253 = n5252 ^ n5247;
  assign n5240 = x28 & x29;
  assign n5239 = x27 & x30;
  assign n5241 = n5240 ^ n5239;
  assign n5238 = x12 & x45;
  assign n5242 = n5241 ^ n5238;
  assign n5254 = n5253 ^ n5242;
  assign n5271 = n5270 ^ n5254;
  assign n5235 = n4997 ^ n4994;
  assign n5236 = n5001 & ~n5235;
  assign n5237 = n5236 ^ n5000;
  assign n5272 = n5271 ^ n5237;
  assign n5232 = n4982 ^ n4960;
  assign n5233 = ~n4961 & ~n5232;
  assign n5234 = n5233 ^ n4982;
  assign n5273 = n5272 ^ n5234;
  assign n5225 = x26 & x31;
  assign n5224 = x25 & x32;
  assign n5226 = n5225 ^ n5224;
  assign n5223 = x24 & x33;
  assign n5227 = n5226 ^ n5223;
  assign n5220 = x23 & x34;
  assign n5219 = x22 & x35;
  assign n5221 = n5220 ^ n5219;
  assign n5218 = x21 & x36;
  assign n5222 = n5221 ^ n5218;
  assign n5228 = n5227 ^ n5222;
  assign n5215 = x16 & x41;
  assign n5214 = x8 & x49;
  assign n5216 = n5215 ^ n5214;
  assign n5213 = x7 & x50;
  assign n5217 = n5216 ^ n5213;
  assign n5229 = n5228 ^ n5217;
  assign n5210 = n4969 ^ n4964;
  assign n5211 = ~n4981 & ~n5210;
  assign n5212 = n5211 ^ n4980;
  assign n5230 = n5229 ^ n5212;
  assign n5205 = n4966 ^ n4965;
  assign n5206 = n4968 & ~n5205;
  assign n5207 = n5206 ^ n4967;
  assign n5202 = n5038 ^ n5037;
  assign n5203 = n5040 & ~n5202;
  assign n5204 = n5203 ^ n5039;
  assign n5208 = n5207 ^ n5204;
  assign n5199 = n5055 ^ n5054;
  assign n5200 = n5057 & ~n5199;
  assign n5201 = n5200 ^ n5056;
  assign n5209 = n5208 ^ n5201;
  assign n5231 = n5230 ^ n5209;
  assign n5274 = n5273 ^ n5231;
  assign n5190 = n5050 ^ n5049;
  assign n5191 = n5052 & ~n5190;
  assign n5192 = n5191 ^ n5051;
  assign n5187 = n5033 ^ n5032;
  assign n5188 = n5035 & ~n5187;
  assign n5189 = n5188 ^ n5034;
  assign n5193 = n5192 ^ n5189;
  assign n5184 = n5028 ^ n5027;
  assign n5185 = n5030 & ~n5184;
  assign n5186 = n5185 ^ n5029;
  assign n5194 = n5193 ^ n5186;
  assign n5180 = ~x2 & ~n1379;
  assign n5181 = x54 & ~n5180;
  assign n5179 = n5071 & ~n5072;
  assign n5182 = n5181 ^ n5179;
  assign n5175 = n5066 ^ n5065;
  assign n5176 = n5068 & ~n5175;
  assign n5177 = n5176 ^ n5067;
  assign n5172 = n5045 ^ n5044;
  assign n5173 = n5047 & ~n5172;
  assign n5174 = n5173 ^ n5046;
  assign n5178 = n5177 ^ n5174;
  assign n5183 = n5182 ^ n5178;
  assign n5195 = n5194 ^ n5183;
  assign n5169 = n5036 ^ n5031;
  assign n5170 = n5042 & ~n5169;
  assign n5171 = n5170 ^ n5041;
  assign n5196 = n5195 ^ n5171;
  assign n5166 = n5075 ^ n5060;
  assign n5167 = ~n5061 & n5166;
  assign n5168 = n5167 ^ n5075;
  assign n5197 = n5196 ^ n5168;
  assign n5161 = n5069 ^ n5064;
  assign n5162 = n5074 & ~n5161;
  assign n5163 = n5162 ^ n5073;
  assign n5158 = n5085 ^ n5082;
  assign n5159 = n5089 & ~n5158;
  assign n5160 = n5159 ^ n5088;
  assign n5164 = n5163 ^ n5160;
  assign n5155 = n5053 ^ n5048;
  assign n5156 = n5059 & ~n5155;
  assign n5157 = n5156 ^ n5058;
  assign n5165 = n5164 ^ n5157;
  assign n5198 = n5197 ^ n5165;
  assign n5275 = n5274 ^ n5198;
  assign n5152 = n4983 ^ n4951;
  assign n5153 = n4984 & n5152;
  assign n5154 = n5153 ^ n4954;
  assign n5276 = n5275 ^ n5154;
  assign n5149 = n5105 ^ n4988;
  assign n5150 = ~n5106 & n5149;
  assign n5151 = n5150 ^ n4988;
  assign n5277 = n5276 ^ n5151;
  assign n5140 = n5096 ^ n5093;
  assign n5141 = n5100 & ~n5140;
  assign n5142 = n5141 ^ n5099;
  assign n5137 = n5014 ^ n5011;
  assign n5138 = n5018 & ~n5137;
  assign n5139 = n5138 ^ n5017;
  assign n5143 = n5142 ^ n5139;
  assign n5133 = x27 & x55;
  assign n5134 = x1 & n5133;
  assign n5135 = x29 & ~n5134;
  assign n5131 = x0 & x57;
  assign n5130 = x1 & x56;
  assign n5132 = n5131 ^ n5130;
  assign n5136 = n5135 ^ n5132;
  assign n5144 = n5143 ^ n5136;
  assign n5127 = n5090 ^ n5079;
  assign n5128 = n5102 & ~n5127;
  assign n5129 = n5128 ^ n5101;
  assign n5145 = n5144 ^ n5129;
  assign n5124 = n5008 ^ n5005;
  assign n5125 = ~n5020 & n5124;
  assign n5126 = n5125 ^ n5005;
  assign n5146 = n5145 ^ n5126;
  assign n5121 = n5002 ^ n4991;
  assign n5122 = n5022 & ~n5121;
  assign n5123 = n5122 ^ n5021;
  assign n5147 = n5146 ^ n5123;
  assign n5118 = n5103 ^ n5026;
  assign n5119 = ~n5104 & n5118;
  assign n5120 = n5119 ^ n5026;
  assign n5148 = n5147 ^ n5120;
  assign n5278 = n5277 ^ n5148;
  assign n5115 = n5107 ^ n4948;
  assign n5116 = ~n5108 & ~n5115;
  assign n5117 = n5116 ^ n4948;
  assign n5279 = n5278 ^ n5117;
  assign n5112 = n4945 ^ n4942;
  assign n5113 = ~n5110 & n5112;
  assign n5114 = n5113 ^ n4942;
  assign n5280 = n5279 ^ n5114;
  assign n5450 = n5148 & ~n5276;
  assign n5451 = n5114 & ~n5450;
  assign n5452 = ~n5117 & n5151;
  assign n5453 = ~n5148 & n5276;
  assign n5454 = ~n5452 & n5453;
  assign n5455 = n5117 & ~n5151;
  assign n5456 = ~n5454 & ~n5455;
  assign n5457 = n5451 & ~n5456;
  assign n5458 = n5450 & ~n5455;
  assign n5459 = n5452 & ~n5453;
  assign n5460 = ~n5458 & ~n5459;
  assign n5461 = ~n5114 & ~n5460;
  assign n5462 = n5151 ^ n5117;
  assign n5463 = n5276 ^ n5148;
  assign n5464 = n5277 & n5463;
  assign n5465 = n5462 & n5464;
  assign n5466 = ~n5461 & ~n5465;
  assign n5467 = ~n5457 & n5466;
  assign n5437 = x18 & x40;
  assign n5436 = x8 & x50;
  assign n5438 = n5437 ^ n5436;
  assign n5435 = x7 & x51;
  assign n5439 = n5438 ^ n5435;
  assign n5432 = x27 & x31;
  assign n5431 = x26 & x32;
  assign n5433 = n5432 ^ n5431;
  assign n5430 = x25 & x33;
  assign n5434 = n5433 ^ n5430;
  assign n5440 = n5439 ^ n5434;
  assign n5427 = x24 & x34;
  assign n5426 = x23 & x35;
  assign n5428 = n5427 ^ n5426;
  assign n5425 = x22 & x36;
  assign n5429 = n5428 ^ n5425;
  assign n5441 = n5440 ^ n5429;
  assign n5422 = n5160 ^ n5157;
  assign n5423 = n5164 & ~n5422;
  assign n5424 = n5423 ^ n5163;
  assign n5442 = n5441 ^ n5424;
  assign n5417 = x17 & x41;
  assign n5416 = x16 & x42;
  assign n5418 = n5417 ^ n5416;
  assign n5415 = x9 & x49;
  assign n5419 = n5418 ^ n5415;
  assign n5412 = x21 & x37;
  assign n5413 = n5412 ^ n2628;
  assign n5411 = x5 & x53;
  assign n5414 = n5413 ^ n5411;
  assign n5420 = n5419 ^ n5414;
  assign n5408 = x4 & x54;
  assign n5407 = x2 & x56;
  assign n5409 = n5408 ^ n5407;
  assign n5406 = x0 & x58;
  assign n5410 = n5409 ^ n5406;
  assign n5421 = n5420 ^ n5410;
  assign n5443 = n5442 ^ n5421;
  assign n5393 = n1493 & n5133;
  assign n5394 = ~n5130 & ~n5393;
  assign n5395 = ~x29 & n5131;
  assign n5396 = x56 & ~n5395;
  assign n5397 = ~n5394 & ~n5396;
  assign n5398 = n5130 & ~n5133;
  assign n5399 = x29 & x57;
  assign n5400 = x0 & n5399;
  assign n5401 = ~n5398 & n5400;
  assign n5402 = ~n5397 & ~n5401;
  assign n5389 = n5214 ^ n5213;
  assign n5390 = n5216 & ~n5389;
  assign n5391 = n5390 ^ n5215;
  assign n5386 = n5244 ^ n5243;
  assign n5387 = n5246 & ~n5386;
  assign n5388 = n5387 ^ n5245;
  assign n5392 = n5391 ^ n5388;
  assign n5403 = n5402 ^ n5392;
  assign n5381 = x19 & x39;
  assign n5380 = x6 & x52;
  assign n5382 = n5381 ^ n5380;
  assign n5379 = x3 & x55;
  assign n5383 = n5382 ^ n5379;
  assign n5376 = x15 & x43;
  assign n5375 = x11 & x47;
  assign n5377 = n5376 ^ n5375;
  assign n5374 = x10 & x48;
  assign n5378 = n5377 ^ n5374;
  assign n5384 = n5383 ^ n5378;
  assign n5371 = x14 & x44;
  assign n5370 = x13 & x45;
  assign n5372 = n5371 ^ n5370;
  assign n5369 = x12 & x46;
  assign n5373 = n5372 ^ n5369;
  assign n5385 = n5384 ^ n5373;
  assign n5404 = n5403 ^ n5385;
  assign n5366 = n5139 ^ n5136;
  assign n5367 = n5143 & ~n5366;
  assign n5368 = n5367 ^ n5142;
  assign n5405 = n5404 ^ n5368;
  assign n5444 = n5443 ^ n5405;
  assign n5363 = n5129 ^ n5126;
  assign n5364 = ~n5145 & n5363;
  assign n5365 = n5364 ^ n5126;
  assign n5445 = n5444 ^ n5365;
  assign n5354 = x29 & x56;
  assign n5355 = n5354 ^ x57;
  assign n5356 = x1 & n5355;
  assign n5353 = x28 & x30;
  assign n5357 = n5356 ^ n5353;
  assign n5350 = n5239 ^ n5238;
  assign n5351 = n5241 & ~n5350;
  assign n5352 = n5351 ^ n5240;
  assign n5358 = n5357 ^ n5352;
  assign n5347 = n5263 ^ n5259;
  assign n5348 = n5269 & ~n5347;
  assign n5349 = n5348 ^ n5268;
  assign n5359 = n5358 ^ n5349;
  assign n5344 = n5247 ^ n5242;
  assign n5345 = n5253 & ~n5344;
  assign n5346 = n5345 ^ n5252;
  assign n5360 = n5359 ^ n5346;
  assign n5337 = n5265 ^ n5264;
  assign n5338 = n5267 & ~n5337;
  assign n5339 = n5338 ^ n5266;
  assign n5334 = n5249 ^ n5248;
  assign n5335 = n5251 & ~n5334;
  assign n5336 = n5335 ^ n5250;
  assign n5340 = n5339 ^ n5336;
  assign n5331 = n5261 ^ n5260;
  assign n5332 = n5262 & ~n5331;
  assign n5333 = n5332 ^ n2445;
  assign n5341 = n5340 ^ n5333;
  assign n5328 = n5222 ^ n5217;
  assign n5329 = n5228 & ~n5328;
  assign n5330 = n5329 ^ n5227;
  assign n5342 = n5341 ^ n5330;
  assign n5323 = n5219 ^ n5218;
  assign n5324 = n5221 & ~n5323;
  assign n5325 = n5324 ^ n5220;
  assign n5320 = n5224 ^ n5223;
  assign n5321 = n5226 & ~n5320;
  assign n5322 = n5321 ^ n5225;
  assign n5326 = n5325 ^ n5322;
  assign n5317 = n5256 ^ n5255;
  assign n5318 = n5258 & ~n5317;
  assign n5319 = n5318 ^ n5257;
  assign n5327 = n5326 ^ n5319;
  assign n5343 = n5342 ^ n5327;
  assign n5361 = n5360 ^ n5343;
  assign n5314 = n5270 ^ n5237;
  assign n5315 = ~n5271 & n5314;
  assign n5316 = n5315 ^ n5237;
  assign n5362 = n5361 ^ n5316;
  assign n5446 = n5445 ^ n5362;
  assign n5311 = n5146 ^ n5120;
  assign n5312 = n5147 & ~n5311;
  assign n5313 = n5312 ^ n5123;
  assign n5447 = n5446 ^ n5313;
  assign n5302 = n5182 ^ n5174;
  assign n5303 = n5178 & ~n5302;
  assign n5304 = n5303 ^ n5177;
  assign n5299 = n5189 ^ n5186;
  assign n5300 = n5193 & ~n5299;
  assign n5301 = n5300 ^ n5192;
  assign n5305 = n5304 ^ n5301;
  assign n5296 = n5204 ^ n5201;
  assign n5297 = n5208 & ~n5296;
  assign n5298 = n5297 ^ n5207;
  assign n5306 = n5305 ^ n5298;
  assign n5293 = n5183 ^ n5171;
  assign n5294 = n5195 & ~n5293;
  assign n5295 = n5294 ^ n5194;
  assign n5307 = n5306 ^ n5295;
  assign n5290 = n5229 ^ n5209;
  assign n5291 = ~n5230 & ~n5290;
  assign n5292 = n5291 ^ n5212;
  assign n5308 = n5307 ^ n5292;
  assign n5287 = n5196 ^ n5165;
  assign n5288 = n5197 & ~n5287;
  assign n5289 = n5288 ^ n5168;
  assign n5309 = n5308 ^ n5289;
  assign n5284 = n5272 ^ n5231;
  assign n5285 = ~n5273 & n5284;
  assign n5286 = n5285 ^ n5234;
  assign n5310 = n5309 ^ n5286;
  assign n5448 = n5447 ^ n5310;
  assign n5281 = n5274 ^ n5154;
  assign n5282 = ~n5275 & ~n5281;
  assign n5283 = n5282 ^ n5154;
  assign n5449 = n5448 ^ n5283;
  assign n5468 = n5467 ^ n5449;
  assign n5645 = n5449 & ~n5454;
  assign n5646 = n5114 & ~n5645;
  assign n5647 = ~n5449 & ~n5450;
  assign n5648 = ~n5455 & ~n5647;
  assign n5649 = ~n5646 & n5648;
  assign n5650 = ~n5449 & ~n5452;
  assign n5651 = ~n5453 & ~n5650;
  assign n5652 = ~n5451 & n5651;
  assign n5653 = ~n5649 & ~n5652;
  assign n5631 = x14 & x45;
  assign n5630 = x12 & x47;
  assign n5632 = n5631 ^ n5630;
  assign n5629 = x11 & x48;
  assign n5633 = n5632 ^ n5629;
  assign n5626 = x17 & x42;
  assign n5625 = x16 & x43;
  assign n5627 = n5626 ^ n5625;
  assign n5624 = x8 & x51;
  assign n5628 = n5627 ^ n5624;
  assign n5634 = n5633 ^ n5628;
  assign n5621 = x29 & x30;
  assign n5620 = x28 & x31;
  assign n5622 = n5621 ^ n5620;
  assign n5619 = x13 & x46;
  assign n5623 = n5622 ^ n5619;
  assign n5635 = n5634 ^ n5623;
  assign n5616 = n5358 ^ n5346;
  assign n5617 = n5359 & ~n5616;
  assign n5618 = n5617 ^ n5349;
  assign n5636 = n5635 ^ n5618;
  assign n5611 = x19 & x40;
  assign n5610 = x5 & x54;
  assign n5612 = n5611 ^ n5610;
  assign n5609 = x4 & x55;
  assign n5613 = n5612 ^ n5609;
  assign n5606 = n5431 ^ n5430;
  assign n5607 = n5433 & ~n5606;
  assign n5608 = n5607 ^ n5432;
  assign n5614 = n5613 ^ n5608;
  assign n5602 = x28 & n1571;
  assign n5603 = n5602 ^ x2;
  assign n5604 = x57 & n5603;
  assign n5601 = x3 & x56;
  assign n5605 = n5604 ^ n5601;
  assign n5615 = n5614 ^ n5605;
  assign n5637 = n5636 ^ n5615;
  assign n5589 = n5353 ^ x57;
  assign n5590 = n5354 & n5589;
  assign n5591 = ~n5352 & ~n5590;
  assign n5592 = ~n5354 & ~n5589;
  assign n5593 = x1 & ~n5592;
  assign n5594 = ~n5591 & n5593;
  assign n5595 = ~x1 & n5353;
  assign n5596 = n5352 & n5595;
  assign n5597 = ~n5594 & ~n5596;
  assign n5585 = x18 & x41;
  assign n5584 = x7 & x52;
  assign n5586 = n5585 ^ n5584;
  assign n5583 = x6 & x53;
  assign n5587 = n5586 ^ n5583;
  assign n5580 = x15 & x44;
  assign n5579 = x10 & x49;
  assign n5581 = n5580 ^ n5579;
  assign n5578 = x9 & x50;
  assign n5582 = n5581 ^ n5578;
  assign n5588 = n5587 ^ n5582;
  assign n5598 = n5597 ^ n5588;
  assign n5573 = x22 & x37;
  assign n5572 = x21 & x38;
  assign n5574 = n5573 ^ n5572;
  assign n5571 = x20 & x39;
  assign n5575 = n5574 ^ n5571;
  assign n5568 = x27 & x32;
  assign n5567 = x26 & x33;
  assign n5569 = n5568 ^ n5567;
  assign n5566 = x0 & x59;
  assign n5570 = n5569 ^ n5566;
  assign n5576 = n5575 ^ n5570;
  assign n5563 = x25 & x34;
  assign n5562 = x24 & x35;
  assign n5564 = n5563 ^ n5562;
  assign n5561 = x23 & x36;
  assign n5565 = n5564 ^ n5561;
  assign n5577 = n5576 ^ n5565;
  assign n5599 = n5598 ^ n5577;
  assign n5558 = n5301 ^ n5298;
  assign n5559 = n5305 & ~n5558;
  assign n5560 = n5559 ^ n5304;
  assign n5600 = n5599 ^ n5560;
  assign n5638 = n5637 ^ n5600;
  assign n5555 = n5295 ^ n5292;
  assign n5556 = ~n5307 & ~n5555;
  assign n5557 = n5556 ^ n5292;
  assign n5639 = n5638 ^ n5557;
  assign n5548 = n5434 ^ n5429;
  assign n5549 = n5440 & ~n5548;
  assign n5550 = n5549 ^ n5439;
  assign n5545 = n5414 ^ n5410;
  assign n5546 = n5420 & ~n5545;
  assign n5547 = n5546 ^ n5419;
  assign n5551 = n5550 ^ n5547;
  assign n5542 = n5378 ^ n5373;
  assign n5543 = n5384 & ~n5542;
  assign n5544 = n5543 ^ n5383;
  assign n5552 = n5551 ^ n5544;
  assign n5535 = n5407 ^ n5406;
  assign n5536 = n5409 & ~n5535;
  assign n5537 = n5536 ^ n5408;
  assign n5532 = n5380 ^ n5379;
  assign n5533 = n5382 & ~n5532;
  assign n5534 = n5533 ^ n5381;
  assign n5538 = n5537 ^ n5534;
  assign n5529 = n5416 ^ n5415;
  assign n5530 = n5418 & ~n5529;
  assign n5531 = n5530 ^ n5417;
  assign n5539 = n5538 ^ n5531;
  assign n5524 = n5375 ^ n5374;
  assign n5525 = n5377 & ~n5524;
  assign n5526 = n5525 ^ n5376;
  assign n5521 = n5370 ^ n5369;
  assign n5522 = n5372 & ~n5521;
  assign n5523 = n5522 ^ n5371;
  assign n5527 = n5526 ^ n5523;
  assign n5519 = x1 & x58;
  assign n5520 = n5519 ^ x30;
  assign n5528 = n5527 ^ n5520;
  assign n5540 = n5539 ^ n5528;
  assign n5514 = n5436 ^ n5435;
  assign n5515 = n5438 & ~n5514;
  assign n5516 = n5515 ^ n5437;
  assign n5511 = n5426 ^ n5425;
  assign n5512 = n5428 & ~n5511;
  assign n5513 = n5512 ^ n5427;
  assign n5517 = n5516 ^ n5513;
  assign n5508 = n5412 ^ n5411;
  assign n5509 = n5413 & ~n5508;
  assign n5510 = n5509 ^ n2628;
  assign n5518 = n5517 ^ n5510;
  assign n5541 = n5540 ^ n5518;
  assign n5553 = n5552 ^ n5541;
  assign n5505 = n5441 ^ n5421;
  assign n5506 = n5442 & ~n5505;
  assign n5507 = n5506 ^ n5424;
  assign n5554 = n5553 ^ n5507;
  assign n5640 = n5639 ^ n5554;
  assign n5502 = n5289 ^ n5286;
  assign n5503 = ~n5309 & n5502;
  assign n5504 = n5503 ^ n5308;
  assign n5641 = n5640 ^ n5504;
  assign n5493 = n5402 ^ n5391;
  assign n5494 = ~n5392 & ~n5493;
  assign n5495 = n5494 ^ n5402;
  assign n5490 = n5322 ^ n5319;
  assign n5491 = n5326 & ~n5490;
  assign n5492 = n5491 ^ n5325;
  assign n5496 = n5495 ^ n5492;
  assign n5487 = n5336 ^ n5333;
  assign n5488 = n5340 & ~n5487;
  assign n5489 = n5488 ^ n5339;
  assign n5497 = n5496 ^ n5489;
  assign n5484 = n5330 ^ n5327;
  assign n5485 = n5342 & ~n5484;
  assign n5486 = n5485 ^ n5341;
  assign n5498 = n5497 ^ n5486;
  assign n5481 = n5403 ^ n5368;
  assign n5482 = n5404 & ~n5481;
  assign n5483 = n5482 ^ n5368;
  assign n5499 = n5498 ^ n5483;
  assign n5478 = n5360 ^ n5316;
  assign n5479 = ~n5361 & n5478;
  assign n5480 = n5479 ^ n5316;
  assign n5500 = n5499 ^ n5480;
  assign n5475 = n5405 ^ n5365;
  assign n5476 = ~n5444 & n5475;
  assign n5477 = n5476 ^ n5443;
  assign n5501 = n5500 ^ n5477;
  assign n5642 = n5641 ^ n5501;
  assign n5472 = n5445 ^ n5313;
  assign n5473 = n5446 & ~n5472;
  assign n5474 = n5473 ^ n5313;
  assign n5643 = n5642 ^ n5474;
  assign n5469 = n5310 ^ n5283;
  assign n5470 = ~n5448 & n5469;
  assign n5471 = n5470 ^ n5447;
  assign n5644 = n5643 ^ n5471;
  assign n5654 = n5653 ^ n5644;
  assign n5818 = x26 & x34;
  assign n5817 = x25 & x35;
  assign n5819 = n5818 ^ n5817;
  assign n5816 = x24 & x36;
  assign n5820 = n5819 ^ n5816;
  assign n5813 = x21 & x39;
  assign n5812 = x22 & x38;
  assign n5814 = n5813 ^ n5812;
  assign n5811 = x20 & x40;
  assign n5815 = n5814 ^ n5811;
  assign n5821 = n5820 ^ n5815;
  assign n5808 = x4 & x56;
  assign n5807 = x3 & x57;
  assign n5809 = n5808 ^ n5807;
  assign n5806 = x2 & x58;
  assign n5810 = n5809 ^ n5806;
  assign n5822 = n5821 ^ n5810;
  assign n5801 = x17 & x43;
  assign n5800 = x16 & x44;
  assign n5802 = n5801 ^ n5800;
  assign n5799 = x9 & x51;
  assign n5803 = n5802 ^ n5799;
  assign n5796 = x15 & x45;
  assign n5795 = x11 & x49;
  assign n5797 = n5796 ^ n5795;
  assign n5794 = x10 & x50;
  assign n5798 = n5797 ^ n5794;
  assign n5804 = n5803 ^ n5798;
  assign n5791 = n5630 ^ n5629;
  assign n5792 = n5632 & ~n5791;
  assign n5793 = n5792 ^ n5631;
  assign n5805 = n5804 ^ n5793;
  assign n5823 = n5822 ^ n5805;
  assign n5788 = n5492 ^ n5489;
  assign n5789 = ~n5496 & ~n5788;
  assign n5790 = n5789 ^ n5495;
  assign n5824 = n5823 ^ n5790;
  assign n5781 = x58 & n1571;
  assign n5779 = x1 & x59;
  assign n5778 = x29 & x31;
  assign n5780 = n5779 ^ n5778;
  assign n5782 = n5781 ^ n5780;
  assign n5777 = x0 & x60;
  assign n5783 = n5782 ^ n5777;
  assign n5774 = x28 & x32;
  assign n5773 = x27 & x33;
  assign n5775 = n5774 ^ n5773;
  assign n5772 = x23 & x37;
  assign n5776 = n5775 ^ n5772;
  assign n5784 = n5783 ^ n5776;
  assign n5769 = n5523 ^ n5520;
  assign n5770 = n5527 & ~n5769;
  assign n5771 = n5770 ^ n5526;
  assign n5785 = n5784 ^ n5771;
  assign n5764 = x14 & x46;
  assign n5763 = x13 & x47;
  assign n5765 = n5764 ^ n5763;
  assign n5762 = x12 & x48;
  assign n5766 = n5765 ^ n5762;
  assign n5759 = x18 & x42;
  assign n5758 = x8 & x52;
  assign n5760 = n5759 ^ n5758;
  assign n5757 = x7 & x53;
  assign n5761 = n5760 ^ n5757;
  assign n5767 = n5766 ^ n5761;
  assign n5754 = x19 & x41;
  assign n5753 = x6 & x54;
  assign n5755 = n5754 ^ n5753;
  assign n5752 = x5 & x55;
  assign n5756 = n5755 ^ n5752;
  assign n5768 = n5767 ^ n5756;
  assign n5786 = n5785 ^ n5768;
  assign n5749 = n5528 ^ n5518;
  assign n5750 = n5540 & ~n5749;
  assign n5751 = n5750 ^ n5539;
  assign n5787 = n5786 ^ n5751;
  assign n5825 = n5824 ^ n5787;
  assign n5746 = n5486 ^ n5483;
  assign n5747 = n5498 & n5746;
  assign n5748 = n5747 ^ n5483;
  assign n5826 = n5825 ^ n5748;
  assign n5737 = n5572 ^ n5571;
  assign n5738 = n5574 & ~n5737;
  assign n5739 = n5738 ^ n5573;
  assign n5734 = n5610 ^ n5609;
  assign n5735 = n5612 & ~n5734;
  assign n5736 = n5735 ^ n5611;
  assign n5740 = n5739 ^ n5736;
  assign n5731 = n5562 ^ n5561;
  assign n5732 = n5564 & ~n5731;
  assign n5733 = n5732 ^ n5563;
  assign n5741 = n5740 ^ n5733;
  assign n5728 = n5597 ^ n5587;
  assign n5729 = ~n5588 & ~n5728;
  assign n5730 = n5729 ^ n5597;
  assign n5742 = n5741 ^ n5730;
  assign n5723 = n5602 ^ n5601;
  assign n5724 = n5603 & ~n5723;
  assign n5725 = n5724 ^ x2;
  assign n5726 = x57 & n5725;
  assign n5719 = n5579 ^ n5578;
  assign n5720 = n5581 & ~n5719;
  assign n5721 = n5720 ^ n5580;
  assign n5716 = n5567 ^ n5566;
  assign n5717 = n5569 & ~n5716;
  assign n5718 = n5717 ^ n5568;
  assign n5722 = n5721 ^ n5718;
  assign n5727 = n5726 ^ n5722;
  assign n5743 = n5742 ^ n5727;
  assign n5713 = n5635 ^ n5615;
  assign n5714 = n5636 & ~n5713;
  assign n5715 = n5714 ^ n5618;
  assign n5744 = n5743 ^ n5715;
  assign n5706 = n5625 ^ n5624;
  assign n5707 = n5627 & ~n5706;
  assign n5708 = n5707 ^ n5626;
  assign n5703 = n5584 ^ n5583;
  assign n5704 = n5586 & ~n5703;
  assign n5705 = n5704 ^ n5585;
  assign n5709 = n5708 ^ n5705;
  assign n5700 = n5620 ^ n5619;
  assign n5701 = n5622 & ~n5700;
  assign n5702 = n5701 ^ n5621;
  assign n5710 = n5709 ^ n5702;
  assign n5697 = n5628 ^ n5623;
  assign n5698 = n5634 & ~n5697;
  assign n5699 = n5698 ^ n5633;
  assign n5711 = n5710 ^ n5699;
  assign n5694 = n5570 ^ n5565;
  assign n5695 = n5576 & ~n5694;
  assign n5696 = n5695 ^ n5575;
  assign n5712 = n5711 ^ n5696;
  assign n5745 = n5744 ^ n5712;
  assign n5827 = n5826 ^ n5745;
  assign n5691 = n5499 ^ n5477;
  assign n5692 = n5500 & ~n5691;
  assign n5693 = n5692 ^ n5477;
  assign n5828 = n5827 ^ n5693;
  assign n5682 = n5513 ^ n5510;
  assign n5683 = n5517 & ~n5682;
  assign n5684 = n5683 ^ n5516;
  assign n5679 = n5534 ^ n5531;
  assign n5680 = n5538 & ~n5679;
  assign n5681 = n5680 ^ n5537;
  assign n5685 = n5684 ^ n5681;
  assign n5676 = n5613 ^ n5605;
  assign n5677 = n5614 & ~n5676;
  assign n5678 = n5677 ^ n5608;
  assign n5686 = n5685 ^ n5678;
  assign n5673 = n5547 ^ n5544;
  assign n5674 = n5551 & ~n5673;
  assign n5675 = n5674 ^ n5550;
  assign n5687 = n5686 ^ n5675;
  assign n5670 = n5598 ^ n5560;
  assign n5671 = n5599 & ~n5670;
  assign n5672 = n5671 ^ n5560;
  assign n5688 = n5687 ^ n5672;
  assign n5667 = n5552 ^ n5507;
  assign n5668 = ~n5553 & n5667;
  assign n5669 = n5668 ^ n5507;
  assign n5689 = n5688 ^ n5669;
  assign n5664 = n5637 ^ n5557;
  assign n5665 = n5638 & ~n5664;
  assign n5666 = n5665 ^ n5557;
  assign n5690 = n5689 ^ n5666;
  assign n5829 = n5828 ^ n5690;
  assign n5661 = n5554 ^ n5504;
  assign n5662 = n5640 & n5661;
  assign n5663 = n5662 ^ n5639;
  assign n5830 = n5829 ^ n5663;
  assign n5658 = n5501 ^ n5474;
  assign n5659 = n5642 & n5658;
  assign n5660 = n5659 ^ n5641;
  assign n5831 = n5830 ^ n5660;
  assign n5655 = n5653 ^ n5471;
  assign n5656 = n5644 & n5655;
  assign n5657 = n5656 ^ n5653;
  assign n5832 = n5831 ^ n5657;
  assign n6004 = n5690 & ~n5828;
  assign n6005 = ~n5663 & n6004;
  assign n6006 = ~n5660 & ~n6005;
  assign n6007 = n5828 ^ n5663;
  assign n6008 = n5829 & n6007;
  assign n6009 = n6008 ^ n5663;
  assign n6010 = ~n6006 & ~n6009;
  assign n6011 = n5657 & n6010;
  assign n6012 = ~n5690 & n5828;
  assign n6013 = n5663 & n6012;
  assign n6014 = ~n5660 & n6013;
  assign n6015 = ~n6011 & ~n6014;
  assign n6016 = n5660 & ~n6013;
  assign n6017 = n6009 & ~n6016;
  assign n6018 = ~n5657 & n6017;
  assign n6019 = n5660 & n6005;
  assign n6020 = ~n6018 & ~n6019;
  assign n6021 = n6015 & n6020;
  assign n5993 = x28 & x33;
  assign n5992 = x27 & x34;
  assign n5994 = n5993 ^ n5992;
  assign n5991 = x26 & x35;
  assign n5995 = n5994 ^ n5991;
  assign n5988 = x19 & x42;
  assign n5987 = x8 & x53;
  assign n5989 = n5988 ^ n5987;
  assign n5986 = x7 & x54;
  assign n5990 = n5989 ^ n5986;
  assign n5996 = n5995 ^ n5990;
  assign n5983 = x18 & x43;
  assign n5982 = x17 & x44;
  assign n5984 = n5983 ^ n5982;
  assign n5981 = x9 & x52;
  assign n5985 = n5984 ^ n5981;
  assign n5997 = n5996 ^ n5985;
  assign n5978 = n5699 ^ n5696;
  assign n5979 = n5711 & ~n5978;
  assign n5980 = n5979 ^ n5710;
  assign n5998 = n5997 ^ n5980;
  assign n5975 = n5741 ^ n5727;
  assign n5976 = ~n5742 & ~n5975;
  assign n5977 = n5976 ^ n5730;
  assign n5999 = n5998 ^ n5977;
  assign n5966 = x29 & x59;
  assign n5967 = x1 & n5966;
  assign n5968 = x31 & ~n5967;
  assign n5965 = x1 & x60;
  assign n5969 = n5968 ^ n5965;
  assign n5962 = n5763 ^ n5762;
  assign n5963 = n5765 & ~n5962;
  assign n5964 = n5963 ^ n5764;
  assign n5970 = n5969 ^ n5964;
  assign n5959 = n5736 ^ n5733;
  assign n5960 = n5740 & ~n5959;
  assign n5961 = n5960 ^ n5739;
  assign n5971 = n5970 ^ n5961;
  assign n5956 = n5803 ^ n5793;
  assign n5957 = ~n5804 & n5956;
  assign n5958 = n5957 ^ n5793;
  assign n5972 = n5971 ^ n5958;
  assign n5951 = x23 & x38;
  assign n5950 = x4 & x57;
  assign n5952 = n5951 ^ n5950;
  assign n5949 = x3 & x58;
  assign n5953 = n5952 ^ n5949;
  assign n5946 = n5705 ^ n5702;
  assign n5947 = n5709 & ~n5946;
  assign n5948 = n5947 ^ n5708;
  assign n5954 = n5953 ^ n5948;
  assign n5943 = n5726 ^ n5721;
  assign n5944 = ~n5722 & n5943;
  assign n5945 = n5944 ^ n5726;
  assign n5955 = n5954 ^ n5945;
  assign n5973 = n5972 ^ n5955;
  assign n5940 = n5822 ^ n5790;
  assign n5941 = ~n5823 & ~n5940;
  assign n5942 = n5941 ^ n5790;
  assign n5974 = n5973 ^ n5942;
  assign n6000 = n5999 ^ n5974;
  assign n5937 = n5824 ^ n5748;
  assign n5938 = n5825 & ~n5937;
  assign n5939 = n5938 ^ n5748;
  assign n6001 = n6000 ^ n5939;
  assign n5934 = n5826 ^ n5693;
  assign n5935 = ~n5827 & ~n5934;
  assign n5936 = n5935 ^ n5693;
  assign n6002 = n6001 ^ n5936;
  assign n5923 = x14 & x47;
  assign n5922 = x12 & x49;
  assign n5924 = n5923 ^ n5922;
  assign n5921 = x11 & x50;
  assign n5925 = n5924 ^ n5921;
  assign n5918 = x16 & x45;
  assign n5917 = x15 & x46;
  assign n5919 = n5918 ^ n5917;
  assign n5916 = x10 & x51;
  assign n5920 = n5919 ^ n5916;
  assign n5926 = n5925 ^ n5920;
  assign n5913 = x30 & x31;
  assign n5912 = x29 & x32;
  assign n5914 = n5913 ^ n5912;
  assign n5911 = x13 & x48;
  assign n5915 = n5914 ^ n5911;
  assign n5927 = n5926 ^ n5915;
  assign n5906 = x5 & x56;
  assign n5905 = x2 & x59;
  assign n5907 = n5906 ^ n5905;
  assign n5904 = x0 & x61;
  assign n5908 = n5907 ^ n5904;
  assign n5901 = x25 & x36;
  assign n5900 = x24 & x37;
  assign n5902 = n5901 ^ n5900;
  assign n5899 = x22 & x39;
  assign n5903 = n5902 ^ n5899;
  assign n5909 = n5908 ^ n5903;
  assign n5897 = n2963 ^ n2856;
  assign n5896 = x6 & x55;
  assign n5898 = n5897 ^ n5896;
  assign n5910 = n5909 ^ n5898;
  assign n5928 = n5927 ^ n5910;
  assign n5893 = n5681 ^ n5678;
  assign n5894 = n5685 & ~n5893;
  assign n5895 = n5894 ^ n5684;
  assign n5929 = n5928 ^ n5895;
  assign n5890 = n5675 ^ n5672;
  assign n5891 = ~n5687 & n5890;
  assign n5892 = n5891 ^ n5672;
  assign n5930 = n5929 ^ n5892;
  assign n5887 = n5743 ^ n5712;
  assign n5888 = ~n5744 & n5887;
  assign n5889 = n5888 ^ n5715;
  assign n5931 = n5930 ^ n5889;
  assign n5878 = n5812 ^ n5811;
  assign n5879 = n5814 & ~n5878;
  assign n5880 = n5879 ^ n5813;
  assign n5875 = n5773 ^ n5772;
  assign n5876 = n5775 & ~n5875;
  assign n5877 = n5876 ^ n5774;
  assign n5881 = n5880 ^ n5877;
  assign n5872 = n5817 ^ n5816;
  assign n5873 = n5819 & ~n5872;
  assign n5874 = n5873 ^ n5818;
  assign n5882 = n5881 ^ n5874;
  assign n5867 = n5753 ^ n5752;
  assign n5868 = n5755 & ~n5867;
  assign n5869 = n5868 ^ n5754;
  assign n5864 = n5807 ^ n5806;
  assign n5865 = n5809 & ~n5864;
  assign n5866 = n5865 ^ n5808;
  assign n5870 = n5869 ^ n5866;
  assign n5861 = n5795 ^ n5794;
  assign n5862 = n5797 & ~n5861;
  assign n5863 = n5862 ^ n5796;
  assign n5871 = n5870 ^ n5863;
  assign n5883 = n5882 ^ n5871;
  assign n5858 = n5815 ^ n5810;
  assign n5859 = n5821 & ~n5858;
  assign n5860 = n5859 ^ n5820;
  assign n5884 = n5883 ^ n5860;
  assign n5855 = n5785 ^ n5751;
  assign n5856 = ~n5786 & n5855;
  assign n5857 = n5856 ^ n5751;
  assign n5885 = n5884 ^ n5857;
  assign n5850 = n5783 ^ n5771;
  assign n5851 = ~n5784 & n5850;
  assign n5852 = n5851 ^ n5771;
  assign n5847 = n5761 ^ n5756;
  assign n5848 = n5767 & ~n5847;
  assign n5849 = n5848 ^ n5766;
  assign n5853 = n5852 ^ n5849;
  assign n5842 = n5800 ^ n5799;
  assign n5843 = n5802 & ~n5842;
  assign n5844 = n5843 ^ n5801;
  assign n5839 = n5758 ^ n5757;
  assign n5840 = n5760 & ~n5839;
  assign n5841 = n5840 ^ n5759;
  assign n5845 = n5844 ^ n5841;
  assign n5836 = n5780 ^ n5777;
  assign n5837 = n5782 & ~n5836;
  assign n5838 = n5837 ^ n5781;
  assign n5846 = n5845 ^ n5838;
  assign n5854 = n5853 ^ n5846;
  assign n5886 = n5885 ^ n5854;
  assign n5932 = n5931 ^ n5886;
  assign n5833 = n5669 ^ n5666;
  assign n5834 = ~n5689 & ~n5833;
  assign n5835 = n5834 ^ n5666;
  assign n5933 = n5932 ^ n5835;
  assign n6003 = n6002 ^ n5933;
  assign n6022 = n6021 ^ n6003;
  assign n6209 = n6003 & ~n6014;
  assign n6210 = ~n6010 & ~n6209;
  assign n6211 = n5657 & ~n6210;
  assign n6212 = n6003 & ~n6017;
  assign n6213 = ~n6019 & ~n6212;
  assign n6214 = ~n6211 & n6213;
  assign n6196 = x0 & x62;
  assign n6194 = n1688 ^ x2;
  assign n6195 = x60 & n6194;
  assign n6197 = n6196 ^ n6195;
  assign n6191 = x17 & x45;
  assign n6190 = x10 & x52;
  assign n6192 = n6191 ^ n6190;
  assign n6189 = x9 & x53;
  assign n6193 = n6192 ^ n6189;
  assign n6198 = n6197 ^ n6193;
  assign n6186 = x26 & x36;
  assign n6185 = x25 & x37;
  assign n6187 = n6186 ^ n6185;
  assign n6184 = x21 & x41;
  assign n6188 = n6187 ^ n6184;
  assign n6199 = n6198 ^ n6188;
  assign n6179 = x19 & x43;
  assign n6178 = x18 & x44;
  assign n6180 = n6179 ^ n6178;
  assign n6177 = x8 & x54;
  assign n6181 = n6180 ^ n6177;
  assign n6174 = x24 & x38;
  assign n6173 = x23 & x39;
  assign n6175 = n6174 ^ n6173;
  assign n6172 = x22 & x40;
  assign n6176 = n6175 ^ n6172;
  assign n6182 = n6181 ^ n6176;
  assign n6169 = x29 & x33;
  assign n6168 = x28 & x34;
  assign n6170 = n6169 ^ n6168;
  assign n6167 = x27 & x35;
  assign n6171 = n6170 ^ n6167;
  assign n6183 = n6182 ^ n6171;
  assign n6200 = n6199 ^ n6183;
  assign n6162 = x14 & x48;
  assign n6161 = x13 & x49;
  assign n6163 = n6162 ^ n6161;
  assign n6160 = x12 & x50;
  assign n6164 = n6163 ^ n6160;
  assign n6157 = x16 & x46;
  assign n6156 = x15 & x47;
  assign n6158 = n6157 ^ n6156;
  assign n6155 = x11 & x51;
  assign n6159 = n6158 ^ n6155;
  assign n6165 = n6164 ^ n6159;
  assign n6152 = x20 & x42;
  assign n6151 = x7 & x55;
  assign n6153 = n6152 ^ n6151;
  assign n6150 = x6 & x56;
  assign n6154 = n6153 ^ n6150;
  assign n6166 = n6165 ^ n6154;
  assign n6201 = n6200 ^ n6166;
  assign n6147 = n5972 ^ n5942;
  assign n6148 = ~n5973 & ~n6147;
  assign n6149 = n6148 ^ n5942;
  assign n6202 = n6201 ^ n6149;
  assign n6144 = n5884 ^ n5854;
  assign n6145 = n5885 & ~n6144;
  assign n6146 = n6145 ^ n5857;
  assign n6203 = n6202 ^ n6146;
  assign n6135 = x5 & x57;
  assign n6134 = x4 & x58;
  assign n6136 = n6135 ^ n6134;
  assign n6133 = x3 & x59;
  assign n6137 = n6136 ^ n6133;
  assign n6130 = n5982 ^ n5981;
  assign n6131 = n5984 & ~n6130;
  assign n6132 = n6131 ^ n5983;
  assign n6138 = n6137 ^ n6132;
  assign n6127 = n5917 ^ n5916;
  assign n6128 = n5919 & ~n6127;
  assign n6129 = n6128 ^ n5918;
  assign n6139 = n6138 ^ n6129;
  assign n6124 = n5953 ^ n5945;
  assign n6125 = n5954 & ~n6124;
  assign n6126 = n6125 ^ n5948;
  assign n6140 = n6139 ^ n6126;
  assign n6121 = n5990 ^ n5985;
  assign n6122 = n5996 & ~n6121;
  assign n6123 = n6122 ^ n5995;
  assign n6141 = n6140 ^ n6123;
  assign n6108 = x60 & n5964;
  assign n6109 = x31 & x59;
  assign n6110 = x29 & n6109;
  assign n6111 = ~n6108 & ~n6110;
  assign n6112 = x31 & x60;
  assign n6113 = x1 & ~n6112;
  assign n6114 = ~n6111 & n6113;
  assign n6115 = n5965 & ~n5966;
  assign n6116 = x31 & ~n6115;
  assign n6117 = n5964 & n6116;
  assign n6118 = ~n6114 & ~n6117;
  assign n6105 = n5844 ^ n5838;
  assign n6106 = ~n5845 & n6105;
  assign n6107 = n6106 ^ n5838;
  assign n6119 = n6118 ^ n6107;
  assign n6102 = n5877 ^ n5874;
  assign n6103 = n5881 & ~n6102;
  assign n6104 = n6103 ^ n5880;
  assign n6120 = n6119 ^ n6104;
  assign n6142 = n6141 ^ n6120;
  assign n6099 = n5927 ^ n5895;
  assign n6100 = ~n5928 & n6099;
  assign n6101 = n6100 ^ n5895;
  assign n6143 = n6142 ^ n6101;
  assign n6204 = n6203 ^ n6143;
  assign n6096 = n5999 ^ n5939;
  assign n6097 = ~n6000 & ~n6096;
  assign n6098 = n6097 ^ n5939;
  assign n6205 = n6204 ^ n6098;
  assign n6087 = n5866 ^ n5863;
  assign n6088 = n5870 & ~n6087;
  assign n6089 = n6088 ^ n5869;
  assign n6084 = n5903 ^ n5898;
  assign n6085 = n5909 & ~n6084;
  assign n6086 = n6085 ^ n5908;
  assign n6090 = n6089 ^ n6086;
  assign n6081 = n5920 ^ n5915;
  assign n6082 = n5926 & ~n6081;
  assign n6083 = n6082 ^ n5925;
  assign n6091 = n6090 ^ n6083;
  assign n6074 = n5912 ^ n5911;
  assign n6075 = n5914 & ~n6074;
  assign n6076 = n6075 ^ n5913;
  assign n6071 = n5922 ^ n5921;
  assign n6072 = n5924 & ~n6071;
  assign n6073 = n6072 ^ n5923;
  assign n6077 = n6076 ^ n6073;
  assign n6069 = x1 & x61;
  assign n6068 = x30 & x32;
  assign n6070 = n6069 ^ n6068;
  assign n6078 = n6077 ^ n6070;
  assign n6063 = n5905 ^ n5904;
  assign n6064 = n5907 & ~n6063;
  assign n6065 = n6064 ^ n5906;
  assign n6060 = n5987 ^ n5986;
  assign n6061 = n5989 & ~n6060;
  assign n6062 = n6061 ^ n5988;
  assign n6066 = n6065 ^ n6062;
  assign n6057 = n5896 ^ n2963;
  assign n6058 = n5897 & ~n6057;
  assign n6059 = n6058 ^ n2856;
  assign n6067 = n6066 ^ n6059;
  assign n6079 = n6078 ^ n6067;
  assign n6052 = n5992 ^ n5991;
  assign n6053 = n5994 & ~n6052;
  assign n6054 = n6053 ^ n5993;
  assign n6049 = n5900 ^ n5899;
  assign n6050 = n5902 & ~n6049;
  assign n6051 = n6050 ^ n5901;
  assign n6055 = n6054 ^ n6051;
  assign n6046 = n5950 ^ n5949;
  assign n6047 = n5952 & ~n6046;
  assign n6048 = n6047 ^ n5951;
  assign n6056 = n6055 ^ n6048;
  assign n6080 = n6079 ^ n6056;
  assign n6092 = n6091 ^ n6080;
  assign n6043 = n5980 ^ n5977;
  assign n6044 = ~n5998 & ~n6043;
  assign n6045 = n6044 ^ n5977;
  assign n6093 = n6092 ^ n6045;
  assign n6038 = n5970 ^ n5958;
  assign n6039 = n5971 & ~n6038;
  assign n6040 = n6039 ^ n5961;
  assign n6035 = n5871 ^ n5860;
  assign n6036 = n5883 & ~n6035;
  assign n6037 = n6036 ^ n5882;
  assign n6041 = n6040 ^ n6037;
  assign n6032 = n5849 ^ n5846;
  assign n6033 = n5853 & ~n6032;
  assign n6034 = n6033 ^ n5852;
  assign n6042 = n6041 ^ n6034;
  assign n6094 = n6093 ^ n6042;
  assign n6029 = n5892 ^ n5889;
  assign n6030 = ~n5930 & n6029;
  assign n6031 = n6030 ^ n5889;
  assign n6095 = n6094 ^ n6031;
  assign n6206 = n6205 ^ n6095;
  assign n6026 = n5931 ^ n5835;
  assign n6027 = ~n5932 & ~n6026;
  assign n6028 = n6027 ^ n5835;
  assign n6207 = n6206 ^ n6028;
  assign n6023 = n6001 ^ n5933;
  assign n6024 = n6002 & n6023;
  assign n6025 = n6024 ^ n5936;
  assign n6208 = n6207 ^ n6025;
  assign n6215 = n6214 ^ n6208;
  assign n6393 = n6086 ^ n6083;
  assign n6394 = n6090 & ~n6393;
  assign n6395 = n6394 ^ n6089;
  assign n6390 = n6067 ^ n6056;
  assign n6391 = n6079 & ~n6390;
  assign n6392 = n6391 ^ n6078;
  assign n6396 = n6395 ^ n6392;
  assign n6387 = n6139 ^ n6123;
  assign n6388 = n6140 & ~n6387;
  assign n6389 = n6388 ^ n6126;
  assign n6397 = n6396 ^ n6389;
  assign n6380 = n6051 ^ n6048;
  assign n6381 = n6055 & ~n6380;
  assign n6382 = n6381 ^ n6054;
  assign n6377 = n6137 ^ n6129;
  assign n6378 = n6138 & ~n6377;
  assign n6379 = n6378 ^ n6132;
  assign n6383 = n6382 ^ n6379;
  assign n6374 = n6073 ^ n6070;
  assign n6375 = n6077 & ~n6374;
  assign n6376 = n6375 ^ n6076;
  assign n6384 = n6383 ^ n6376;
  assign n6367 = ~x2 & ~n1688;
  assign n6368 = x60 & ~n6367;
  assign n6366 = n6195 & ~n6196;
  assign n6369 = n6368 ^ n6366;
  assign n6363 = n6134 ^ n6133;
  assign n6364 = n6136 & ~n6363;
  assign n6365 = n6364 ^ n6135;
  assign n6370 = n6369 ^ n6365;
  assign n6360 = n6185 ^ n6184;
  assign n6361 = n6187 & ~n6360;
  assign n6362 = n6361 ^ n6186;
  assign n6371 = n6370 ^ n6362;
  assign n6355 = n6161 ^ n6160;
  assign n6356 = n6163 & ~n6355;
  assign n6357 = n6356 ^ n6162;
  assign n6352 = n6173 ^ n6172;
  assign n6353 = n6175 & ~n6352;
  assign n6354 = n6353 ^ n6174;
  assign n6358 = n6357 ^ n6354;
  assign n6349 = n6151 ^ n6150;
  assign n6350 = n6153 & ~n6349;
  assign n6351 = n6350 ^ n6152;
  assign n6359 = n6358 ^ n6351;
  assign n6372 = n6371 ^ n6359;
  assign n6346 = n6062 ^ n6059;
  assign n6347 = n6066 & ~n6346;
  assign n6348 = n6347 ^ n6065;
  assign n6373 = n6372 ^ n6348;
  assign n6385 = n6384 ^ n6373;
  assign n6343 = n6183 ^ n6166;
  assign n6344 = n6200 & ~n6343;
  assign n6345 = n6344 ^ n6199;
  assign n6386 = n6385 ^ n6345;
  assign n6398 = n6397 ^ n6386;
  assign n6340 = n6201 ^ n6146;
  assign n6341 = ~n6202 & ~n6340;
  assign n6342 = n6341 ^ n6149;
  assign n6399 = n6398 ^ n6342;
  assign n6337 = n6203 ^ n6098;
  assign n6338 = ~n6204 & ~n6337;
  assign n6339 = n6338 ^ n6098;
  assign n6400 = n6399 ^ n6339;
  assign n6326 = x31 & x32;
  assign n6325 = x30 & x33;
  assign n6327 = n6326 ^ n6325;
  assign n6324 = x14 & x49;
  assign n6328 = n6327 ^ n6324;
  assign n6321 = x23 & x40;
  assign n6320 = x20 & x43;
  assign n6322 = n6321 ^ n6320;
  assign n6319 = x6 & x57;
  assign n6323 = n6322 ^ n6319;
  assign n6329 = n6328 ^ n6323;
  assign n6316 = x19 & x44;
  assign n6315 = x8 & x55;
  assign n6317 = n6316 ^ n6315;
  assign n6314 = x7 & x56;
  assign n6318 = n6317 ^ n6314;
  assign n6330 = n6329 ^ n6318;
  assign n6309 = x15 & x48;
  assign n6308 = x13 & x50;
  assign n6310 = n6309 ^ n6308;
  assign n6307 = x12 & x51;
  assign n6311 = n6310 ^ n6307;
  assign n6304 = x18 & x45;
  assign n6303 = x17 & x46;
  assign n6305 = n6304 ^ n6303;
  assign n6302 = x9 & x54;
  assign n6306 = n6305 ^ n6302;
  assign n6312 = n6311 ^ n6306;
  assign n6299 = x16 & x47;
  assign n6298 = x11 & x52;
  assign n6300 = n6299 ^ n6298;
  assign n6297 = x10 & x53;
  assign n6301 = n6300 ^ n6297;
  assign n6313 = n6312 ^ n6301;
  assign n6331 = n6330 ^ n6313;
  assign n6292 = x4 & x59;
  assign n6291 = x3 & x60;
  assign n6293 = n6292 ^ n6291;
  assign n6290 = x2 & x61;
  assign n6294 = n6293 ^ n6290;
  assign n6287 = x22 & x41;
  assign n6286 = x21 & x42;
  assign n6288 = n6287 ^ n6286;
  assign n6285 = x5 & x58;
  assign n6289 = n6288 ^ n6285;
  assign n6295 = n6294 ^ n6289;
  assign n6282 = n6156 ^ n6155;
  assign n6283 = n6158 & ~n6282;
  assign n6284 = n6283 ^ n6157;
  assign n6296 = n6295 ^ n6284;
  assign n6332 = n6331 ^ n6296;
  assign n6279 = n6120 ^ n6101;
  assign n6280 = ~n6142 & n6279;
  assign n6281 = n6280 ^ n6141;
  assign n6333 = n6332 ^ n6281;
  assign n6276 = n6091 ^ n6045;
  assign n6277 = ~n6092 & ~n6276;
  assign n6278 = n6277 ^ n6045;
  assign n6334 = n6333 ^ n6278;
  assign n6267 = x29 & x34;
  assign n6266 = x28 & x35;
  assign n6268 = n6267 ^ n6266;
  assign n6265 = x27 & x36;
  assign n6269 = n6268 ^ n6265;
  assign n6262 = x26 & x37;
  assign n6261 = x25 & x38;
  assign n6263 = n6262 ^ n6261;
  assign n6260 = x24 & x39;
  assign n6264 = n6263 ^ n6260;
  assign n6270 = n6269 ^ n6264;
  assign n6256 = x30 & x61;
  assign n6257 = x1 & n6256;
  assign n6258 = x32 & ~n6257;
  assign n6254 = x0 & x63;
  assign n6253 = x1 & x62;
  assign n6255 = n6254 ^ n6253;
  assign n6259 = n6258 ^ n6255;
  assign n6271 = n6270 ^ n6259;
  assign n6250 = n6193 ^ n6188;
  assign n6251 = n6198 & ~n6250;
  assign n6252 = n6251 ^ n6197;
  assign n6272 = n6271 ^ n6252;
  assign n6247 = n6107 ^ n6104;
  assign n6248 = ~n6119 & ~n6247;
  assign n6249 = n6248 ^ n6118;
  assign n6273 = n6272 ^ n6249;
  assign n6240 = n6178 ^ n6177;
  assign n6241 = n6180 & ~n6240;
  assign n6242 = n6241 ^ n6179;
  assign n6237 = n6190 ^ n6189;
  assign n6238 = n6192 & ~n6237;
  assign n6239 = n6238 ^ n6191;
  assign n6243 = n6242 ^ n6239;
  assign n6234 = n6168 ^ n6167;
  assign n6235 = n6170 & ~n6234;
  assign n6236 = n6235 ^ n6169;
  assign n6244 = n6243 ^ n6236;
  assign n6231 = n6159 ^ n6154;
  assign n6232 = n6165 & ~n6231;
  assign n6233 = n6232 ^ n6164;
  assign n6245 = n6244 ^ n6233;
  assign n6228 = n6176 ^ n6171;
  assign n6229 = n6182 & ~n6228;
  assign n6230 = n6229 ^ n6181;
  assign n6246 = n6245 ^ n6230;
  assign n6274 = n6273 ^ n6246;
  assign n6225 = n6040 ^ n6034;
  assign n6226 = ~n6041 & n6225;
  assign n6227 = n6226 ^ n6034;
  assign n6275 = n6274 ^ n6227;
  assign n6335 = n6334 ^ n6275;
  assign n6222 = n6093 ^ n6031;
  assign n6223 = n6094 & ~n6222;
  assign n6224 = n6223 ^ n6031;
  assign n6336 = n6335 ^ n6224;
  assign n6401 = n6400 ^ n6336;
  assign n6219 = n6205 ^ n6028;
  assign n6220 = n6206 & ~n6219;
  assign n6221 = n6220 ^ n6028;
  assign n6402 = n6401 ^ n6221;
  assign n6216 = n6214 ^ n6207;
  assign n6217 = ~n6208 & n6216;
  assign n6218 = n6217 ^ n6214;
  assign n6403 = n6402 ^ n6218;
  assign n6590 = x32 & x62;
  assign n6591 = ~x63 & ~n6590;
  assign n6592 = x1 & ~n6591;
  assign n6521 = x32 & x63;
  assign n6593 = x62 & n6521;
  assign n6594 = n6592 & ~n6593;
  assign n6587 = n6325 ^ n6324;
  assign n6588 = n6327 & ~n6587;
  assign n6589 = n6588 ^ n6326;
  assign n6595 = n6594 ^ n6589;
  assign n6583 = x13 & x51;
  assign n6582 = x12 & x52;
  assign n6584 = n6583 ^ n6582;
  assign n6581 = x11 & x53;
  assign n6585 = n6584 ^ n6581;
  assign n6578 = x15 & x49;
  assign n6577 = x10 & x54;
  assign n6579 = n6578 ^ n6577;
  assign n6576 = x9 & x55;
  assign n6580 = n6579 ^ n6576;
  assign n6586 = n6585 ^ n6580;
  assign n6596 = n6595 ^ n6586;
  assign n6573 = n6379 ^ n6376;
  assign n6574 = n6383 & ~n6573;
  assign n6575 = n6574 ^ n6382;
  assign n6597 = n6596 ^ n6575;
  assign n6570 = n6294 ^ n6284;
  assign n6571 = ~n6295 & n6570;
  assign n6572 = n6571 ^ n6284;
  assign n6598 = n6597 ^ n6572;
  assign n6563 = n6298 ^ n6297;
  assign n6564 = n6300 & ~n6563;
  assign n6565 = n6564 ^ n6299;
  assign n6560 = n6308 ^ n6307;
  assign n6561 = n6310 & ~n6560;
  assign n6562 = n6561 ^ n6309;
  assign n6566 = n6565 ^ n6562;
  assign n6557 = n6261 ^ n6260;
  assign n6558 = n6263 & ~n6557;
  assign n6559 = n6558 ^ n6262;
  assign n6567 = n6566 ^ n6559;
  assign n6554 = n6323 ^ n6318;
  assign n6555 = n6329 & ~n6554;
  assign n6556 = n6555 ^ n6328;
  assign n6568 = n6567 ^ n6556;
  assign n6551 = n6306 ^ n6301;
  assign n6552 = n6312 & ~n6551;
  assign n6553 = n6552 ^ n6311;
  assign n6569 = n6568 ^ n6553;
  assign n6599 = n6598 ^ n6569;
  assign n6548 = n6395 ^ n6389;
  assign n6549 = ~n6396 & n6548;
  assign n6550 = n6549 ^ n6389;
  assign n6600 = n6599 ^ n6550;
  assign n6539 = n6354 ^ n6351;
  assign n6540 = n6358 & ~n6539;
  assign n6541 = n6540 ^ n6357;
  assign n6536 = n6239 ^ n6236;
  assign n6537 = n6243 & ~n6536;
  assign n6538 = n6537 ^ n6242;
  assign n6542 = n6541 ^ n6538;
  assign n6533 = n6365 ^ n6362;
  assign n6534 = n6370 & ~n6533;
  assign n6535 = n6534 ^ n6369;
  assign n6543 = n6542 ^ n6535;
  assign n6530 = n6371 ^ n6348;
  assign n6531 = ~n6372 & n6530;
  assign n6532 = n6531 ^ n6348;
  assign n6544 = n6543 ^ n6532;
  assign n6527 = n6233 ^ n6230;
  assign n6528 = n6245 & ~n6527;
  assign n6529 = n6528 ^ n6244;
  assign n6545 = n6544 ^ n6529;
  assign n6514 = x32 & x61;
  assign n6515 = n1571 & n6514;
  assign n6516 = ~n6253 & ~n6515;
  assign n6517 = ~x32 & n6254;
  assign n6518 = x62 & ~n6517;
  assign n6519 = ~n6516 & ~n6518;
  assign n6520 = n6253 & ~n6256;
  assign n6522 = x0 & n6521;
  assign n6523 = ~n6520 & n6522;
  assign n6524 = ~n6519 & ~n6523;
  assign n6510 = x19 & x45;
  assign n6509 = x18 & x46;
  assign n6511 = n6510 ^ n6509;
  assign n6508 = x5 & x59;
  assign n6512 = n6511 ^ n6508;
  assign n6505 = x4 & x60;
  assign n6504 = x3 & x61;
  assign n6506 = n6505 ^ n6504;
  assign n6503 = x2 & x62;
  assign n6507 = n6506 ^ n6503;
  assign n6513 = n6512 ^ n6507;
  assign n6525 = n6524 ^ n6513;
  assign n6497 = x17 & x47;
  assign n6496 = x7 & x57;
  assign n6498 = n6497 ^ n6496;
  assign n6495 = x6 & x58;
  assign n6499 = n6498 ^ n6495;
  assign n6492 = x25 & x39;
  assign n6491 = x24 & x40;
  assign n6493 = n6492 ^ n6491;
  assign n6490 = x23 & x41;
  assign n6494 = n6493 ^ n6490;
  assign n6500 = n6499 ^ n6494;
  assign n6488 = n3238 ^ n3200;
  assign n6487 = x20 & x44;
  assign n6489 = n6488 ^ n6487;
  assign n6501 = n6500 ^ n6489;
  assign n6482 = x29 & x35;
  assign n6481 = x28 & x36;
  assign n6483 = n6482 ^ n6481;
  assign n6480 = x27 & x37;
  assign n6484 = n6483 ^ n6480;
  assign n6477 = x26 & x38;
  assign n6476 = x16 & x48;
  assign n6478 = n6477 ^ n6476;
  assign n6475 = x8 & x56;
  assign n6479 = n6478 ^ n6475;
  assign n6485 = n6484 ^ n6479;
  assign n6472 = x31 & x33;
  assign n6471 = x30 & x34;
  assign n6473 = n6472 ^ n6471;
  assign n6470 = x14 & x50;
  assign n6474 = n6473 ^ n6470;
  assign n6486 = n6485 ^ n6474;
  assign n6502 = n6501 ^ n6486;
  assign n6526 = n6525 ^ n6502;
  assign n6546 = n6545 ^ n6526;
  assign n6467 = n6384 ^ n6345;
  assign n6468 = ~n6385 & n6467;
  assign n6469 = n6468 ^ n6345;
  assign n6547 = n6546 ^ n6469;
  assign n6601 = n6600 ^ n6547;
  assign n6464 = n6397 ^ n6342;
  assign n6465 = ~n6398 & ~n6464;
  assign n6466 = n6465 ^ n6342;
  assign n6602 = n6601 ^ n6466;
  assign n6453 = n6266 ^ n6265;
  assign n6454 = n6268 & ~n6453;
  assign n6455 = n6454 ^ n6267;
  assign n6450 = n6303 ^ n6302;
  assign n6451 = n6305 & ~n6450;
  assign n6452 = n6451 ^ n6304;
  assign n6456 = n6455 ^ n6452;
  assign n6447 = n6320 ^ n6319;
  assign n6448 = n6322 & ~n6447;
  assign n6449 = n6448 ^ n6321;
  assign n6457 = n6456 ^ n6449;
  assign n6442 = n6291 ^ n6290;
  assign n6443 = n6293 & ~n6442;
  assign n6444 = n6443 ^ n6292;
  assign n6439 = n6315 ^ n6314;
  assign n6440 = n6317 & ~n6439;
  assign n6441 = n6440 ^ n6316;
  assign n6445 = n6444 ^ n6441;
  assign n6436 = n6286 ^ n6285;
  assign n6437 = n6288 & ~n6436;
  assign n6438 = n6437 ^ n6287;
  assign n6446 = n6445 ^ n6438;
  assign n6458 = n6457 ^ n6446;
  assign n6433 = n6264 ^ n6259;
  assign n6434 = n6270 & ~n6433;
  assign n6435 = n6434 ^ n6269;
  assign n6459 = n6458 ^ n6435;
  assign n6430 = n6313 ^ n6296;
  assign n6431 = n6331 & ~n6430;
  assign n6432 = n6431 ^ n6330;
  assign n6460 = n6459 ^ n6432;
  assign n6427 = n6252 ^ n6249;
  assign n6428 = ~n6272 & ~n6427;
  assign n6429 = n6428 ^ n6249;
  assign n6461 = n6460 ^ n6429;
  assign n6424 = n6273 ^ n6227;
  assign n6425 = n6274 & ~n6424;
  assign n6426 = n6425 ^ n6227;
  assign n6462 = n6461 ^ n6426;
  assign n6421 = n6332 ^ n6278;
  assign n6422 = n6333 & n6421;
  assign n6423 = n6422 ^ n6281;
  assign n6463 = n6462 ^ n6423;
  assign n6603 = n6602 ^ n6463;
  assign n6418 = n6334 ^ n6224;
  assign n6419 = ~n6335 & ~n6418;
  assign n6420 = n6419 ^ n6224;
  assign n6604 = n6603 ^ n6420;
  assign n6404 = ~n6221 & n6339;
  assign n6405 = n6336 & ~n6399;
  assign n6406 = n6404 & n6405;
  assign n6407 = n6221 & ~n6339;
  assign n6408 = ~n6336 & n6399;
  assign n6409 = n6407 & n6408;
  assign n6410 = ~n6406 & ~n6409;
  assign n6412 = ~n6407 & ~n6408;
  assign n6411 = ~n6404 & ~n6405;
  assign n6413 = n6412 ^ n6411;
  assign n6414 = n6411 ^ n6218;
  assign n6415 = n6413 & n6414;
  assign n6416 = n6410 & n6415;
  assign n6417 = n6416 ^ n6410;
  assign n6605 = n6604 ^ n6417;
  assign n6786 = n6411 & ~n6412;
  assign n6787 = ~n6406 & n6604;
  assign n6788 = ~n6786 & ~n6787;
  assign n6789 = ~n6218 & ~n6788;
  assign n6790 = ~n6411 & n6412;
  assign n6791 = ~n6409 & ~n6604;
  assign n6792 = ~n6790 & ~n6791;
  assign n6793 = ~n6789 & ~n6792;
  assign n6773 = n6452 ^ n6449;
  assign n6774 = n6456 & ~n6773;
  assign n6775 = n6774 ^ n6455;
  assign n6770 = n6562 ^ n6559;
  assign n6771 = n6566 & ~n6770;
  assign n6772 = n6771 ^ n6565;
  assign n6776 = n6775 ^ n6772;
  assign n6767 = n6441 ^ n6438;
  assign n6768 = n6445 & ~n6767;
  assign n6769 = n6768 ^ n6444;
  assign n6777 = n6776 ^ n6769;
  assign n6764 = n6446 ^ n6435;
  assign n6765 = n6458 & ~n6764;
  assign n6766 = n6765 ^ n6457;
  assign n6778 = n6777 ^ n6766;
  assign n6761 = n6556 ^ n6553;
  assign n6762 = n6568 & ~n6761;
  assign n6763 = n6762 ^ n6567;
  assign n6779 = n6778 ^ n6763;
  assign n6754 = x22 & x43;
  assign n6753 = x21 & x44;
  assign n6755 = n6754 ^ n6753;
  assign n6752 = x8 & x57;
  assign n6756 = n6755 ^ n6752;
  assign n6749 = x7 & x58;
  assign n6748 = x6 & x59;
  assign n6750 = n6749 ^ n6748;
  assign n6747 = x5 & x60;
  assign n6751 = n6750 ^ n6747;
  assign n6757 = n6756 ^ n6751;
  assign n6745 = ~n6589 & n6594;
  assign n6746 = n6745 ^ n6592;
  assign n6758 = n6757 ^ n6746;
  assign n6740 = x29 & x36;
  assign n6739 = x19 & x46;
  assign n6741 = n6740 ^ n6739;
  assign n6738 = x11 & x54;
  assign n6742 = n6741 ^ n6738;
  assign n6735 = x3 & x62;
  assign n6734 = x17 & x48;
  assign n6736 = n6735 ^ n6734;
  assign n6737 = n6736 ^ x33;
  assign n6743 = n6742 ^ n6737;
  assign n6731 = x32 & x33;
  assign n6730 = x31 & x34;
  assign n6732 = n6731 ^ n6730;
  assign n6729 = x30 & x35;
  assign n6733 = n6732 ^ n6729;
  assign n6744 = n6743 ^ n6733;
  assign n6759 = n6758 ^ n6744;
  assign n6724 = x28 & x37;
  assign n6723 = x27 & x38;
  assign n6725 = n6724 ^ n6723;
  assign n6722 = x26 & x39;
  assign n6726 = n6725 ^ n6722;
  assign n6719 = x25 & x40;
  assign n6718 = x24 & x41;
  assign n6720 = n6719 ^ n6718;
  assign n6721 = n6720 ^ n3436;
  assign n6727 = n6726 ^ n6721;
  assign n6715 = x20 & x45;
  assign n6714 = x10 & x55;
  assign n6716 = n6715 ^ n6714;
  assign n6713 = x9 & x56;
  assign n6717 = n6716 ^ n6713;
  assign n6728 = n6727 ^ n6717;
  assign n6760 = n6759 ^ n6728;
  assign n6780 = n6779 ^ n6760;
  assign n6710 = n6459 ^ n6429;
  assign n6711 = ~n6460 & ~n6710;
  assign n6712 = n6711 ^ n6429;
  assign n6781 = n6780 ^ n6712;
  assign n6702 = x2 & x63;
  assign n6701 = x4 & x61;
  assign n6703 = n6702 ^ n6701;
  assign n6698 = n6471 ^ n6470;
  assign n6699 = n6473 & ~n6698;
  assign n6700 = n6699 ^ n6472;
  assign n6704 = n6703 ^ n6700;
  assign n6694 = x18 & x47;
  assign n6693 = x13 & x52;
  assign n6695 = n6694 ^ n6693;
  assign n6692 = x12 & x53;
  assign n6696 = n6695 ^ n6692;
  assign n6689 = x16 & x49;
  assign n6688 = x15 & x50;
  assign n6690 = n6689 ^ n6688;
  assign n6687 = x14 & x51;
  assign n6691 = n6690 ^ n6687;
  assign n6697 = n6696 ^ n6691;
  assign n6705 = n6704 ^ n6697;
  assign n6684 = n6524 ^ n6512;
  assign n6685 = ~n6513 & ~n6684;
  assign n6686 = n6685 ^ n6524;
  assign n6706 = n6705 ^ n6686;
  assign n6681 = n6538 ^ n6535;
  assign n6682 = n6542 & ~n6681;
  assign n6683 = n6682 ^ n6541;
  assign n6707 = n6706 ^ n6683;
  assign n6674 = n6582 ^ n6581;
  assign n6675 = n6584 & ~n6674;
  assign n6676 = n6675 ^ n6583;
  assign n6671 = n6481 ^ n6480;
  assign n6672 = n6483 & ~n6671;
  assign n6673 = n6672 ^ n6482;
  assign n6677 = n6676 ^ n6673;
  assign n6668 = n6487 ^ n3238;
  assign n6669 = n6488 & ~n6668;
  assign n6670 = n6669 ^ n3200;
  assign n6678 = n6677 ^ n6670;
  assign n6665 = n6494 ^ n6489;
  assign n6666 = n6500 & ~n6665;
  assign n6667 = n6666 ^ n6499;
  assign n6679 = n6678 ^ n6667;
  assign n6662 = n6479 ^ n6474;
  assign n6663 = n6485 & ~n6662;
  assign n6664 = n6663 ^ n6484;
  assign n6680 = n6679 ^ n6664;
  assign n6708 = n6707 ^ n6680;
  assign n6659 = n6543 ^ n6529;
  assign n6660 = n6544 & ~n6659;
  assign n6661 = n6660 ^ n6532;
  assign n6709 = n6708 ^ n6661;
  assign n6782 = n6781 ^ n6709;
  assign n6656 = n6461 ^ n6423;
  assign n6657 = ~n6462 & n6656;
  assign n6658 = n6657 ^ n6426;
  assign n6783 = n6782 ^ n6658;
  assign n6653 = n6602 ^ n6420;
  assign n6654 = n6603 & n6653;
  assign n6655 = n6654 ^ n6420;
  assign n6784 = n6783 ^ n6655;
  assign n6641 = n6509 ^ n6508;
  assign n6642 = n6511 & ~n6641;
  assign n6643 = n6642 ^ n6510;
  assign n6638 = n6504 ^ n6503;
  assign n6639 = n6506 & ~n6638;
  assign n6640 = n6639 ^ n6505;
  assign n6644 = n6643 ^ n6640;
  assign n6635 = n6476 ^ n6475;
  assign n6636 = n6478 & ~n6635;
  assign n6637 = n6636 ^ n6477;
  assign n6645 = n6644 ^ n6637;
  assign n6632 = n6595 ^ n6585;
  assign n6633 = ~n6586 & n6632;
  assign n6634 = n6633 ^ n6595;
  assign n6646 = n6645 ^ n6634;
  assign n6627 = n6577 ^ n6576;
  assign n6628 = n6579 & ~n6627;
  assign n6629 = n6628 ^ n6578;
  assign n6624 = n6496 ^ n6495;
  assign n6625 = n6498 & ~n6624;
  assign n6626 = n6625 ^ n6497;
  assign n6630 = n6629 ^ n6626;
  assign n6621 = n6491 ^ n6490;
  assign n6622 = n6493 & ~n6621;
  assign n6623 = n6622 ^ n6492;
  assign n6631 = n6630 ^ n6623;
  assign n6647 = n6646 ^ n6631;
  assign n6618 = n6525 ^ n6501;
  assign n6619 = ~n6502 & ~n6618;
  assign n6620 = n6619 ^ n6525;
  assign n6648 = n6647 ^ n6620;
  assign n6615 = n6596 ^ n6572;
  assign n6616 = n6597 & ~n6615;
  assign n6617 = n6616 ^ n6575;
  assign n6649 = n6648 ^ n6617;
  assign n6612 = n6545 ^ n6469;
  assign n6613 = n6546 & n6612;
  assign n6614 = n6613 ^ n6469;
  assign n6650 = n6649 ^ n6614;
  assign n6609 = n6598 ^ n6550;
  assign n6610 = ~n6599 & n6609;
  assign n6611 = n6610 ^ n6550;
  assign n6651 = n6650 ^ n6611;
  assign n6606 = n6600 ^ n6466;
  assign n6607 = n6601 & ~n6606;
  assign n6608 = n6607 ^ n6466;
  assign n6652 = n6651 ^ n6608;
  assign n6785 = n6784 ^ n6652;
  assign n6794 = n6793 ^ n6785;
  assign n6972 = n6655 & n6783;
  assign n6973 = n6608 & n6651;
  assign n6974 = ~n6972 & n6973;
  assign n6975 = ~n6655 & ~n6783;
  assign n6976 = ~n6608 & ~n6651;
  assign n6977 = n6975 & ~n6976;
  assign n6978 = ~n6974 & ~n6977;
  assign n6979 = ~n6793 & ~n6978;
  assign n6980 = n6783 ^ n6608;
  assign n6981 = ~n6652 & n6980;
  assign n6982 = ~n6784 & n6981;
  assign n6983 = ~n6979 & ~n6982;
  assign n6984 = n6972 & ~n6973;
  assign n6985 = ~n6975 & n6976;
  assign n6986 = ~n6984 & ~n6985;
  assign n6987 = n6793 & ~n6986;
  assign n6988 = n6983 & ~n6987;
  assign n6959 = n6640 ^ n6637;
  assign n6960 = n6644 & ~n6959;
  assign n6961 = n6960 ^ n6643;
  assign n6956 = n6673 ^ n6670;
  assign n6957 = n6677 & ~n6956;
  assign n6958 = n6957 ^ n6676;
  assign n6962 = n6961 ^ n6958;
  assign n6953 = n6626 ^ n6623;
  assign n6954 = n6630 & ~n6953;
  assign n6955 = n6954 ^ n6629;
  assign n6963 = n6962 ^ n6955;
  assign n6950 = n6667 ^ n6664;
  assign n6951 = n6679 & ~n6950;
  assign n6952 = n6951 ^ n6678;
  assign n6964 = n6963 ^ n6952;
  assign n6947 = n6645 ^ n6631;
  assign n6948 = n6646 & ~n6947;
  assign n6949 = n6948 ^ n6634;
  assign n6965 = n6964 ^ n6949;
  assign n6940 = x18 & x48;
  assign n6939 = x15 & x51;
  assign n6941 = n6940 ^ n6939;
  assign n6938 = x13 & x53;
  assign n6942 = n6941 ^ n6938;
  assign n6935 = x31 & x35;
  assign n6934 = x30 & x36;
  assign n6936 = n6935 ^ n6934;
  assign n6933 = x14 & x52;
  assign n6937 = n6936 ^ n6933;
  assign n6943 = n6942 ^ n6937;
  assign n6930 = x32 & x34;
  assign n6929 = x17 & x49;
  assign n6931 = n6930 ^ n6929;
  assign n6928 = x16 & x50;
  assign n6932 = n6931 ^ n6928;
  assign n6944 = n6943 ^ n6932;
  assign n6923 = x19 & x47;
  assign n6922 = x12 & x54;
  assign n6924 = n6923 ^ n6922;
  assign n6921 = x11 & x55;
  assign n6925 = n6924 ^ n6921;
  assign n6918 = x29 & x37;
  assign n6917 = x28 & x38;
  assign n6919 = n6918 ^ n6917;
  assign n6916 = x27 & x39;
  assign n6920 = n6919 ^ n6916;
  assign n6926 = n6925 ^ n6920;
  assign n6913 = x5 & x61;
  assign n6912 = x4 & x62;
  assign n6914 = n6913 ^ n6912;
  assign n6911 = x3 & x63;
  assign n6915 = n6914 ^ n6911;
  assign n6927 = n6926 ^ n6915;
  assign n6945 = n6944 ^ n6927;
  assign n6906 = x22 & x44;
  assign n6905 = x21 & x45;
  assign n6907 = n6906 ^ n6905;
  assign n6904 = x20 & x46;
  assign n6908 = n6907 ^ n6904;
  assign n6901 = x26 & x40;
  assign n6900 = x25 & x41;
  assign n6902 = n6901 ^ n6900;
  assign n6899 = x10 & x56;
  assign n6903 = n6902 ^ n6899;
  assign n6909 = n6908 ^ n6903;
  assign n6896 = x23 & x43;
  assign n6895 = x24 & x42;
  assign n6897 = n6896 ^ n6895;
  assign n6894 = x9 & x57;
  assign n6898 = n6897 ^ n6894;
  assign n6910 = n6909 ^ n6898;
  assign n6946 = n6945 ^ n6910;
  assign n6966 = n6965 ^ n6946;
  assign n6891 = n6647 ^ n6617;
  assign n6892 = n6648 & n6891;
  assign n6893 = n6892 ^ n6617;
  assign n6967 = n6966 ^ n6893;
  assign n6888 = n6779 ^ n6712;
  assign n6889 = ~n6780 & ~n6888;
  assign n6890 = n6889 ^ n6712;
  assign n6968 = n6967 ^ n6890;
  assign n6885 = n6649 ^ n6611;
  assign n6886 = n6650 & ~n6885;
  assign n6887 = n6886 ^ n6611;
  assign n6969 = n6968 ^ n6887;
  assign n6874 = n6714 ^ n6713;
  assign n6875 = n6716 & ~n6874;
  assign n6876 = n6875 ^ n6715;
  assign n6871 = n6693 ^ n6692;
  assign n6872 = n6695 & ~n6871;
  assign n6873 = n6872 ^ n6694;
  assign n6877 = n6876 ^ n6873;
  assign n6868 = n6719 ^ n3436;
  assign n6869 = ~n6720 & n6868;
  assign n6870 = n6869 ^ n3436;
  assign n6878 = n6877 ^ n6870;
  assign n6865 = n6721 ^ n6717;
  assign n6866 = n6727 & ~n6865;
  assign n6867 = n6866 ^ n6726;
  assign n6879 = n6878 ^ n6867;
  assign n6862 = n6756 ^ n6746;
  assign n6863 = ~n6757 & n6862;
  assign n6864 = n6863 ^ n6746;
  assign n6880 = n6879 ^ n6864;
  assign n6859 = n6744 ^ n6728;
  assign n6860 = n6759 & ~n6859;
  assign n6861 = n6860 ^ n6758;
  assign n6881 = n6880 ^ n6861;
  assign n6856 = n6686 ^ n6683;
  assign n6857 = n6706 & ~n6856;
  assign n6858 = n6857 ^ n6683;
  assign n6882 = n6881 ^ n6858;
  assign n6847 = n6700 & n6703;
  assign n6848 = x4 & x63;
  assign n6849 = n6290 & n6848;
  assign n6850 = ~n6847 & ~n6849;
  assign n6843 = x8 & x58;
  assign n6842 = x7 & x59;
  assign n6844 = n6843 ^ n6842;
  assign n6841 = x6 & x60;
  assign n6845 = n6844 ^ n6841;
  assign n6838 = n6723 ^ n6722;
  assign n6839 = n6725 & ~n6838;
  assign n6840 = n6839 ^ n6724;
  assign n6846 = n6845 ^ n6840;
  assign n6851 = n6850 ^ n6846;
  assign n6835 = n6704 ^ n6696;
  assign n6836 = ~n6697 & n6835;
  assign n6837 = n6836 ^ n6704;
  assign n6852 = n6851 ^ n6837;
  assign n6832 = n6772 ^ n6769;
  assign n6833 = n6776 & ~n6832;
  assign n6834 = n6833 ^ n6775;
  assign n6853 = n6852 ^ n6834;
  assign n6825 = n6688 ^ n6687;
  assign n6826 = n6690 & ~n6825;
  assign n6827 = n6826 ^ n6689;
  assign n6822 = n6730 ^ n6729;
  assign n6823 = n6732 & ~n6822;
  assign n6824 = n6823 ^ n6731;
  assign n6828 = n6827 ^ n6824;
  assign n6818 = x48 & n3990;
  assign n6819 = ~n6735 & ~n6818;
  assign n6820 = ~x33 & ~n6734;
  assign n6821 = ~n6819 & ~n6820;
  assign n6829 = n6828 ^ n6821;
  assign n6813 = n6739 ^ n6738;
  assign n6814 = n6741 & ~n6813;
  assign n6815 = n6814 ^ n6740;
  assign n6810 = n6753 ^ n6752;
  assign n6811 = n6755 & ~n6810;
  assign n6812 = n6811 ^ n6754;
  assign n6816 = n6815 ^ n6812;
  assign n6807 = n6748 ^ n6747;
  assign n6808 = n6750 & ~n6807;
  assign n6809 = n6808 ^ n6749;
  assign n6817 = n6816 ^ n6809;
  assign n6830 = n6829 ^ n6817;
  assign n6804 = n6737 ^ n6733;
  assign n6805 = n6743 & ~n6804;
  assign n6806 = n6805 ^ n6742;
  assign n6831 = n6830 ^ n6806;
  assign n6854 = n6853 ^ n6831;
  assign n6801 = n6777 ^ n6763;
  assign n6802 = n6778 & ~n6801;
  assign n6803 = n6802 ^ n6766;
  assign n6855 = n6854 ^ n6803;
  assign n6883 = n6882 ^ n6855;
  assign n6798 = n6707 ^ n6661;
  assign n6799 = n6708 & ~n6798;
  assign n6800 = n6799 ^ n6661;
  assign n6884 = n6883 ^ n6800;
  assign n6970 = n6969 ^ n6884;
  assign n6795 = n6781 ^ n6658;
  assign n6796 = ~n6782 & ~n6795;
  assign n6797 = n6796 ^ n6658;
  assign n6971 = n6970 ^ n6797;
  assign n6989 = n6988 ^ n6971;
  assign n7164 = ~n6971 & ~n6972;
  assign n7165 = ~n6985 & n7164;
  assign n7166 = n6971 & ~n6975;
  assign n7167 = n6973 & ~n7166;
  assign n7168 = ~n7165 & ~n7167;
  assign n7169 = n6793 & n7168;
  assign n7170 = n6976 & ~n7164;
  assign n7171 = ~n6974 & n7166;
  assign n7172 = ~n7170 & ~n7171;
  assign n7173 = ~n7169 & n7172;
  assign n7150 = n6873 ^ n6870;
  assign n7151 = n6877 & ~n7150;
  assign n7152 = n7151 ^ n6876;
  assign n7147 = n6812 ^ n6809;
  assign n7148 = n6816 & ~n7147;
  assign n7149 = n7148 ^ n6815;
  assign n7153 = n7152 ^ n7149;
  assign n7144 = n6824 ^ n6821;
  assign n7145 = n6828 & ~n7144;
  assign n7146 = n7145 ^ n6827;
  assign n7154 = n7153 ^ n7146;
  assign n7141 = n6817 ^ n6806;
  assign n7142 = n6830 & ~n7141;
  assign n7143 = n7142 ^ n6829;
  assign n7155 = n7154 ^ n7143;
  assign n7138 = n6867 ^ n6864;
  assign n7139 = ~n6879 & n7138;
  assign n7140 = n7139 ^ n6864;
  assign n7156 = n7155 ^ n7140;
  assign n7131 = x26 & x41;
  assign n7130 = x25 & x42;
  assign n7132 = n7131 ^ n7130;
  assign n7129 = x21 & x46;
  assign n7133 = n7132 ^ n7129;
  assign n7126 = x19 & x48;
  assign n7125 = x17 & x50;
  assign n7127 = n7126 ^ n7125;
  assign n7124 = x14 & x53;
  assign n7128 = n7127 ^ n7124;
  assign n7134 = n7133 ^ n7128;
  assign n7121 = x28 & x39;
  assign n7120 = x27 & x40;
  assign n7122 = n7121 ^ n7120;
  assign n7123 = n7122 ^ n6848;
  assign n7135 = n7134 ^ n7123;
  assign n7115 = x33 & x34;
  assign n7114 = x32 & x35;
  assign n7116 = n7115 ^ n7114;
  assign n7113 = x31 & x36;
  assign n7117 = n7116 ^ n7113;
  assign n7110 = x5 & x62;
  assign n7109 = x18 & x49;
  assign n7111 = n7110 ^ n7109;
  assign n7112 = n7111 ^ x34;
  assign n7118 = n7117 ^ n7112;
  assign n7106 = x29 & x38;
  assign n7105 = x13 & x54;
  assign n7107 = n7106 ^ n7105;
  assign n7104 = x12 & x55;
  assign n7108 = n7107 ^ n7104;
  assign n7119 = n7118 ^ n7108;
  assign n7136 = n7135 ^ n7119;
  assign n7099 = x9 & x58;
  assign n7098 = x8 & x59;
  assign n7100 = n7099 ^ n7098;
  assign n7097 = x7 & x60;
  assign n7101 = n7100 ^ n7097;
  assign n7094 = x24 & x43;
  assign n7095 = n7094 ^ n3432;
  assign n7093 = x22 & x45;
  assign n7096 = n7095 ^ n7093;
  assign n7102 = n7101 ^ n7096;
  assign n7090 = x30 & x37;
  assign n7089 = x16 & x51;
  assign n7091 = n7090 ^ n7089;
  assign n7088 = x15 & x52;
  assign n7092 = n7091 ^ n7088;
  assign n7103 = n7102 ^ n7092;
  assign n7137 = n7136 ^ n7103;
  assign n7157 = n7156 ^ n7137;
  assign n7085 = n6861 ^ n6858;
  assign n7086 = ~n6881 & n7085;
  assign n7087 = n7086 ^ n6858;
  assign n7158 = n7157 ^ n7087;
  assign n7082 = n6965 ^ n6893;
  assign n7083 = ~n6966 & n7082;
  assign n7084 = n7083 ^ n6893;
  assign n7159 = n7158 ^ n7084;
  assign n7079 = n6882 ^ n6800;
  assign n7080 = n6883 & n7079;
  assign n7081 = n7080 ^ n6800;
  assign n7160 = n7159 ^ n7081;
  assign n7070 = n6850 ^ n6840;
  assign n7071 = ~n6846 & ~n7070;
  assign n7072 = n7071 ^ n6850;
  assign n7067 = n6920 ^ n6915;
  assign n7068 = n6926 & ~n7067;
  assign n7069 = n7068 ^ n6925;
  assign n7073 = n7072 ^ n7069;
  assign n7064 = n6903 ^ n6898;
  assign n7065 = n6909 & ~n7064;
  assign n7066 = n7065 ^ n6908;
  assign n7074 = n7073 ^ n7066;
  assign n7057 = n6917 ^ n6916;
  assign n7058 = n6919 & ~n7057;
  assign n7059 = n7058 ^ n6918;
  assign n7054 = n6912 ^ n6911;
  assign n7055 = n6914 & ~n7054;
  assign n7056 = n7055 ^ n6913;
  assign n7060 = n7059 ^ n7056;
  assign n7051 = n6842 ^ n6841;
  assign n7052 = n6844 & ~n7051;
  assign n7053 = n7052 ^ n6843;
  assign n7061 = n7060 ^ n7053;
  assign n7048 = x6 & x61;
  assign n7045 = n6929 ^ n6928;
  assign n7046 = n6931 & ~n7045;
  assign n7047 = n7046 ^ n6930;
  assign n7049 = n7048 ^ n7047;
  assign n7042 = n6934 ^ n6933;
  assign n7043 = n6936 & ~n7042;
  assign n7044 = n7043 ^ n6935;
  assign n7050 = n7049 ^ n7044;
  assign n7062 = n7061 ^ n7050;
  assign n7037 = n6905 ^ n6904;
  assign n7038 = n6907 & ~n7037;
  assign n7039 = n7038 ^ n6906;
  assign n7034 = n6895 ^ n6894;
  assign n7035 = n6897 & ~n7034;
  assign n7036 = n7035 ^ n6896;
  assign n7040 = n7039 ^ n7036;
  assign n7031 = n6900 ^ n6899;
  assign n7032 = n6902 & ~n7031;
  assign n7033 = n7032 ^ n6901;
  assign n7041 = n7040 ^ n7033;
  assign n7063 = n7062 ^ n7041;
  assign n7075 = n7074 ^ n7063;
  assign n7028 = n6952 ^ n6949;
  assign n7029 = ~n6964 & n7028;
  assign n7030 = n7029 ^ n6949;
  assign n7076 = n7075 ^ n7030;
  assign n7019 = x20 & x47;
  assign n7018 = x11 & x56;
  assign n7020 = n7019 ^ n7018;
  assign n7017 = x10 & x57;
  assign n7021 = n7020 ^ n7017;
  assign n7014 = n6922 ^ n6921;
  assign n7015 = n6924 & ~n7014;
  assign n7016 = n7015 ^ n6923;
  assign n7022 = n7021 ^ n7016;
  assign n7011 = n6939 ^ n6938;
  assign n7012 = n6941 & ~n7011;
  assign n7013 = n7012 ^ n6940;
  assign n7023 = n7022 ^ n7013;
  assign n7008 = n6937 ^ n6932;
  assign n7009 = n6943 & ~n7008;
  assign n7010 = n7009 ^ n6942;
  assign n7024 = n7023 ^ n7010;
  assign n7005 = n6958 ^ n6955;
  assign n7006 = n6962 & ~n7005;
  assign n7007 = n7006 ^ n6961;
  assign n7025 = n7024 ^ n7007;
  assign n7002 = n6927 ^ n6910;
  assign n7003 = n6945 & ~n7002;
  assign n7004 = n7003 ^ n6944;
  assign n7026 = n7025 ^ n7004;
  assign n6999 = n6837 ^ n6834;
  assign n7000 = n6852 & n6999;
  assign n7001 = n7000 ^ n6834;
  assign n7027 = n7026 ^ n7001;
  assign n7077 = n7076 ^ n7027;
  assign n6996 = n6831 ^ n6803;
  assign n6997 = ~n6854 & ~n6996;
  assign n6998 = n6997 ^ n6853;
  assign n7078 = n7077 ^ n6998;
  assign n7161 = n7160 ^ n7078;
  assign n6993 = n6890 ^ n6887;
  assign n6994 = n6968 & ~n6993;
  assign n6995 = n6994 ^ n6887;
  assign n7162 = n7161 ^ n6995;
  assign n6990 = n6969 ^ n6797;
  assign n6991 = ~n6970 & ~n6990;
  assign n6992 = n6991 ^ n6797;
  assign n7163 = n7162 ^ n6992;
  assign n7174 = n7173 ^ n7163;
  assign n7340 = n7069 ^ n7066;
  assign n7341 = ~n7073 & ~n7340;
  assign n7342 = n7341 ^ n7072;
  assign n7337 = n7050 ^ n7041;
  assign n7338 = n7062 & ~n7337;
  assign n7339 = n7338 ^ n7061;
  assign n7343 = n7342 ^ n7339;
  assign n7334 = n7010 ^ n7007;
  assign n7335 = ~n7024 & n7334;
  assign n7336 = n7335 ^ n7007;
  assign n7344 = n7343 ^ n7336;
  assign n7327 = x33 & x35;
  assign n7326 = x19 & x49;
  assign n7328 = n7327 ^ n7326;
  assign n7325 = x18 & x50;
  assign n7329 = n7328 ^ n7325;
  assign n7322 = x17 & x51;
  assign n7321 = x13 & x55;
  assign n7323 = n7322 ^ n7321;
  assign n7320 = x12 & x56;
  assign n7324 = n7323 ^ n7320;
  assign n7330 = n7329 ^ n7324;
  assign n7317 = x32 & x36;
  assign n7316 = x31 & x37;
  assign n7318 = n7317 ^ n7316;
  assign n7315 = x30 & x38;
  assign n7319 = n7318 ^ n7315;
  assign n7331 = n7330 ^ n7319;
  assign n7310 = x16 & x52;
  assign n7309 = x15 & x53;
  assign n7311 = n7310 ^ n7309;
  assign n7308 = x14 & x54;
  assign n7312 = n7311 ^ n7308;
  assign n7305 = x26 & x42;
  assign n7304 = x25 & x43;
  assign n7306 = n7305 ^ n7304;
  assign n7303 = x24 & x44;
  assign n7307 = n7306 ^ n7303;
  assign n7313 = n7312 ^ n7307;
  assign n7300 = x23 & x45;
  assign n7299 = x22 & x46;
  assign n7301 = n7300 ^ n7299;
  assign n7298 = x20 & x48;
  assign n7302 = n7301 ^ n7298;
  assign n7314 = n7313 ^ n7302;
  assign n7332 = n7331 ^ n7314;
  assign n7293 = x29 & x39;
  assign n7292 = x28 & x40;
  assign n7294 = n7293 ^ n7292;
  assign n7291 = x27 & x41;
  assign n7295 = n7294 ^ n7291;
  assign n7288 = x21 & x47;
  assign n7287 = x6 & x62;
  assign n7289 = n7288 ^ n7287;
  assign n7286 = x5 & x63;
  assign n7290 = n7289 ^ n7286;
  assign n7296 = n7295 ^ n7290;
  assign n7283 = x11 & x57;
  assign n7282 = x10 & x58;
  assign n7284 = n7283 ^ n7282;
  assign n7281 = x9 & x59;
  assign n7285 = n7284 ^ n7281;
  assign n7297 = n7296 ^ n7285;
  assign n7333 = n7332 ^ n7297;
  assign n7345 = n7344 ^ n7333;
  assign n7278 = n7004 ^ n7001;
  assign n7279 = n7026 & ~n7278;
  assign n7280 = n7279 ^ n7025;
  assign n7346 = n7345 ^ n7280;
  assign n7275 = n7156 ^ n7087;
  assign n7276 = ~n7157 & n7275;
  assign n7277 = n7276 ^ n7087;
  assign n7347 = n7346 ^ n7277;
  assign n7272 = n7027 ^ n6998;
  assign n7273 = ~n7077 & n7272;
  assign n7274 = n7273 ^ n7076;
  assign n7348 = n7347 ^ n7274;
  assign n7261 = n7098 ^ n7097;
  assign n7262 = n7100 & ~n7261;
  assign n7263 = n7262 ^ n7099;
  assign n7258 = n7094 ^ n7093;
  assign n7259 = n7095 & ~n7258;
  assign n7260 = n7259 ^ n3432;
  assign n7264 = n7263 ^ n7260;
  assign n7255 = n7018 ^ n7017;
  assign n7256 = n7020 & ~n7255;
  assign n7257 = n7256 ^ n7019;
  assign n7265 = n7264 ^ n7257;
  assign n7250 = n7089 ^ n7088;
  assign n7251 = n7091 & ~n7250;
  assign n7252 = n7251 ^ n7090;
  assign n7247 = n7114 ^ n7113;
  assign n7248 = n7116 & ~n7247;
  assign n7249 = n7248 ^ n7115;
  assign n7253 = n7252 ^ n7249;
  assign n7244 = n7121 ^ n6848;
  assign n7245 = ~n7122 & n7244;
  assign n7246 = n7245 ^ n6848;
  assign n7254 = n7253 ^ n7246;
  assign n7266 = n7265 ^ n7254;
  assign n7241 = n7149 ^ n7146;
  assign n7242 = n7153 & ~n7241;
  assign n7243 = n7242 ^ n7152;
  assign n7267 = n7266 ^ n7243;
  assign n7234 = n7105 ^ n7104;
  assign n7235 = n7107 & ~n7234;
  assign n7236 = n7235 ^ n7106;
  assign n7231 = n7130 ^ n7129;
  assign n7232 = n7132 & ~n7231;
  assign n7233 = n7232 ^ n7131;
  assign n7237 = n7236 ^ n7233;
  assign n7228 = n7125 ^ n7124;
  assign n7229 = n7127 & ~n7228;
  assign n7230 = n7229 ^ n7126;
  assign n7238 = n7237 ^ n7230;
  assign n7225 = n7112 ^ n7108;
  assign n7226 = n7118 & ~n7225;
  assign n7227 = n7226 ^ n7117;
  assign n7239 = n7238 ^ n7227;
  assign n7222 = n7128 ^ n7123;
  assign n7223 = n7134 & ~n7222;
  assign n7224 = n7223 ^ n7133;
  assign n7240 = n7239 ^ n7224;
  assign n7268 = n7267 ^ n7240;
  assign n7219 = n7154 ^ n7140;
  assign n7220 = ~n7155 & n7219;
  assign n7221 = n7220 ^ n7140;
  assign n7269 = n7268 ^ n7221;
  assign n7212 = n7021 ^ n7013;
  assign n7213 = n7022 & ~n7212;
  assign n7214 = n7213 ^ n7016;
  assign n7209 = n7096 ^ n7092;
  assign n7210 = n7102 & ~n7209;
  assign n7211 = n7210 ^ n7101;
  assign n7215 = n7214 ^ n7211;
  assign n7206 = n7036 ^ n7033;
  assign n7207 = n7040 & ~n7206;
  assign n7208 = n7207 ^ n7039;
  assign n7216 = n7215 ^ n7208;
  assign n7203 = n7119 ^ n7103;
  assign n7204 = n7136 & ~n7203;
  assign n7205 = n7204 ^ n7135;
  assign n7217 = n7216 ^ n7205;
  assign n7196 = x49 & n4296;
  assign n7197 = ~n7110 & ~n7196;
  assign n7198 = ~x34 & ~n7109;
  assign n7199 = ~n7197 & ~n7198;
  assign n7194 = x7 & x61;
  assign n7193 = x8 & x60;
  assign n7195 = n7194 ^ n7193;
  assign n7200 = n7199 ^ n7195;
  assign n7190 = n7056 ^ n7053;
  assign n7191 = n7060 & ~n7190;
  assign n7192 = n7191 ^ n7059;
  assign n7201 = n7200 ^ n7192;
  assign n7187 = n7048 ^ n7044;
  assign n7188 = n7049 & ~n7187;
  assign n7189 = n7188 ^ n7047;
  assign n7202 = n7201 ^ n7189;
  assign n7218 = n7217 ^ n7202;
  assign n7270 = n7269 ^ n7218;
  assign n7184 = n7074 ^ n7030;
  assign n7185 = n7075 & ~n7184;
  assign n7186 = n7185 ^ n7030;
  assign n7271 = n7270 ^ n7186;
  assign n7349 = n7348 ^ n7271;
  assign n7181 = n7084 ^ n7081;
  assign n7182 = ~n7159 & n7181;
  assign n7183 = n7182 ^ n7081;
  assign n7350 = n7349 ^ n7183;
  assign n7178 = n7160 ^ n6995;
  assign n7179 = ~n7161 & n7178;
  assign n7180 = n7179 ^ n6995;
  assign n7351 = n7350 ^ n7180;
  assign n7175 = n7173 ^ n6992;
  assign n7176 = ~n7163 & ~n7175;
  assign n7177 = n7176 ^ n7173;
  assign n7352 = n7351 ^ n7177;
  assign n7519 = ~n7271 & ~n7348;
  assign n7520 = ~n7183 & n7519;
  assign n7521 = ~n7180 & n7520;
  assign n7522 = ~n7177 & ~n7521;
  assign n7523 = n7348 ^ n7183;
  assign n7524 = ~n7349 & n7523;
  assign n7525 = n7524 ^ n7183;
  assign n7526 = ~n7180 & ~n7525;
  assign n7527 = ~n7520 & ~n7526;
  assign n7528 = ~n7522 & ~n7527;
  assign n7529 = n7271 & n7348;
  assign n7530 = n7183 & n7529;
  assign n7531 = ~n7180 & ~n7530;
  assign n7532 = n7525 & ~n7531;
  assign n7533 = ~n7177 & n7532;
  assign n7534 = n7180 & n7530;
  assign n7535 = ~n7533 & ~n7534;
  assign n7536 = ~n7528 & n7535;
  assign n7508 = n7233 ^ n7230;
  assign n7509 = n7237 & ~n7508;
  assign n7510 = n7509 ^ n7236;
  assign n7505 = n7249 ^ n7246;
  assign n7506 = n7253 & ~n7505;
  assign n7507 = n7506 ^ n7252;
  assign n7511 = n7510 ^ n7507;
  assign n7500 = n7292 ^ n7291;
  assign n7501 = n7294 & ~n7500;
  assign n7502 = n7501 ^ n7293;
  assign n7497 = n7321 ^ n7320;
  assign n7498 = n7323 & ~n7497;
  assign n7499 = n7498 ^ n7322;
  assign n7503 = n7502 ^ n7499;
  assign n7494 = n7304 ^ n7303;
  assign n7495 = n7306 & ~n7494;
  assign n7496 = n7495 ^ n7305;
  assign n7504 = n7503 ^ n7496;
  assign n7512 = n7511 ^ n7504;
  assign n7491 = n7314 ^ n7297;
  assign n7492 = n7332 & ~n7491;
  assign n7493 = n7492 ^ n7331;
  assign n7513 = n7512 ^ n7493;
  assign n7488 = n7265 ^ n7243;
  assign n7489 = ~n7266 & n7488;
  assign n7490 = n7489 ^ n7243;
  assign n7514 = n7513 ^ n7490;
  assign n7485 = n7267 ^ n7221;
  assign n7486 = ~n7268 & n7485;
  assign n7487 = n7486 ^ n7221;
  assign n7515 = n7514 ^ n7487;
  assign n7478 = n7324 ^ n7319;
  assign n7479 = n7330 & ~n7478;
  assign n7480 = n7479 ^ n7329;
  assign n7475 = n7307 ^ n7302;
  assign n7476 = n7313 & ~n7475;
  assign n7477 = n7476 ^ n7312;
  assign n7481 = n7480 ^ n7477;
  assign n7472 = n7200 ^ n7189;
  assign n7473 = n7201 & ~n7472;
  assign n7474 = n7473 ^ n7192;
  assign n7482 = n7481 ^ n7474;
  assign n7465 = n7287 ^ n7286;
  assign n7466 = n7289 & ~n7465;
  assign n7467 = n7466 ^ n7288;
  assign n7462 = n7282 ^ n7281;
  assign n7463 = n7284 & ~n7462;
  assign n7464 = n7463 ^ n7283;
  assign n7468 = n7467 ^ n7464;
  assign n7459 = n7299 ^ n7298;
  assign n7460 = n7301 & ~n7459;
  assign n7461 = n7460 ^ n7300;
  assign n7469 = n7468 ^ n7461;
  assign n7454 = n7316 ^ n7315;
  assign n7455 = n7318 & ~n7454;
  assign n7456 = n7455 ^ n7317;
  assign n7451 = n7326 ^ n7325;
  assign n7452 = n7328 & ~n7451;
  assign n7453 = n7452 ^ n7327;
  assign n7457 = n7456 ^ n7453;
  assign n7448 = n7309 ^ n7308;
  assign n7449 = n7311 & ~n7448;
  assign n7450 = n7449 ^ n7310;
  assign n7458 = n7457 ^ n7450;
  assign n7470 = n7469 ^ n7458;
  assign n7445 = n7290 ^ n7285;
  assign n7446 = n7296 & ~n7445;
  assign n7447 = n7446 ^ n7295;
  assign n7471 = n7470 ^ n7447;
  assign n7483 = n7482 ^ n7471;
  assign n7442 = n7339 ^ n7336;
  assign n7443 = ~n7343 & ~n7442;
  assign n7444 = n7443 ^ n7342;
  assign n7484 = n7483 ^ n7444;
  assign n7516 = n7515 ^ n7484;
  assign n7439 = n7346 ^ n7274;
  assign n7440 = ~n7347 & ~n7439;
  assign n7441 = n7440 ^ n7277;
  assign n7517 = n7516 ^ n7441;
  assign n7428 = x10 & x59;
  assign n7427 = x9 & x60;
  assign n7429 = n7428 ^ n7427;
  assign n7426 = x8 & x61;
  assign n7430 = n7429 ^ n7426;
  assign n7423 = x25 & x44;
  assign n7422 = x24 & x45;
  assign n7424 = n7423 ^ n7422;
  assign n7421 = x23 & x46;
  assign n7425 = n7424 ^ n7421;
  assign n7431 = n7430 ^ n7425;
  assign n7418 = x27 & x42;
  assign n7417 = x26 & x43;
  assign n7419 = n7418 ^ n7417;
  assign n7416 = x6 & x63;
  assign n7420 = n7419 ^ n7416;
  assign n7432 = n7431 ^ n7420;
  assign n7413 = n7211 ^ n7208;
  assign n7414 = n7215 & ~n7413;
  assign n7415 = n7414 ^ n7214;
  assign n7433 = n7432 ^ n7415;
  assign n7408 = n7195 & n7199;
  assign n7409 = x60 & x61;
  assign n7410 = n388 & n7409;
  assign n7411 = ~n7408 & ~n7410;
  assign n7404 = x22 & x47;
  assign n7403 = x21 & x48;
  assign n7405 = n7404 ^ n7403;
  assign n7402 = x14 & x55;
  assign n7406 = n7405 ^ n7402;
  assign n7399 = x13 & x56;
  assign n7398 = x12 & x57;
  assign n7400 = n7399 ^ n7398;
  assign n7397 = x11 & x58;
  assign n7401 = n7400 ^ n7397;
  assign n7407 = n7406 ^ n7401;
  assign n7412 = n7411 ^ n7407;
  assign n7434 = n7433 ^ n7412;
  assign n7390 = x30 & x39;
  assign n7389 = x29 & x40;
  assign n7391 = n7390 ^ n7389;
  assign n7388 = x28 & x41;
  assign n7392 = n7391 ^ n7388;
  assign n7385 = x19 & x50;
  assign n7384 = x18 & x51;
  assign n7386 = n7385 ^ n7384;
  assign n7383 = x17 & x52;
  assign n7387 = n7386 ^ n7383;
  assign n7393 = n7392 ^ n7387;
  assign n7380 = n7260 ^ n7257;
  assign n7381 = n7264 & ~n7380;
  assign n7382 = n7381 ^ n7263;
  assign n7394 = n7393 ^ n7382;
  assign n7375 = x20 & x49;
  assign n7374 = x16 & x53;
  assign n7376 = n7375 ^ n7374;
  assign n7373 = x15 & x54;
  assign n7377 = n7376 ^ n7373;
  assign n7370 = x33 & x36;
  assign n7369 = x32 & x37;
  assign n7371 = n7370 ^ n7369;
  assign n7368 = x31 & x38;
  assign n7372 = n7371 ^ n7368;
  assign n7378 = n7377 ^ n7372;
  assign n7366 = x7 & x62;
  assign n7365 = ~x34 & x35;
  assign n7367 = n7366 ^ n7365;
  assign n7379 = n7378 ^ n7367;
  assign n7395 = n7394 ^ n7379;
  assign n7362 = n7227 ^ n7224;
  assign n7363 = n7239 & ~n7362;
  assign n7364 = n7363 ^ n7238;
  assign n7396 = n7395 ^ n7364;
  assign n7435 = n7434 ^ n7396;
  assign n7359 = n7205 ^ n7202;
  assign n7360 = n7217 & ~n7359;
  assign n7361 = n7360 ^ n7216;
  assign n7436 = n7435 ^ n7361;
  assign n7356 = n7333 ^ n7280;
  assign n7357 = ~n7345 & ~n7356;
  assign n7358 = n7357 ^ n7344;
  assign n7437 = n7436 ^ n7358;
  assign n7353 = n7269 ^ n7186;
  assign n7354 = ~n7270 & n7353;
  assign n7355 = n7354 ^ n7186;
  assign n7438 = n7437 ^ n7355;
  assign n7518 = n7517 ^ n7438;
  assign n7537 = n7536 ^ n7518;
  assign n7703 = n7518 & ~n7534;
  assign n7704 = n7527 & ~n7703;
  assign n7705 = n7177 & ~n7704;
  assign n7706 = n7518 & ~n7532;
  assign n7707 = ~n7521 & ~n7706;
  assign n7708 = ~n7705 & n7707;
  assign n7689 = n7384 ^ n7383;
  assign n7690 = n7386 & ~n7689;
  assign n7691 = n7690 ^ n7385;
  assign n7686 = n7374 ^ n7373;
  assign n7687 = n7376 & ~n7686;
  assign n7688 = n7687 ^ n7375;
  assign n7692 = n7691 ^ n7688;
  assign n7683 = x34 & x36;
  assign n7682 = x33 & x37;
  assign n7684 = n7683 ^ n7682;
  assign n7681 = x32 & x38;
  assign n7685 = n7684 ^ n7681;
  assign n7693 = n7692 ^ n7685;
  assign n7678 = n7507 ^ n7504;
  assign n7679 = n7511 & ~n7678;
  assign n7680 = n7679 ^ n7510;
  assign n7694 = n7693 ^ n7680;
  assign n7673 = x11 & x59;
  assign n7672 = x10 & x60;
  assign n7674 = n7673 ^ n7672;
  assign n7671 = x9 & x61;
  assign n7675 = n7674 ^ n7671;
  assign n7668 = x18 & x52;
  assign n7667 = x17 & x53;
  assign n7669 = n7668 ^ n7667;
  assign n7666 = x16 & x54;
  assign n7670 = n7669 ^ n7666;
  assign n7676 = n7675 ^ n7670;
  assign n7663 = x24 & x46;
  assign n7662 = x13 & x57;
  assign n7664 = n7663 ^ n7662;
  assign n7661 = x12 & x58;
  assign n7665 = n7664 ^ n7661;
  assign n7677 = n7676 ^ n7665;
  assign n7695 = n7694 ^ n7677;
  assign n7654 = x28 & x42;
  assign n7655 = n7654 ^ n3924;
  assign n7653 = x7 & x63;
  assign n7656 = n7655 ^ n7653;
  assign n7650 = x31 & x39;
  assign n7649 = x30 & x40;
  assign n7651 = n7650 ^ n7649;
  assign n7648 = x29 & x41;
  assign n7652 = n7651 ^ n7648;
  assign n7657 = n7656 ^ n7652;
  assign n7645 = n7453 ^ n7450;
  assign n7646 = n7457 & ~n7645;
  assign n7647 = n7646 ^ n7456;
  assign n7658 = n7657 ^ n7647;
  assign n7640 = x27 & x43;
  assign n7639 = x26 & x44;
  assign n7641 = n7640 ^ n7639;
  assign n7638 = x25 & x45;
  assign n7642 = n7641 ^ n7638;
  assign n7635 = x21 & x49;
  assign n7634 = x20 & x50;
  assign n7636 = n7635 ^ n7634;
  assign n7633 = x19 & x51;
  assign n7637 = n7636 ^ n7633;
  assign n7643 = n7642 ^ n7637;
  assign n7630 = x22 & x48;
  assign n7629 = x15 & x55;
  assign n7631 = n7630 ^ n7629;
  assign n7628 = x14 & x56;
  assign n7632 = n7631 ^ n7628;
  assign n7644 = n7643 ^ n7632;
  assign n7659 = n7658 ^ n7644;
  assign n7625 = n7458 ^ n7447;
  assign n7626 = n7470 & ~n7625;
  assign n7627 = n7626 ^ n7469;
  assign n7660 = n7659 ^ n7627;
  assign n7696 = n7695 ^ n7660;
  assign n7622 = n7512 ^ n7490;
  assign n7623 = ~n7513 & n7622;
  assign n7624 = n7623 ^ n7490;
  assign n7697 = n7696 ^ n7624;
  assign n7614 = ~x34 & ~n7366;
  assign n7615 = x35 & ~n7614;
  assign n7613 = x8 & x62;
  assign n7616 = n7615 ^ n7613;
  assign n7610 = n7369 ^ n7368;
  assign n7611 = n7371 & ~n7610;
  assign n7612 = n7611 ^ n7370;
  assign n7617 = n7616 ^ n7612;
  assign n7607 = n7392 ^ n7382;
  assign n7608 = ~n7393 & n7607;
  assign n7609 = n7608 ^ n7382;
  assign n7618 = n7617 ^ n7609;
  assign n7602 = n7422 ^ n7421;
  assign n7603 = n7424 & ~n7602;
  assign n7604 = n7603 ^ n7423;
  assign n7599 = n7417 ^ n7416;
  assign n7600 = n7419 & ~n7599;
  assign n7601 = n7600 ^ n7418;
  assign n7605 = n7604 ^ n7601;
  assign n7596 = n7389 ^ n7388;
  assign n7597 = n7391 & ~n7596;
  assign n7598 = n7597 ^ n7390;
  assign n7606 = n7605 ^ n7598;
  assign n7619 = n7618 ^ n7606;
  assign n7591 = n7425 ^ n7420;
  assign n7592 = n7431 & ~n7591;
  assign n7593 = n7592 ^ n7430;
  assign n7588 = n7372 ^ n7367;
  assign n7589 = n7378 & ~n7588;
  assign n7590 = n7589 ^ n7377;
  assign n7594 = n7593 ^ n7590;
  assign n7585 = n7411 ^ n7406;
  assign n7586 = ~n7407 & ~n7585;
  assign n7587 = n7586 ^ n7411;
  assign n7595 = n7594 ^ n7587;
  assign n7620 = n7619 ^ n7595;
  assign n7582 = n7394 ^ n7364;
  assign n7583 = ~n7395 & n7582;
  assign n7584 = n7583 ^ n7364;
  assign n7621 = n7620 ^ n7584;
  assign n7698 = n7697 ^ n7621;
  assign n7579 = n7514 ^ n7484;
  assign n7580 = n7515 & n7579;
  assign n7581 = n7580 ^ n7487;
  assign n7699 = n7698 ^ n7581;
  assign n7570 = n7499 ^ n7496;
  assign n7571 = n7503 & ~n7570;
  assign n7572 = n7571 ^ n7502;
  assign n7567 = n7464 ^ n7461;
  assign n7568 = n7468 & ~n7567;
  assign n7569 = n7568 ^ n7467;
  assign n7573 = n7572 ^ n7569;
  assign n7562 = n7398 ^ n7397;
  assign n7563 = n7400 & ~n7562;
  assign n7564 = n7563 ^ n7399;
  assign n7559 = n7403 ^ n7402;
  assign n7560 = n7405 & ~n7559;
  assign n7561 = n7560 ^ n7404;
  assign n7565 = n7564 ^ n7561;
  assign n7556 = n7427 ^ n7426;
  assign n7557 = n7429 & ~n7556;
  assign n7558 = n7557 ^ n7428;
  assign n7566 = n7565 ^ n7558;
  assign n7574 = n7573 ^ n7566;
  assign n7553 = n7480 ^ n7474;
  assign n7554 = ~n7481 & n7553;
  assign n7555 = n7554 ^ n7474;
  assign n7575 = n7574 ^ n7555;
  assign n7550 = n7432 ^ n7412;
  assign n7551 = n7433 & n7550;
  assign n7552 = n7551 ^ n7415;
  assign n7576 = n7575 ^ n7552;
  assign n7547 = n7396 ^ n7361;
  assign n7548 = ~n7435 & ~n7547;
  assign n7549 = n7548 ^ n7434;
  assign n7577 = n7576 ^ n7549;
  assign n7544 = n7482 ^ n7444;
  assign n7545 = ~n7483 & ~n7544;
  assign n7546 = n7545 ^ n7444;
  assign n7578 = n7577 ^ n7546;
  assign n7700 = n7699 ^ n7578;
  assign n7541 = n7436 ^ n7355;
  assign n7542 = n7437 & n7541;
  assign n7543 = n7542 ^ n7358;
  assign n7701 = n7700 ^ n7543;
  assign n7538 = n7516 ^ n7438;
  assign n7539 = ~n7517 & n7538;
  assign n7540 = n7539 ^ n7441;
  assign n7702 = n7701 ^ n7540;
  assign n7709 = n7708 ^ n7702;
  assign n7865 = n7601 ^ n7598;
  assign n7866 = n7605 & ~n7865;
  assign n7867 = n7866 ^ n7604;
  assign n7862 = n7615 ^ n7612;
  assign n7863 = ~n7616 & n7862;
  assign n7864 = n7863 ^ n7612;
  assign n7868 = n7867 ^ n7864;
  assign n7859 = n7688 ^ n7685;
  assign n7860 = n7692 & ~n7859;
  assign n7861 = n7860 ^ n7691;
  assign n7869 = n7868 ^ n7861;
  assign n7856 = n7617 ^ n7606;
  assign n7857 = n7618 & ~n7856;
  assign n7858 = n7857 ^ n7609;
  assign n7870 = n7869 ^ n7858;
  assign n7853 = n7693 ^ n7677;
  assign n7854 = n7694 & ~n7853;
  assign n7855 = n7854 ^ n7680;
  assign n7871 = n7870 ^ n7855;
  assign n7850 = n7595 ^ n7584;
  assign n7851 = ~n7620 & n7850;
  assign n7852 = n7851 ^ n7619;
  assign n7872 = n7871 ^ n7852;
  assign n7847 = n7695 ^ n7624;
  assign n7848 = ~n7696 & n7847;
  assign n7849 = n7848 ^ n7624;
  assign n7873 = n7872 ^ n7849;
  assign n7844 = n7697 ^ n7581;
  assign n7845 = n7698 & n7844;
  assign n7846 = n7845 ^ n7581;
  assign n7874 = n7873 ^ n7846;
  assign n7834 = x12 & x59;
  assign n7833 = x13 & x58;
  assign n7835 = n7834 ^ n7833;
  assign n7830 = n7634 ^ n7633;
  assign n7831 = n7636 & ~n7830;
  assign n7832 = n7831 ^ n7635;
  assign n7836 = n7835 ^ n7832;
  assign n7826 = x16 & x55;
  assign n7825 = x15 & x56;
  assign n7827 = n7826 ^ n7825;
  assign n7824 = x14 & x57;
  assign n7828 = n7827 ^ n7824;
  assign n7821 = x26 & x45;
  assign n7820 = x25 & x46;
  assign n7822 = n7821 ^ n7820;
  assign n7819 = x24 & x47;
  assign n7823 = n7822 ^ n7819;
  assign n7829 = n7828 ^ n7823;
  assign n7837 = n7836 ^ n7829;
  assign n7816 = n7593 ^ n7587;
  assign n7817 = ~n7594 & ~n7816;
  assign n7818 = n7817 ^ n7587;
  assign n7838 = n7837 ^ n7818;
  assign n7811 = x32 & x39;
  assign n7810 = x31 & x40;
  assign n7812 = n7811 ^ n7810;
  assign n7809 = x30 & x41;
  assign n7813 = n7812 ^ n7809;
  assign n7806 = x29 & x42;
  assign n7805 = x28 & x43;
  assign n7807 = n7806 ^ n7805;
  assign n7804 = x27 & x44;
  assign n7808 = n7807 ^ n7804;
  assign n7814 = n7813 ^ n7808;
  assign n7801 = x23 & x48;
  assign n7800 = x18 & x53;
  assign n7802 = n7801 ^ n7800;
  assign n7799 = x17 & x54;
  assign n7803 = n7802 ^ n7799;
  assign n7815 = n7814 ^ n7803;
  assign n7839 = n7838 ^ n7815;
  assign n7792 = x11 & x60;
  assign n7791 = x10 & x61;
  assign n7793 = n7792 ^ n7791;
  assign n7790 = x8 & x63;
  assign n7794 = n7793 ^ n7790;
  assign n7787 = n7667 ^ n7666;
  assign n7788 = n7669 & ~n7787;
  assign n7789 = n7788 ^ n7668;
  assign n7795 = n7794 ^ n7789;
  assign n7784 = n7682 ^ n7681;
  assign n7785 = n7684 & ~n7784;
  assign n7786 = n7785 ^ n7683;
  assign n7796 = n7795 ^ n7786;
  assign n7779 = x21 & x50;
  assign n7778 = x20 & x51;
  assign n7780 = n7779 ^ n7778;
  assign n7777 = x19 & x52;
  assign n7781 = n7780 ^ n7777;
  assign n7774 = x35 & x36;
  assign n7773 = x34 & x37;
  assign n7775 = n7774 ^ n7773;
  assign n7772 = x33 & x38;
  assign n7776 = n7775 ^ n7772;
  assign n7782 = n7781 ^ n7776;
  assign n7769 = x9 & x62;
  assign n7768 = x22 & x49;
  assign n7770 = n7769 ^ n7768;
  assign n7771 = n7770 ^ x36;
  assign n7783 = n7782 ^ n7771;
  assign n7797 = n7796 ^ n7783;
  assign n7765 = n7569 ^ n7566;
  assign n7766 = n7573 & ~n7765;
  assign n7767 = n7766 ^ n7572;
  assign n7798 = n7797 ^ n7767;
  assign n7840 = n7839 ^ n7798;
  assign n7762 = n7555 ^ n7552;
  assign n7763 = ~n7575 & n7762;
  assign n7764 = n7763 ^ n7552;
  assign n7841 = n7840 ^ n7764;
  assign n7753 = n7662 ^ n7661;
  assign n7754 = n7664 & ~n7753;
  assign n7755 = n7754 ^ n7663;
  assign n7750 = n7672 ^ n7671;
  assign n7751 = n7674 & ~n7750;
  assign n7752 = n7751 ^ n7673;
  assign n7756 = n7755 ^ n7752;
  assign n7747 = n7639 ^ n7638;
  assign n7748 = n7641 & ~n7747;
  assign n7749 = n7748 ^ n7640;
  assign n7757 = n7756 ^ n7749;
  assign n7744 = n7656 ^ n7647;
  assign n7745 = ~n7657 & n7744;
  assign n7746 = n7745 ^ n7647;
  assign n7758 = n7757 ^ n7746;
  assign n7739 = n7629 ^ n7628;
  assign n7740 = n7631 & ~n7739;
  assign n7741 = n7740 ^ n7630;
  assign n7736 = n7649 ^ n7648;
  assign n7737 = n7651 & ~n7736;
  assign n7738 = n7737 ^ n7650;
  assign n7742 = n7741 ^ n7738;
  assign n7733 = n7654 ^ n7653;
  assign n7734 = n7655 & ~n7733;
  assign n7735 = n7734 ^ n3924;
  assign n7743 = n7742 ^ n7735;
  assign n7759 = n7758 ^ n7743;
  assign n7728 = n7561 ^ n7558;
  assign n7729 = n7565 & ~n7728;
  assign n7730 = n7729 ^ n7564;
  assign n7725 = n7637 ^ n7632;
  assign n7726 = n7643 & ~n7725;
  assign n7727 = n7726 ^ n7642;
  assign n7731 = n7730 ^ n7727;
  assign n7722 = n7670 ^ n7665;
  assign n7723 = n7676 & ~n7722;
  assign n7724 = n7723 ^ n7675;
  assign n7732 = n7731 ^ n7724;
  assign n7760 = n7759 ^ n7732;
  assign n7719 = n7658 ^ n7627;
  assign n7720 = ~n7659 & n7719;
  assign n7721 = n7720 ^ n7627;
  assign n7761 = n7760 ^ n7721;
  assign n7842 = n7841 ^ n7761;
  assign n7716 = n7576 ^ n7546;
  assign n7717 = ~n7577 & n7716;
  assign n7718 = n7717 ^ n7549;
  assign n7843 = n7842 ^ n7718;
  assign n7875 = n7874 ^ n7843;
  assign n7713 = n7699 ^ n7543;
  assign n7714 = n7700 & n7713;
  assign n7715 = n7714 ^ n7543;
  assign n7876 = n7875 ^ n7715;
  assign n7710 = n7708 ^ n7540;
  assign n7711 = ~n7702 & n7710;
  assign n7712 = n7711 ^ n7708;
  assign n7877 = n7876 ^ n7712;
  assign n8036 = x20 & x52;
  assign n8035 = x18 & x54;
  assign n8037 = n8036 ^ n8035;
  assign n8034 = x17 & x55;
  assign n8038 = n8037 ^ n8034;
  assign n8031 = x35 & x37;
  assign n8030 = x22 & x50;
  assign n8032 = n8031 ^ n8030;
  assign n8029 = x21 & x51;
  assign n8033 = n8032 ^ n8029;
  assign n8039 = n8038 ^ n8033;
  assign n8026 = x32 & x40;
  assign n8025 = x23 & x49;
  assign n8027 = n8026 ^ n8025;
  assign n8024 = x16 & x56;
  assign n8028 = n8027 ^ n8024;
  assign n8040 = n8039 ^ n8028;
  assign n8021 = n7727 ^ n7724;
  assign n8022 = n7731 & ~n8021;
  assign n8023 = n8022 ^ n7730;
  assign n8041 = n8040 ^ n8023;
  assign n8017 = n7832 & n7835;
  assign n7982 = x13 & x59;
  assign n8018 = n7661 & n7982;
  assign n8019 = ~n8017 & ~n8018;
  assign n8013 = x11 & x61;
  assign n8012 = x10 & x62;
  assign n8014 = n8013 ^ n8012;
  assign n8011 = x9 & x63;
  assign n8015 = n8014 ^ n8011;
  assign n8008 = x24 & x48;
  assign n8009 = n8008 ^ n4012;
  assign n8007 = x12 & x60;
  assign n8010 = n8009 ^ n8007;
  assign n8016 = n8015 ^ n8010;
  assign n8020 = n8019 ^ n8016;
  assign n8042 = n8041 ^ n8020;
  assign n8000 = n7791 ^ n7790;
  assign n8001 = n7793 & ~n8000;
  assign n8002 = n8001 ^ n7792;
  assign n7997 = n7820 ^ n7819;
  assign n7998 = n7822 & ~n7997;
  assign n7999 = n7998 ^ n7821;
  assign n8003 = n8002 ^ n7999;
  assign n7994 = n7825 ^ n7824;
  assign n7995 = n7827 & ~n7994;
  assign n7996 = n7995 ^ n7826;
  assign n8004 = n8003 ^ n7996;
  assign n7991 = n7864 ^ n7861;
  assign n7992 = n7868 & ~n7991;
  assign n7993 = n7992 ^ n7867;
  assign n8005 = n8004 ^ n7993;
  assign n7986 = x34 & x38;
  assign n7985 = x33 & x39;
  assign n7987 = n7986 ^ n7985;
  assign n7984 = x19 & x53;
  assign n7988 = n7987 ^ n7984;
  assign n7980 = x15 & x57;
  assign n7979 = x14 & x58;
  assign n7981 = n7980 ^ n7979;
  assign n7983 = n7982 ^ n7981;
  assign n7989 = n7988 ^ n7983;
  assign n7976 = x28 & x44;
  assign n7975 = x27 & x45;
  assign n7977 = n7976 ^ n7975;
  assign n7974 = x26 & x46;
  assign n7978 = n7977 ^ n7974;
  assign n7990 = n7989 ^ n7978;
  assign n8006 = n8005 ^ n7990;
  assign n8043 = n8042 ^ n8006;
  assign n7971 = n7858 ^ n7855;
  assign n7972 = ~n7870 & n7971;
  assign n7973 = n7972 ^ n7855;
  assign n8044 = n8043 ^ n7973;
  assign n7962 = n7778 ^ n7777;
  assign n7963 = n7780 & ~n7962;
  assign n7964 = n7963 ^ n7779;
  assign n7959 = n7773 ^ n7772;
  assign n7960 = n7775 & ~n7959;
  assign n7961 = n7960 ^ n7774;
  assign n7965 = n7964 ^ n7961;
  assign n7955 = x49 & n5425;
  assign n7956 = ~n7769 & ~n7955;
  assign n7957 = ~x36 & ~n7768;
  assign n7958 = ~n7956 & ~n7957;
  assign n7966 = n7965 ^ n7958;
  assign n7952 = n7836 ^ n7828;
  assign n7953 = ~n7829 & n7952;
  assign n7954 = n7953 ^ n7836;
  assign n7967 = n7966 ^ n7954;
  assign n7947 = n7805 ^ n7804;
  assign n7948 = n7807 & ~n7947;
  assign n7949 = n7948 ^ n7806;
  assign n7944 = n7800 ^ n7799;
  assign n7945 = n7802 & ~n7944;
  assign n7946 = n7945 ^ n7801;
  assign n7950 = n7949 ^ n7946;
  assign n7941 = n7810 ^ n7809;
  assign n7942 = n7812 & ~n7941;
  assign n7943 = n7942 ^ n7811;
  assign n7951 = n7950 ^ n7943;
  assign n7968 = n7967 ^ n7951;
  assign n7936 = n7776 ^ n7771;
  assign n7937 = n7782 & ~n7936;
  assign n7938 = n7937 ^ n7781;
  assign n7933 = n7808 ^ n7803;
  assign n7934 = n7814 & ~n7933;
  assign n7935 = n7934 ^ n7813;
  assign n7939 = n7938 ^ n7935;
  assign n7930 = n7752 ^ n7749;
  assign n7931 = n7756 & ~n7930;
  assign n7932 = n7931 ^ n7755;
  assign n7940 = n7939 ^ n7932;
  assign n7969 = n7968 ^ n7940;
  assign n7927 = n7837 ^ n7815;
  assign n7928 = ~n7838 & ~n7927;
  assign n7929 = n7928 ^ n7818;
  assign n7970 = n7969 ^ n7929;
  assign n8045 = n8044 ^ n7970;
  assign n7924 = n7852 ^ n7849;
  assign n7925 = ~n7872 & n7924;
  assign n7926 = n7925 ^ n7849;
  assign n8046 = n8045 ^ n7926;
  assign n7915 = x31 & x41;
  assign n7914 = x30 & x42;
  assign n7916 = n7915 ^ n7914;
  assign n7913 = x29 & x43;
  assign n7917 = n7916 ^ n7913;
  assign n7910 = n7738 ^ n7735;
  assign n7911 = n7742 & ~n7910;
  assign n7912 = n7911 ^ n7741;
  assign n7918 = n7917 ^ n7912;
  assign n7907 = n7794 ^ n7786;
  assign n7908 = n7795 & ~n7907;
  assign n7909 = n7908 ^ n7789;
  assign n7919 = n7918 ^ n7909;
  assign n7904 = n7757 ^ n7743;
  assign n7905 = n7758 & ~n7904;
  assign n7906 = n7905 ^ n7746;
  assign n7920 = n7919 ^ n7906;
  assign n7901 = n7796 ^ n7767;
  assign n7902 = ~n7797 & n7901;
  assign n7903 = n7902 ^ n7767;
  assign n7921 = n7920 ^ n7903;
  assign n7898 = n7732 ^ n7721;
  assign n7899 = n7760 & ~n7898;
  assign n7900 = n7899 ^ n7759;
  assign n7922 = n7921 ^ n7900;
  assign n7895 = n7839 ^ n7764;
  assign n7896 = n7840 & ~n7895;
  assign n7897 = n7896 ^ n7764;
  assign n7923 = n7922 ^ n7897;
  assign n8047 = n8046 ^ n7923;
  assign n7892 = n7841 ^ n7718;
  assign n7893 = n7842 & n7892;
  assign n7894 = n7893 ^ n7718;
  assign n8048 = n8047 ^ n7894;
  assign n7878 = n7715 & ~n7846;
  assign n7879 = ~n7843 & ~n7873;
  assign n7880 = n7878 & n7879;
  assign n7881 = ~n7715 & n7846;
  assign n7882 = n7843 & n7873;
  assign n7883 = n7881 & n7882;
  assign n7884 = ~n7880 & ~n7883;
  assign n7885 = ~n7878 & ~n7879;
  assign n7886 = n7885 ^ n7712;
  assign n7887 = ~n7881 & ~n7882;
  assign n7888 = n7887 ^ n7885;
  assign n7889 = ~n7886 & n7888;
  assign n7890 = n7884 & n7889;
  assign n7891 = n7890 ^ n7884;
  assign n8049 = n8048 ^ n7891;
  assign n8206 = ~n7878 & ~n8048;
  assign n8207 = ~n7882 & ~n8206;
  assign n8208 = ~n7879 & ~n8048;
  assign n8209 = ~n7881 & ~n8208;
  assign n8210 = ~n8207 & ~n8209;
  assign n8211 = ~n7712 & ~n8210;
  assign n8212 = n7885 & ~n7887;
  assign n8213 = ~n7880 & ~n8048;
  assign n8214 = ~n8212 & ~n8213;
  assign n8215 = ~n8211 & ~n8214;
  assign n8194 = x33 & x40;
  assign n8193 = x32 & x41;
  assign n8195 = n8194 ^ n8193;
  assign n8192 = x31 & x42;
  assign n8196 = n8195 ^ n8192;
  assign n8189 = n7999 ^ n7996;
  assign n8190 = n8003 & ~n8189;
  assign n8191 = n8190 ^ n8002;
  assign n8197 = n8196 ^ n8191;
  assign n8186 = n7946 ^ n7943;
  assign n8187 = n7950 & ~n8186;
  assign n8188 = n8187 ^ n7949;
  assign n8198 = n8197 ^ n8188;
  assign n8183 = n8004 ^ n7990;
  assign n8184 = n8005 & ~n8183;
  assign n8185 = n8184 ^ n7993;
  assign n8199 = n8198 ^ n8185;
  assign n8180 = n7966 ^ n7951;
  assign n8181 = n7967 & ~n8180;
  assign n8182 = n8181 ^ n7954;
  assign n8200 = n8199 ^ n8182;
  assign n8177 = n7968 ^ n7929;
  assign n8178 = ~n7969 & ~n8177;
  assign n8179 = n8178 ^ n7929;
  assign n8201 = n8200 ^ n8179;
  assign n8174 = n8042 ^ n7973;
  assign n8175 = n8043 & ~n8174;
  assign n8176 = n8175 ^ n7973;
  assign n8202 = n8201 ^ n8176;
  assign n8171 = n8044 ^ n7926;
  assign n8172 = ~n8045 & ~n8171;
  assign n8173 = n8172 ^ n7926;
  assign n8203 = n8202 ^ n8173;
  assign n8160 = x30 & x43;
  assign n8159 = x29 & x44;
  assign n8161 = n8160 ^ n8159;
  assign n8158 = x28 & x45;
  assign n8162 = n8161 ^ n8158;
  assign n8155 = x12 & x61;
  assign n8156 = n8155 ^ n4015;
  assign n8154 = x10 & x63;
  assign n8157 = n8156 ^ n8154;
  assign n8163 = n8162 ^ n8157;
  assign n8151 = x36 & x37;
  assign n8150 = x35 & x38;
  assign n8152 = n8151 ^ n8150;
  assign n8149 = x34 & x39;
  assign n8153 = n8152 ^ n8149;
  assign n8164 = n8163 ^ n8153;
  assign n8146 = n7917 ^ n7909;
  assign n8147 = n7918 & ~n8146;
  assign n8148 = n8147 ^ n7912;
  assign n8165 = n8164 ^ n8148;
  assign n8141 = n7914 ^ n7913;
  assign n8142 = n7916 & ~n8141;
  assign n8143 = n8142 ^ n7915;
  assign n8138 = n7982 ^ n7980;
  assign n8139 = ~n7981 & n8138;
  assign n8140 = n8139 ^ n7982;
  assign n8144 = n8143 ^ n8140;
  assign n8135 = n7975 ^ n7974;
  assign n8136 = n7977 & ~n8135;
  assign n8137 = n8136 ^ n7976;
  assign n8145 = n8144 ^ n8137;
  assign n8166 = n8165 ^ n8145;
  assign n8128 = x22 & x51;
  assign n8127 = x21 & x52;
  assign n8129 = n8128 ^ n8127;
  assign n8126 = x20 & x53;
  assign n8130 = n8129 ^ n8126;
  assign n8123 = x19 & x54;
  assign n8124 = n8123 ^ n4255;
  assign n8122 = x18 & x55;
  assign n8125 = n8124 ^ n8122;
  assign n8131 = n8130 ^ n8125;
  assign n8119 = x11 & x62;
  assign n8118 = x23 & x50;
  assign n8120 = n8119 ^ n8118;
  assign n8121 = n8120 ^ x37;
  assign n8132 = n8131 ^ n8121;
  assign n8115 = n7938 ^ n7932;
  assign n8116 = ~n7939 & n8115;
  assign n8117 = n8116 ^ n7932;
  assign n8133 = n8132 ^ n8117;
  assign n8110 = x27 & x46;
  assign n8109 = x26 & x47;
  assign n8111 = n8110 ^ n8109;
  assign n8108 = x17 & x56;
  assign n8112 = n8111 ^ n8108;
  assign n8105 = n8025 ^ n8024;
  assign n8106 = n8027 & ~n8105;
  assign n8107 = n8106 ^ n8026;
  assign n8113 = n8112 ^ n8107;
  assign n8102 = x16 & x57;
  assign n8101 = x15 & x58;
  assign n8103 = n8102 ^ n8101;
  assign n8100 = x14 & x59;
  assign n8104 = n8103 ^ n8100;
  assign n8114 = n8113 ^ n8104;
  assign n8134 = n8133 ^ n8114;
  assign n8167 = n8166 ^ n8134;
  assign n8097 = n7919 ^ n7903;
  assign n8098 = n7920 & ~n8097;
  assign n8099 = n8098 ^ n7906;
  assign n8168 = n8167 ^ n8099;
  assign n8090 = x13 & x60;
  assign n8087 = n8030 ^ n8029;
  assign n8088 = n8032 & ~n8087;
  assign n8089 = n8088 ^ n8031;
  assign n8091 = n8090 ^ n8089;
  assign n8084 = n7985 ^ n7984;
  assign n8085 = n7987 & ~n8084;
  assign n8086 = n8085 ^ n7986;
  assign n8092 = n8091 ^ n8086;
  assign n8081 = n8033 ^ n8028;
  assign n8082 = n8039 & ~n8081;
  assign n8083 = n8082 ^ n8038;
  assign n8093 = n8092 ^ n8083;
  assign n8076 = n8035 ^ n8034;
  assign n8077 = n8037 & ~n8076;
  assign n8078 = n8077 ^ n8036;
  assign n8073 = n8012 ^ n8011;
  assign n8074 = n8014 & ~n8073;
  assign n8075 = n8074 ^ n8013;
  assign n8079 = n8078 ^ n8075;
  assign n8070 = n8008 ^ n8007;
  assign n8071 = n8009 & ~n8070;
  assign n8072 = n8071 ^ n4012;
  assign n8080 = n8079 ^ n8072;
  assign n8094 = n8093 ^ n8080;
  assign n8067 = n8040 ^ n8020;
  assign n8068 = n8041 & n8067;
  assign n8069 = n8068 ^ n8023;
  assign n8095 = n8094 ^ n8069;
  assign n8062 = n8019 ^ n8015;
  assign n8063 = ~n8016 & ~n8062;
  assign n8064 = n8063 ^ n8019;
  assign n8059 = n7961 ^ n7958;
  assign n8060 = n7965 & ~n8059;
  assign n8061 = n8060 ^ n7964;
  assign n8065 = n8064 ^ n8061;
  assign n8056 = n7983 ^ n7978;
  assign n8057 = n7989 & ~n8056;
  assign n8058 = n8057 ^ n7988;
  assign n8066 = n8065 ^ n8058;
  assign n8096 = n8095 ^ n8066;
  assign n8169 = n8168 ^ n8096;
  assign n8053 = n7900 ^ n7897;
  assign n8054 = ~n7922 & n8053;
  assign n8055 = n8054 ^ n7897;
  assign n8170 = n8169 ^ n8055;
  assign n8204 = n8203 ^ n8170;
  assign n8050 = n8046 ^ n7894;
  assign n8051 = ~n8047 & ~n8050;
  assign n8052 = n8051 ^ n7894;
  assign n8205 = n8204 ^ n8052;
  assign n8216 = n8215 ^ n8205;
  assign n8369 = n8052 & n8170;
  assign n8370 = n8215 & ~n8369;
  assign n8371 = ~n8052 & ~n8170;
  assign n8372 = n8173 & ~n8202;
  assign n8373 = ~n8371 & ~n8372;
  assign n8374 = ~n8173 & n8202;
  assign n8375 = ~n8373 & ~n8374;
  assign n8376 = n8370 & n8375;
  assign n8377 = ~n8369 & ~n8374;
  assign n8378 = n8373 & ~n8377;
  assign n8379 = ~n8215 & n8378;
  assign n8380 = n8173 ^ n8052;
  assign n8381 = n8202 ^ n8170;
  assign n8382 = n8203 & ~n8381;
  assign n8383 = n8380 & n8382;
  assign n8384 = ~n8379 & ~n8383;
  assign n8385 = ~n8376 & n8384;
  assign n8360 = n8164 ^ n8145;
  assign n8361 = n8165 & ~n8360;
  assign n8362 = n8361 ^ n8148;
  assign n8357 = n8132 ^ n8114;
  assign n8358 = n8133 & ~n8357;
  assign n8359 = n8358 ^ n8117;
  assign n8363 = n8362 ^ n8359;
  assign n8350 = x16 & x58;
  assign n8349 = x15 & x59;
  assign n8351 = n8350 ^ n8349;
  assign n8348 = x14 & x60;
  assign n8352 = n8351 ^ n8348;
  assign n8345 = n8150 ^ n8149;
  assign n8346 = n8152 & ~n8345;
  assign n8347 = n8346 ^ n8151;
  assign n8353 = n8352 ^ n8347;
  assign n8342 = n8193 ^ n8192;
  assign n8343 = n8195 & ~n8342;
  assign n8344 = n8343 ^ n8194;
  assign n8354 = n8353 ^ n8344;
  assign n8339 = n8196 ^ n8188;
  assign n8340 = n8197 & ~n8339;
  assign n8341 = n8340 ^ n8191;
  assign n8355 = n8354 ^ n8341;
  assign n8336 = n8125 ^ n8121;
  assign n8337 = n8131 & ~n8336;
  assign n8338 = n8337 ^ n8130;
  assign n8356 = n8355 ^ n8338;
  assign n8364 = n8363 ^ n8356;
  assign n8333 = n8179 ^ n8176;
  assign n8334 = n8201 & ~n8333;
  assign n8335 = n8334 ^ n8176;
  assign n8365 = n8364 ^ n8335;
  assign n8323 = x50 & n5772;
  assign n8324 = ~n8119 & ~n8323;
  assign n8325 = ~x37 & ~n8118;
  assign n8326 = ~n8324 & ~n8325;
  assign n8321 = x12 & x62;
  assign n8320 = x13 & x61;
  assign n8322 = n8321 ^ n8320;
  assign n8327 = n8326 ^ n8322;
  assign n8317 = x30 & x44;
  assign n8316 = x29 & x45;
  assign n8318 = n8317 ^ n8316;
  assign n8315 = x17 & x57;
  assign n8319 = n8318 ^ n8315;
  assign n8328 = n8327 ^ n8319;
  assign n8312 = n8140 ^ n8137;
  assign n8313 = n8144 & ~n8312;
  assign n8314 = n8313 ^ n8143;
  assign n8329 = n8328 ^ n8314;
  assign n8306 = x33 & x41;
  assign n8305 = x25 & x49;
  assign n8307 = n8306 ^ n8305;
  assign n8304 = x18 & x56;
  assign n8308 = n8307 ^ n8304;
  assign n8301 = x32 & x42;
  assign n8300 = x31 & x43;
  assign n8302 = n8301 ^ n8300;
  assign n8299 = x11 & x63;
  assign n8303 = n8302 ^ n8299;
  assign n8309 = n8308 ^ n8303;
  assign n8296 = x28 & x46;
  assign n8295 = x27 & x47;
  assign n8297 = n8296 ^ n8295;
  assign n8294 = x26 & x48;
  assign n8298 = n8297 ^ n8294;
  assign n8310 = n8309 ^ n8298;
  assign n8289 = x22 & x52;
  assign n8288 = x21 & x53;
  assign n8290 = n8289 ^ n8288;
  assign n8287 = x19 & x55;
  assign n8291 = n8290 ^ n8287;
  assign n8284 = x35 & x39;
  assign n8283 = x34 & x40;
  assign n8285 = n8284 ^ n8283;
  assign n8282 = x20 & x54;
  assign n8286 = n8285 ^ n8282;
  assign n8292 = n8291 ^ n8286;
  assign n8279 = x36 & x38;
  assign n8278 = x24 & x50;
  assign n8280 = n8279 ^ n8278;
  assign n8277 = x23 & x51;
  assign n8281 = n8280 ^ n8277;
  assign n8293 = n8292 ^ n8281;
  assign n8311 = n8310 ^ n8293;
  assign n8330 = n8329 ^ n8311;
  assign n8270 = n8159 ^ n8158;
  assign n8271 = n8161 & ~n8270;
  assign n8272 = n8271 ^ n8160;
  assign n8267 = n8109 ^ n8108;
  assign n8268 = n8111 & ~n8267;
  assign n8269 = n8268 ^ n8110;
  assign n8273 = n8272 ^ n8269;
  assign n8264 = n8101 ^ n8100;
  assign n8265 = n8103 & ~n8264;
  assign n8266 = n8265 ^ n8102;
  assign n8274 = n8273 ^ n8266;
  assign n8261 = n8157 ^ n8153;
  assign n8262 = n8163 & ~n8261;
  assign n8263 = n8262 ^ n8162;
  assign n8275 = n8274 ^ n8263;
  assign n8256 = n8127 ^ n8126;
  assign n8257 = n8129 & ~n8256;
  assign n8258 = n8257 ^ n8128;
  assign n8253 = n8123 ^ n8122;
  assign n8254 = n8124 & ~n8253;
  assign n8255 = n8254 ^ n4255;
  assign n8259 = n8258 ^ n8255;
  assign n8250 = n8155 ^ n8154;
  assign n8251 = n8156 & ~n8250;
  assign n8252 = n8251 ^ n4015;
  assign n8260 = n8259 ^ n8252;
  assign n8276 = n8275 ^ n8260;
  assign n8331 = n8330 ^ n8276;
  assign n8247 = n8198 ^ n8182;
  assign n8248 = n8199 & ~n8247;
  assign n8249 = n8248 ^ n8185;
  assign n8332 = n8331 ^ n8249;
  assign n8366 = n8365 ^ n8332;
  assign n8238 = n8112 ^ n8104;
  assign n8239 = n8113 & ~n8238;
  assign n8240 = n8239 ^ n8107;
  assign n8235 = n8090 ^ n8086;
  assign n8236 = n8091 & ~n8235;
  assign n8237 = n8236 ^ n8089;
  assign n8241 = n8240 ^ n8237;
  assign n8232 = n8075 ^ n8072;
  assign n8233 = n8079 & ~n8232;
  assign n8234 = n8233 ^ n8078;
  assign n8242 = n8241 ^ n8234;
  assign n8229 = n8061 ^ n8058;
  assign n8230 = ~n8065 & ~n8229;
  assign n8231 = n8230 ^ n8064;
  assign n8243 = n8242 ^ n8231;
  assign n8226 = n8083 ^ n8080;
  assign n8227 = n8093 & ~n8226;
  assign n8228 = n8227 ^ n8092;
  assign n8244 = n8243 ^ n8228;
  assign n8223 = n8094 ^ n8066;
  assign n8224 = n8095 & n8223;
  assign n8225 = n8224 ^ n8069;
  assign n8245 = n8244 ^ n8225;
  assign n8220 = n8166 ^ n8099;
  assign n8221 = ~n8167 & n8220;
  assign n8222 = n8221 ^ n8099;
  assign n8246 = n8245 ^ n8222;
  assign n8367 = n8366 ^ n8246;
  assign n8217 = n8168 ^ n8055;
  assign n8218 = n8169 & n8217;
  assign n8219 = n8218 ^ n8055;
  assign n8368 = n8367 ^ n8219;
  assign n8386 = n8385 ^ n8368;
  assign n8539 = ~n8368 & ~n8374;
  assign n8540 = ~n8371 & ~n8539;
  assign n8541 = ~n8370 & n8540;
  assign n8542 = ~n8368 & ~n8369;
  assign n8543 = ~n8372 & ~n8542;
  assign n8544 = ~n8215 & n8543;
  assign n8545 = n8368 & ~n8375;
  assign n8546 = ~n8544 & ~n8545;
  assign n8547 = ~n8541 & n8546;
  assign n8529 = n8354 ^ n8338;
  assign n8530 = n8355 & ~n8529;
  assign n8531 = n8530 ^ n8341;
  assign n8526 = n8263 ^ n8260;
  assign n8527 = n8275 & ~n8526;
  assign n8528 = n8527 ^ n8274;
  assign n8532 = n8531 ^ n8528;
  assign n8521 = x33 & x42;
  assign n8520 = x32 & x43;
  assign n8522 = n8521 ^ n8520;
  assign n8519 = x31 & x44;
  assign n8523 = n8522 ^ n8519;
  assign n8516 = x24 & x51;
  assign n8515 = x22 & x53;
  assign n8517 = n8516 ^ n8515;
  assign n8514 = x21 & x54;
  assign n8518 = n8517 ^ n8514;
  assign n8524 = n8523 ^ n8518;
  assign n8511 = x34 & x41;
  assign n8510 = x25 & x50;
  assign n8512 = n8511 ^ n8510;
  assign n8509 = x20 & x55;
  assign n8513 = n8512 ^ n8509;
  assign n8525 = n8524 ^ n8513;
  assign n8533 = n8532 ^ n8525;
  assign n8506 = n8330 ^ n8249;
  assign n8507 = ~n8331 & n8506;
  assign n8508 = n8507 ^ n8249;
  assign n8534 = n8533 ^ n8508;
  assign n8503 = n8359 ^ n8356;
  assign n8504 = n8363 & ~n8503;
  assign n8505 = n8504 ^ n8362;
  assign n8535 = n8534 ^ n8505;
  assign n8492 = n8316 ^ n8315;
  assign n8493 = n8318 & ~n8492;
  assign n8494 = n8493 ^ n8317;
  assign n8489 = n8295 ^ n8294;
  assign n8490 = n8297 & ~n8489;
  assign n8491 = n8490 ^ n8296;
  assign n8495 = n8494 ^ n8491;
  assign n8486 = n8349 ^ n8348;
  assign n8487 = n8351 & ~n8486;
  assign n8488 = n8487 ^ n8350;
  assign n8496 = n8495 ^ n8488;
  assign n8483 = n8303 ^ n8298;
  assign n8484 = n8309 & ~n8483;
  assign n8485 = n8484 ^ n8308;
  assign n8497 = n8496 ^ n8485;
  assign n8480 = n8286 ^ n8281;
  assign n8481 = n8292 & ~n8480;
  assign n8482 = n8481 ^ n8291;
  assign n8498 = n8497 ^ n8482;
  assign n8477 = n8242 ^ n8228;
  assign n8478 = ~n8243 & ~n8477;
  assign n8479 = n8478 ^ n8231;
  assign n8499 = n8498 ^ n8479;
  assign n8470 = x16 & x59;
  assign n8469 = x15 & x60;
  assign n8471 = n8470 ^ n8469;
  assign n8468 = x14 & x61;
  assign n8472 = n8471 ^ n8468;
  assign n8465 = x26 & x49;
  assign n8464 = x18 & x57;
  assign n8466 = n8465 ^ n8464;
  assign n8463 = x17 & x58;
  assign n8467 = n8466 ^ n8463;
  assign n8473 = n8472 ^ n8467;
  assign n8460 = x29 & x46;
  assign n8459 = x28 & x47;
  assign n8461 = n8460 ^ n8459;
  assign n8458 = x27 & x48;
  assign n8462 = n8461 ^ n8458;
  assign n8474 = n8473 ^ n8462;
  assign n8453 = x36 & x39;
  assign n8452 = x35 & x40;
  assign n8454 = n8453 ^ n8452;
  assign n8451 = x23 & x52;
  assign n8455 = n8454 ^ n8451;
  assign n8448 = x30 & x45;
  assign n8447 = x19 & x56;
  assign n8449 = n8448 ^ n8447;
  assign n8446 = x12 & x63;
  assign n8450 = n8449 ^ n8446;
  assign n8456 = n8455 ^ n8450;
  assign n8444 = x13 & x62;
  assign n8443 = ~x37 & x38;
  assign n8445 = n8444 ^ n8443;
  assign n8457 = n8456 ^ n8445;
  assign n8475 = n8474 ^ n8457;
  assign n8440 = n8237 ^ n8234;
  assign n8441 = n8241 & ~n8440;
  assign n8442 = n8441 ^ n8240;
  assign n8476 = n8475 ^ n8442;
  assign n8500 = n8499 ^ n8476;
  assign n8431 = n8322 & n8326;
  assign n8432 = x61 & x62;
  assign n8433 = n1046 & n8432;
  assign n8434 = ~n8431 & ~n8433;
  assign n8427 = n8305 ^ n8304;
  assign n8428 = n8307 & ~n8427;
  assign n8429 = n8428 ^ n8306;
  assign n8424 = n8300 ^ n8299;
  assign n8425 = n8302 & ~n8424;
  assign n8426 = n8425 ^ n8301;
  assign n8430 = n8429 ^ n8426;
  assign n8435 = n8434 ^ n8430;
  assign n8419 = n8278 ^ n8277;
  assign n8420 = n8280 & ~n8419;
  assign n8421 = n8420 ^ n8279;
  assign n8416 = n8288 ^ n8287;
  assign n8417 = n8290 & ~n8416;
  assign n8418 = n8417 ^ n8289;
  assign n8422 = n8421 ^ n8418;
  assign n8413 = n8283 ^ n8282;
  assign n8414 = n8285 & ~n8413;
  assign n8415 = n8414 ^ n8284;
  assign n8423 = n8422 ^ n8415;
  assign n8436 = n8435 ^ n8423;
  assign n8410 = n8327 ^ n8314;
  assign n8411 = ~n8328 & n8410;
  assign n8412 = n8411 ^ n8314;
  assign n8437 = n8436 ^ n8412;
  assign n8405 = n8255 ^ n8252;
  assign n8406 = n8259 & ~n8405;
  assign n8407 = n8406 ^ n8258;
  assign n8402 = n8269 ^ n8266;
  assign n8403 = n8273 & ~n8402;
  assign n8404 = n8403 ^ n8272;
  assign n8408 = n8407 ^ n8404;
  assign n8399 = n8352 ^ n8344;
  assign n8400 = n8353 & ~n8399;
  assign n8401 = n8400 ^ n8347;
  assign n8409 = n8408 ^ n8401;
  assign n8438 = n8437 ^ n8409;
  assign n8396 = n8329 ^ n8310;
  assign n8397 = ~n8311 & n8396;
  assign n8398 = n8397 ^ n8329;
  assign n8439 = n8438 ^ n8398;
  assign n8501 = n8500 ^ n8439;
  assign n8393 = n8244 ^ n8222;
  assign n8394 = ~n8245 & n8393;
  assign n8395 = n8394 ^ n8225;
  assign n8502 = n8501 ^ n8395;
  assign n8536 = n8535 ^ n8502;
  assign n8390 = n8364 ^ n8332;
  assign n8391 = n8365 & ~n8390;
  assign n8392 = n8391 ^ n8335;
  assign n8537 = n8536 ^ n8392;
  assign n8387 = n8246 ^ n8219;
  assign n8388 = ~n8367 & n8387;
  assign n8389 = n8388 ^ n8366;
  assign n8538 = n8537 ^ n8389;
  assign n8548 = n8547 ^ n8538;
  assign n8692 = ~n8389 & ~n8392;
  assign n8693 = ~n8502 & ~n8535;
  assign n8695 = n8389 & n8392;
  assign n8696 = n8502 & n8535;
  assign n8697 = ~n8695 & ~n8696;
  assign n8700 = ~n8693 & ~n8697;
  assign n8701 = ~n8692 & n8700;
  assign n8694 = ~n8692 & ~n8693;
  assign n8698 = n8697 ^ n8694;
  assign n8699 = ~n8547 & n8698;
  assign n8702 = n8701 ^ n8699;
  assign n8703 = n8392 ^ n8389;
  assign n8704 = n8535 ^ n8392;
  assign n8705 = ~n8536 & ~n8704;
  assign n8706 = ~n8703 & n8705;
  assign n8707 = ~n8702 & ~n8706;
  assign n8683 = n8435 ^ n8412;
  assign n8684 = n8436 & ~n8683;
  assign n8685 = n8684 ^ n8412;
  assign n8680 = n8496 ^ n8482;
  assign n8681 = n8497 & ~n8680;
  assign n8682 = n8681 ^ n8485;
  assign n8686 = n8685 ^ n8682;
  assign n8675 = x32 & x44;
  assign n8674 = x31 & x45;
  assign n8676 = n8675 ^ n8674;
  assign n8673 = x13 & x63;
  assign n8677 = n8676 ^ n8673;
  assign n8670 = x33 & x43;
  assign n8669 = x23 & x53;
  assign n8671 = n8670 ^ n8669;
  assign n8668 = x19 & x57;
  assign n8672 = n8671 ^ n8668;
  assign n8678 = n8677 ^ n8672;
  assign n8665 = x22 & x54;
  assign n8664 = x21 & x55;
  assign n8666 = n8665 ^ n8664;
  assign n8663 = x20 & x56;
  assign n8667 = n8666 ^ n8663;
  assign n8679 = n8678 ^ n8667;
  assign n8687 = n8686 ^ n8679;
  assign n8660 = n8498 ^ n8476;
  assign n8661 = ~n8499 & ~n8660;
  assign n8662 = n8661 ^ n8479;
  assign n8688 = n8687 ^ n8662;
  assign n8657 = n8409 ^ n8398;
  assign n8658 = ~n8438 & ~n8657;
  assign n8659 = n8658 ^ n8437;
  assign n8689 = n8688 ^ n8659;
  assign n8654 = n8500 ^ n8395;
  assign n8655 = ~n8501 & ~n8654;
  assign n8656 = n8655 ^ n8395;
  assign n8690 = n8689 ^ n8656;
  assign n8645 = n8450 ^ n8445;
  assign n8646 = n8456 & ~n8645;
  assign n8647 = n8646 ^ n8455;
  assign n8642 = n8467 ^ n8462;
  assign n8643 = n8473 & ~n8642;
  assign n8644 = n8643 ^ n8472;
  assign n8648 = n8647 ^ n8644;
  assign n8637 = n8520 ^ n8519;
  assign n8638 = n8522 & ~n8637;
  assign n8639 = n8638 ^ n8521;
  assign n8634 = n8464 ^ n8463;
  assign n8635 = n8466 & ~n8634;
  assign n8636 = n8635 ^ n8465;
  assign n8640 = n8639 ^ n8636;
  assign n8631 = n8469 ^ n8468;
  assign n8632 = n8471 & ~n8631;
  assign n8633 = n8632 ^ n8470;
  assign n8641 = n8640 ^ n8633;
  assign n8649 = n8648 ^ n8641;
  assign n8628 = n8528 ^ n8525;
  assign n8629 = n8532 & ~n8628;
  assign n8630 = n8629 ^ n8531;
  assign n8650 = n8649 ^ n8630;
  assign n8621 = x36 & x40;
  assign n8620 = x35 & x41;
  assign n8622 = n8621 ^ n8620;
  assign n8619 = x34 & x42;
  assign n8623 = n8622 ^ n8619;
  assign n8616 = x37 & x39;
  assign n8615 = x25 & x51;
  assign n8617 = n8616 ^ n8615;
  assign n8614 = x24 & x52;
  assign n8618 = n8617 ^ n8614;
  assign n8624 = n8623 ^ n8618;
  assign n8611 = x30 & x46;
  assign n8610 = x29 & x47;
  assign n8612 = n8611 ^ n8610;
  assign n8609 = x28 & x48;
  assign n8613 = n8612 ^ n8609;
  assign n8625 = n8624 ^ n8613;
  assign n8606 = n8404 ^ n8401;
  assign n8607 = n8408 & ~n8606;
  assign n8608 = n8607 ^ n8407;
  assign n8626 = n8625 ^ n8608;
  assign n8601 = x27 & x49;
  assign n8602 = n8601 ^ n4353;
  assign n8600 = x18 & x58;
  assign n8603 = n8602 ^ n8600;
  assign n8597 = n8515 ^ n8514;
  assign n8598 = n8517 & ~n8597;
  assign n8599 = n8598 ^ n8516;
  assign n8604 = n8603 ^ n8599;
  assign n8594 = x17 & x59;
  assign n8593 = x16 & x60;
  assign n8595 = n8594 ^ n8593;
  assign n8592 = x15 & x61;
  assign n8596 = n8595 ^ n8592;
  assign n8605 = n8604 ^ n8596;
  assign n8627 = n8626 ^ n8605;
  assign n8651 = n8650 ^ n8627;
  assign n8585 = n8434 ^ n8429;
  assign n8586 = ~n8430 & ~n8585;
  assign n8587 = n8586 ^ n8434;
  assign n8582 = n8491 ^ n8488;
  assign n8583 = n8495 & ~n8582;
  assign n8584 = n8583 ^ n8494;
  assign n8588 = n8587 ^ n8584;
  assign n8579 = n8418 ^ n8415;
  assign n8580 = n8422 & ~n8579;
  assign n8581 = n8580 ^ n8421;
  assign n8589 = n8588 ^ n8581;
  assign n8572 = n8510 ^ n8509;
  assign n8573 = n8512 & ~n8572;
  assign n8574 = n8573 ^ n8511;
  assign n8569 = n8459 ^ n8458;
  assign n8570 = n8461 & ~n8569;
  assign n8571 = n8570 ^ n8460;
  assign n8575 = n8574 ^ n8571;
  assign n8566 = n8447 ^ n8446;
  assign n8567 = n8449 & ~n8566;
  assign n8568 = n8567 ^ n8448;
  assign n8576 = n8575 ^ n8568;
  assign n8562 = ~x37 & ~n8444;
  assign n8563 = x38 & ~n8562;
  assign n8561 = x14 & x62;
  assign n8564 = n8563 ^ n8561;
  assign n8558 = n8452 ^ n8451;
  assign n8559 = n8454 & ~n8558;
  assign n8560 = n8559 ^ n8453;
  assign n8565 = n8564 ^ n8560;
  assign n8577 = n8576 ^ n8565;
  assign n8555 = n8518 ^ n8513;
  assign n8556 = n8524 & ~n8555;
  assign n8557 = n8556 ^ n8523;
  assign n8578 = n8577 ^ n8557;
  assign n8590 = n8589 ^ n8578;
  assign n8552 = n8474 ^ n8442;
  assign n8553 = ~n8475 & n8552;
  assign n8554 = n8553 ^ n8442;
  assign n8591 = n8590 ^ n8554;
  assign n8652 = n8651 ^ n8591;
  assign n8549 = n8533 ^ n8505;
  assign n8550 = n8534 & ~n8549;
  assign n8551 = n8550 ^ n8508;
  assign n8653 = n8652 ^ n8551;
  assign n8691 = n8690 ^ n8653;
  assign n8708 = n8707 ^ n8691;
  assign n8853 = n8547 & ~n8692;
  assign n8854 = ~n8691 & ~n8693;
  assign n8855 = ~n8695 & ~n8854;
  assign n8856 = ~n8853 & n8855;
  assign n8857 = ~n8691 & ~n8692;
  assign n8858 = ~n8696 & ~n8857;
  assign n8859 = ~n8547 & n8858;
  assign n8860 = n8691 & ~n8700;
  assign n8861 = ~n8859 & ~n8860;
  assign n8862 = ~n8856 & n8861;
  assign n8841 = n8563 ^ n8560;
  assign n8842 = ~n8564 & n8841;
  assign n8843 = n8842 ^ n8560;
  assign n8838 = n8618 ^ n8613;
  assign n8839 = n8624 & ~n8838;
  assign n8840 = n8839 ^ n8623;
  assign n8844 = n8843 ^ n8840;
  assign n8835 = n8603 ^ n8596;
  assign n8836 = n8604 & ~n8835;
  assign n8837 = n8836 ^ n8599;
  assign n8845 = n8844 ^ n8837;
  assign n8832 = n8682 ^ n8679;
  assign n8833 = n8686 & ~n8832;
  assign n8834 = n8833 ^ n8685;
  assign n8846 = n8845 ^ n8834;
  assign n8825 = x21 & x56;
  assign n8824 = x20 & x57;
  assign n8826 = n8825 ^ n8824;
  assign n8823 = x19 & x58;
  assign n8827 = n8826 ^ n8823;
  assign n8820 = x29 & x48;
  assign n8819 = x28 & x49;
  assign n8821 = n8820 ^ n8819;
  assign n8818 = x27 & x50;
  assign n8822 = n8821 ^ n8818;
  assign n8828 = n8827 ^ n8822;
  assign n8815 = n8620 ^ n8619;
  assign n8816 = n8622 & ~n8815;
  assign n8817 = n8816 ^ n8621;
  assign n8829 = n8828 ^ n8817;
  assign n8810 = x31 & x46;
  assign n8809 = x30 & x47;
  assign n8811 = n8810 ^ n8809;
  assign n8808 = x14 & x63;
  assign n8812 = n8811 ^ n8808;
  assign n8805 = x37 & x40;
  assign n8804 = x36 & x41;
  assign n8806 = n8805 ^ n8804;
  assign n8803 = x35 & x42;
  assign n8807 = n8806 ^ n8803;
  assign n8813 = n8812 ^ n8807;
  assign n8801 = x15 & x62;
  assign n8800 = ~x38 & x39;
  assign n8802 = n8801 ^ n8800;
  assign n8814 = n8813 ^ n8802;
  assign n8830 = n8829 ^ n8814;
  assign n8797 = n8584 ^ n8581;
  assign n8798 = ~n8588 & ~n8797;
  assign n8799 = n8798 ^ n8587;
  assign n8831 = n8830 ^ n8799;
  assign n8847 = n8846 ^ n8831;
  assign n8790 = x17 & x60;
  assign n8789 = x18 & x59;
  assign n8791 = n8790 ^ n8789;
  assign n8786 = n8615 ^ n8614;
  assign n8787 = n8617 & ~n8786;
  assign n8788 = n8787 ^ n8616;
  assign n8792 = n8791 ^ n8788;
  assign n8783 = n8571 ^ n8568;
  assign n8784 = n8575 & ~n8783;
  assign n8785 = n8784 ^ n8574;
  assign n8793 = n8792 ^ n8785;
  assign n8780 = n8636 ^ n8633;
  assign n8781 = n8640 & ~n8780;
  assign n8782 = n8781 ^ n8639;
  assign n8794 = n8793 ^ n8782;
  assign n8773 = n8669 ^ n8668;
  assign n8774 = n8671 & ~n8773;
  assign n8775 = n8774 ^ n8670;
  assign n8770 = n8593 ^ n8592;
  assign n8771 = n8595 & ~n8770;
  assign n8772 = n8771 ^ n8594;
  assign n8776 = n8775 ^ n8772;
  assign n8767 = n8601 ^ n8600;
  assign n8768 = n8602 & ~n8767;
  assign n8769 = n8768 ^ n4353;
  assign n8777 = n8776 ^ n8769;
  assign n8764 = n8672 ^ n8667;
  assign n8765 = n8678 & ~n8764;
  assign n8766 = n8765 ^ n8677;
  assign n8778 = n8777 ^ n8766;
  assign n8759 = n8664 ^ n8663;
  assign n8760 = n8666 & ~n8759;
  assign n8761 = n8760 ^ n8665;
  assign n8756 = n8674 ^ n8673;
  assign n8757 = n8676 & ~n8756;
  assign n8758 = n8757 ^ n8675;
  assign n8762 = n8761 ^ n8758;
  assign n8753 = n8610 ^ n8609;
  assign n8754 = n8612 & ~n8753;
  assign n8755 = n8754 ^ n8611;
  assign n8763 = n8762 ^ n8755;
  assign n8779 = n8778 ^ n8763;
  assign n8795 = n8794 ^ n8779;
  assign n8750 = n8625 ^ n8605;
  assign n8751 = n8626 & ~n8750;
  assign n8752 = n8751 ^ n8608;
  assign n8796 = n8795 ^ n8752;
  assign n8848 = n8847 ^ n8796;
  assign n8747 = n8687 ^ n8659;
  assign n8748 = ~n8688 & n8747;
  assign n8749 = n8748 ^ n8662;
  assign n8849 = n8848 ^ n8749;
  assign n8738 = x34 & x43;
  assign n8739 = n8738 ^ n4357;
  assign n8737 = x22 & x55;
  assign n8740 = n8739 ^ n8737;
  assign n8734 = x33 & x44;
  assign n8733 = x32 & x45;
  assign n8735 = n8734 ^ n8733;
  assign n8732 = x16 & x61;
  assign n8736 = n8735 ^ n8732;
  assign n8741 = n8740 ^ n8736;
  assign n8729 = x25 & x52;
  assign n8728 = x24 & x53;
  assign n8730 = n8729 ^ n8728;
  assign n8727 = x23 & x54;
  assign n8731 = n8730 ^ n8727;
  assign n8742 = n8741 ^ n8731;
  assign n8724 = n8644 ^ n8641;
  assign n8725 = n8648 & ~n8724;
  assign n8726 = n8725 ^ n8647;
  assign n8743 = n8742 ^ n8726;
  assign n8721 = n8565 ^ n8557;
  assign n8722 = n8577 & ~n8721;
  assign n8723 = n8722 ^ n8576;
  assign n8744 = n8743 ^ n8723;
  assign n8718 = n8589 ^ n8554;
  assign n8719 = n8590 & ~n8718;
  assign n8720 = n8719 ^ n8554;
  assign n8745 = n8744 ^ n8720;
  assign n8715 = n8649 ^ n8627;
  assign n8716 = n8650 & ~n8715;
  assign n8717 = n8716 ^ n8630;
  assign n8746 = n8745 ^ n8717;
  assign n8850 = n8849 ^ n8746;
  assign n8712 = n8651 ^ n8551;
  assign n8713 = n8652 & n8712;
  assign n8714 = n8713 ^ n8551;
  assign n8851 = n8850 ^ n8714;
  assign n8709 = n8689 ^ n8653;
  assign n8710 = n8690 & n8709;
  assign n8711 = n8710 ^ n8656;
  assign n8852 = n8851 ^ n8711;
  assign n8863 = n8862 ^ n8852;
  assign n9003 = n8711 & n8714;
  assign n9004 = n8746 & n8849;
  assign n9005 = ~n9003 & ~n9004;
  assign n9006 = n9005 ^ n8862;
  assign n9007 = ~n8711 & ~n8714;
  assign n9008 = ~n8746 & ~n8849;
  assign n9009 = ~n9007 & ~n9008;
  assign n9010 = n9009 ^ n9005;
  assign n9011 = n9006 & n9010;
  assign n9012 = n8714 ^ n8711;
  assign n9013 = n8849 ^ n8714;
  assign n9014 = ~n8850 & ~n9013;
  assign n9015 = ~n9012 & n9014;
  assign n9016 = ~n9011 & ~n9015;
  assign n8990 = x36 & x42;
  assign n8989 = x35 & x43;
  assign n8991 = n8990 ^ n8989;
  assign n8988 = x23 & x55;
  assign n8992 = n8991 ^ n8988;
  assign n8985 = x38 & x40;
  assign n8984 = x37 & x41;
  assign n8986 = n8985 ^ n8984;
  assign n8983 = x26 & x52;
  assign n8987 = n8986 ^ n8983;
  assign n8993 = n8992 ^ n8987;
  assign n8980 = n8758 ^ n8755;
  assign n8981 = n8762 & ~n8980;
  assign n8982 = n8981 ^ n8761;
  assign n8994 = n8993 ^ n8982;
  assign n8975 = n8788 & n8791;
  assign n8976 = x59 & x60;
  assign n8977 = n2037 & n8976;
  assign n8978 = ~n8975 & ~n8977;
  assign n8971 = n8824 ^ n8823;
  assign n8972 = n8826 & ~n8971;
  assign n8973 = n8972 ^ n8825;
  assign n8968 = n8738 ^ n8737;
  assign n8969 = n8739 & ~n8968;
  assign n8970 = n8969 ^ n4357;
  assign n8974 = n8973 ^ n8970;
  assign n8979 = n8978 ^ n8974;
  assign n8995 = n8994 ^ n8979;
  assign n8965 = n8792 ^ n8782;
  assign n8966 = n8793 & ~n8965;
  assign n8967 = n8966 ^ n8785;
  assign n8996 = n8995 ^ n8967;
  assign n8962 = n8742 ^ n8723;
  assign n8963 = n8743 & ~n8962;
  assign n8964 = n8963 ^ n8726;
  assign n8997 = n8996 ^ n8964;
  assign n8959 = n8829 ^ n8799;
  assign n8960 = ~n8830 & ~n8959;
  assign n8961 = n8960 ^ n8799;
  assign n8998 = n8997 ^ n8961;
  assign n8950 = n8728 ^ n8727;
  assign n8951 = n8730 & ~n8950;
  assign n8952 = n8951 ^ n8729;
  assign n8947 = n8804 ^ n8803;
  assign n8948 = n8806 & ~n8947;
  assign n8949 = n8948 ^ n8805;
  assign n8953 = n8952 ^ n8949;
  assign n8945 = ~x38 & ~n8801;
  assign n8946 = x39 & ~n8945;
  assign n8954 = n8953 ^ n8946;
  assign n8942 = n8772 ^ n8769;
  assign n8943 = n8776 & ~n8942;
  assign n8944 = n8943 ^ n8775;
  assign n8955 = n8954 ^ n8944;
  assign n8937 = n8809 ^ n8808;
  assign n8938 = n8811 & ~n8937;
  assign n8939 = n8938 ^ n8810;
  assign n8934 = n8819 ^ n8818;
  assign n8935 = n8821 & ~n8934;
  assign n8936 = n8935 ^ n8820;
  assign n8940 = n8939 ^ n8936;
  assign n8931 = n8733 ^ n8732;
  assign n8932 = n8735 & ~n8931;
  assign n8933 = n8932 ^ n8734;
  assign n8941 = n8940 ^ n8933;
  assign n8956 = n8955 ^ n8941;
  assign n8926 = n8736 ^ n8731;
  assign n8927 = n8741 & ~n8926;
  assign n8928 = n8927 ^ n8740;
  assign n8923 = n8807 ^ n8802;
  assign n8924 = n8813 & ~n8923;
  assign n8925 = n8924 ^ n8812;
  assign n8929 = n8928 ^ n8925;
  assign n8920 = n8827 ^ n8817;
  assign n8921 = ~n8828 & n8920;
  assign n8922 = n8921 ^ n8817;
  assign n8930 = n8929 ^ n8922;
  assign n8957 = n8956 ^ n8930;
  assign n8917 = n8777 ^ n8763;
  assign n8918 = n8778 & ~n8917;
  assign n8919 = n8918 ^ n8766;
  assign n8958 = n8957 ^ n8919;
  assign n8999 = n8998 ^ n8958;
  assign n8914 = n8720 ^ n8717;
  assign n8915 = ~n8745 & n8914;
  assign n8916 = n8915 ^ n8717;
  assign n9000 = n8999 ^ n8916;
  assign n8909 = n8845 ^ n8831;
  assign n8910 = n8846 & n8909;
  assign n8911 = n8910 ^ n8834;
  assign n8906 = n8794 ^ n8752;
  assign n8907 = ~n8795 & n8906;
  assign n8908 = n8907 ^ n8752;
  assign n8912 = n8911 ^ n8908;
  assign n8899 = x34 & x44;
  assign n8898 = x33 & x45;
  assign n8900 = n8899 ^ n8898;
  assign n8897 = x32 & x46;
  assign n8901 = n8900 ^ n8897;
  assign n8894 = x31 & x47;
  assign n8893 = x30 & x48;
  assign n8895 = n8894 ^ n8893;
  assign n8892 = x20 & x58;
  assign n8896 = n8895 ^ n8892;
  assign n8902 = n8901 ^ n8896;
  assign n8889 = x25 & x53;
  assign n8888 = x24 & x54;
  assign n8890 = n8889 ^ n8888;
  assign n8887 = x22 & x56;
  assign n8891 = n8890 ^ n8887;
  assign n8903 = n8902 ^ n8891;
  assign n8882 = x21 & x57;
  assign n8881 = x19 & x59;
  assign n8883 = n8882 ^ n8881;
  assign n8880 = x18 & x60;
  assign n8884 = n8883 ^ n8880;
  assign n8877 = x17 & x61;
  assign n8876 = x16 & x62;
  assign n8878 = n8877 ^ n8876;
  assign n8875 = x15 & x63;
  assign n8879 = n8878 ^ n8875;
  assign n8885 = n8884 ^ n8879;
  assign n8872 = x29 & x49;
  assign n8871 = x28 & x50;
  assign n8873 = n8872 ^ n8871;
  assign n8870 = x27 & x51;
  assign n8874 = n8873 ^ n8870;
  assign n8886 = n8885 ^ n8874;
  assign n8904 = n8903 ^ n8886;
  assign n8867 = n8843 ^ n8837;
  assign n8868 = ~n8844 & n8867;
  assign n8869 = n8868 ^ n8837;
  assign n8905 = n8904 ^ n8869;
  assign n8913 = n8912 ^ n8905;
  assign n9001 = n9000 ^ n8913;
  assign n8864 = n8847 ^ n8749;
  assign n8865 = n8848 & n8864;
  assign n8866 = n8865 ^ n8749;
  assign n9002 = n9001 ^ n8866;
  assign n9017 = n9016 ^ n9002;
  assign n9156 = n8862 & ~n9007;
  assign n9157 = ~n9002 & ~n9008;
  assign n9158 = ~n9003 & ~n9157;
  assign n9159 = ~n9156 & n9158;
  assign n9160 = ~n9002 & ~n9007;
  assign n9161 = ~n9004 & ~n9160;
  assign n9162 = ~n8862 & n9161;
  assign n9163 = ~n9005 & ~n9008;
  assign n9164 = n9002 & ~n9163;
  assign n9165 = ~n9162 & ~n9164;
  assign n9166 = ~n9159 & n9165;
  assign n9142 = n8881 ^ n8880;
  assign n9143 = n8883 & ~n9142;
  assign n9144 = n9143 ^ n8882;
  assign n9139 = n8871 ^ n8870;
  assign n9140 = n8873 & ~n9139;
  assign n9141 = n9140 ^ n8872;
  assign n9145 = n9144 ^ n9141;
  assign n9136 = n8888 ^ n8887;
  assign n9137 = n8890 & ~n9136;
  assign n9138 = n9137 ^ n8889;
  assign n9146 = n9145 ^ n9138;
  assign n9133 = n8992 ^ n8982;
  assign n9134 = ~n8993 & n9133;
  assign n9135 = n9134 ^ n8982;
  assign n9147 = n9146 ^ n9135;
  assign n9128 = x36 & x43;
  assign n9129 = n9128 ^ n4755;
  assign n9127 = x23 & x56;
  assign n9130 = n9129 ^ n9127;
  assign n9124 = x35 & x44;
  assign n9123 = x34 & x45;
  assign n9125 = n9124 ^ n9123;
  assign n9122 = x16 & x63;
  assign n9126 = n9125 ^ n9122;
  assign n9131 = n9130 ^ n9126;
  assign n9119 = n8978 ^ n8973;
  assign n9120 = ~n8974 & ~n9119;
  assign n9121 = n9120 ^ n8978;
  assign n9132 = n9131 ^ n9121;
  assign n9148 = n9147 ^ n9132;
  assign n9114 = x18 & x61;
  assign n9111 = n8984 ^ n8983;
  assign n9112 = n8986 & ~n9111;
  assign n9113 = n9112 ^ n8985;
  assign n9115 = n9114 ^ n9113;
  assign n9108 = n8989 ^ n8988;
  assign n9109 = n8991 & ~n9108;
  assign n9110 = n9109 ^ n8990;
  assign n9116 = n9115 ^ n9110;
  assign n9105 = n8896 ^ n8891;
  assign n9106 = n8902 & ~n9105;
  assign n9107 = n9106 ^ n8901;
  assign n9117 = n9116 ^ n9107;
  assign n9100 = n8893 ^ n8892;
  assign n9101 = n8895 & ~n9100;
  assign n9102 = n9101 ^ n8894;
  assign n9097 = n8898 ^ n8897;
  assign n9098 = n8900 & ~n9097;
  assign n9099 = n9098 ^ n8899;
  assign n9103 = n9102 ^ n9099;
  assign n9094 = n8876 ^ n8875;
  assign n9095 = n8878 & ~n9094;
  assign n9096 = n9095 ^ n8877;
  assign n9104 = n9103 ^ n9096;
  assign n9118 = n9117 ^ n9104;
  assign n9149 = n9148 ^ n9118;
  assign n9091 = n8903 ^ n8869;
  assign n9092 = ~n8904 & n9091;
  assign n9093 = n9092 ^ n8869;
  assign n9150 = n9149 ^ n9093;
  assign n9088 = n8964 ^ n8961;
  assign n9089 = n8997 & ~n9088;
  assign n9090 = n9089 ^ n8961;
  assign n9151 = n9150 ^ n9090;
  assign n9085 = n8908 ^ n8905;
  assign n9086 = n8912 & ~n9085;
  assign n9087 = n9086 ^ n8911;
  assign n9152 = n9151 ^ n9087;
  assign n9082 = n8998 ^ n8916;
  assign n9083 = ~n8999 & n9082;
  assign n9084 = n9083 ^ n8916;
  assign n9153 = n9152 ^ n9084;
  assign n9073 = x30 & x49;
  assign n9072 = x29 & x50;
  assign n9074 = n9073 ^ n9072;
  assign n9071 = x22 & x57;
  assign n9075 = n9074 ^ n9071;
  assign n9068 = x33 & x46;
  assign n9067 = x32 & x47;
  assign n9069 = n9068 ^ n9067;
  assign n9066 = x31 & x48;
  assign n9070 = n9069 ^ n9066;
  assign n9076 = n9075 ^ n9070;
  assign n9063 = x21 & x58;
  assign n9062 = x20 & x59;
  assign n9064 = n9063 ^ n9062;
  assign n9061 = x19 & x60;
  assign n9065 = n9064 ^ n9061;
  assign n9077 = n9076 ^ n9065;
  assign n9058 = n8954 ^ n8941;
  assign n9059 = n8955 & ~n9058;
  assign n9060 = n9059 ^ n8944;
  assign n9078 = n9077 ^ n9060;
  assign n9053 = x39 & x40;
  assign n9052 = x38 & x41;
  assign n9054 = n9053 ^ n9052;
  assign n9051 = x37 & x42;
  assign n9055 = n9054 ^ n9051;
  assign n9048 = x17 & x62;
  assign n9047 = x28 & x51;
  assign n9049 = n9048 ^ n9047;
  assign n9050 = n9049 ^ x40;
  assign n9056 = n9055 ^ n9050;
  assign n9044 = x25 & x54;
  assign n9045 = n9044 ^ n4926;
  assign n9043 = x24 & x55;
  assign n9046 = n9045 ^ n9043;
  assign n9057 = n9056 ^ n9046;
  assign n9079 = n9078 ^ n9057;
  assign n9040 = n8930 ^ n8919;
  assign n9041 = n8957 & ~n9040;
  assign n9042 = n9041 ^ n8956;
  assign n9080 = n9079 ^ n9042;
  assign n9033 = n8949 ^ n8946;
  assign n9034 = n8953 & ~n9033;
  assign n9035 = n9034 ^ n8952;
  assign n9030 = n8879 ^ n8874;
  assign n9031 = n8885 & ~n9030;
  assign n9032 = n9031 ^ n8884;
  assign n9036 = n9035 ^ n9032;
  assign n9027 = n8936 ^ n8933;
  assign n9028 = n8940 & ~n9027;
  assign n9029 = n9028 ^ n8939;
  assign n9037 = n9036 ^ n9029;
  assign n9024 = n8925 ^ n8922;
  assign n9025 = n8929 & ~n9024;
  assign n9026 = n9025 ^ n8928;
  assign n9038 = n9037 ^ n9026;
  assign n9021 = n8994 ^ n8967;
  assign n9022 = n8995 & n9021;
  assign n9023 = n9022 ^ n8967;
  assign n9039 = n9038 ^ n9023;
  assign n9081 = n9080 ^ n9039;
  assign n9154 = n9153 ^ n9081;
  assign n9018 = n8913 ^ n8866;
  assign n9019 = n9001 & n9018;
  assign n9020 = n9019 ^ n9000;
  assign n9155 = n9154 ^ n9020;
  assign n9167 = n9166 ^ n9155;
  assign n9306 = n9020 & n9154;
  assign n9307 = ~n9166 & ~n9306;
  assign n9308 = ~n9020 & ~n9154;
  assign n9309 = ~n9307 & ~n9308;
  assign n9294 = n9130 ^ n9121;
  assign n9295 = ~n9131 & ~n9294;
  assign n9296 = n9295 ^ n9121;
  assign n9291 = n9032 ^ n9029;
  assign n9292 = n9036 & ~n9291;
  assign n9293 = n9292 ^ n9035;
  assign n9297 = n9296 ^ n9293;
  assign n9286 = n9044 ^ n9043;
  assign n9287 = n9045 & ~n9286;
  assign n9288 = n9287 ^ n4926;
  assign n9283 = n9123 ^ n9122;
  assign n9284 = n9125 & ~n9283;
  assign n9285 = n9284 ^ n9124;
  assign n9289 = n9288 ^ n9285;
  assign n9280 = n9128 ^ n9127;
  assign n9281 = n9129 & ~n9280;
  assign n9282 = n9281 ^ n4755;
  assign n9290 = n9289 ^ n9282;
  assign n9298 = n9297 ^ n9290;
  assign n9273 = n9072 ^ n9071;
  assign n9274 = n9074 & ~n9273;
  assign n9275 = n9274 ^ n9073;
  assign n9270 = n9067 ^ n9066;
  assign n9271 = n9069 & ~n9270;
  assign n9272 = n9271 ^ n9068;
  assign n9276 = n9275 ^ n9272;
  assign n9267 = n9062 ^ n9061;
  assign n9268 = n9064 & ~n9267;
  assign n9269 = n9268 ^ n9063;
  assign n9277 = n9276 ^ n9269;
  assign n9264 = n9050 ^ n9046;
  assign n9265 = n9056 & ~n9264;
  assign n9266 = n9265 ^ n9055;
  assign n9278 = n9277 ^ n9266;
  assign n9261 = n9070 ^ n9065;
  assign n9262 = n9076 & ~n9261;
  assign n9263 = n9262 ^ n9075;
  assign n9279 = n9278 ^ n9263;
  assign n9299 = n9298 ^ n9279;
  assign n9258 = n9077 ^ n9057;
  assign n9259 = n9078 & ~n9258;
  assign n9260 = n9259 ^ n9060;
  assign n9300 = n9299 ^ n9260;
  assign n9251 = n9141 ^ n9138;
  assign n9252 = n9145 & ~n9251;
  assign n9253 = n9252 ^ n9144;
  assign n9248 = n9099 ^ n9096;
  assign n9249 = n9103 & ~n9248;
  assign n9250 = n9249 ^ n9102;
  assign n9254 = n9253 ^ n9250;
  assign n9245 = n9114 ^ n9110;
  assign n9246 = n9115 & ~n9245;
  assign n9247 = n9246 ^ n9113;
  assign n9255 = n9254 ^ n9247;
  assign n9242 = n9107 ^ n9104;
  assign n9243 = n9117 & ~n9242;
  assign n9244 = n9243 ^ n9116;
  assign n9256 = n9255 ^ n9244;
  assign n9239 = n9146 ^ n9132;
  assign n9240 = n9147 & n9239;
  assign n9241 = n9240 ^ n9135;
  assign n9257 = n9256 ^ n9241;
  assign n9301 = n9300 ^ n9257;
  assign n9236 = n9079 ^ n9039;
  assign n9237 = n9080 & ~n9236;
  assign n9238 = n9237 ^ n9042;
  assign n9302 = n9301 ^ n9238;
  assign n9226 = x51 & n7292;
  assign n9227 = ~n9048 & ~n9226;
  assign n9228 = ~x40 & ~n9047;
  assign n9229 = ~n9227 & ~n9228;
  assign n9224 = x18 & x62;
  assign n9223 = x19 & x61;
  assign n9225 = n9224 ^ n9223;
  assign n9230 = n9229 ^ n9225;
  assign n9219 = x36 & x44;
  assign n9218 = x35 & x45;
  assign n9220 = n9219 ^ n9218;
  assign n9217 = x34 & x46;
  assign n9221 = n9220 ^ n9217;
  assign n9214 = x33 & x47;
  assign n9213 = x29 & x51;
  assign n9215 = n9214 ^ n9213;
  assign n9212 = x17 & x63;
  assign n9216 = n9215 ^ n9212;
  assign n9222 = n9221 ^ n9216;
  assign n9231 = n9230 ^ n9222;
  assign n9207 = x39 & x41;
  assign n9206 = x28 & x52;
  assign n9208 = n9207 ^ n9206;
  assign n9205 = x27 & x53;
  assign n9209 = n9208 ^ n9205;
  assign n9202 = x38 & x42;
  assign n9201 = x37 & x43;
  assign n9203 = n9202 ^ n9201;
  assign n9200 = x25 & x55;
  assign n9204 = n9203 ^ n9200;
  assign n9210 = n9209 ^ n9204;
  assign n9197 = x26 & x54;
  assign n9196 = x24 & x56;
  assign n9198 = n9197 ^ n9196;
  assign n9195 = x23 & x57;
  assign n9199 = n9198 ^ n9195;
  assign n9211 = n9210 ^ n9199;
  assign n9232 = n9231 ^ n9211;
  assign n9190 = x22 & x58;
  assign n9189 = x21 & x59;
  assign n9191 = n9190 ^ n9189;
  assign n9188 = x20 & x60;
  assign n9192 = n9191 ^ n9188;
  assign n9185 = x32 & x48;
  assign n9184 = x31 & x49;
  assign n9186 = n9185 ^ n9184;
  assign n9183 = x30 & x50;
  assign n9187 = n9186 ^ n9183;
  assign n9193 = n9192 ^ n9187;
  assign n9180 = n9052 ^ n9051;
  assign n9181 = n9054 & ~n9180;
  assign n9182 = n9181 ^ n9053;
  assign n9194 = n9193 ^ n9182;
  assign n9233 = n9232 ^ n9194;
  assign n9177 = n9118 ^ n9093;
  assign n9178 = ~n9149 & ~n9177;
  assign n9179 = n9178 ^ n9148;
  assign n9234 = n9233 ^ n9179;
  assign n9174 = n9026 ^ n9023;
  assign n9175 = ~n9038 & n9174;
  assign n9176 = n9175 ^ n9023;
  assign n9235 = n9234 ^ n9176;
  assign n9303 = n9302 ^ n9235;
  assign n9171 = n9090 ^ n9087;
  assign n9172 = ~n9151 & ~n9171;
  assign n9173 = n9172 ^ n9087;
  assign n9304 = n9303 ^ n9173;
  assign n9168 = n9152 ^ n9081;
  assign n9169 = n9153 & ~n9168;
  assign n9170 = n9169 ^ n9084;
  assign n9305 = n9304 ^ n9170;
  assign n9310 = n9309 ^ n9305;
  assign n9439 = ~n9235 & ~n9302;
  assign n9440 = ~n9173 & ~n9439;
  assign n9441 = ~n9170 & n9440;
  assign n9442 = n9235 & n9302;
  assign n9443 = ~n9441 & ~n9442;
  assign n9444 = n9170 & n9173;
  assign n9445 = ~n9443 & ~n9444;
  assign n9446 = ~n9309 & n9445;
  assign n9448 = ~n9173 & n9442;
  assign n9447 = n9173 & n9439;
  assign n9449 = n9448 ^ n9447;
  assign n9450 = n9170 & n9449;
  assign n9451 = n9450 ^ n9448;
  assign n9452 = ~n9446 & ~n9451;
  assign n9453 = ~n9170 & ~n9447;
  assign n9454 = ~n9440 & ~n9442;
  assign n9455 = ~n9453 & n9454;
  assign n9456 = n9309 & n9455;
  assign n9457 = n9452 & ~n9456;
  assign n9426 = n9196 ^ n9195;
  assign n9427 = n9198 & ~n9426;
  assign n9428 = n9427 ^ n9197;
  assign n9423 = n9206 ^ n9205;
  assign n9424 = n9208 & ~n9423;
  assign n9425 = n9424 ^ n9207;
  assign n9429 = n9428 ^ n9425;
  assign n9420 = n9201 ^ n9200;
  assign n9421 = n9203 & ~n9420;
  assign n9422 = n9421 ^ n9202;
  assign n9430 = n9429 ^ n9422;
  assign n9417 = n9192 ^ n9182;
  assign n9418 = ~n9193 & n9417;
  assign n9419 = n9418 ^ n9182;
  assign n9431 = n9430 ^ n9419;
  assign n9414 = n9204 ^ n9199;
  assign n9415 = n9210 & ~n9414;
  assign n9416 = n9415 ^ n9209;
  assign n9432 = n9431 ^ n9416;
  assign n9411 = n9211 ^ n9194;
  assign n9412 = n9232 & ~n9411;
  assign n9413 = n9412 ^ n9231;
  assign n9433 = n9432 ^ n9413;
  assign n9405 = n9225 & n9229;
  assign n9406 = n2253 & n8432;
  assign n9407 = ~n9405 & ~n9406;
  assign n9401 = x32 & x49;
  assign n9400 = x31 & x50;
  assign n9402 = n9401 ^ n9400;
  assign n9399 = x30 & x51;
  assign n9403 = n9402 ^ n9399;
  assign n9396 = n9218 ^ n9217;
  assign n9397 = n9220 & ~n9396;
  assign n9398 = n9397 ^ n9219;
  assign n9404 = n9403 ^ n9398;
  assign n9408 = n9407 ^ n9404;
  assign n9393 = n9230 ^ n9221;
  assign n9394 = ~n9222 & n9393;
  assign n9395 = n9394 ^ n9230;
  assign n9409 = n9408 ^ n9395;
  assign n9388 = n9213 ^ n9212;
  assign n9389 = n9215 & ~n9388;
  assign n9390 = n9389 ^ n9214;
  assign n9385 = n9189 ^ n9188;
  assign n9386 = n9191 & ~n9385;
  assign n9387 = n9386 ^ n9190;
  assign n9391 = n9390 ^ n9387;
  assign n9382 = n9184 ^ n9183;
  assign n9383 = n9186 & ~n9382;
  assign n9384 = n9383 ^ n9185;
  assign n9392 = n9391 ^ n9384;
  assign n9410 = n9409 ^ n9392;
  assign n9434 = n9433 ^ n9410;
  assign n9379 = n9179 ^ n9176;
  assign n9380 = n9234 & ~n9379;
  assign n9381 = n9380 ^ n9176;
  assign n9435 = n9434 ^ n9381;
  assign n9372 = x39 & x42;
  assign n9371 = x38 & x43;
  assign n9373 = n9372 ^ n9371;
  assign n9370 = x27 & x54;
  assign n9374 = n9373 ^ n9370;
  assign n9367 = n9272 ^ n9269;
  assign n9368 = n9276 & ~n9367;
  assign n9369 = n9368 ^ n9275;
  assign n9375 = n9374 ^ n9369;
  assign n9364 = n9285 ^ n9282;
  assign n9365 = n9289 & ~n9364;
  assign n9366 = n9365 ^ n9288;
  assign n9376 = n9375 ^ n9366;
  assign n9361 = n9266 ^ n9263;
  assign n9362 = n9278 & ~n9361;
  assign n9363 = n9362 ^ n9277;
  assign n9377 = n9376 ^ n9363;
  assign n9358 = n9293 ^ n9290;
  assign n9359 = ~n9297 & ~n9358;
  assign n9360 = n9359 ^ n9296;
  assign n9378 = n9377 ^ n9360;
  assign n9436 = n9435 ^ n9378;
  assign n9355 = n9300 ^ n9238;
  assign n9356 = n9301 & ~n9355;
  assign n9357 = n9356 ^ n9238;
  assign n9437 = n9436 ^ n9357;
  assign n9346 = x29 & x52;
  assign n9347 = n9346 ^ n4971;
  assign n9345 = x26 & x55;
  assign n9348 = n9347 ^ n9345;
  assign n9342 = x37 & x44;
  assign n9341 = x36 & x45;
  assign n9343 = n9342 ^ n9341;
  assign n9340 = x35 & x46;
  assign n9344 = n9343 ^ n9340;
  assign n9349 = n9348 ^ n9344;
  assign n9337 = x21 & x60;
  assign n9336 = x20 & x61;
  assign n9338 = n9337 ^ n9336;
  assign n9335 = x18 & x63;
  assign n9339 = n9338 ^ n9335;
  assign n9350 = n9349 ^ n9339;
  assign n9332 = n9250 ^ n9247;
  assign n9333 = n9254 & ~n9332;
  assign n9334 = n9333 ^ n9253;
  assign n9351 = n9350 ^ n9334;
  assign n9327 = x34 & x47;
  assign n9326 = x33 & x48;
  assign n9328 = n9327 ^ n9326;
  assign n9325 = x24 & x57;
  assign n9329 = n9328 ^ n9325;
  assign n9322 = x25 & x56;
  assign n9321 = x23 & x58;
  assign n9323 = n9322 ^ n9321;
  assign n9320 = x22 & x59;
  assign n9324 = n9323 ^ n9320;
  assign n9330 = n9329 ^ n9324;
  assign n9318 = x19 & x62;
  assign n9317 = ~x40 & x41;
  assign n9319 = n9318 ^ n9317;
  assign n9331 = n9330 ^ n9319;
  assign n9352 = n9351 ^ n9331;
  assign n9314 = n9298 ^ n9260;
  assign n9315 = n9299 & ~n9314;
  assign n9316 = n9315 ^ n9260;
  assign n9353 = n9352 ^ n9316;
  assign n9311 = n9244 ^ n9241;
  assign n9312 = ~n9256 & n9311;
  assign n9313 = n9312 ^ n9241;
  assign n9354 = n9353 ^ n9313;
  assign n9438 = n9437 ^ n9354;
  assign n9458 = n9457 ^ n9438;
  assign n9587 = ~n9170 & ~n9173;
  assign n9588 = ~n9308 & ~n9587;
  assign n9589 = ~n9307 & n9588;
  assign n9590 = ~n9444 & ~n9589;
  assign n9591 = ~n9438 & ~n9439;
  assign n9592 = ~n9590 & ~n9591;
  assign n9593 = ~n9438 & ~n9444;
  assign n9594 = ~n9442 & ~n9593;
  assign n9595 = n9309 & n9594;
  assign n9596 = n9438 & n9443;
  assign n9597 = ~n9595 & ~n9596;
  assign n9598 = ~n9592 & n9597;
  assign n9575 = x19 & x63;
  assign n9572 = n9371 ^ n9370;
  assign n9573 = n9373 & ~n9572;
  assign n9574 = n9573 ^ n9372;
  assign n9576 = n9575 ^ n9574;
  assign n9570 = ~x40 & ~n9318;
  assign n9571 = x41 & ~n9570;
  assign n9577 = n9576 ^ n9571;
  assign n9567 = n9324 ^ n9319;
  assign n9568 = n9330 & ~n9567;
  assign n9569 = n9568 ^ n9329;
  assign n9578 = n9577 ^ n9569;
  assign n9564 = n9407 ^ n9398;
  assign n9565 = ~n9404 & ~n9564;
  assign n9566 = n9565 ^ n9407;
  assign n9579 = n9578 ^ n9566;
  assign n9561 = n9350 ^ n9331;
  assign n9562 = n9351 & ~n9561;
  assign n9563 = n9562 ^ n9334;
  assign n9580 = n9579 ^ n9563;
  assign n9554 = n9321 ^ n9320;
  assign n9555 = n9323 & ~n9554;
  assign n9556 = n9555 ^ n9322;
  assign n9551 = n9336 ^ n9335;
  assign n9552 = n9338 & ~n9551;
  assign n9553 = n9552 ^ n9337;
  assign n9557 = n9556 ^ n9553;
  assign n9548 = n9341 ^ n9340;
  assign n9549 = n9343 & ~n9548;
  assign n9550 = n9549 ^ n9342;
  assign n9558 = n9557 ^ n9550;
  assign n9545 = n9344 ^ n9339;
  assign n9546 = n9349 & ~n9545;
  assign n9547 = n9546 ^ n9348;
  assign n9559 = n9558 ^ n9547;
  assign n9540 = n9346 ^ n9345;
  assign n9541 = n9347 & ~n9540;
  assign n9542 = n9541 ^ n4971;
  assign n9537 = n9326 ^ n9325;
  assign n9538 = n9328 & ~n9537;
  assign n9539 = n9538 ^ n9327;
  assign n9543 = n9542 ^ n9539;
  assign n9534 = n9400 ^ n9399;
  assign n9535 = n9402 & ~n9534;
  assign n9536 = n9535 ^ n9401;
  assign n9544 = n9543 ^ n9536;
  assign n9560 = n9559 ^ n9544;
  assign n9581 = n9580 ^ n9560;
  assign n9528 = n5133 ^ n4974;
  assign n9527 = x25 & x57;
  assign n9529 = n9528 ^ n9527;
  assign n9524 = n9425 ^ n9422;
  assign n9525 = n9429 & ~n9524;
  assign n9526 = n9525 ^ n9428;
  assign n9530 = n9529 ^ n9526;
  assign n9521 = n9387 ^ n9384;
  assign n9522 = n9391 & ~n9521;
  assign n9523 = n9522 ^ n9390;
  assign n9531 = n9530 ^ n9523;
  assign n9518 = n9430 ^ n9416;
  assign n9519 = n9431 & ~n9518;
  assign n9520 = n9519 ^ n9419;
  assign n9532 = n9531 ^ n9520;
  assign n9515 = n9395 ^ n9392;
  assign n9516 = ~n9409 & ~n9515;
  assign n9517 = n9516 ^ n9408;
  assign n9533 = n9532 ^ n9517;
  assign n9582 = n9581 ^ n9533;
  assign n9512 = n9352 ^ n9313;
  assign n9513 = n9353 & ~n9512;
  assign n9514 = n9513 ^ n9316;
  assign n9583 = n9582 ^ n9514;
  assign n9503 = x40 & x42;
  assign n9502 = x30 & x52;
  assign n9504 = n9503 ^ n9502;
  assign n9501 = x29 & x53;
  assign n9505 = n9504 ^ n9501;
  assign n9498 = x37 & x45;
  assign n9497 = x36 & x46;
  assign n9499 = n9498 ^ n9497;
  assign n9496 = x35 & x47;
  assign n9500 = n9499 ^ n9496;
  assign n9506 = n9505 ^ n9500;
  assign n9493 = x39 & x43;
  assign n9492 = x38 & x44;
  assign n9494 = n9493 ^ n9492;
  assign n9491 = x26 & x56;
  assign n9495 = n9494 ^ n9491;
  assign n9507 = n9506 ^ n9495;
  assign n9486 = x31 & x51;
  assign n9485 = x21 & x61;
  assign n9487 = n9486 ^ n9485;
  assign n9484 = x20 & x62;
  assign n9488 = n9487 ^ n9484;
  assign n9481 = x24 & x58;
  assign n9480 = x23 & x59;
  assign n9482 = n9481 ^ n9480;
  assign n9479 = x22 & x60;
  assign n9483 = n9482 ^ n9479;
  assign n9489 = n9488 ^ n9483;
  assign n9476 = x34 & x48;
  assign n9475 = x33 & x49;
  assign n9477 = n9476 ^ n9475;
  assign n9474 = x32 & x50;
  assign n9478 = n9477 ^ n9474;
  assign n9490 = n9489 ^ n9478;
  assign n9508 = n9507 ^ n9490;
  assign n9471 = n9374 ^ n9366;
  assign n9472 = n9375 & ~n9471;
  assign n9473 = n9472 ^ n9369;
  assign n9509 = n9508 ^ n9473;
  assign n9468 = n9363 ^ n9360;
  assign n9469 = ~n9377 & ~n9468;
  assign n9470 = n9469 ^ n9360;
  assign n9510 = n9509 ^ n9470;
  assign n9465 = n9432 ^ n9410;
  assign n9466 = n9433 & n9465;
  assign n9467 = n9466 ^ n9413;
  assign n9511 = n9510 ^ n9467;
  assign n9584 = n9583 ^ n9511;
  assign n9462 = n9434 ^ n9378;
  assign n9463 = ~n9435 & ~n9462;
  assign n9464 = n9463 ^ n9381;
  assign n9585 = n9584 ^ n9464;
  assign n9459 = n9357 ^ n9354;
  assign n9460 = n9437 & ~n9459;
  assign n9461 = n9460 ^ n9436;
  assign n9586 = n9585 ^ n9461;
  assign n9599 = n9598 ^ n9586;
  assign n9723 = ~n9464 & n9511;
  assign n9724 = ~n9583 & n9723;
  assign n9725 = n9461 & ~n9724;
  assign n9726 = n9583 ^ n9464;
  assign n9727 = n9584 & n9726;
  assign n9728 = n9727 ^ n9464;
  assign n9729 = ~n9725 & ~n9728;
  assign n9730 = n9598 & n9729;
  assign n9731 = n9464 & ~n9511;
  assign n9732 = n9583 & n9731;
  assign n9733 = n9732 ^ n9724;
  assign n9734 = n9461 & n9733;
  assign n9735 = n9734 ^ n9724;
  assign n9736 = ~n9730 & ~n9735;
  assign n9737 = ~n9461 & ~n9732;
  assign n9738 = n9728 & ~n9737;
  assign n9739 = ~n9598 & n9738;
  assign n9740 = n9736 & ~n9739;
  assign n9710 = n9485 ^ n9484;
  assign n9711 = n9487 & ~n9710;
  assign n9712 = n9711 ^ n9486;
  assign n9707 = n9475 ^ n9474;
  assign n9708 = n9477 & ~n9707;
  assign n9709 = n9708 ^ n9476;
  assign n9713 = n9712 ^ n9709;
  assign n9704 = n9527 ^ n5133;
  assign n9705 = n9528 & ~n9704;
  assign n9706 = n9705 ^ n4974;
  assign n9714 = n9713 ^ n9706;
  assign n9699 = n9497 ^ n9496;
  assign n9700 = n9499 & ~n9699;
  assign n9701 = n9700 ^ n9498;
  assign n9696 = n9492 ^ n9491;
  assign n9697 = n9494 & ~n9696;
  assign n9698 = n9697 ^ n9493;
  assign n9702 = n9701 ^ n9698;
  assign n9693 = n9480 ^ n9479;
  assign n9694 = n9482 & ~n9693;
  assign n9695 = n9694 ^ n9481;
  assign n9703 = n9702 ^ n9695;
  assign n9715 = n9714 ^ n9703;
  assign n9690 = n9500 ^ n9495;
  assign n9691 = n9506 & ~n9690;
  assign n9692 = n9691 ^ n9505;
  assign n9716 = n9715 ^ n9692;
  assign n9687 = n9547 ^ n9544;
  assign n9688 = n9559 & ~n9687;
  assign n9689 = n9688 ^ n9558;
  assign n9717 = n9716 ^ n9689;
  assign n9684 = n9507 ^ n9473;
  assign n9685 = ~n9508 & n9684;
  assign n9686 = n9685 ^ n9473;
  assign n9718 = n9717 ^ n9686;
  assign n9677 = n9539 ^ n9536;
  assign n9678 = n9543 & ~n9677;
  assign n9679 = n9678 ^ n9542;
  assign n9674 = n9483 ^ n9478;
  assign n9675 = n9489 & ~n9674;
  assign n9676 = n9675 ^ n9488;
  assign n9680 = n9679 ^ n9676;
  assign n9671 = n9553 ^ n9550;
  assign n9672 = n9557 & ~n9671;
  assign n9673 = n9672 ^ n9556;
  assign n9681 = n9680 ^ n9673;
  assign n9668 = n9577 ^ n9566;
  assign n9669 = ~n9578 & ~n9668;
  assign n9670 = n9669 ^ n9566;
  assign n9682 = n9681 ^ n9670;
  assign n9663 = x23 & x60;
  assign n9662 = x24 & x59;
  assign n9664 = n9663 ^ n9662;
  assign n9659 = n9502 ^ n9501;
  assign n9660 = n9504 & ~n9659;
  assign n9661 = n9660 ^ n9503;
  assign n9665 = n9664 ^ n9661;
  assign n9656 = x31 & x52;
  assign n9655 = x30 & x53;
  assign n9657 = n9656 ^ n9655;
  assign n9654 = x28 & x55;
  assign n9658 = n9657 ^ n9654;
  assign n9666 = n9665 ^ n9658;
  assign n9651 = n9575 ^ n9571;
  assign n9652 = n9576 & ~n9651;
  assign n9653 = n9652 ^ n9574;
  assign n9667 = n9666 ^ n9653;
  assign n9683 = n9682 ^ n9667;
  assign n9719 = n9718 ^ n9683;
  assign n9648 = n9509 ^ n9467;
  assign n9649 = ~n9510 & ~n9648;
  assign n9650 = n9649 ^ n9470;
  assign n9720 = n9719 ^ n9650;
  assign n9645 = n9581 ^ n9514;
  assign n9646 = ~n9582 & ~n9645;
  assign n9647 = n9646 ^ n9514;
  assign n9721 = n9720 ^ n9647;
  assign n9636 = x32 & x51;
  assign n9635 = x26 & x57;
  assign n9637 = n9636 ^ n9635;
  assign n9634 = x25 & x58;
  assign n9638 = n9637 ^ n9634;
  assign n9631 = x38 & x45;
  assign n9630 = x37 & x46;
  assign n9632 = n9631 ^ n9630;
  assign n9629 = x36 & x47;
  assign n9633 = n9632 ^ n9629;
  assign n9639 = n9638 ^ n9633;
  assign n9626 = x27 & x56;
  assign n9625 = x22 & x61;
  assign n9627 = n9626 ^ n9625;
  assign n9624 = x20 & x63;
  assign n9628 = n9627 ^ n9624;
  assign n9640 = n9639 ^ n9628;
  assign n9619 = x40 & x43;
  assign n9618 = x39 & x44;
  assign n9620 = n9619 ^ n9618;
  assign n9617 = x29 & x54;
  assign n9621 = n9620 ^ n9617;
  assign n9614 = x35 & x48;
  assign n9613 = x34 & x49;
  assign n9615 = n9614 ^ n9613;
  assign n9612 = x33 & x50;
  assign n9616 = n9615 ^ n9612;
  assign n9622 = n9621 ^ n9616;
  assign n9610 = x21 & x62;
  assign n9609 = ~x41 & x42;
  assign n9611 = n9610 ^ n9609;
  assign n9623 = n9622 ^ n9611;
  assign n9641 = n9640 ^ n9623;
  assign n9606 = n9529 ^ n9523;
  assign n9607 = n9530 & ~n9606;
  assign n9608 = n9607 ^ n9526;
  assign n9642 = n9641 ^ n9608;
  assign n9603 = n9520 ^ n9517;
  assign n9604 = ~n9532 & ~n9603;
  assign n9605 = n9604 ^ n9517;
  assign n9643 = n9642 ^ n9605;
  assign n9600 = n9579 ^ n9560;
  assign n9601 = ~n9580 & n9600;
  assign n9602 = n9601 ^ n9563;
  assign n9644 = n9643 ^ n9602;
  assign n9722 = n9721 ^ n9644;
  assign n9741 = n9740 ^ n9722;
  assign n9866 = n9461 & n9583;
  assign n9867 = n9598 & ~n9866;
  assign n9868 = ~n9461 & ~n9583;
  assign n9869 = n9722 & ~n9731;
  assign n9870 = ~n9868 & ~n9869;
  assign n9871 = ~n9867 & n9870;
  assign n9872 = ~n9731 & n9868;
  assign n9873 = ~n9722 & ~n9872;
  assign n9874 = n9598 & ~n9873;
  assign n9875 = n9722 & ~n9866;
  assign n9876 = ~n9723 & ~n9875;
  assign n9877 = ~n9874 & n9876;
  assign n9878 = ~n9871 & ~n9877;
  assign n9856 = n9676 ^ n9673;
  assign n9857 = n9680 & ~n9856;
  assign n9858 = n9857 ^ n9679;
  assign n9853 = n9665 ^ n9653;
  assign n9854 = ~n9666 & n9853;
  assign n9855 = n9854 ^ n9653;
  assign n9859 = n9858 ^ n9855;
  assign n9849 = n9661 & n9664;
  assign n9850 = n3520 & n8976;
  assign n9851 = ~n9849 & ~n9850;
  assign n9845 = x32 & x52;
  assign n9844 = x31 & x53;
  assign n9846 = n9845 ^ n9844;
  assign n9843 = x26 & x58;
  assign n9847 = n9846 ^ n9843;
  assign n9840 = n9625 ^ n9624;
  assign n9841 = n9627 & ~n9840;
  assign n9842 = n9841 ^ n9626;
  assign n9848 = n9847 ^ n9842;
  assign n9852 = n9851 ^ n9848;
  assign n9860 = n9859 ^ n9852;
  assign n9837 = n9681 ^ n9667;
  assign n9838 = ~n9682 & ~n9837;
  assign n9839 = n9838 ^ n9670;
  assign n9861 = n9860 ^ n9839;
  assign n9829 = n9635 ^ n9634;
  assign n9830 = n9637 & ~n9829;
  assign n9831 = n9830 ^ n9636;
  assign n9826 = n9613 ^ n9612;
  assign n9827 = n9615 & ~n9826;
  assign n9828 = n9827 ^ n9614;
  assign n9832 = n9831 ^ n9828;
  assign n9823 = n9630 ^ n9629;
  assign n9824 = n9632 & ~n9823;
  assign n9825 = n9824 ^ n9631;
  assign n9833 = n9832 ^ n9825;
  assign n9820 = n9698 ^ n9695;
  assign n9821 = n9702 & ~n9820;
  assign n9822 = n9821 ^ n9701;
  assign n9834 = n9833 ^ n9822;
  assign n9817 = n9709 ^ n9706;
  assign n9818 = n9713 & ~n9817;
  assign n9819 = n9818 ^ n9712;
  assign n9835 = n9834 ^ n9819;
  assign n9811 = x41 & x43;
  assign n9810 = x40 & x44;
  assign n9812 = n9811 ^ n9810;
  assign n9809 = x39 & x45;
  assign n9813 = n9812 ^ n9809;
  assign n9806 = x38 & x46;
  assign n9805 = x29 & x55;
  assign n9807 = n9806 ^ n9805;
  assign n9804 = x28 & x56;
  assign n9808 = n9807 ^ n9804;
  assign n9814 = n9813 ^ n9808;
  assign n9801 = x37 & x47;
  assign n9800 = x30 & x54;
  assign n9802 = n9801 ^ n9800;
  assign n9799 = x27 & x57;
  assign n9803 = n9802 ^ n9799;
  assign n9815 = n9814 ^ n9803;
  assign n9794 = x36 & x48;
  assign n9793 = x35 & x49;
  assign n9795 = n9794 ^ n9793;
  assign n9792 = x34 & x50;
  assign n9796 = n9795 ^ n9792;
  assign n9789 = x33 & x51;
  assign n9788 = x25 & x59;
  assign n9790 = n9789 ^ n9788;
  assign n9787 = x24 & x60;
  assign n9791 = n9790 ^ n9787;
  assign n9797 = n9796 ^ n9791;
  assign n9784 = x23 & x61;
  assign n9783 = x22 & x62;
  assign n9785 = n9784 ^ n9783;
  assign n9782 = x21 & x63;
  assign n9786 = n9785 ^ n9782;
  assign n9798 = n9797 ^ n9786;
  assign n9816 = n9815 ^ n9798;
  assign n9836 = n9835 ^ n9816;
  assign n9862 = n9861 ^ n9836;
  assign n9779 = n9718 ^ n9650;
  assign n9780 = n9719 & ~n9779;
  assign n9781 = n9780 ^ n9650;
  assign n9863 = n9862 ^ n9781;
  assign n9774 = n9605 ^ n9602;
  assign n9775 = n9643 & ~n9774;
  assign n9776 = n9775 ^ n9602;
  assign n9771 = n9689 ^ n9686;
  assign n9772 = ~n9717 & n9771;
  assign n9773 = n9772 ^ n9686;
  assign n9777 = n9776 ^ n9773;
  assign n9762 = n9618 ^ n9617;
  assign n9763 = n9620 & ~n9762;
  assign n9764 = n9763 ^ n9619;
  assign n9759 = n9655 ^ n9654;
  assign n9760 = n9657 & ~n9759;
  assign n9761 = n9760 ^ n9656;
  assign n9765 = n9764 ^ n9761;
  assign n9757 = ~x41 & ~n9610;
  assign n9758 = x42 & ~n9757;
  assign n9766 = n9765 ^ n9758;
  assign n9754 = n9616 ^ n9611;
  assign n9755 = n9622 & ~n9754;
  assign n9756 = n9755 ^ n9621;
  assign n9767 = n9766 ^ n9756;
  assign n9751 = n9633 ^ n9628;
  assign n9752 = n9639 & ~n9751;
  assign n9753 = n9752 ^ n9638;
  assign n9768 = n9767 ^ n9753;
  assign n9748 = n9703 ^ n9692;
  assign n9749 = n9715 & ~n9748;
  assign n9750 = n9749 ^ n9714;
  assign n9769 = n9768 ^ n9750;
  assign n9745 = n9640 ^ n9608;
  assign n9746 = ~n9641 & n9745;
  assign n9747 = n9746 ^ n9608;
  assign n9770 = n9769 ^ n9747;
  assign n9778 = n9777 ^ n9770;
  assign n9864 = n9863 ^ n9778;
  assign n9742 = n9720 ^ n9644;
  assign n9743 = n9721 & n9742;
  assign n9744 = n9743 ^ n9647;
  assign n9865 = n9864 ^ n9744;
  assign n9879 = n9878 ^ n9865;
  assign n10000 = n9744 & ~n9864;
  assign n10001 = n9878 & ~n10000;
  assign n10002 = ~n9744 & n9864;
  assign n10003 = ~n10001 & ~n10002;
  assign n9988 = n9761 ^ n9758;
  assign n9989 = n9765 & ~n9988;
  assign n9990 = n9989 ^ n9764;
  assign n9985 = n9828 ^ n9825;
  assign n9986 = n9832 & ~n9985;
  assign n9987 = n9986 ^ n9831;
  assign n9991 = n9990 ^ n9987;
  assign n9982 = n9851 ^ n9842;
  assign n9983 = ~n9848 & ~n9982;
  assign n9984 = n9983 ^ n9851;
  assign n9992 = n9991 ^ n9984;
  assign n9979 = n9855 ^ n9852;
  assign n9980 = n9859 & n9979;
  assign n9981 = n9980 ^ n9858;
  assign n9993 = n9992 ^ n9981;
  assign n9976 = n9835 ^ n9815;
  assign n9977 = ~n9816 & n9976;
  assign n9978 = n9977 ^ n9835;
  assign n9994 = n9993 ^ n9978;
  assign n9973 = n9860 ^ n9836;
  assign n9974 = n9861 & n9973;
  assign n9975 = n9974 ^ n9839;
  assign n9995 = n9994 ^ n9975;
  assign n9970 = n9750 ^ n9747;
  assign n9971 = ~n9769 & n9970;
  assign n9972 = n9971 ^ n9747;
  assign n9996 = n9995 ^ n9972;
  assign n9963 = x24 & x61;
  assign n9960 = n9810 ^ n9809;
  assign n9961 = n9812 & ~n9960;
  assign n9962 = n9961 ^ n9811;
  assign n9964 = n9963 ^ n9962;
  assign n9957 = n9805 ^ n9804;
  assign n9958 = n9807 & ~n9957;
  assign n9959 = n9958 ^ n9806;
  assign n9965 = n9964 ^ n9959;
  assign n9952 = x27 & x58;
  assign n9951 = x26 & x59;
  assign n9953 = n9952 ^ n9951;
  assign n9950 = x25 & x60;
  assign n9954 = n9953 ^ n9950;
  assign n9947 = n9844 ^ n9843;
  assign n9948 = n9846 & ~n9947;
  assign n9949 = n9948 ^ n9845;
  assign n9955 = n9954 ^ n9949;
  assign n9944 = n9800 ^ n9799;
  assign n9945 = n9802 & ~n9944;
  assign n9946 = n9945 ^ n9801;
  assign n9956 = n9955 ^ n9946;
  assign n9966 = n9965 ^ n9956;
  assign n9941 = n9833 ^ n9819;
  assign n9942 = n9834 & ~n9941;
  assign n9943 = n9942 ^ n9822;
  assign n9967 = n9966 ^ n9943;
  assign n9936 = n9791 ^ n9786;
  assign n9937 = n9797 & ~n9936;
  assign n9938 = n9937 ^ n9796;
  assign n9933 = n9808 ^ n9803;
  assign n9934 = n9814 & ~n9933;
  assign n9935 = n9934 ^ n9813;
  assign n9939 = n9938 ^ n9935;
  assign n9928 = n9788 ^ n9787;
  assign n9929 = n9790 & ~n9928;
  assign n9930 = n9929 ^ n9789;
  assign n9925 = n9783 ^ n9782;
  assign n9926 = n9785 & ~n9925;
  assign n9927 = n9926 ^ n9784;
  assign n9931 = n9930 ^ n9927;
  assign n9922 = n9793 ^ n9792;
  assign n9923 = n9795 & ~n9922;
  assign n9924 = n9923 ^ n9794;
  assign n9932 = n9931 ^ n9924;
  assign n9940 = n9939 ^ n9932;
  assign n9968 = n9967 ^ n9940;
  assign n9915 = x31 & x54;
  assign n9916 = n9915 ^ n5354;
  assign n9914 = x30 & x55;
  assign n9917 = n9916 ^ n9914;
  assign n9911 = x38 & x47;
  assign n9910 = x37 & x48;
  assign n9912 = n9911 ^ n9910;
  assign n9909 = x36 & x49;
  assign n9913 = n9912 ^ n9909;
  assign n9918 = n9917 ^ n9913;
  assign n9907 = x23 & x62;
  assign n9906 = ~x42 & x43;
  assign n9908 = n9907 ^ n9906;
  assign n9919 = n9918 ^ n9908;
  assign n9903 = n9766 ^ n9753;
  assign n9904 = n9767 & ~n9903;
  assign n9905 = n9904 ^ n9756;
  assign n9920 = n9919 ^ n9905;
  assign n9898 = x35 & x50;
  assign n9897 = x28 & x57;
  assign n9899 = n9898 ^ n9897;
  assign n9896 = x22 & x63;
  assign n9900 = n9899 ^ n9896;
  assign n9893 = x34 & x51;
  assign n9892 = x33 & x52;
  assign n9894 = n9893 ^ n9892;
  assign n9891 = x32 & x53;
  assign n9895 = n9894 ^ n9891;
  assign n9901 = n9900 ^ n9895;
  assign n9888 = x41 & x44;
  assign n9887 = x40 & x45;
  assign n9889 = n9888 ^ n9887;
  assign n9886 = x39 & x46;
  assign n9890 = n9889 ^ n9886;
  assign n9902 = n9901 ^ n9890;
  assign n9921 = n9920 ^ n9902;
  assign n9969 = n9968 ^ n9921;
  assign n9997 = n9996 ^ n9969;
  assign n9883 = n9773 ^ n9770;
  assign n9884 = n9777 & ~n9883;
  assign n9885 = n9884 ^ n9776;
  assign n9998 = n9997 ^ n9885;
  assign n9880 = n9862 ^ n9778;
  assign n9881 = ~n9863 & ~n9880;
  assign n9882 = n9881 ^ n9781;
  assign n9999 = n9998 ^ n9882;
  assign n10004 = n10003 ^ n9999;
  assign n10118 = n9882 & ~n9885;
  assign n10119 = n9969 & ~n10118;
  assign n10120 = ~n9882 & n9885;
  assign n10121 = ~n10119 & ~n10120;
  assign n10122 = ~n9969 & n10118;
  assign n10123 = n9996 & ~n10122;
  assign n10124 = n10121 & ~n10123;
  assign n10125 = ~n10003 & n10124;
  assign n10126 = n9969 & n10120;
  assign n10127 = ~n10122 & ~n10126;
  assign n10128 = ~n9997 & ~n10127;
  assign n10129 = ~n10125 & ~n10128;
  assign n10130 = ~n9996 & ~n10126;
  assign n10131 = ~n10121 & ~n10130;
  assign n10132 = n10003 & n10131;
  assign n10133 = n10129 & ~n10132;
  assign n10108 = n9897 ^ n9896;
  assign n10109 = n9899 & ~n10108;
  assign n10110 = n10109 ^ n9898;
  assign n10105 = n9951 ^ n9950;
  assign n10106 = n9953 & ~n10105;
  assign n10107 = n10106 ^ n9952;
  assign n10111 = n10110 ^ n10107;
  assign n10102 = n9892 ^ n9891;
  assign n10103 = n9894 & ~n10102;
  assign n10104 = n10103 ^ n9893;
  assign n10112 = n10111 ^ n10104;
  assign n10099 = n9990 ^ n9984;
  assign n10100 = ~n9991 & ~n10099;
  assign n10101 = n10100 ^ n9984;
  assign n10113 = n10112 ^ n10101;
  assign n10094 = n9910 ^ n9909;
  assign n10095 = n9912 & ~n10094;
  assign n10096 = n10095 ^ n9911;
  assign n10091 = n9887 ^ n9886;
  assign n10092 = n9889 & ~n10091;
  assign n10093 = n10092 ^ n9888;
  assign n10097 = n10096 ^ n10093;
  assign n10088 = n9915 ^ n9914;
  assign n10089 = n9916 & ~n10088;
  assign n10090 = n10089 ^ n5354;
  assign n10098 = n10097 ^ n10090;
  assign n10114 = n10113 ^ n10098;
  assign n10080 = x38 & x48;
  assign n10079 = x31 & x55;
  assign n10081 = n10080 ^ n10079;
  assign n10082 = n10081 ^ n5399;
  assign n10076 = x37 & x49;
  assign n10075 = x36 & x50;
  assign n10077 = n10076 ^ n10075;
  assign n10074 = x23 & x63;
  assign n10078 = n10077 ^ n10074;
  assign n10083 = n10082 ^ n10078;
  assign n10071 = x35 & x51;
  assign n10070 = x34 & x52;
  assign n10072 = n10071 ^ n10070;
  assign n10069 = x33 & x53;
  assign n10073 = n10072 ^ n10069;
  assign n10084 = n10083 ^ n10073;
  assign n10064 = x40 & x46;
  assign n10063 = x39 & x47;
  assign n10065 = n10064 ^ n10063;
  assign n10062 = x30 & x56;
  assign n10066 = n10065 ^ n10062;
  assign n10059 = x28 & x58;
  assign n10058 = x27 & x59;
  assign n10060 = n10059 ^ n10058;
  assign n10057 = x26 & x60;
  assign n10061 = n10060 ^ n10057;
  assign n10067 = n10066 ^ n10061;
  assign n10054 = x42 & x44;
  assign n10053 = x41 & x45;
  assign n10055 = n10054 ^ n10053;
  assign n10052 = x32 & x54;
  assign n10056 = n10055 ^ n10052;
  assign n10068 = n10067 ^ n10056;
  assign n10085 = n10084 ^ n10068;
  assign n10049 = n9935 ^ n9932;
  assign n10050 = n9939 & ~n10049;
  assign n10051 = n10050 ^ n9938;
  assign n10086 = n10085 ^ n10051;
  assign n10044 = n9954 ^ n9946;
  assign n10045 = n9955 & ~n10044;
  assign n10046 = n10045 ^ n9949;
  assign n10041 = n9913 ^ n9908;
  assign n10042 = n9918 & ~n10041;
  assign n10043 = n10042 ^ n9917;
  assign n10047 = n10046 ^ n10043;
  assign n10038 = n9895 ^ n9890;
  assign n10039 = n9901 & ~n10038;
  assign n10040 = n10039 ^ n9900;
  assign n10048 = n10047 ^ n10040;
  assign n10087 = n10086 ^ n10048;
  assign n10115 = n10114 ^ n10087;
  assign n10035 = n9994 ^ n9972;
  assign n10036 = n9995 & n10035;
  assign n10037 = n10036 ^ n9975;
  assign n10116 = n10115 ^ n10037;
  assign n10028 = n9965 ^ n9943;
  assign n10029 = ~n9966 & n10028;
  assign n10030 = n10029 ^ n9943;
  assign n10025 = n9919 ^ n9902;
  assign n10026 = n9920 & ~n10025;
  assign n10027 = n10026 ^ n9905;
  assign n10031 = n10030 ^ n10027;
  assign n10020 = ~x42 & ~n9907;
  assign n10021 = x43 & ~n10020;
  assign n10018 = x25 & x61;
  assign n10017 = x24 & x62;
  assign n10019 = n10018 ^ n10017;
  assign n10022 = n10021 ^ n10019;
  assign n10014 = n9927 ^ n9924;
  assign n10015 = n9931 & ~n10014;
  assign n10016 = n10015 ^ n9930;
  assign n10023 = n10022 ^ n10016;
  assign n10011 = n9963 ^ n9959;
  assign n10012 = n9964 & ~n10011;
  assign n10013 = n10012 ^ n9962;
  assign n10024 = n10023 ^ n10013;
  assign n10032 = n10031 ^ n10024;
  assign n10008 = n9992 ^ n9978;
  assign n10009 = ~n9993 & n10008;
  assign n10010 = n10009 ^ n9981;
  assign n10033 = n10032 ^ n10010;
  assign n10005 = n9940 ^ n9921;
  assign n10006 = n9968 & ~n10005;
  assign n10007 = n10006 ^ n9967;
  assign n10034 = n10033 ^ n10007;
  assign n10117 = n10116 ^ n10034;
  assign n10134 = n10133 ^ n10117;
  assign n10266 = ~n10002 & ~n10118;
  assign n10267 = ~n10001 & n10266;
  assign n10268 = ~n10120 & ~n10267;
  assign n10269 = n9969 & n9996;
  assign n10270 = ~n10117 & ~n10269;
  assign n10271 = ~n10268 & ~n10270;
  assign n10272 = ~n10117 & ~n10120;
  assign n10273 = ~n9969 & ~n9996;
  assign n10274 = ~n10272 & ~n10273;
  assign n10275 = n10003 & n10274;
  assign n10276 = ~n10119 & ~n10123;
  assign n10277 = n10117 & ~n10276;
  assign n10278 = ~n10275 & ~n10277;
  assign n10279 = ~n10271 & n10278;
  assign n10256 = n10112 ^ n10098;
  assign n10257 = ~n10113 & ~n10256;
  assign n10258 = n10257 ^ n10101;
  assign n10253 = n10043 ^ n10040;
  assign n10254 = n10047 & ~n10253;
  assign n10255 = n10254 ^ n10046;
  assign n10259 = n10258 ^ n10255;
  assign n10246 = n10058 ^ n10057;
  assign n10247 = n10060 & ~n10246;
  assign n10248 = n10247 ^ n10059;
  assign n10243 = n10075 ^ n10074;
  assign n10244 = n10077 & ~n10243;
  assign n10245 = n10244 ^ n10076;
  assign n10249 = n10248 ^ n10245;
  assign n10240 = n10070 ^ n10069;
  assign n10241 = n10072 & ~n10240;
  assign n10242 = n10241 ^ n10071;
  assign n10250 = n10249 ^ n10242;
  assign n10237 = n10022 ^ n10013;
  assign n10238 = n10023 & ~n10237;
  assign n10239 = n10238 ^ n10016;
  assign n10251 = n10250 ^ n10239;
  assign n10232 = n10080 ^ n5399;
  assign n10233 = ~n10081 & n10232;
  assign n10234 = n10233 ^ n5399;
  assign n10229 = n10063 ^ n10062;
  assign n10230 = n10065 & ~n10229;
  assign n10231 = n10230 ^ n10064;
  assign n10235 = n10234 ^ n10231;
  assign n10226 = n10053 ^ n10052;
  assign n10227 = n10055 & ~n10226;
  assign n10228 = n10227 ^ n10054;
  assign n10236 = n10235 ^ n10228;
  assign n10252 = n10251 ^ n10236;
  assign n10260 = n10259 ^ n10252;
  assign n10223 = n10114 ^ n10086;
  assign n10224 = ~n10087 & ~n10223;
  assign n10225 = n10224 ^ n10114;
  assign n10261 = n10260 ^ n10225;
  assign n10216 = x40 & x47;
  assign n10215 = x33 & x54;
  assign n10217 = n10216 ^ n10215;
  assign n10214 = x31 & x56;
  assign n10218 = n10217 ^ n10214;
  assign n10212 = x25 & x62;
  assign n10211 = ~x43 & x44;
  assign n10213 = n10212 ^ n10211;
  assign n10219 = n10218 ^ n10213;
  assign n10208 = n10107 ^ n10104;
  assign n10209 = n10111 & ~n10208;
  assign n10210 = n10209 ^ n10110;
  assign n10220 = n10219 ^ n10210;
  assign n10203 = x42 & x45;
  assign n10202 = x41 & x46;
  assign n10204 = n10203 ^ n10202;
  assign n10201 = x32 & x55;
  assign n10205 = n10204 ^ n10201;
  assign n10198 = x27 & x60;
  assign n10197 = x26 & x61;
  assign n10199 = n10198 ^ n10197;
  assign n10196 = x24 & x63;
  assign n10200 = n10199 ^ n10196;
  assign n10206 = n10205 ^ n10200;
  assign n10193 = x39 & x48;
  assign n10192 = x38 & x49;
  assign n10194 = n10193 ^ n10192;
  assign n10191 = x37 & x50;
  assign n10195 = n10194 ^ n10191;
  assign n10207 = n10206 ^ n10195;
  assign n10221 = n10220 ^ n10207;
  assign n10180 = ~n6895 & ~n6896;
  assign n10181 = ~x24 & ~n10018;
  assign n10182 = x43 & x62;
  assign n10183 = ~n10181 & n10182;
  assign n10184 = ~n10180 & n10183;
  assign n10185 = n10017 & n10018;
  assign n10186 = x42 & x61;
  assign n10187 = n7304 & n10186;
  assign n10188 = ~n10185 & ~n10187;
  assign n10189 = ~n10184 & n10188;
  assign n10176 = x36 & x51;
  assign n10175 = x35 & x52;
  assign n10177 = n10176 ^ n10175;
  assign n10174 = x29 & x58;
  assign n10178 = n10177 ^ n10174;
  assign n10171 = x34 & x53;
  assign n10170 = x30 & x57;
  assign n10172 = n10171 ^ n10170;
  assign n10169 = x28 & x59;
  assign n10173 = n10172 ^ n10169;
  assign n10179 = n10178 ^ n10173;
  assign n10190 = n10189 ^ n10179;
  assign n10222 = n10221 ^ n10190;
  assign n10262 = n10261 ^ n10222;
  assign n10151 = n10061 ^ n10056;
  assign n10152 = n10067 & ~n10151;
  assign n10153 = n10152 ^ n10066;
  assign n10154 = n10085 & n10153;
  assign n10155 = n10051 & n10154;
  assign n10156 = n10061 & n10066;
  assign n10157 = n10056 & n10156;
  assign n10158 = n10084 & n10157;
  assign n10159 = ~n10155 & ~n10158;
  assign n10160 = ~n10061 & ~n10066;
  assign n10161 = ~n10056 & n10160;
  assign n10162 = ~n10051 & n10161;
  assign n10163 = n10159 & ~n10162;
  assign n10164 = ~n10084 & ~n10153;
  assign n10165 = n10086 & n10164;
  assign n10166 = n10163 & ~n10165;
  assign n10147 = n10093 ^ n10090;
  assign n10148 = n10097 & ~n10147;
  assign n10149 = n10148 ^ n10096;
  assign n10144 = n10078 ^ n10073;
  assign n10145 = n10083 & ~n10144;
  assign n10146 = n10145 ^ n10082;
  assign n10150 = n10149 ^ n10146;
  assign n10167 = n10166 ^ n10150;
  assign n10141 = n10027 ^ n10024;
  assign n10142 = n10031 & ~n10141;
  assign n10143 = n10142 ^ n10030;
  assign n10168 = n10167 ^ n10143;
  assign n10263 = n10262 ^ n10168;
  assign n10138 = n10032 ^ n10007;
  assign n10139 = n10033 & ~n10138;
  assign n10140 = n10139 ^ n10010;
  assign n10264 = n10263 ^ n10140;
  assign n10135 = n10115 ^ n10034;
  assign n10136 = n10116 & n10135;
  assign n10137 = n10136 ^ n10037;
  assign n10265 = n10264 ^ n10137;
  assign n10280 = n10279 ^ n10265;
  assign n10399 = n10137 & n10264;
  assign n10400 = ~n10279 & ~n10399;
  assign n10401 = ~n10137 & ~n10264;
  assign n10402 = ~n10400 & ~n10401;
  assign n10391 = n10255 ^ n10252;
  assign n10392 = ~n10259 & ~n10391;
  assign n10393 = n10392 ^ n10258;
  assign n10388 = n10207 ^ n10190;
  assign n10389 = n10221 & n10388;
  assign n10390 = n10389 ^ n10220;
  assign n10394 = n10393 ^ n10390;
  assign n10383 = n10189 ^ n10178;
  assign n10384 = ~n10179 & ~n10383;
  assign n10385 = n10384 ^ n10189;
  assign n10380 = n10245 ^ n10242;
  assign n10381 = n10249 & ~n10380;
  assign n10382 = n10381 ^ n10248;
  assign n10386 = n10385 ^ n10382;
  assign n10377 = n10200 ^ n10195;
  assign n10378 = n10206 & ~n10377;
  assign n10379 = n10378 ^ n10205;
  assign n10387 = n10386 ^ n10379;
  assign n10395 = n10394 ^ n10387;
  assign n10374 = n10225 ^ n10222;
  assign n10375 = n10261 & ~n10374;
  assign n10376 = n10375 ^ n10260;
  assign n10396 = n10395 ^ n10376;
  assign n10365 = x40 & x48;
  assign n10364 = x32 & x56;
  assign n10366 = n10365 ^ n10364;
  assign n10363 = x30 & x58;
  assign n10367 = n10366 ^ n10363;
  assign n10360 = x39 & x49;
  assign n10359 = x38 & x50;
  assign n10361 = n10360 ^ n10359;
  assign n10362 = n10361 ^ n5966;
  assign n10368 = n10367 ^ n10362;
  assign n10356 = n10231 ^ n10228;
  assign n10357 = n10235 & ~n10356;
  assign n10358 = n10357 ^ n10234;
  assign n10369 = n10368 ^ n10358;
  assign n10346 = ~x43 & ~n10212;
  assign n10347 = x44 & ~n10346;
  assign n10348 = x25 & x63;
  assign n10349 = ~n10347 & ~n10348;
  assign n10350 = x62 & x63;
  assign n10351 = x43 & x63;
  assign n10352 = ~n10350 & ~n10351;
  assign n10353 = n7423 & ~n10352;
  assign n10354 = ~n10349 & ~n10353;
  assign n10343 = n10202 ^ n10201;
  assign n10344 = n10204 & ~n10343;
  assign n10345 = n10344 ^ n10203;
  assign n10355 = n10354 ^ n10345;
  assign n10370 = n10369 ^ n10355;
  assign n10338 = x42 & x46;
  assign n10337 = x41 & x47;
  assign n10339 = n10338 ^ n10337;
  assign n10336 = x31 & x57;
  assign n10340 = n10339 ^ n10336;
  assign n10333 = x28 & x60;
  assign n10332 = x27 & x61;
  assign n10334 = n10333 ^ n10332;
  assign n10331 = x26 & x62;
  assign n10335 = n10334 ^ n10331;
  assign n10341 = n10340 ^ n10335;
  assign n10328 = x37 & x51;
  assign n10327 = x36 & x52;
  assign n10329 = n10328 ^ n10327;
  assign n10326 = x35 & x53;
  assign n10330 = n10329 ^ n10326;
  assign n10342 = n10341 ^ n10330;
  assign n10371 = n10370 ^ n10342;
  assign n10321 = n10150 & ~n10153;
  assign n10322 = n10159 & ~n10321;
  assign n10323 = n10322 ^ n10143;
  assign n10324 = ~n10167 & ~n10323;
  assign n10325 = n10324 ^ n10143;
  assign n10372 = n10371 ^ n10325;
  assign n10316 = n10250 ^ n10236;
  assign n10317 = n10251 & ~n10316;
  assign n10318 = n10317 ^ n10239;
  assign n10313 = n10153 ^ n10149;
  assign n10314 = ~n10150 & n10313;
  assign n10315 = n10314 ^ n10153;
  assign n10319 = n10318 ^ n10315;
  assign n10306 = x43 & x45;
  assign n10305 = x34 & x54;
  assign n10307 = n10306 ^ n10305;
  assign n10304 = x33 & x55;
  assign n10308 = n10307 ^ n10304;
  assign n10301 = n10215 ^ n10214;
  assign n10302 = n10217 & ~n10301;
  assign n10303 = n10302 ^ n10216;
  assign n10309 = n10308 ^ n10303;
  assign n10298 = n10175 ^ n10174;
  assign n10299 = n10177 & ~n10298;
  assign n10300 = n10299 ^ n10176;
  assign n10310 = n10309 ^ n10300;
  assign n10295 = n10218 ^ n10210;
  assign n10296 = ~n10219 & n10295;
  assign n10297 = n10296 ^ n10210;
  assign n10311 = n10310 ^ n10297;
  assign n10290 = n10197 ^ n10196;
  assign n10291 = n10199 & ~n10290;
  assign n10292 = n10291 ^ n10198;
  assign n10287 = n10192 ^ n10191;
  assign n10288 = n10194 & ~n10287;
  assign n10289 = n10288 ^ n10193;
  assign n10293 = n10292 ^ n10289;
  assign n10284 = n10170 ^ n10169;
  assign n10285 = n10172 & ~n10284;
  assign n10286 = n10285 ^ n10171;
  assign n10294 = n10293 ^ n10286;
  assign n10312 = n10311 ^ n10294;
  assign n10320 = n10319 ^ n10312;
  assign n10373 = n10372 ^ n10320;
  assign n10397 = n10396 ^ n10373;
  assign n10281 = n10262 ^ n10140;
  assign n10282 = n10263 & ~n10281;
  assign n10283 = n10282 ^ n10140;
  assign n10398 = n10397 ^ n10283;
  assign n10403 = n10402 ^ n10398;
  assign n10512 = n10283 & ~n10397;
  assign n10513 = ~n10401 & ~n10512;
  assign n10514 = ~n10400 & n10513;
  assign n10515 = ~n10283 & n10397;
  assign n10516 = ~n10514 & ~n10515;
  assign n10501 = n10345 & n10354;
  assign n10502 = n10501 ^ n10353;
  assign n10498 = n10308 ^ n10300;
  assign n10499 = n10309 & ~n10498;
  assign n10500 = n10499 ^ n10303;
  assign n10503 = n10502 ^ n10500;
  assign n10495 = n10289 ^ n10286;
  assign n10496 = n10293 & ~n10495;
  assign n10497 = n10496 ^ n10292;
  assign n10504 = n10503 ^ n10497;
  assign n10492 = n10382 ^ n10379;
  assign n10493 = ~n10386 & ~n10492;
  assign n10494 = n10493 ^ n10385;
  assign n10505 = n10504 ^ n10494;
  assign n10489 = n10310 ^ n10294;
  assign n10490 = n10311 & ~n10489;
  assign n10491 = n10490 ^ n10297;
  assign n10506 = n10505 ^ n10491;
  assign n10486 = n10390 ^ n10387;
  assign n10487 = ~n10394 & n10486;
  assign n10488 = n10487 ^ n10393;
  assign n10507 = n10506 ^ n10488;
  assign n10479 = x28 & x61;
  assign n10478 = x29 & x60;
  assign n10480 = n10479 ^ n10478;
  assign n10475 = n10305 ^ n10304;
  assign n10476 = n10307 & ~n10475;
  assign n10477 = n10476 ^ n10306;
  assign n10481 = n10480 ^ n10477;
  assign n10472 = x43 & x46;
  assign n10471 = x42 & x47;
  assign n10473 = n10472 ^ n10471;
  assign n10470 = x34 & x55;
  assign n10474 = n10473 ^ n10470;
  assign n10482 = n10481 ^ n10474;
  assign n10468 = x27 & x62;
  assign n10467 = ~x44 & x45;
  assign n10469 = n10468 ^ n10467;
  assign n10483 = n10482 ^ n10469;
  assign n10462 = x32 & x57;
  assign n10461 = x31 & x58;
  assign n10463 = n10462 ^ n10461;
  assign n10460 = x30 & x59;
  assign n10464 = n10463 ^ n10460;
  assign n10457 = x38 & x51;
  assign n10456 = x37 & x52;
  assign n10458 = n10457 ^ n10456;
  assign n10455 = x36 & x53;
  assign n10459 = n10458 ^ n10455;
  assign n10465 = n10464 ^ n10459;
  assign n10452 = x41 & x48;
  assign n10451 = x35 & x54;
  assign n10453 = n10452 ^ n10451;
  assign n10450 = x33 & x56;
  assign n10454 = n10453 ^ n10450;
  assign n10466 = n10465 ^ n10454;
  assign n10484 = n10483 ^ n10466;
  assign n10445 = n10364 ^ n10363;
  assign n10446 = n10366 & ~n10445;
  assign n10447 = n10446 ^ n10365;
  assign n10442 = n10327 ^ n10326;
  assign n10443 = n10329 & ~n10442;
  assign n10444 = n10443 ^ n10328;
  assign n10448 = n10447 ^ n10444;
  assign n10439 = n10332 ^ n10331;
  assign n10440 = n10334 & ~n10439;
  assign n10441 = n10440 ^ n10333;
  assign n10449 = n10448 ^ n10441;
  assign n10485 = n10484 ^ n10449;
  assign n10508 = n10507 ^ n10485;
  assign n10434 = n10315 ^ n10312;
  assign n10435 = n10319 & ~n10434;
  assign n10436 = n10435 ^ n10318;
  assign n10431 = n10355 ^ n10342;
  assign n10432 = n10370 & ~n10431;
  assign n10433 = n10432 ^ n10369;
  assign n10437 = n10436 ^ n10433;
  assign n10424 = x40 & x49;
  assign n10423 = x39 & x50;
  assign n10425 = n10424 ^ n10423;
  assign n10422 = x26 & x63;
  assign n10426 = n10425 ^ n10422;
  assign n10419 = n10360 ^ n5966;
  assign n10420 = ~n10361 & n10419;
  assign n10421 = n10420 ^ n5966;
  assign n10427 = n10426 ^ n10421;
  assign n10416 = n10337 ^ n10336;
  assign n10417 = n10339 & ~n10416;
  assign n10418 = n10417 ^ n10338;
  assign n10428 = n10427 ^ n10418;
  assign n10413 = n10367 ^ n10358;
  assign n10414 = ~n10368 & n10413;
  assign n10415 = n10414 ^ n10358;
  assign n10429 = n10428 ^ n10415;
  assign n10410 = n10335 ^ n10330;
  assign n10411 = n10341 & ~n10410;
  assign n10412 = n10411 ^ n10340;
  assign n10430 = n10429 ^ n10412;
  assign n10438 = n10437 ^ n10430;
  assign n10509 = n10508 ^ n10438;
  assign n10407 = n10371 ^ n10320;
  assign n10408 = n10372 & ~n10407;
  assign n10409 = n10408 ^ n10325;
  assign n10510 = n10509 ^ n10409;
  assign n10404 = n10376 ^ n10373;
  assign n10405 = ~n10396 & n10404;
  assign n10406 = n10405 ^ n10395;
  assign n10511 = n10510 ^ n10406;
  assign n10517 = n10516 ^ n10511;
  assign n10615 = n10477 & n10480;
  assign n10616 = n5240 & n7409;
  assign n10617 = ~n10615 & ~n10616;
  assign n10611 = x32 & x58;
  assign n10612 = n10611 ^ n6109;
  assign n10610 = x30 & x60;
  assign n10613 = n10612 ^ n10610;
  assign n10607 = x29 & x61;
  assign n10606 = x28 & x62;
  assign n10608 = n10607 ^ n10606;
  assign n10605 = x27 & x63;
  assign n10609 = n10608 ^ n10605;
  assign n10614 = n10613 ^ n10609;
  assign n10618 = n10617 ^ n10614;
  assign n10602 = n10428 ^ n10412;
  assign n10603 = n10429 & ~n10602;
  assign n10604 = n10603 ^ n10415;
  assign n10619 = n10618 ^ n10604;
  assign n10597 = x41 & x49;
  assign n10596 = x40 & x50;
  assign n10598 = n10597 ^ n10596;
  assign n10595 = x39 & x51;
  assign n10599 = n10598 ^ n10595;
  assign n10592 = n10426 ^ n10418;
  assign n10593 = n10427 & ~n10592;
  assign n10594 = n10593 ^ n10421;
  assign n10600 = n10599 ^ n10594;
  assign n10589 = n10444 ^ n10441;
  assign n10590 = n10448 & ~n10589;
  assign n10591 = n10590 ^ n10447;
  assign n10601 = n10600 ^ n10591;
  assign n10620 = n10619 ^ n10601;
  assign n10586 = n10433 ^ n10430;
  assign n10587 = n10437 & ~n10586;
  assign n10588 = n10587 ^ n10436;
  assign n10621 = n10620 ^ n10588;
  assign n10579 = n10461 ^ n10460;
  assign n10580 = n10463 & ~n10579;
  assign n10581 = n10580 ^ n10462;
  assign n10576 = n10423 ^ n10422;
  assign n10577 = n10425 & ~n10576;
  assign n10578 = n10577 ^ n10424;
  assign n10582 = n10581 ^ n10578;
  assign n10573 = n10456 ^ n10455;
  assign n10574 = n10458 & ~n10573;
  assign n10575 = n10574 ^ n10457;
  assign n10583 = n10582 ^ n10575;
  assign n10568 = x35 & x55;
  assign n10567 = x34 & x56;
  assign n10569 = n10568 ^ n10567;
  assign n10566 = x33 & x57;
  assign n10570 = n10569 ^ n10566;
  assign n10563 = x38 & x52;
  assign n10562 = x37 & x53;
  assign n10564 = n10563 ^ n10562;
  assign n10561 = x36 & x54;
  assign n10565 = n10564 ^ n10561;
  assign n10571 = n10570 ^ n10565;
  assign n10558 = x44 & x46;
  assign n10557 = x43 & x47;
  assign n10559 = n10558 ^ n10557;
  assign n10556 = x42 & x48;
  assign n10560 = n10559 ^ n10556;
  assign n10572 = n10571 ^ n10560;
  assign n10584 = n10583 ^ n10572;
  assign n10553 = n10502 ^ n10497;
  assign n10554 = n10503 & ~n10553;
  assign n10555 = n10554 ^ n10500;
  assign n10585 = n10584 ^ n10555;
  assign n10622 = n10621 ^ n10585;
  assign n10550 = n10506 ^ n10485;
  assign n10551 = n10507 & n10550;
  assign n10552 = n10551 ^ n10488;
  assign n10623 = n10622 ^ n10552;
  assign n10541 = n10471 ^ n10470;
  assign n10542 = n10473 & ~n10541;
  assign n10543 = n10542 ^ n10472;
  assign n10538 = n10451 ^ n10450;
  assign n10539 = n10453 & ~n10538;
  assign n10540 = n10539 ^ n10452;
  assign n10544 = n10543 ^ n10540;
  assign n10536 = ~x44 & ~n10468;
  assign n10537 = x45 & ~n10536;
  assign n10545 = n10544 ^ n10537;
  assign n10533 = n10474 ^ n10469;
  assign n10534 = n10482 & ~n10533;
  assign n10535 = n10534 ^ n10481;
  assign n10546 = n10545 ^ n10535;
  assign n10530 = n10459 ^ n10454;
  assign n10531 = n10465 & ~n10530;
  assign n10532 = n10531 ^ n10464;
  assign n10547 = n10546 ^ n10532;
  assign n10527 = n10466 ^ n10449;
  assign n10528 = n10484 & ~n10527;
  assign n10529 = n10528 ^ n10483;
  assign n10548 = n10547 ^ n10529;
  assign n10524 = n10494 ^ n10491;
  assign n10525 = n10505 & ~n10524;
  assign n10526 = n10525 ^ n10491;
  assign n10549 = n10548 ^ n10526;
  assign n10624 = n10623 ^ n10549;
  assign n10521 = n10438 ^ n10409;
  assign n10522 = n10509 & ~n10521;
  assign n10523 = n10522 ^ n10508;
  assign n10625 = n10624 ^ n10523;
  assign n10518 = n10516 ^ n10510;
  assign n10519 = ~n10511 & n10518;
  assign n10520 = n10519 ^ n10516;
  assign n10626 = n10625 ^ n10520;
  assign n10719 = x44 & x47;
  assign n10718 = x43 & x48;
  assign n10720 = n10719 ^ n10718;
  assign n10717 = x35 & x56;
  assign n10721 = n10720 ^ n10717;
  assign n10714 = x41 & x50;
  assign n10713 = x40 & x51;
  assign n10715 = n10714 ^ n10713;
  assign n10712 = x28 & x63;
  assign n10716 = n10715 ^ n10712;
  assign n10722 = n10721 ^ n10716;
  assign n10710 = x29 & x62;
  assign n10709 = ~x45 & x46;
  assign n10711 = n10710 ^ n10709;
  assign n10723 = n10722 ^ n10711;
  assign n10706 = n10599 ^ n10591;
  assign n10707 = n10600 & ~n10706;
  assign n10708 = n10707 ^ n10594;
  assign n10724 = n10723 ^ n10708;
  assign n10701 = n10611 ^ n10610;
  assign n10702 = n10612 & ~n10701;
  assign n10703 = n10702 ^ n6109;
  assign n10698 = n10562 ^ n10561;
  assign n10699 = n10564 & ~n10698;
  assign n10700 = n10699 ^ n10563;
  assign n10704 = n10703 ^ n10700;
  assign n10695 = n10606 ^ n10605;
  assign n10696 = n10608 & ~n10695;
  assign n10697 = n10696 ^ n10607;
  assign n10705 = n10704 ^ n10697;
  assign n10725 = n10724 ^ n10705;
  assign n10692 = n10529 ^ n10526;
  assign n10693 = ~n10548 & n10692;
  assign n10694 = n10693 ^ n10526;
  assign n10726 = n10725 ^ n10694;
  assign n10685 = x42 & x49;
  assign n10684 = x36 & x55;
  assign n10686 = n10685 ^ n10684;
  assign n10683 = x34 & x57;
  assign n10687 = n10686 ^ n10683;
  assign n10680 = n10540 ^ n10537;
  assign n10681 = n10544 & ~n10680;
  assign n10682 = n10681 ^ n10543;
  assign n10688 = n10687 ^ n10682;
  assign n10677 = n10578 ^ n10575;
  assign n10678 = n10582 & ~n10677;
  assign n10679 = n10678 ^ n10581;
  assign n10689 = n10688 ^ n10679;
  assign n10674 = n10545 ^ n10532;
  assign n10675 = n10546 & ~n10674;
  assign n10676 = n10675 ^ n10535;
  assign n10690 = n10689 ^ n10676;
  assign n10669 = x33 & x58;
  assign n10668 = x32 & x59;
  assign n10670 = n10669 ^ n10668;
  assign n10671 = n10670 ^ n6112;
  assign n10665 = x39 & x52;
  assign n10664 = x38 & x53;
  assign n10666 = n10665 ^ n10664;
  assign n10663 = x37 & x54;
  assign n10667 = n10666 ^ n10663;
  assign n10672 = n10671 ^ n10667;
  assign n10660 = n10596 ^ n10595;
  assign n10661 = n10598 & ~n10660;
  assign n10662 = n10661 ^ n10597;
  assign n10673 = n10672 ^ n10662;
  assign n10691 = n10690 ^ n10673;
  assign n10727 = n10726 ^ n10691;
  assign n10651 = n10557 ^ n10556;
  assign n10652 = n10559 & ~n10651;
  assign n10653 = n10652 ^ n10558;
  assign n10648 = n10567 ^ n10566;
  assign n10649 = n10569 & ~n10648;
  assign n10650 = n10649 ^ n10568;
  assign n10654 = n10653 ^ n10650;
  assign n10655 = n10654 ^ n6256;
  assign n10645 = n10565 ^ n10560;
  assign n10646 = n10571 & ~n10645;
  assign n10647 = n10646 ^ n10570;
  assign n10656 = n10655 ^ n10647;
  assign n10642 = n10617 ^ n10613;
  assign n10643 = ~n10614 & ~n10642;
  assign n10644 = n10643 ^ n10617;
  assign n10657 = n10656 ^ n10644;
  assign n10639 = n10618 ^ n10601;
  assign n10640 = ~n10619 & n10639;
  assign n10641 = n10640 ^ n10604;
  assign n10658 = n10657 ^ n10641;
  assign n10636 = n10583 ^ n10555;
  assign n10637 = ~n10584 & n10636;
  assign n10638 = n10637 ^ n10555;
  assign n10659 = n10658 ^ n10638;
  assign n10728 = n10727 ^ n10659;
  assign n10633 = n10620 ^ n10585;
  assign n10634 = ~n10621 & n10633;
  assign n10635 = n10634 ^ n10588;
  assign n10729 = n10728 ^ n10635;
  assign n10630 = n10622 ^ n10549;
  assign n10631 = n10623 & n10630;
  assign n10632 = n10631 ^ n10552;
  assign n10730 = n10729 ^ n10632;
  assign n10627 = n10523 ^ n10520;
  assign n10628 = ~n10625 & n10627;
  assign n10629 = n10628 ^ n10520;
  assign n10731 = n10730 ^ n10629;
  assign n10834 = ~n10659 & n10727;
  assign n10835 = n10659 & ~n10727;
  assign n10836 = n10635 & ~n10835;
  assign n10837 = ~n10632 & n10836;
  assign n10838 = ~n10834 & ~n10837;
  assign n10839 = n10632 & ~n10635;
  assign n10840 = ~n10838 & ~n10839;
  assign n10828 = n10635 ^ n10632;
  assign n10829 = n10659 ^ n10635;
  assign n10830 = n10828 & n10829;
  assign n10831 = ~n10730 & n10830;
  assign n10832 = n10831 ^ n10730;
  assign n10833 = ~n10629 & n10832;
  assign n10841 = n10840 ^ n10833;
  assign n10842 = n10728 & n10830;
  assign n10843 = ~n10841 & ~n10842;
  assign n10821 = n10657 ^ n10638;
  assign n10822 = ~n10658 & n10821;
  assign n10823 = n10822 ^ n10641;
  assign n10818 = n10689 ^ n10673;
  assign n10819 = n10690 & ~n10818;
  assign n10820 = n10819 ^ n10676;
  assign n10824 = n10823 ^ n10820;
  assign n10811 = ~x45 & ~n10710;
  assign n10812 = x46 & ~n10811;
  assign n10809 = x31 & x61;
  assign n10808 = x30 & x62;
  assign n10810 = n10809 ^ n10808;
  assign n10813 = n10812 ^ n10810;
  assign n10805 = x41 & x51;
  assign n10804 = x40 & x52;
  assign n10806 = n10805 ^ n10804;
  assign n10803 = x39 & x53;
  assign n10807 = n10806 ^ n10803;
  assign n10814 = n10813 ^ n10807;
  assign n10800 = n10653 ^ n6256;
  assign n10801 = ~n10654 & n10800;
  assign n10802 = n10801 ^ n6256;
  assign n10815 = n10814 ^ n10802;
  assign n10795 = x42 & x50;
  assign n10794 = x35 & x57;
  assign n10796 = n10795 ^ n10794;
  assign n10793 = x34 & x58;
  assign n10797 = n10796 ^ n10793;
  assign n10790 = x45 & x47;
  assign n10789 = x44 & x48;
  assign n10791 = n10790 ^ n10789;
  assign n10788 = x43 & x49;
  assign n10792 = n10791 ^ n10788;
  assign n10798 = n10797 ^ n10792;
  assign n10785 = x36 & x56;
  assign n10784 = x33 & x59;
  assign n10786 = n10785 ^ n10784;
  assign n10783 = x29 & x63;
  assign n10787 = n10786 ^ n10783;
  assign n10799 = n10798 ^ n10787;
  assign n10816 = n10815 ^ n10799;
  assign n10780 = n10647 ^ n10644;
  assign n10781 = ~n10656 & ~n10780;
  assign n10782 = n10781 ^ n10644;
  assign n10817 = n10816 ^ n10782;
  assign n10825 = n10824 ^ n10817;
  assign n10777 = n10725 ^ n10691;
  assign n10778 = n10726 & ~n10777;
  assign n10779 = n10778 ^ n10694;
  assign n10826 = n10825 ^ n10779;
  assign n10768 = n10664 ^ n10663;
  assign n10769 = n10666 & ~n10768;
  assign n10770 = n10769 ^ n10665;
  assign n10765 = n10713 ^ n10712;
  assign n10766 = n10715 & ~n10765;
  assign n10767 = n10766 ^ n10714;
  assign n10771 = n10770 ^ n10767;
  assign n10762 = n10669 ^ n6112;
  assign n10763 = ~n10670 & n10762;
  assign n10764 = n10763 ^ n6112;
  assign n10772 = n10771 ^ n10764;
  assign n10759 = n10687 ^ n10679;
  assign n10760 = n10688 & ~n10759;
  assign n10761 = n10760 ^ n10682;
  assign n10773 = n10772 ^ n10761;
  assign n10754 = x38 & x54;
  assign n10753 = x37 & x55;
  assign n10755 = n10754 ^ n10753;
  assign n10752 = x32 & x60;
  assign n10756 = n10755 ^ n10752;
  assign n10749 = n10718 ^ n10717;
  assign n10750 = n10720 & ~n10749;
  assign n10751 = n10750 ^ n10719;
  assign n10757 = n10756 ^ n10751;
  assign n10746 = n10684 ^ n10683;
  assign n10747 = n10686 & ~n10746;
  assign n10748 = n10747 ^ n10685;
  assign n10758 = n10757 ^ n10748;
  assign n10774 = n10773 ^ n10758;
  assign n10741 = n10716 ^ n10711;
  assign n10742 = n10722 & ~n10741;
  assign n10743 = n10742 ^ n10721;
  assign n10738 = n10671 ^ n10662;
  assign n10739 = ~n10672 & n10738;
  assign n10740 = n10739 ^ n10662;
  assign n10744 = n10743 ^ n10740;
  assign n10735 = n10700 ^ n10697;
  assign n10736 = n10704 & ~n10735;
  assign n10737 = n10736 ^ n10703;
  assign n10745 = n10744 ^ n10737;
  assign n10775 = n10774 ^ n10745;
  assign n10732 = n10723 ^ n10705;
  assign n10733 = n10724 & ~n10732;
  assign n10734 = n10733 ^ n10708;
  assign n10776 = n10775 ^ n10734;
  assign n10827 = n10826 ^ n10776;
  assign n10844 = n10843 ^ n10827;
  assign n10947 = n10629 & ~n10839;
  assign n10948 = ~n10632 & n10635;
  assign n10949 = ~n10827 & ~n10835;
  assign n10950 = ~n10948 & ~n10949;
  assign n10951 = ~n10947 & n10950;
  assign n10952 = ~n10827 & ~n10839;
  assign n10953 = ~n10834 & ~n10952;
  assign n10954 = ~n10629 & n10953;
  assign n10955 = n10827 & n10838;
  assign n10956 = ~n10954 & ~n10955;
  assign n10957 = ~n10951 & n10956;
  assign n10935 = n10794 ^ n10793;
  assign n10936 = n10796 & ~n10935;
  assign n10937 = n10936 ^ n10795;
  assign n10932 = n10789 ^ n10788;
  assign n10933 = n10791 & ~n10932;
  assign n10934 = n10933 ^ n10790;
  assign n10938 = n10937 ^ n10934;
  assign n10929 = n10804 ^ n10803;
  assign n10930 = n10806 & ~n10929;
  assign n10931 = n10930 ^ n10805;
  assign n10939 = n10938 ^ n10931;
  assign n10926 = n10813 ^ n10802;
  assign n10927 = ~n10814 & n10926;
  assign n10928 = n10927 ^ n10802;
  assign n10940 = n10939 ^ n10928;
  assign n10921 = n10784 ^ n10783;
  assign n10922 = n10786 & ~n10921;
  assign n10923 = n10922 ^ n10785;
  assign n10918 = n10753 ^ n10752;
  assign n10919 = n10755 & ~n10918;
  assign n10920 = n10919 ^ n10754;
  assign n10924 = n10923 ^ n10920;
  assign n10909 = x45 & x46;
  assign n10910 = ~n10808 & ~n10909;
  assign n10911 = n10809 & ~n10910;
  assign n10912 = ~x29 & ~n8448;
  assign n10913 = x46 & x62;
  assign n10914 = ~n10912 & n10913;
  assign n10915 = ~n10911 & ~n10914;
  assign n10916 = ~x30 & ~n10809;
  assign n10917 = ~n10915 & ~n10916;
  assign n10925 = n10924 ^ n10917;
  assign n10941 = n10940 ^ n10925;
  assign n10904 = n10767 ^ n10764;
  assign n10905 = n10771 & ~n10904;
  assign n10906 = n10905 ^ n10770;
  assign n10901 = n10792 ^ n10787;
  assign n10902 = n10798 & ~n10901;
  assign n10903 = n10902 ^ n10797;
  assign n10907 = n10906 ^ n10903;
  assign n10898 = n10756 ^ n10748;
  assign n10899 = n10757 & ~n10898;
  assign n10900 = n10899 ^ n10751;
  assign n10908 = n10907 ^ n10900;
  assign n10942 = n10941 ^ n10908;
  assign n10895 = n10772 ^ n10758;
  assign n10896 = n10773 & ~n10895;
  assign n10897 = n10896 ^ n10761;
  assign n10943 = n10942 ^ n10897;
  assign n10892 = n10820 ^ n10817;
  assign n10893 = n10824 & n10892;
  assign n10894 = n10893 ^ n10823;
  assign n10944 = n10943 ^ n10894;
  assign n10883 = x45 & x48;
  assign n10882 = x38 & x55;
  assign n10884 = n10883 ^ n10882;
  assign n10881 = x37 & x56;
  assign n10885 = n10884 ^ n10881;
  assign n10878 = x44 & x49;
  assign n10877 = x43 & x50;
  assign n10879 = n10878 ^ n10877;
  assign n10876 = x42 & x51;
  assign n10880 = n10879 ^ n10876;
  assign n10886 = n10885 ^ n10880;
  assign n10874 = x31 & x62;
  assign n10873 = ~x46 & x47;
  assign n10875 = n10874 ^ n10873;
  assign n10887 = n10886 ^ n10875;
  assign n10868 = x39 & x54;
  assign n10867 = x36 & x57;
  assign n10869 = n10868 ^ n10867;
  assign n10866 = x35 & x58;
  assign n10870 = n10869 ^ n10866;
  assign n10863 = x33 & x60;
  assign n10864 = n10863 ^ n6514;
  assign n10862 = x30 & x63;
  assign n10865 = n10864 ^ n10862;
  assign n10871 = n10870 ^ n10865;
  assign n10859 = x41 & x52;
  assign n10858 = x40 & x53;
  assign n10860 = n10859 ^ n10858;
  assign n10857 = x34 & x59;
  assign n10861 = n10860 ^ n10857;
  assign n10872 = n10871 ^ n10861;
  assign n10888 = n10887 ^ n10872;
  assign n10854 = n10743 ^ n10737;
  assign n10855 = ~n10744 & n10854;
  assign n10856 = n10855 ^ n10737;
  assign n10889 = n10888 ^ n10856;
  assign n10851 = n10815 ^ n10782;
  assign n10852 = ~n10816 & ~n10851;
  assign n10853 = n10852 ^ n10782;
  assign n10890 = n10889 ^ n10853;
  assign n10848 = n10774 ^ n10734;
  assign n10849 = ~n10775 & n10848;
  assign n10850 = n10849 ^ n10734;
  assign n10891 = n10890 ^ n10850;
  assign n10945 = n10944 ^ n10891;
  assign n10845 = n10825 ^ n10776;
  assign n10846 = ~n10826 & n10845;
  assign n10847 = n10846 ^ n10779;
  assign n10946 = n10945 ^ n10847;
  assign n10958 = n10957 ^ n10946;
  assign n11035 = ~n10850 & n10853;
  assign n11045 = n10920 ^ n10917;
  assign n11046 = n10924 & ~n11045;
  assign n11047 = n11046 ^ n10923;
  assign n11042 = n10865 ^ n10861;
  assign n11043 = n10871 & ~n11042;
  assign n11044 = n11043 ^ n10870;
  assign n11048 = n11047 ^ n11044;
  assign n11039 = n10934 ^ n10931;
  assign n11040 = n10938 & ~n11039;
  assign n11041 = n11040 ^ n10937;
  assign n11049 = n11048 ^ n11041;
  assign n11036 = n10939 ^ n10925;
  assign n11037 = n10940 & ~n11036;
  assign n11038 = n11037 ^ n10928;
  assign n11050 = n11049 ^ n11038;
  assign n11051 = n10872 & n10887;
  assign n11052 = ~n11050 & ~n11051;
  assign n11053 = ~n11035 & ~n11052;
  assign n11054 = ~n10872 & ~n10887;
  assign n11055 = ~n11050 & ~n11054;
  assign n11056 = ~n10856 & ~n11051;
  assign n11057 = n11055 & ~n11056;
  assign n11058 = n11050 & n11054;
  assign n11059 = ~n11057 & ~n11058;
  assign n11060 = n11059 ^ n10888;
  assign n11061 = n10856 & ~n11060;
  assign n11062 = n11061 ^ n10888;
  assign n11063 = n11053 & n11062;
  assign n11064 = n10850 & ~n10853;
  assign n11065 = ~n11059 & n11064;
  assign n11066 = ~n11063 & ~n11065;
  assign n11067 = ~n10889 & ~n11055;
  assign n11068 = n11050 & n11056;
  assign n11069 = n11067 & ~n11068;
  assign n11070 = ~n11064 & n11069;
  assign n11071 = n11050 & ~n11051;
  assign n11072 = ~n11057 & ~n11071;
  assign n11073 = n11035 & n11072;
  assign n11074 = ~n11070 & ~n11073;
  assign n11075 = n11066 & n11074;
  assign n11026 = x44 & x50;
  assign n11025 = x43 & x51;
  assign n11027 = n11026 ^ n11025;
  assign n11024 = x36 & x58;
  assign n11028 = n11027 ^ n11024;
  assign n11021 = x42 & x52;
  assign n11020 = x41 & x53;
  assign n11022 = n11021 ^ n11020;
  assign n11019 = x40 & x54;
  assign n11023 = n11022 ^ n11019;
  assign n11029 = n11028 ^ n11023;
  assign n11016 = x46 & x48;
  assign n11015 = x45 & x49;
  assign n11017 = n11016 ^ n11015;
  assign n11014 = x38 & x56;
  assign n11018 = n11017 ^ n11014;
  assign n11030 = n11029 ^ n11018;
  assign n11011 = n10903 ^ n10900;
  assign n11012 = n10907 & ~n11011;
  assign n11013 = n11012 ^ n10906;
  assign n11031 = n11030 ^ n11013;
  assign n11006 = x39 & x55;
  assign n11005 = x37 & x57;
  assign n11007 = n11006 ^ n11005;
  assign n11004 = x34 & x60;
  assign n11008 = n11007 ^ n11004;
  assign n11001 = n10877 ^ n10876;
  assign n11002 = n10879 & ~n11001;
  assign n11003 = n11002 ^ n10878;
  assign n11009 = n11008 ^ n11003;
  assign n10998 = x35 & x59;
  assign n10999 = n10998 ^ n6590;
  assign n10997 = x33 & x61;
  assign n11000 = n10999 ^ n10997;
  assign n11010 = n11009 ^ n11000;
  assign n11032 = n11031 ^ n11010;
  assign n10985 = x47 & x62;
  assign n10986 = ~x63 & ~n10985;
  assign n10987 = x31 & ~n10986;
  assign n10988 = x46 & x47;
  assign n10989 = ~n10987 & ~n10988;
  assign n10990 = x46 & x63;
  assign n10991 = ~n10350 & ~n10990;
  assign n10992 = n8894 & ~n10991;
  assign n10993 = ~n10989 & ~n10992;
  assign n10982 = n10882 ^ n10881;
  assign n10983 = n10884 & ~n10982;
  assign n10984 = n10983 ^ n10883;
  assign n10994 = n10993 ^ n10984;
  assign n10979 = n10880 ^ n10875;
  assign n10980 = n10886 & ~n10979;
  assign n10981 = n10980 ^ n10885;
  assign n10995 = n10994 ^ n10981;
  assign n10974 = n10863 ^ n10862;
  assign n10975 = n10864 & ~n10974;
  assign n10976 = n10975 ^ n6514;
  assign n10971 = n10867 ^ n10866;
  assign n10972 = n10869 & ~n10971;
  assign n10973 = n10972 ^ n10868;
  assign n10977 = n10976 ^ n10973;
  assign n10968 = n10858 ^ n10857;
  assign n10969 = n10860 & ~n10968;
  assign n10970 = n10969 ^ n10859;
  assign n10978 = n10977 ^ n10970;
  assign n10996 = n10995 ^ n10978;
  assign n11033 = n11032 ^ n10996;
  assign n10965 = n10941 ^ n10897;
  assign n10966 = ~n10942 & n10965;
  assign n10967 = n10966 ^ n10897;
  assign n11034 = n11033 ^ n10967;
  assign n11076 = n11075 ^ n11034;
  assign n10962 = n10943 ^ n10891;
  assign n10963 = n10944 & n10962;
  assign n10964 = n10963 ^ n10894;
  assign n11077 = n11076 ^ n10964;
  assign n10959 = n10957 ^ n10945;
  assign n10960 = n10946 & ~n10959;
  assign n10961 = n10960 ^ n10957;
  assign n11078 = n11077 ^ n10961;
  assign n11079 = ~n10961 & ~n10964;
  assign n11158 = n11056 ^ n11049;
  assign n11159 = n11050 & n11158;
  assign n11160 = n11159 ^ n11038;
  assign n11161 = ~n11058 & n11160;
  assign n11151 = x44 & x51;
  assign n11150 = x43 & x52;
  assign n11152 = n11151 ^ n11150;
  assign n11149 = x42 & x53;
  assign n11153 = n11152 ^ n11149;
  assign n11146 = x46 & x49;
  assign n11145 = x45 & x50;
  assign n11147 = n11146 ^ n11145;
  assign n11144 = x39 & x56;
  assign n11148 = n11147 ^ n11144;
  assign n11154 = n11153 ^ n11148;
  assign n11142 = x33 & x62;
  assign n11141 = ~x47 & x48;
  assign n11143 = n11142 ^ n11141;
  assign n11155 = n11154 ^ n11143;
  assign n11138 = n11044 ^ n11041;
  assign n11139 = n11048 & ~n11138;
  assign n11140 = n11139 ^ n11047;
  assign n11156 = n11155 ^ n11140;
  assign n11133 = x41 & x54;
  assign n11132 = x34 & x61;
  assign n11134 = n11133 ^ n11132;
  assign n11135 = n11134 ^ n6521;
  assign n11129 = x40 & x55;
  assign n11128 = x38 & x57;
  assign n11130 = n11129 ^ n11128;
  assign n11127 = x37 & x58;
  assign n11131 = n11130 ^ n11127;
  assign n11136 = n11135 ^ n11131;
  assign n11124 = n11025 ^ n11024;
  assign n11125 = n11027 & ~n11124;
  assign n11126 = n11125 ^ n11026;
  assign n11137 = n11136 ^ n11126;
  assign n11157 = n11156 ^ n11137;
  assign n11162 = n11161 ^ n11157;
  assign n11117 = n11005 ^ n11004;
  assign n11118 = n11007 & ~n11117;
  assign n11119 = n11118 ^ n11006;
  assign n11114 = n11020 ^ n11019;
  assign n11115 = n11022 & ~n11114;
  assign n11116 = n11115 ^ n11021;
  assign n11120 = n11119 ^ n11116;
  assign n11111 = n10998 ^ n10997;
  assign n11112 = n10999 & ~n11111;
  assign n11113 = n11112 ^ n6590;
  assign n11121 = n11120 ^ n11113;
  assign n11108 = n11008 ^ n11000;
  assign n11109 = n11009 & ~n11108;
  assign n11110 = n11109 ^ n11003;
  assign n11122 = n11121 ^ n11110;
  assign n11105 = n11023 ^ n11018;
  assign n11106 = n11029 & ~n11105;
  assign n11107 = n11106 ^ n11028;
  assign n11123 = n11122 ^ n11107;
  assign n11163 = n11162 ^ n11123;
  assign n11102 = n11032 ^ n10967;
  assign n11103 = ~n11033 & n11102;
  assign n11104 = n11103 ^ n10967;
  assign n11164 = n11163 ^ n11104;
  assign n11096 = ~n10984 & n10993;
  assign n11097 = n11096 ^ n10989;
  assign n11093 = x35 & x60;
  assign n11092 = x36 & x59;
  assign n11094 = n11093 ^ n11092;
  assign n11089 = n11015 ^ n11014;
  assign n11090 = n11017 & ~n11089;
  assign n11091 = n11090 ^ n11016;
  assign n11095 = n11094 ^ n11091;
  assign n11098 = n11097 ^ n11095;
  assign n11086 = n10973 ^ n10970;
  assign n11087 = n10977 & ~n11086;
  assign n11088 = n11087 ^ n10976;
  assign n11099 = n11098 ^ n11088;
  assign n11083 = n10994 ^ n10978;
  assign n11084 = n10995 & ~n11083;
  assign n11085 = n11084 ^ n10981;
  assign n11100 = n11099 ^ n11085;
  assign n11080 = n11030 ^ n11010;
  assign n11081 = n11031 & ~n11080;
  assign n11082 = n11081 ^ n11013;
  assign n11101 = n11100 ^ n11082;
  assign n11165 = n11164 ^ n11101;
  assign n11166 = n11079 & n11165;
  assign n11167 = n10961 & n10964;
  assign n11168 = ~n11165 & n11167;
  assign n11169 = ~n11166 & ~n11168;
  assign n11170 = ~n11066 & ~n11169;
  assign n11171 = n10964 ^ n10961;
  assign n11172 = n11165 ^ n10964;
  assign n11173 = ~n11171 & ~n11172;
  assign n11174 = ~n11074 & n11173;
  assign n11175 = ~n11170 & ~n11174;
  assign n11176 = ~n11034 & n11066;
  assign n11177 = ~n11165 & n11176;
  assign n11178 = n11079 & n11177;
  assign n11179 = n11034 & n11074;
  assign n11180 = n11168 & n11179;
  assign n11181 = ~n11178 & ~n11180;
  assign n11182 = n11074 ^ n11066;
  assign n11183 = ~n11165 & n11182;
  assign n11184 = n11183 ^ n11066;
  assign n11185 = n11076 & n11184;
  assign n11186 = ~n11177 & n11185;
  assign n11187 = ~n11079 & n11186;
  assign n11188 = n11066 & n11165;
  assign n11189 = ~n11034 & ~n11184;
  assign n11190 = ~n11188 & ~n11189;
  assign n11191 = ~n11167 & ~n11190;
  assign n11192 = ~n11179 & ~n11189;
  assign n11193 = n11191 & ~n11192;
  assign n11194 = ~n11187 & ~n11193;
  assign n11195 = n11181 & n11194;
  assign n11196 = n11175 & n11195;
  assign n11285 = ~n11079 & ~n11165;
  assign n11286 = n11074 & ~n11176;
  assign n11287 = ~n11285 & ~n11286;
  assign n11288 = ~n11166 & ~n11191;
  assign n11289 = ~n11287 & n11288;
  assign n11273 = x35 & x61;
  assign n11272 = x34 & x62;
  assign n11274 = n11273 ^ n11272;
  assign n11271 = x33 & x63;
  assign n11275 = n11274 ^ n11271;
  assign n11268 = x43 & x53;
  assign n11267 = x42 & x54;
  assign n11269 = n11268 ^ n11267;
  assign n11266 = x41 & x55;
  assign n11270 = n11269 ^ n11266;
  assign n11276 = n11275 ^ n11270;
  assign n11263 = n11116 ^ n11113;
  assign n11264 = n11120 & ~n11263;
  assign n11265 = n11264 ^ n11119;
  assign n11277 = n11276 ^ n11265;
  assign n11260 = n11097 ^ n11088;
  assign n11261 = n11098 & ~n11260;
  assign n11262 = n11261 ^ n11088;
  assign n11278 = n11277 ^ n11262;
  assign n11256 = n11091 & n11094;
  assign n11257 = n7774 & n8976;
  assign n11258 = ~n11256 & ~n11257;
  assign n11252 = n11128 ^ n11127;
  assign n11253 = n11130 & ~n11252;
  assign n11254 = n11253 ^ n11129;
  assign n11249 = n11133 ^ n6521;
  assign n11250 = ~n11134 & n11249;
  assign n11251 = n11250 ^ n6521;
  assign n11255 = n11254 ^ n11251;
  assign n11259 = n11258 ^ n11255;
  assign n11279 = n11278 ^ n11259;
  assign n11242 = n11150 ^ n11149;
  assign n11243 = n11152 & ~n11242;
  assign n11244 = n11243 ^ n11151;
  assign n11239 = n11145 ^ n11144;
  assign n11240 = n11147 & ~n11239;
  assign n11241 = n11240 ^ n11146;
  assign n11245 = n11244 ^ n11241;
  assign n11237 = ~x47 & ~n11142;
  assign n11238 = x48 & ~n11237;
  assign n11246 = n11245 ^ n11238;
  assign n11234 = n11148 ^ n11143;
  assign n11235 = n11154 & ~n11234;
  assign n11236 = n11235 ^ n11153;
  assign n11247 = n11246 ^ n11236;
  assign n11231 = n11135 ^ n11126;
  assign n11232 = ~n11136 & n11231;
  assign n11233 = n11232 ^ n11126;
  assign n11248 = n11247 ^ n11233;
  assign n11280 = n11279 ^ n11248;
  assign n11228 = n11085 ^ n11082;
  assign n11229 = n11100 & n11228;
  assign n11230 = n11229 ^ n11082;
  assign n11281 = n11280 ^ n11230;
  assign n11221 = x47 & x49;
  assign n11220 = x46 & x50;
  assign n11222 = n11221 ^ n11220;
  assign n11219 = x45 & x51;
  assign n11223 = n11222 ^ n11219;
  assign n11216 = x44 & x52;
  assign n11215 = x39 & x57;
  assign n11217 = n11216 ^ n11215;
  assign n11214 = x38 & x58;
  assign n11218 = n11217 ^ n11214;
  assign n11224 = n11223 ^ n11218;
  assign n11211 = x40 & x56;
  assign n11210 = x37 & x59;
  assign n11212 = n11211 ^ n11210;
  assign n11209 = x36 & x60;
  assign n11213 = n11212 ^ n11209;
  assign n11225 = n11224 ^ n11213;
  assign n11206 = n11121 ^ n11107;
  assign n11207 = n11122 & ~n11206;
  assign n11208 = n11207 ^ n11110;
  assign n11226 = n11225 ^ n11208;
  assign n11203 = n11155 ^ n11137;
  assign n11204 = n11156 & ~n11203;
  assign n11205 = n11204 ^ n11140;
  assign n11227 = n11226 ^ n11205;
  assign n11282 = n11281 ^ n11227;
  assign n11200 = n11157 ^ n11123;
  assign n11201 = n11162 & ~n11200;
  assign n11202 = n11201 ^ n11161;
  assign n11283 = n11282 ^ n11202;
  assign n11197 = n11104 ^ n11101;
  assign n11198 = n11164 & n11197;
  assign n11199 = n11198 ^ n11163;
  assign n11284 = n11283 ^ n11199;
  assign n11290 = n11289 ^ n11284;
  assign n11372 = ~n11227 & n11281;
  assign n11373 = n11202 & ~n11372;
  assign n11374 = n11227 & ~n11281;
  assign n11375 = ~n11373 & ~n11374;
  assign n11379 = n11199 & ~n11375;
  assign n11380 = n11202 & n11374;
  assign n11381 = ~n11379 & ~n11380;
  assign n11376 = ~n11199 & n11375;
  assign n11377 = ~n11202 & n11372;
  assign n11378 = ~n11376 & ~n11377;
  assign n11382 = n11381 ^ n11378;
  assign n11383 = ~n11289 & n11382;
  assign n11384 = n11383 ^ n11381;
  assign n11385 = n11380 ^ n11377;
  assign n11386 = ~n11199 & n11385;
  assign n11387 = n11386 ^ n11380;
  assign n11388 = n11384 & ~n11387;
  assign n11361 = x47 & x50;
  assign n11360 = x46 & x51;
  assign n11362 = n11361 ^ n11360;
  assign n11359 = x40 & x57;
  assign n11363 = n11362 ^ n11359;
  assign n11356 = n11241 ^ n11238;
  assign n11357 = n11245 & ~n11356;
  assign n11358 = n11357 ^ n11244;
  assign n11364 = n11363 ^ n11358;
  assign n11354 = x35 & x62;
  assign n11353 = ~x48 & x49;
  assign n11355 = n11354 ^ n11353;
  assign n11365 = n11364 ^ n11355;
  assign n11350 = n11275 ^ n11265;
  assign n11351 = ~n11276 & n11350;
  assign n11352 = n11351 ^ n11265;
  assign n11366 = n11365 ^ n11352;
  assign n11345 = n11210 ^ n11209;
  assign n11346 = n11212 & ~n11345;
  assign n11347 = n11346 ^ n11211;
  assign n11342 = n11272 ^ n11271;
  assign n11343 = n11274 & ~n11342;
  assign n11344 = n11343 ^ n11273;
  assign n11348 = n11347 ^ n11344;
  assign n11339 = n11267 ^ n11266;
  assign n11340 = n11269 & ~n11339;
  assign n11341 = n11340 ^ n11268;
  assign n11349 = n11348 ^ n11341;
  assign n11367 = n11366 ^ n11349;
  assign n11334 = x36 & x61;
  assign n11331 = n11215 ^ n11214;
  assign n11332 = n11217 & ~n11331;
  assign n11333 = n11332 ^ n11216;
  assign n11335 = n11334 ^ n11333;
  assign n11328 = n11220 ^ n11219;
  assign n11329 = n11222 & ~n11328;
  assign n11330 = n11329 ^ n11221;
  assign n11336 = n11335 ^ n11330;
  assign n11325 = n11258 ^ n11254;
  assign n11326 = ~n11255 & ~n11325;
  assign n11327 = n11326 ^ n11258;
  assign n11337 = n11336 ^ n11327;
  assign n11322 = n11218 ^ n11213;
  assign n11323 = n11224 & ~n11322;
  assign n11324 = n11323 ^ n11223;
  assign n11338 = n11337 ^ n11324;
  assign n11368 = n11367 ^ n11338;
  assign n11319 = n11208 ^ n11205;
  assign n11320 = ~n11226 & n11319;
  assign n11321 = n11320 ^ n11205;
  assign n11369 = n11368 ^ n11321;
  assign n11316 = n11279 ^ n11230;
  assign n11317 = n11280 & ~n11316;
  assign n11318 = n11317 ^ n11230;
  assign n11370 = n11369 ^ n11318;
  assign n11311 = n11277 ^ n11259;
  assign n11312 = n11278 & n11311;
  assign n11313 = n11312 ^ n11262;
  assign n11308 = n11246 ^ n11233;
  assign n11309 = n11247 & ~n11308;
  assign n11310 = n11309 ^ n11236;
  assign n11314 = n11313 ^ n11310;
  assign n11303 = x42 & x55;
  assign n11302 = x41 & x56;
  assign n11304 = n11303 ^ n11302;
  assign n11301 = x34 & x63;
  assign n11305 = n11304 ^ n11301;
  assign n11298 = x39 & x58;
  assign n11297 = x38 & x59;
  assign n11299 = n11298 ^ n11297;
  assign n11296 = x37 & x60;
  assign n11300 = n11299 ^ n11296;
  assign n11306 = n11305 ^ n11300;
  assign n11293 = x43 & x54;
  assign n11292 = x44 & x53;
  assign n11294 = n11293 ^ n11292;
  assign n11291 = x45 & x52;
  assign n11295 = n11294 ^ n11291;
  assign n11307 = n11306 ^ n11295;
  assign n11315 = n11314 ^ n11307;
  assign n11371 = n11370 ^ n11315;
  assign n11389 = n11388 ^ n11371;
  assign n11472 = ~n11199 & ~n11202;
  assign n11473 = n11288 & ~n11472;
  assign n11474 = ~n11287 & n11473;
  assign n11475 = n11199 & n11202;
  assign n11476 = ~n11474 & ~n11475;
  assign n11477 = n11371 & ~n11374;
  assign n11478 = ~n11476 & ~n11477;
  assign n11479 = ~n11371 & ~n11372;
  assign n11480 = ~n11376 & n11479;
  assign n11481 = ~n11289 & ~n11480;
  assign n11482 = n11199 & n11373;
  assign n11483 = ~n11479 & ~n11482;
  assign n11484 = ~n11481 & ~n11483;
  assign n11485 = ~n11478 & ~n11484;
  assign n11460 = n11297 ^ n11296;
  assign n11461 = n11299 & ~n11460;
  assign n11462 = n11461 ^ n11298;
  assign n11457 = n11302 ^ n11301;
  assign n11458 = n11304 & ~n11457;
  assign n11459 = n11458 ^ n11303;
  assign n11463 = n11462 ^ n11459;
  assign n11454 = n11291 & n11294;
  assign n11401 = x44 & x54;
  assign n11455 = n11268 & n11401;
  assign n11456 = ~n11454 & ~n11455;
  assign n11464 = n11463 ^ n11456;
  assign n11451 = n11363 ^ n11355;
  assign n11452 = n11364 & ~n11451;
  assign n11453 = n11452 ^ n11358;
  assign n11465 = n11464 ^ n11453;
  assign n11446 = x48 & x50;
  assign n11445 = x47 & x51;
  assign n11447 = n11446 ^ n11445;
  assign n11444 = x46 & x52;
  assign n11448 = n11447 ^ n11444;
  assign n11441 = x45 & x53;
  assign n11440 = x40 & x58;
  assign n11442 = n11441 ^ n11440;
  assign n11439 = x39 & x59;
  assign n11443 = n11442 ^ n11439;
  assign n11449 = n11448 ^ n11443;
  assign n11436 = ~x48 & ~n11354;
  assign n11437 = x49 & ~n11436;
  assign n11434 = x37 & x61;
  assign n11433 = x36 & x62;
  assign n11435 = n11434 ^ n11433;
  assign n11438 = n11437 ^ n11435;
  assign n11450 = n11449 ^ n11438;
  assign n11466 = n11465 ^ n11450;
  assign n11428 = n11334 ^ n11330;
  assign n11429 = n11335 & ~n11428;
  assign n11430 = n11429 ^ n11333;
  assign n11425 = n11300 ^ n11295;
  assign n11426 = n11306 & ~n11425;
  assign n11427 = n11426 ^ n11305;
  assign n11431 = n11430 ^ n11427;
  assign n11422 = n11344 ^ n11341;
  assign n11423 = n11348 & ~n11422;
  assign n11424 = n11423 ^ n11347;
  assign n11432 = n11431 ^ n11424;
  assign n11467 = n11466 ^ n11432;
  assign n11419 = n11310 ^ n11307;
  assign n11420 = n11314 & ~n11419;
  assign n11421 = n11420 ^ n11313;
  assign n11468 = n11467 ^ n11421;
  assign n11414 = n11365 ^ n11349;
  assign n11415 = n11366 & ~n11414;
  assign n11416 = n11415 ^ n11352;
  assign n11411 = n11336 ^ n11324;
  assign n11412 = ~n11337 & ~n11411;
  assign n11413 = n11412 ^ n11327;
  assign n11417 = n11416 ^ n11413;
  assign n11406 = x42 & x56;
  assign n11405 = x41 & x57;
  assign n11407 = n11406 ^ n11405;
  assign n11404 = x38 & x60;
  assign n11408 = n11407 ^ n11404;
  assign n11400 = x43 & x55;
  assign n11402 = n11401 ^ n11400;
  assign n11399 = x35 & x63;
  assign n11403 = n11402 ^ n11399;
  assign n11409 = n11408 ^ n11403;
  assign n11396 = n11360 ^ n11359;
  assign n11397 = n11362 & ~n11396;
  assign n11398 = n11397 ^ n11361;
  assign n11410 = n11409 ^ n11398;
  assign n11418 = n11417 ^ n11410;
  assign n11469 = n11468 ^ n11418;
  assign n11393 = n11367 ^ n11321;
  assign n11394 = n11368 & n11393;
  assign n11395 = n11394 ^ n11321;
  assign n11470 = n11469 ^ n11395;
  assign n11390 = n11369 ^ n11315;
  assign n11391 = ~n11370 & n11390;
  assign n11392 = n11391 ^ n11318;
  assign n11471 = n11470 ^ n11392;
  assign n11486 = n11485 ^ n11471;
  assign n11558 = ~x35 & ~n9794;
  assign n11559 = x49 & x62;
  assign n11560 = ~n11558 & n11559;
  assign n11561 = ~x36 & ~n11434;
  assign n11562 = n11560 & ~n11561;
  assign n11563 = x48 & x49;
  assign n11564 = ~n11433 & ~n11563;
  assign n11565 = n11434 & ~n11564;
  assign n11566 = ~n11562 & ~n11565;
  assign n11554 = x39 & x60;
  assign n11553 = x38 & x61;
  assign n11555 = n11554 ^ n11553;
  assign n11552 = x36 & x63;
  assign n11556 = n11555 ^ n11552;
  assign n11549 = n11405 ^ n11404;
  assign n11550 = n11407 & ~n11549;
  assign n11551 = n11550 ^ n11406;
  assign n11557 = n11556 ^ n11551;
  assign n11567 = n11566 ^ n11557;
  assign n11546 = n11443 ^ n11438;
  assign n11547 = n11449 & ~n11546;
  assign n11548 = n11547 ^ n11448;
  assign n11568 = n11567 ^ n11548;
  assign n11541 = n11440 ^ n11439;
  assign n11542 = n11442 & ~n11541;
  assign n11543 = n11542 ^ n11441;
  assign n11538 = n11400 ^ n11399;
  assign n11539 = n11402 & ~n11538;
  assign n11540 = n11539 ^ n11401;
  assign n11544 = n11543 ^ n11540;
  assign n11535 = n11445 ^ n11444;
  assign n11536 = n11447 & ~n11535;
  assign n11537 = n11536 ^ n11446;
  assign n11545 = n11544 ^ n11537;
  assign n11569 = n11568 ^ n11545;
  assign n11531 = x37 & x62;
  assign n11530 = ~x49 & x50;
  assign n11532 = n11531 ^ n11530;
  assign n11527 = n11408 ^ n11398;
  assign n11528 = ~n11409 & n11527;
  assign n11529 = n11528 ^ n11398;
  assign n11533 = n11532 ^ n11529;
  assign n11524 = n11459 ^ n11456;
  assign n11525 = n11463 & n11524;
  assign n11526 = n11525 ^ n11462;
  assign n11534 = n11533 ^ n11526;
  assign n11570 = n11569 ^ n11534;
  assign n11521 = n11413 ^ n11410;
  assign n11522 = ~n11417 & n11521;
  assign n11523 = n11522 ^ n11416;
  assign n11571 = n11570 ^ n11523;
  assign n11514 = x48 & x51;
  assign n11513 = x43 & x56;
  assign n11515 = n11514 ^ n11513;
  assign n11512 = x42 & x57;
  assign n11516 = n11515 ^ n11512;
  assign n11509 = x44 & x55;
  assign n11508 = x41 & x58;
  assign n11510 = n11509 ^ n11508;
  assign n11507 = x40 & x59;
  assign n11511 = n11510 ^ n11507;
  assign n11517 = n11516 ^ n11511;
  assign n11504 = x47 & x52;
  assign n11503 = x46 & x53;
  assign n11505 = n11504 ^ n11503;
  assign n11502 = x45 & x54;
  assign n11506 = n11505 ^ n11502;
  assign n11518 = n11517 ^ n11506;
  assign n11499 = n11464 ^ n11450;
  assign n11500 = ~n11465 & n11499;
  assign n11501 = n11500 ^ n11453;
  assign n11519 = n11518 ^ n11501;
  assign n11496 = n11427 ^ n11424;
  assign n11497 = n11431 & ~n11496;
  assign n11498 = n11497 ^ n11430;
  assign n11520 = n11519 ^ n11498;
  assign n11572 = n11571 ^ n11520;
  assign n11493 = n11466 ^ n11421;
  assign n11494 = n11467 & ~n11493;
  assign n11495 = n11494 ^ n11421;
  assign n11573 = n11572 ^ n11495;
  assign n11490 = n11468 ^ n11395;
  assign n11491 = ~n11469 & ~n11490;
  assign n11492 = n11491 ^ n11395;
  assign n11574 = n11573 ^ n11492;
  assign n11487 = n11485 ^ n11392;
  assign n11488 = ~n11471 & ~n11487;
  assign n11489 = n11488 ^ n11485;
  assign n11575 = n11574 ^ n11489;
  assign n11652 = n11492 & n11495;
  assign n11653 = n11489 & ~n11652;
  assign n11654 = ~n11492 & ~n11495;
  assign n11655 = n11654 ^ n11520;
  assign n11656 = ~n11572 & n11655;
  assign n11657 = n11656 ^ n11571;
  assign n11658 = n11653 & n11657;
  assign n11659 = n11492 & n11520;
  assign n11660 = n11573 & n11659;
  assign n11661 = ~n11492 & ~n11520;
  assign n11662 = n11495 & ~n11571;
  assign n11663 = ~n11661 & n11662;
  assign n11664 = ~n11660 & ~n11663;
  assign n11665 = ~n11489 & ~n11664;
  assign n11666 = n11520 ^ n11495;
  assign n11667 = n11495 ^ n11492;
  assign n11668 = ~n11666 & ~n11667;
  assign n11669 = n11572 & n11668;
  assign n11670 = ~n11665 & ~n11669;
  assign n11671 = ~n11658 & n11670;
  assign n11643 = x49 & x51;
  assign n11642 = x48 & x52;
  assign n11644 = n11643 ^ n11642;
  assign n11641 = x47 & x53;
  assign n11645 = n11644 ^ n11641;
  assign n11638 = n11540 ^ n11537;
  assign n11639 = n11544 & ~n11638;
  assign n11640 = n11639 ^ n11543;
  assign n11646 = n11645 ^ n11640;
  assign n11635 = n11566 ^ n11551;
  assign n11636 = ~n11557 & ~n11635;
  assign n11637 = n11636 ^ n11566;
  assign n11647 = n11646 ^ n11637;
  assign n11624 = ~x49 & ~n11531;
  assign n11625 = x50 & ~n11624;
  assign n11626 = x37 & x63;
  assign n11627 = ~n11625 & ~n11626;
  assign n11628 = x49 & x63;
  assign n11629 = ~n10350 & ~n11628;
  assign n11630 = n10191 & ~n11629;
  assign n11631 = ~n11627 & ~n11630;
  assign n11621 = n11513 ^ n11512;
  assign n11622 = n11515 & ~n11621;
  assign n11623 = n11622 ^ n11514;
  assign n11632 = n11631 ^ n11623;
  assign n11618 = n11511 ^ n11506;
  assign n11619 = n11517 & ~n11618;
  assign n11620 = n11619 ^ n11516;
  assign n11633 = n11632 ^ n11620;
  assign n11613 = n11503 ^ n11502;
  assign n11614 = n11505 & ~n11613;
  assign n11615 = n11614 ^ n11504;
  assign n11610 = n11508 ^ n11507;
  assign n11611 = n11510 & ~n11610;
  assign n11612 = n11611 ^ n11509;
  assign n11616 = n11615 ^ n11612;
  assign n11607 = n11553 ^ n11552;
  assign n11608 = n11555 & ~n11607;
  assign n11609 = n11608 ^ n11554;
  assign n11617 = n11616 ^ n11609;
  assign n11634 = n11633 ^ n11617;
  assign n11648 = n11647 ^ n11634;
  assign n11604 = n11518 ^ n11498;
  assign n11605 = n11519 & ~n11604;
  assign n11606 = n11605 ^ n11501;
  assign n11649 = n11648 ^ n11606;
  assign n11601 = n11569 ^ n11523;
  assign n11602 = n11570 & ~n11601;
  assign n11603 = n11602 ^ n11523;
  assign n11650 = n11649 ^ n11603;
  assign n11594 = x45 & x55;
  assign n11593 = x44 & x56;
  assign n11595 = n11594 ^ n11593;
  assign n11592 = x43 & x57;
  assign n11596 = n11595 ^ n11592;
  assign n11589 = x46 & x54;
  assign n11588 = x42 & x58;
  assign n11590 = n11589 ^ n11588;
  assign n11587 = x41 & x59;
  assign n11591 = n11590 ^ n11587;
  assign n11597 = n11596 ^ n11591;
  assign n11584 = x40 & x60;
  assign n11583 = x39 & x61;
  assign n11585 = n11584 ^ n11583;
  assign n11582 = x38 & x62;
  assign n11586 = n11585 ^ n11582;
  assign n11598 = n11597 ^ n11586;
  assign n11579 = n11529 ^ n11526;
  assign n11580 = ~n11533 & n11579;
  assign n11581 = n11580 ^ n11526;
  assign n11599 = n11598 ^ n11581;
  assign n11576 = n11567 ^ n11545;
  assign n11577 = ~n11568 & n11576;
  assign n11578 = n11577 ^ n11548;
  assign n11600 = n11599 ^ n11578;
  assign n11651 = n11650 ^ n11600;
  assign n11672 = n11671 ^ n11651;
  assign n11745 = n11520 & ~n11571;
  assign n11746 = n11651 & ~n11745;
  assign n11747 = ~n11654 & ~n11746;
  assign n11748 = ~n11653 & n11747;
  assign n11749 = ~n11520 & n11571;
  assign n11750 = n11651 & ~n11652;
  assign n11751 = ~n11749 & ~n11750;
  assign n11752 = ~n11489 & n11751;
  assign n11753 = ~n11651 & ~n11657;
  assign n11754 = ~n11752 & ~n11753;
  assign n11755 = ~n11748 & n11754;
  assign n11733 = n11588 ^ n11587;
  assign n11734 = n11590 & ~n11733;
  assign n11735 = n11734 ^ n11589;
  assign n11730 = n11583 ^ n11582;
  assign n11731 = n11585 & ~n11730;
  assign n11732 = n11731 ^ n11584;
  assign n11736 = n11735 ^ n11732;
  assign n11727 = n11593 ^ n11592;
  assign n11728 = n11595 & ~n11727;
  assign n11729 = n11728 ^ n11594;
  assign n11737 = n11736 ^ n11729;
  assign n11724 = n11591 ^ n11586;
  assign n11725 = n11597 & ~n11724;
  assign n11726 = n11725 ^ n11596;
  assign n11738 = n11737 ^ n11726;
  assign n11721 = n11612 ^ n11609;
  assign n11722 = n11616 & ~n11721;
  assign n11723 = n11722 ^ n11615;
  assign n11739 = n11738 ^ n11723;
  assign n11718 = n11632 ^ n11617;
  assign n11719 = n11633 & ~n11718;
  assign n11720 = n11719 ^ n11620;
  assign n11740 = n11739 ^ n11720;
  assign n11715 = n11598 ^ n11578;
  assign n11716 = n11599 & ~n11715;
  assign n11717 = n11716 ^ n11581;
  assign n11741 = n11740 ^ n11717;
  assign n11708 = x49 & x52;
  assign n11707 = x48 & x53;
  assign n11709 = n11708 ^ n11707;
  assign n11706 = x44 & x57;
  assign n11710 = n11709 ^ n11706;
  assign n11703 = x47 & x54;
  assign n11702 = x46 & x55;
  assign n11704 = n11703 ^ n11702;
  assign n11701 = x38 & x63;
  assign n11705 = n11704 ^ n11701;
  assign n11711 = n11710 ^ n11705;
  assign n11698 = x45 & x56;
  assign n11697 = x43 & x58;
  assign n11699 = n11698 ^ n11697;
  assign n11696 = x42 & x59;
  assign n11700 = n11699 ^ n11696;
  assign n11712 = n11711 ^ n11700;
  assign n11693 = n11645 ^ n11637;
  assign n11694 = n11646 & n11693;
  assign n11695 = n11694 ^ n11640;
  assign n11713 = n11712 ^ n11695;
  assign n11689 = ~n11623 & n11631;
  assign n11690 = n11689 ^ n11627;
  assign n11686 = x40 & x61;
  assign n11685 = x41 & x60;
  assign n11687 = n11686 ^ n11685;
  assign n11682 = n11642 ^ n11641;
  assign n11683 = n11644 & ~n11682;
  assign n11684 = n11683 ^ n11643;
  assign n11688 = n11687 ^ n11684;
  assign n11691 = n11690 ^ n11688;
  assign n11680 = x39 & x62;
  assign n11679 = ~x50 & x51;
  assign n11681 = n11680 ^ n11679;
  assign n11692 = n11691 ^ n11681;
  assign n11714 = n11713 ^ n11692;
  assign n11742 = n11741 ^ n11714;
  assign n11676 = n11647 ^ n11606;
  assign n11677 = n11648 & ~n11676;
  assign n11678 = n11677 ^ n11606;
  assign n11743 = n11742 ^ n11678;
  assign n11673 = n11649 ^ n11600;
  assign n11674 = ~n11650 & n11673;
  assign n11675 = n11674 ^ n11603;
  assign n11744 = n11743 ^ n11675;
  assign n11756 = n11755 ^ n11744;
  assign n11823 = n11741 ^ n11678;
  assign n11824 = n11742 & n11823;
  assign n11825 = n11824 ^ n11678;
  assign n11826 = ~n11675 & ~n11825;
  assign n11827 = n11714 & ~n11741;
  assign n11828 = ~n11678 & n11827;
  assign n11829 = ~n11826 & ~n11828;
  assign n11830 = n11755 & ~n11829;
  assign n11831 = ~n11714 & n11741;
  assign n11832 = n11678 & n11831;
  assign n11833 = n11832 ^ n11828;
  assign n11834 = n11675 & n11833;
  assign n11835 = n11834 ^ n11828;
  assign n11836 = ~n11830 & ~n11835;
  assign n11837 = n11675 & n11825;
  assign n11838 = ~n11832 & ~n11837;
  assign n11839 = ~n11755 & ~n11838;
  assign n11840 = n11836 & ~n11839;
  assign n11816 = n11712 ^ n11692;
  assign n11817 = n11713 & n11816;
  assign n11818 = n11817 ^ n11695;
  assign n11813 = n11726 ^ n11723;
  assign n11814 = ~n11738 & n11813;
  assign n11815 = n11814 ^ n11723;
  assign n11819 = n11818 ^ n11815;
  assign n11808 = n11732 ^ n11729;
  assign n11809 = n11736 & ~n11808;
  assign n11810 = n11809 ^ n11735;
  assign n11805 = n11705 ^ n11700;
  assign n11806 = n11711 & ~n11805;
  assign n11807 = n11806 ^ n11710;
  assign n11811 = n11810 ^ n11807;
  assign n11800 = n11702 ^ n11701;
  assign n11801 = n11704 & ~n11800;
  assign n11802 = n11801 ^ n11703;
  assign n11797 = n11707 ^ n11706;
  assign n11798 = n11709 & ~n11797;
  assign n11799 = n11798 ^ n11708;
  assign n11803 = n11802 ^ n11799;
  assign n11795 = ~x50 & ~n11680;
  assign n11796 = x51 & ~n11795;
  assign n11804 = n11803 ^ n11796;
  assign n11812 = n11811 ^ n11804;
  assign n11820 = n11819 ^ n11812;
  assign n11789 = n11684 & n11687;
  assign n11785 = x41 & x61;
  assign n11790 = n11584 & n11785;
  assign n11791 = ~n11789 & ~n11790;
  assign n11784 = x42 & x60;
  assign n11786 = n11785 ^ n11784;
  assign n11783 = x39 & x63;
  assign n11787 = n11786 ^ n11783;
  assign n11780 = n11697 ^ n11696;
  assign n11781 = n11699 & ~n11780;
  assign n11782 = n11781 ^ n11698;
  assign n11788 = n11787 ^ n11782;
  assign n11792 = n11791 ^ n11788;
  assign n11775 = x50 & x52;
  assign n11774 = x49 & x53;
  assign n11776 = n11775 ^ n11774;
  assign n11773 = x48 & x54;
  assign n11777 = n11776 ^ n11773;
  assign n11770 = x44 & x58;
  assign n11769 = x43 & x59;
  assign n11771 = n11770 ^ n11769;
  assign n11768 = x40 & x62;
  assign n11772 = n11771 ^ n11768;
  assign n11778 = n11777 ^ n11772;
  assign n11765 = x47 & x55;
  assign n11764 = x46 & x56;
  assign n11766 = n11765 ^ n11764;
  assign n11763 = x45 & x57;
  assign n11767 = n11766 ^ n11763;
  assign n11779 = n11778 ^ n11767;
  assign n11793 = n11792 ^ n11779;
  assign n11760 = n11688 ^ n11681;
  assign n11761 = ~n11691 & ~n11760;
  assign n11762 = n11761 ^ n11690;
  assign n11794 = n11793 ^ n11762;
  assign n11821 = n11820 ^ n11794;
  assign n11757 = n11720 ^ n11717;
  assign n11758 = ~n11740 & n11757;
  assign n11759 = n11758 ^ n11717;
  assign n11822 = n11821 ^ n11759;
  assign n11841 = n11840 ^ n11822;
  assign n11908 = n11822 & ~n11828;
  assign n11909 = ~n11832 & ~n11908;
  assign n11910 = n11675 & ~n11909;
  assign n11911 = n11822 & n11825;
  assign n11912 = ~n11910 & ~n11911;
  assign n11913 = n11755 & n11912;
  assign n11914 = ~n11675 & n11909;
  assign n11915 = ~n11822 & ~n11825;
  assign n11916 = ~n11914 & ~n11915;
  assign n11917 = ~n11913 & n11916;
  assign n11898 = n11799 ^ n11796;
  assign n11899 = n11803 & ~n11898;
  assign n11900 = n11899 ^ n11802;
  assign n11895 = n11772 ^ n11767;
  assign n11896 = n11778 & ~n11895;
  assign n11897 = n11896 ^ n11777;
  assign n11901 = n11900 ^ n11897;
  assign n11892 = n11791 ^ n11782;
  assign n11893 = ~n11788 & ~n11892;
  assign n11894 = n11893 ^ n11791;
  assign n11902 = n11901 ^ n11894;
  assign n11889 = n11807 ^ n11804;
  assign n11890 = n11811 & ~n11889;
  assign n11891 = n11890 ^ n11810;
  assign n11903 = n11902 ^ n11891;
  assign n11886 = n11792 ^ n11762;
  assign n11887 = n11793 & n11886;
  assign n11888 = n11887 ^ n11762;
  assign n11904 = n11903 ^ n11888;
  assign n11881 = x40 & x63;
  assign n11878 = n11764 ^ n11763;
  assign n11879 = n11766 & ~n11878;
  assign n11880 = n11879 ^ n11765;
  assign n11882 = n11881 ^ n11880;
  assign n11875 = n11774 ^ n11773;
  assign n11876 = n11776 & ~n11875;
  assign n11877 = n11876 ^ n11775;
  assign n11883 = n11882 ^ n11877;
  assign n11870 = x50 & x53;
  assign n11869 = x49 & x54;
  assign n11871 = n11870 ^ n11869;
  assign n11868 = x48 & x55;
  assign n11872 = n11871 ^ n11868;
  assign n11865 = x47 & x56;
  assign n11864 = x46 & x57;
  assign n11866 = n11865 ^ n11864;
  assign n11863 = x43 & x60;
  assign n11867 = n11866 ^ n11863;
  assign n11873 = n11872 ^ n11867;
  assign n11861 = x41 & x62;
  assign n11860 = ~x51 & x52;
  assign n11862 = n11861 ^ n11860;
  assign n11874 = n11873 ^ n11862;
  assign n11884 = n11883 ^ n11874;
  assign n11855 = x45 & x58;
  assign n11854 = x44 & x59;
  assign n11856 = n11855 ^ n11854;
  assign n11857 = n11856 ^ n10186;
  assign n11851 = n11769 ^ n11768;
  assign n11852 = n11771 & ~n11851;
  assign n11853 = n11852 ^ n11770;
  assign n11858 = n11857 ^ n11853;
  assign n11848 = n11784 ^ n11783;
  assign n11849 = n11786 & ~n11848;
  assign n11850 = n11849 ^ n11785;
  assign n11859 = n11858 ^ n11850;
  assign n11885 = n11884 ^ n11859;
  assign n11905 = n11904 ^ n11885;
  assign n11845 = n11815 ^ n11812;
  assign n11846 = n11819 & ~n11845;
  assign n11847 = n11846 ^ n11818;
  assign n11906 = n11905 ^ n11847;
  assign n11842 = n11794 ^ n11759;
  assign n11843 = n11821 & ~n11842;
  assign n11844 = n11843 ^ n11820;
  assign n11907 = n11906 ^ n11844;
  assign n11918 = n11917 ^ n11907;
  assign n11997 = ~n11844 & ~n11906;
  assign n11998 = n11916 & ~n11997;
  assign n11999 = ~n11913 & n11998;
  assign n12000 = n11844 & n11906;
  assign n12001 = ~n11999 & ~n12000;
  assign n11992 = n11904 ^ n11847;
  assign n11993 = ~n11905 & n11992;
  assign n11994 = n11993 ^ n11847;
  assign n11989 = n11891 ^ n11888;
  assign n11990 = n11903 & ~n11989;
  assign n11991 = n11990 ^ n11888;
  assign n11995 = n11994 ^ n11991;
  assign n11964 = x51 & x52;
  assign n11966 = x42 & x62;
  assign n11965 = ~x62 & x63;
  assign n11967 = n11966 ^ n11965;
  assign n11968 = x41 & n11967;
  assign n11969 = n11968 ^ n11966;
  assign n11970 = ~n11964 & n11969;
  assign n11971 = x63 ^ x42;
  assign n11972 = x52 & x62;
  assign n11973 = x41 & n11972;
  assign n11974 = ~n11971 & n11973;
  assign n11975 = ~n11970 & ~n11974;
  assign n11976 = ~x41 & ~n11966;
  assign n11977 = ~x62 & ~x63;
  assign n11978 = ~n11976 & ~n11977;
  assign n11979 = ~x52 & n11971;
  assign n11980 = n11979 ^ n11964;
  assign n11981 = n11978 & n11980;
  assign n11982 = n11981 ^ n11964;
  assign n11983 = n11975 & ~n11982;
  assign n11961 = n11881 ^ n11877;
  assign n11962 = n11882 & ~n11961;
  assign n11963 = n11962 ^ n11880;
  assign n11984 = n11983 ^ n11963;
  assign n11958 = n11857 ^ n11850;
  assign n11959 = n11858 & ~n11958;
  assign n11960 = n11959 ^ n11853;
  assign n11985 = n11984 ^ n11960;
  assign n11955 = n11874 ^ n11859;
  assign n11956 = n11884 & ~n11955;
  assign n11957 = n11956 ^ n11883;
  assign n11986 = n11985 ^ n11957;
  assign n11952 = n11900 ^ n11894;
  assign n11953 = ~n11901 & ~n11952;
  assign n11954 = n11953 ^ n11894;
  assign n11987 = n11986 ^ n11954;
  assign n11945 = x45 & x59;
  assign n11944 = x44 & x60;
  assign n11946 = n11945 ^ n11944;
  assign n11943 = x43 & x61;
  assign n11947 = n11946 ^ n11943;
  assign n11940 = x51 & x53;
  assign n11939 = x50 & x54;
  assign n11941 = n11940 ^ n11939;
  assign n11938 = x49 & x55;
  assign n11942 = n11941 ^ n11938;
  assign n11948 = n11947 ^ n11942;
  assign n11935 = x48 & x56;
  assign n11934 = x47 & x57;
  assign n11936 = n11935 ^ n11934;
  assign n11933 = x46 & x58;
  assign n11937 = n11936 ^ n11933;
  assign n11949 = n11948 ^ n11937;
  assign n11930 = n11867 ^ n11862;
  assign n11931 = n11873 & ~n11930;
  assign n11932 = n11931 ^ n11872;
  assign n11950 = n11949 ^ n11932;
  assign n11925 = n11855 ^ n10186;
  assign n11926 = ~n11856 & n11925;
  assign n11927 = n11926 ^ n10186;
  assign n11922 = n11864 ^ n11863;
  assign n11923 = n11866 & ~n11922;
  assign n11924 = n11923 ^ n11865;
  assign n11928 = n11927 ^ n11924;
  assign n11919 = n11869 ^ n11868;
  assign n11920 = n11871 & ~n11919;
  assign n11921 = n11920 ^ n11870;
  assign n11929 = n11928 ^ n11921;
  assign n11951 = n11950 ^ n11929;
  assign n11988 = n11987 ^ n11951;
  assign n11996 = n11995 ^ n11988;
  assign n12002 = n12001 ^ n11996;
  assign n12065 = ~n11951 & ~n11987;
  assign n12066 = n11991 & n12065;
  assign n12067 = n11951 & n11987;
  assign n12068 = ~n11991 & n12067;
  assign n12069 = ~n12066 & ~n12068;
  assign n12070 = n11995 & ~n12069;
  assign n12071 = n11991 ^ n11987;
  assign n12072 = ~n11988 & ~n12071;
  assign n12073 = n12072 ^ n11991;
  assign n12076 = ~n11994 & n12073;
  assign n12077 = ~n12066 & ~n12076;
  assign n12074 = ~n11994 & ~n12068;
  assign n12075 = ~n12073 & ~n12074;
  assign n12078 = n12077 ^ n12075;
  assign n12079 = ~n12001 & ~n12078;
  assign n12080 = n12079 ^ n12077;
  assign n12081 = ~n12070 & n12080;
  assign n12058 = n11983 ^ n11960;
  assign n12059 = ~n11984 & n12058;
  assign n12060 = n12059 ^ n11963;
  assign n12055 = n11942 ^ n11937;
  assign n12056 = n11948 & ~n12055;
  assign n12057 = n12056 ^ n11947;
  assign n12061 = n12060 ^ n12057;
  assign n12050 = n11934 ^ n11933;
  assign n12051 = n11936 & ~n12050;
  assign n12052 = n12051 ^ n11935;
  assign n12047 = n11939 ^ n11938;
  assign n12048 = n11941 & ~n12047;
  assign n12049 = n12048 ^ n11940;
  assign n12053 = n12052 ^ n12049;
  assign n12044 = n11944 ^ n11943;
  assign n12045 = n11946 & ~n12044;
  assign n12046 = n12045 ^ n11945;
  assign n12054 = n12053 ^ n12046;
  assign n12062 = n12061 ^ n12054;
  assign n12032 = ~x41 & ~n10876;
  assign n12033 = ~x42 & ~x63;
  assign n12034 = n11972 & ~n12033;
  assign n12035 = ~n12032 & n12034;
  assign n12036 = x52 & x63;
  assign n12037 = n10805 & n12036;
  assign n12024 = x42 & x63;
  assign n12038 = n11861 & n12024;
  assign n12039 = ~n12037 & ~n12038;
  assign n12040 = ~n12035 & n12039;
  assign n12028 = x48 & x57;
  assign n12027 = x47 & x58;
  assign n12029 = n12028 ^ n12027;
  assign n12026 = x46 & x59;
  assign n12030 = n12029 ^ n12026;
  assign n12022 = x45 & x60;
  assign n12021 = x44 & x61;
  assign n12023 = n12022 ^ n12021;
  assign n12025 = n12024 ^ n12023;
  assign n12031 = n12030 ^ n12025;
  assign n12041 = n12040 ^ n12031;
  assign n12018 = n11949 ^ n11929;
  assign n12019 = n11950 & ~n12018;
  assign n12020 = n12019 ^ n11932;
  assign n12042 = n12041 ^ n12020;
  assign n12013 = x51 & x54;
  assign n12012 = x50 & x55;
  assign n12014 = n12013 ^ n12012;
  assign n12011 = x49 & x56;
  assign n12015 = n12014 ^ n12011;
  assign n12008 = n11924 ^ n11921;
  assign n12009 = n11928 & ~n12008;
  assign n12010 = n12009 ^ n11927;
  assign n12016 = n12015 ^ n12010;
  assign n12006 = ~x52 & x53;
  assign n12007 = n12006 ^ n10182;
  assign n12017 = n12016 ^ n12007;
  assign n12043 = n12042 ^ n12017;
  assign n12063 = n12062 ^ n12043;
  assign n12003 = n11957 ^ n11954;
  assign n12004 = n11986 & ~n12003;
  assign n12005 = n12004 ^ n11954;
  assign n12064 = n12063 ^ n12005;
  assign n12082 = n12081 ^ n12064;
  assign n12140 = n12064 & ~n12070;
  assign n12141 = ~n12075 & ~n12140;
  assign n12142 = ~n12001 & ~n12141;
  assign n12143 = n12064 & n12077;
  assign n12144 = n11994 & n12068;
  assign n12145 = ~n12143 & ~n12144;
  assign n12146 = ~n12142 & n12145;
  assign n12131 = x52 & x54;
  assign n12130 = x51 & x55;
  assign n12132 = n12131 ^ n12130;
  assign n12129 = x50 & x56;
  assign n12133 = n12132 ^ n12129;
  assign n12126 = x49 & x57;
  assign n12125 = x48 & x58;
  assign n12127 = n12126 ^ n12125;
  assign n12124 = x47 & x59;
  assign n12128 = n12127 ^ n12124;
  assign n12134 = n12133 ^ n12128;
  assign n12121 = n12049 ^ n12046;
  assign n12122 = n12053 & ~n12121;
  assign n12123 = n12122 ^ n12052;
  assign n12135 = n12134 ^ n12123;
  assign n12118 = n12057 ^ n12054;
  assign n12119 = n12061 & ~n12118;
  assign n12120 = n12119 ^ n12060;
  assign n12136 = n12135 ^ n12120;
  assign n12113 = x46 & x60;
  assign n12112 = x45 & x61;
  assign n12114 = n12113 ^ n12112;
  assign n12111 = x44 & x62;
  assign n12115 = n12114 ^ n12111;
  assign n12108 = n12027 ^ n12026;
  assign n12109 = n12029 & ~n12108;
  assign n12110 = n12109 ^ n12028;
  assign n12116 = n12115 ^ n12110;
  assign n12105 = n12024 ^ n12022;
  assign n12106 = ~n12023 & n12105;
  assign n12107 = n12106 ^ n12024;
  assign n12117 = n12116 ^ n12107;
  assign n12137 = n12136 ^ n12117;
  assign n12099 = n12015 ^ n12007;
  assign n12100 = n12016 & ~n12099;
  assign n12101 = n12100 ^ n12010;
  assign n12096 = n12040 ^ n12030;
  assign n12097 = ~n12031 & ~n12096;
  assign n12098 = n12097 ^ n12040;
  assign n12102 = n12101 ^ n12098;
  assign n12092 = ~x52 & ~n10182;
  assign n12093 = x53 & ~n12092;
  assign n12094 = n12093 ^ n10351;
  assign n12089 = n12012 ^ n12011;
  assign n12090 = n12014 & ~n12089;
  assign n12091 = n12090 ^ n12013;
  assign n12095 = n12094 ^ n12091;
  assign n12103 = n12102 ^ n12095;
  assign n12086 = n12041 ^ n12017;
  assign n12087 = ~n12042 & n12086;
  assign n12088 = n12087 ^ n12020;
  assign n12104 = n12103 ^ n12088;
  assign n12138 = n12137 ^ n12104;
  assign n12083 = n12043 ^ n12005;
  assign n12084 = ~n12063 & ~n12083;
  assign n12085 = n12084 ^ n12062;
  assign n12139 = n12138 ^ n12085;
  assign n12147 = n12146 ^ n12139;
  assign n12207 = n12085 & ~n12138;
  assign n12208 = n12145 & ~n12207;
  assign n12209 = ~n12142 & n12208;
  assign n12210 = ~n12085 & n12138;
  assign n12211 = ~n12209 & ~n12210;
  assign n12197 = x46 & x61;
  assign n12196 = x47 & x60;
  assign n12198 = n12197 ^ n12196;
  assign n12193 = n12130 ^ n12129;
  assign n12194 = n12132 & ~n12193;
  assign n12195 = n12194 ^ n12131;
  assign n12199 = n12198 ^ n12195;
  assign n12190 = x52 & x55;
  assign n12189 = x51 & x56;
  assign n12191 = n12190 ^ n12189;
  assign n12188 = x50 & x57;
  assign n12192 = n12191 ^ n12188;
  assign n12200 = n12199 ^ n12192;
  assign n12186 = x45 & x62;
  assign n12185 = ~x53 & x54;
  assign n12187 = n12186 ^ n12185;
  assign n12201 = n12200 ^ n12187;
  assign n12180 = n12112 ^ n12111;
  assign n12181 = n12114 & ~n12180;
  assign n12182 = n12181 ^ n12113;
  assign n12177 = n12125 ^ n12124;
  assign n12178 = n12127 & ~n12177;
  assign n12179 = n12178 ^ n12126;
  assign n12183 = n12182 ^ n12179;
  assign n12174 = x49 & x58;
  assign n12173 = x48 & x59;
  assign n12175 = n12174 ^ n12173;
  assign n12172 = x44 & x63;
  assign n12176 = n12175 ^ n12172;
  assign n12184 = n12183 ^ n12176;
  assign n12202 = n12201 ^ n12184;
  assign n12169 = n12098 ^ n12095;
  assign n12170 = ~n12102 & n12169;
  assign n12171 = n12170 ^ n12101;
  assign n12203 = n12202 ^ n12171;
  assign n12160 = n12091 & n12093;
  assign n12161 = ~n10351 & ~n12160;
  assign n12162 = x52 & x53;
  assign n12163 = x53 & x62;
  assign n12164 = ~n12162 & ~n12163;
  assign n12165 = ~n12091 & n12164;
  assign n12166 = ~n12161 & ~n12165;
  assign n12157 = n12115 ^ n12107;
  assign n12158 = n12116 & ~n12157;
  assign n12159 = n12158 ^ n12110;
  assign n12167 = n12166 ^ n12159;
  assign n12154 = n12133 ^ n12123;
  assign n12155 = ~n12134 & n12154;
  assign n12156 = n12155 ^ n12123;
  assign n12168 = n12167 ^ n12156;
  assign n12204 = n12203 ^ n12168;
  assign n12151 = n12135 ^ n12117;
  assign n12152 = n12136 & ~n12151;
  assign n12153 = n12152 ^ n12120;
  assign n12205 = n12204 ^ n12153;
  assign n12148 = n12137 ^ n12088;
  assign n12149 = n12104 & n12148;
  assign n12150 = n12149 ^ n12137;
  assign n12206 = n12205 ^ n12150;
  assign n12212 = n12211 ^ n12206;
  assign n12260 = ~n12168 & ~n12203;
  assign n12261 = ~n12150 & ~n12153;
  assign n12263 = n12150 & n12153;
  assign n12264 = n12168 & n12203;
  assign n12265 = ~n12263 & ~n12264;
  assign n12268 = ~n12261 & ~n12265;
  assign n12269 = ~n12260 & n12268;
  assign n12262 = ~n12260 & ~n12261;
  assign n12266 = n12265 ^ n12262;
  assign n12267 = ~n12211 & n12266;
  assign n12270 = n12269 ^ n12267;
  assign n12271 = n12153 ^ n12150;
  assign n12272 = n12203 ^ n12153;
  assign n12273 = ~n12204 & ~n12272;
  assign n12274 = ~n12271 & n12273;
  assign n12275 = ~n12270 & ~n12274;
  assign n12251 = n12173 ^ n12172;
  assign n12252 = n12175 & ~n12251;
  assign n12253 = n12252 ^ n12174;
  assign n12248 = n12189 ^ n12188;
  assign n12249 = n12191 & ~n12248;
  assign n12250 = n12249 ^ n12190;
  assign n12254 = n12253 ^ n12250;
  assign n12246 = ~x53 & ~n12186;
  assign n12247 = x54 & ~n12246;
  assign n12255 = n12254 ^ n12247;
  assign n12243 = n12166 ^ n12156;
  assign n12244 = ~n12167 & n12243;
  assign n12245 = n12244 ^ n12156;
  assign n12256 = n12255 ^ n12245;
  assign n12238 = x47 & x61;
  assign n12239 = n12238 ^ n10913;
  assign n12237 = x45 & x63;
  assign n12240 = n12239 ^ n12237;
  assign n12234 = x50 & x58;
  assign n12233 = x49 & x59;
  assign n12235 = n12234 ^ n12233;
  assign n12232 = x48 & x60;
  assign n12236 = n12235 ^ n12232;
  assign n12241 = n12240 ^ n12236;
  assign n12229 = n12197 ^ n12195;
  assign n12230 = ~n12198 & n12229;
  assign n12231 = n12230 ^ n12195;
  assign n12242 = n12241 ^ n12231;
  assign n12257 = n12256 ^ n12242;
  assign n12226 = n12201 ^ n12171;
  assign n12227 = ~n12202 & n12226;
  assign n12228 = n12227 ^ n12171;
  assign n12258 = n12257 ^ n12228;
  assign n12221 = x53 & x55;
  assign n12220 = x52 & x56;
  assign n12222 = n12221 ^ n12220;
  assign n12219 = x51 & x57;
  assign n12223 = n12222 ^ n12219;
  assign n12216 = n12179 ^ n12176;
  assign n12217 = n12183 & ~n12216;
  assign n12218 = n12217 ^ n12182;
  assign n12224 = n12223 ^ n12218;
  assign n12213 = n12192 ^ n12187;
  assign n12214 = n12200 & ~n12213;
  assign n12215 = n12214 ^ n12199;
  assign n12225 = n12224 ^ n12215;
  assign n12259 = n12258 ^ n12225;
  assign n12276 = n12275 ^ n12259;
  assign n12324 = n12259 & ~n12261;
  assign n12325 = ~n12264 & ~n12324;
  assign n12326 = n12259 & ~n12260;
  assign n12327 = ~n12263 & ~n12326;
  assign n12328 = ~n12325 & ~n12327;
  assign n12329 = ~n12211 & ~n12328;
  assign n12330 = ~n12259 & ~n12268;
  assign n12331 = n12260 & ~n12324;
  assign n12332 = ~n12330 & ~n12331;
  assign n12333 = ~n12329 & n12332;
  assign n12319 = n12257 ^ n12225;
  assign n12320 = n12258 & ~n12319;
  assign n12321 = n12320 ^ n12228;
  assign n12316 = n12255 ^ n12242;
  assign n12317 = n12256 & ~n12316;
  assign n12318 = n12317 ^ n12245;
  assign n12322 = n12321 ^ n12318;
  assign n12308 = n12233 ^ n12232;
  assign n12309 = n12235 & ~n12308;
  assign n12310 = n12309 ^ n12234;
  assign n12311 = n12310 ^ n10990;
  assign n12305 = n12220 ^ n12219;
  assign n12306 = n12222 & ~n12305;
  assign n12307 = n12306 ^ n12221;
  assign n12312 = n12311 ^ n12307;
  assign n12300 = x53 & x56;
  assign n12299 = x52 & x57;
  assign n12301 = n12300 ^ n12299;
  assign n12298 = x51 & x58;
  assign n12302 = n12301 ^ n12298;
  assign n12295 = x50 & x59;
  assign n12294 = x49 & x60;
  assign n12296 = n12295 ^ n12294;
  assign n12293 = x48 & x61;
  assign n12297 = n12296 ^ n12293;
  assign n12303 = n12302 ^ n12297;
  assign n12290 = n12238 ^ n12237;
  assign n12291 = n12239 & ~n12290;
  assign n12292 = n12291 ^ n10913;
  assign n12304 = n12303 ^ n12292;
  assign n12313 = n12312 ^ n12304;
  assign n12287 = n12218 ^ n12215;
  assign n12288 = ~n12224 & n12287;
  assign n12289 = n12288 ^ n12215;
  assign n12314 = n12313 ^ n12289;
  assign n12283 = ~x54 & x55;
  assign n12284 = n12283 ^ n10985;
  assign n12280 = n12250 ^ n12247;
  assign n12281 = n12254 & ~n12280;
  assign n12282 = n12281 ^ n12253;
  assign n12285 = n12284 ^ n12282;
  assign n12277 = n12240 ^ n12231;
  assign n12278 = ~n12241 & n12277;
  assign n12279 = n12278 ^ n12231;
  assign n12286 = n12285 ^ n12279;
  assign n12315 = n12314 ^ n12286;
  assign n12323 = n12322 ^ n12315;
  assign n12334 = n12333 ^ n12323;
  assign n12387 = ~n12286 & ~n12314;
  assign n12388 = ~n12318 & n12387;
  assign n12389 = n12321 & ~n12388;
  assign n12390 = n12286 & n12314;
  assign n12391 = ~n12318 & ~n12390;
  assign n12392 = ~n12387 & ~n12391;
  assign n12393 = ~n12389 & ~n12392;
  assign n12394 = ~n12333 & n12393;
  assign n12395 = n12318 & n12390;
  assign n12396 = ~n12388 & ~n12395;
  assign n12397 = ~n12322 & ~n12396;
  assign n12398 = ~n12394 & ~n12397;
  assign n12399 = n12321 & n12392;
  assign n12400 = ~n12395 & ~n12399;
  assign n12401 = n12333 & ~n12400;
  assign n12402 = n12398 & ~n12401;
  assign n12378 = x51 & x59;
  assign n12377 = x50 & x60;
  assign n12379 = n12378 ^ n12377;
  assign n12376 = x49 & x61;
  assign n12380 = n12379 ^ n12376;
  assign n12373 = n12299 ^ n12298;
  assign n12374 = n12301 & ~n12373;
  assign n12375 = n12374 ^ n12300;
  assign n12381 = n12380 ^ n12375;
  assign n12370 = n12294 ^ n12293;
  assign n12371 = n12296 & ~n12370;
  assign n12372 = n12371 ^ n12295;
  assign n12382 = n12381 ^ n12372;
  assign n12367 = n12282 ^ n12279;
  assign n12368 = ~n12285 & n12367;
  assign n12369 = n12368 ^ n12279;
  assign n12383 = n12382 ^ n12369;
  assign n12364 = n12302 ^ n12292;
  assign n12365 = ~n12303 & n12364;
  assign n12366 = n12365 ^ n12292;
  assign n12384 = n12383 ^ n12366;
  assign n12361 = n12312 ^ n12289;
  assign n12362 = ~n12313 & n12361;
  assign n12363 = n12362 ^ n12289;
  assign n12385 = n12384 ^ n12363;
  assign n12343 = x48 & x63;
  assign n12344 = ~x55 & ~n12343;
  assign n12345 = n10985 & ~n12344;
  assign n12346 = x48 & x62;
  assign n12347 = x47 & x63;
  assign n12348 = ~n12346 & ~n12347;
  assign n12349 = x54 & x55;
  assign n12350 = ~n12348 & ~n12349;
  assign n12351 = ~n12345 & n12350;
  assign n12352 = n12348 & n12349;
  assign n12353 = x63 ^ x48;
  assign n12354 = x55 & x62;
  assign n12355 = ~n12353 & n12354;
  assign n12356 = x47 & n12355;
  assign n12357 = ~n12352 & ~n12356;
  assign n12358 = ~n12351 & n12357;
  assign n12340 = x54 & x56;
  assign n12339 = x53 & x57;
  assign n12341 = n12340 ^ n12339;
  assign n12338 = x52 & x58;
  assign n12342 = n12341 ^ n12338;
  assign n12359 = n12358 ^ n12342;
  assign n12335 = n12310 ^ n12307;
  assign n12336 = n12311 & ~n12335;
  assign n12337 = n12336 ^ n10990;
  assign n12360 = n12359 ^ n12337;
  assign n12386 = n12385 ^ n12360;
  assign n12403 = n12402 ^ n12386;
  assign n12449 = n12318 & n12321;
  assign n12450 = ~n12333 & ~n12449;
  assign n12451 = ~n12318 & ~n12321;
  assign n12452 = n12386 & ~n12390;
  assign n12453 = ~n12451 & ~n12452;
  assign n12454 = ~n12450 & n12453;
  assign n12455 = ~n12321 & n12391;
  assign n12456 = ~n12386 & ~n12455;
  assign n12457 = ~n12333 & ~n12456;
  assign n12458 = n12386 & ~n12449;
  assign n12459 = ~n12387 & ~n12458;
  assign n12460 = ~n12457 & n12459;
  assign n12461 = ~n12454 & ~n12460;
  assign n12439 = n12339 ^ n12338;
  assign n12440 = n12341 & ~n12439;
  assign n12441 = n12440 ^ n12340;
  assign n12436 = n12377 ^ n12376;
  assign n12437 = n12379 & ~n12436;
  assign n12438 = n12437 ^ n12378;
  assign n12442 = n12441 ^ n12438;
  assign n12429 = ~n12346 & ~n12349;
  assign n12430 = n12347 & ~n12429;
  assign n12431 = ~x47 & ~n11773;
  assign n12432 = ~x48 & ~x63;
  assign n12433 = n12354 & ~n12432;
  assign n12434 = ~n12431 & n12433;
  assign n12435 = ~n12430 & ~n12434;
  assign n12443 = n12442 ^ n12435;
  assign n12426 = n12358 ^ n12337;
  assign n12427 = n12359 & ~n12426;
  assign n12428 = n12427 ^ n12337;
  assign n12444 = n12443 ^ n12428;
  assign n12423 = n12380 ^ n12372;
  assign n12424 = n12381 & ~n12423;
  assign n12425 = n12424 ^ n12375;
  assign n12445 = n12444 ^ n12425;
  assign n12418 = x54 & x57;
  assign n12417 = x53 & x58;
  assign n12419 = n12418 ^ n12417;
  assign n12416 = x52 & x59;
  assign n12420 = n12419 ^ n12416;
  assign n12413 = x51 & x60;
  assign n12412 = x50 & x61;
  assign n12414 = n12413 ^ n12412;
  assign n12415 = n12414 ^ n12343;
  assign n12421 = n12420 ^ n12415;
  assign n12410 = ~x55 & x56;
  assign n12411 = n12410 ^ n11559;
  assign n12422 = n12421 ^ n12411;
  assign n12446 = n12445 ^ n12422;
  assign n12407 = n12382 ^ n12366;
  assign n12408 = n12383 & ~n12407;
  assign n12409 = n12408 ^ n12369;
  assign n12447 = n12446 ^ n12409;
  assign n12404 = n12363 ^ n12360;
  assign n12405 = n12385 & n12404;
  assign n12406 = n12405 ^ n12384;
  assign n12448 = n12447 ^ n12406;
  assign n12462 = n12461 ^ n12448;
  assign n12498 = ~n12422 & n12445;
  assign n12499 = n12409 & ~n12498;
  assign n12500 = n12422 & ~n12445;
  assign n12501 = ~n12499 & ~n12500;
  assign n12505 = ~n12409 & n12498;
  assign n12506 = n12406 & ~n12505;
  assign n12507 = n12501 & ~n12506;
  assign n12502 = n12406 & ~n12501;
  assign n12503 = n12409 & n12500;
  assign n12504 = ~n12502 & ~n12503;
  assign n12508 = n12507 ^ n12504;
  assign n12509 = ~n12461 & ~n12508;
  assign n12510 = n12509 ^ n12507;
  assign n12511 = n12505 ^ n12503;
  assign n12512 = n12406 & n12511;
  assign n12513 = n12512 ^ n12505;
  assign n12514 = ~n12510 & ~n12513;
  assign n12491 = x52 & x60;
  assign n12490 = x51 & x61;
  assign n12492 = n12491 ^ n12490;
  assign n12493 = n12492 ^ n11628;
  assign n12487 = n12413 ^ n12343;
  assign n12488 = ~n12414 & n12487;
  assign n12489 = n12488 ^ n12343;
  assign n12494 = n12493 ^ n12489;
  assign n12484 = x55 & x57;
  assign n12483 = x54 & x58;
  assign n12485 = n12484 ^ n12483;
  assign n12482 = x53 & x59;
  assign n12486 = n12485 ^ n12482;
  assign n12495 = n12494 ^ n12486;
  assign n12479 = n12443 ^ n12425;
  assign n12480 = ~n12444 & n12479;
  assign n12481 = n12480 ^ n12428;
  assign n12496 = n12495 ^ n12481;
  assign n12473 = ~x55 & ~n11559;
  assign n12474 = x56 & ~n12473;
  assign n12472 = x50 & x62;
  assign n12475 = n12474 ^ n12472;
  assign n12469 = n12417 ^ n12416;
  assign n12470 = n12419 & ~n12469;
  assign n12471 = n12470 ^ n12418;
  assign n12476 = n12475 ^ n12471;
  assign n12466 = n12415 ^ n12411;
  assign n12467 = n12421 & ~n12466;
  assign n12468 = n12467 ^ n12420;
  assign n12477 = n12476 ^ n12468;
  assign n12463 = n12438 ^ n12435;
  assign n12464 = n12442 & n12463;
  assign n12465 = n12464 ^ n12441;
  assign n12478 = n12477 ^ n12465;
  assign n12497 = n12496 ^ n12478;
  assign n12515 = n12514 ^ n12497;
  assign n12553 = ~n12406 & ~n12409;
  assign n12554 = ~n12461 & ~n12553;
  assign n12555 = n12406 & n12409;
  assign n12556 = n12497 & ~n12498;
  assign n12557 = ~n12555 & ~n12556;
  assign n12558 = ~n12554 & n12557;
  assign n12559 = n12406 & n12499;
  assign n12560 = ~n12497 & ~n12559;
  assign n12561 = ~n12461 & ~n12560;
  assign n12562 = n12497 & ~n12553;
  assign n12563 = ~n12500 & ~n12562;
  assign n12564 = ~n12561 & n12563;
  assign n12565 = ~n12558 & ~n12564;
  assign n12545 = x52 & x61;
  assign n12544 = x53 & x60;
  assign n12546 = n12545 ^ n12544;
  assign n12541 = n12483 ^ n12482;
  assign n12542 = n12485 & ~n12541;
  assign n12543 = n12542 ^ n12484;
  assign n12547 = n12546 ^ n12543;
  assign n12538 = n12474 ^ n12471;
  assign n12539 = ~n12475 & n12538;
  assign n12540 = n12539 ^ n12471;
  assign n12548 = n12547 ^ n12540;
  assign n12535 = n12493 ^ n12486;
  assign n12536 = n12494 & ~n12535;
  assign n12537 = n12536 ^ n12489;
  assign n12549 = n12548 ^ n12537;
  assign n12530 = x55 & x58;
  assign n12529 = x54 & x59;
  assign n12531 = n12530 ^ n12529;
  assign n12528 = x50 & x63;
  assign n12532 = n12531 ^ n12528;
  assign n12525 = n12491 ^ n11628;
  assign n12526 = ~n12492 & n12525;
  assign n12527 = n12526 ^ n11628;
  assign n12533 = n12532 ^ n12527;
  assign n12523 = x51 & x62;
  assign n12522 = ~x56 & x57;
  assign n12524 = n12523 ^ n12522;
  assign n12534 = n12533 ^ n12524;
  assign n12550 = n12549 ^ n12534;
  assign n12519 = n12468 ^ n12465;
  assign n12520 = ~n12477 & n12519;
  assign n12521 = n12520 ^ n12465;
  assign n12551 = n12550 ^ n12521;
  assign n12516 = n12495 ^ n12478;
  assign n12517 = n12496 & ~n12516;
  assign n12518 = n12517 ^ n12481;
  assign n12552 = n12551 ^ n12518;
  assign n12566 = n12565 ^ n12552;
  assign n12596 = ~n12518 & ~n12521;
  assign n12597 = ~n12534 & ~n12549;
  assign n12598 = ~n12596 & ~n12597;
  assign n12599 = n12518 & n12521;
  assign n12600 = n12534 & n12549;
  assign n12601 = ~n12599 & ~n12600;
  assign n12602 = ~n12598 & n12601;
  assign n12603 = ~n12565 & n12602;
  assign n12604 = n12549 ^ n12518;
  assign n12605 = n12534 ^ n12521;
  assign n12606 = ~n12550 & ~n12605;
  assign n12607 = ~n12604 & n12606;
  assign n12608 = ~n12603 & ~n12607;
  assign n12609 = ~n12597 & n12599;
  assign n12610 = ~n12596 & n12600;
  assign n12611 = ~n12609 & ~n12610;
  assign n12612 = n12565 & ~n12611;
  assign n12613 = n12608 & ~n12612;
  assign n12589 = x53 & x61;
  assign n12590 = n12589 ^ n11972;
  assign n12588 = x51 & x63;
  assign n12591 = n12590 ^ n12588;
  assign n12585 = x56 & x58;
  assign n12584 = x55 & x59;
  assign n12586 = n12585 ^ n12584;
  assign n12583 = x54 & x60;
  assign n12587 = n12586 ^ n12583;
  assign n12592 = n12591 ^ n12587;
  assign n12580 = n12532 ^ n12524;
  assign n12581 = n12533 & ~n12580;
  assign n12582 = n12581 ^ n12527;
  assign n12593 = n12592 ^ n12582;
  assign n12577 = n12540 ^ n12537;
  assign n12578 = ~n12548 & n12577;
  assign n12579 = n12578 ^ n12537;
  assign n12594 = n12593 ^ n12579;
  assign n12572 = n12543 & n12546;
  assign n12573 = n7409 & n12162;
  assign n12574 = ~n12572 & ~n12573;
  assign n12569 = n12529 ^ n12528;
  assign n12570 = n12531 & ~n12569;
  assign n12571 = n12570 ^ n12530;
  assign n12575 = n12574 ^ n12571;
  assign n12567 = ~x56 & ~n12523;
  assign n12568 = x57 & ~n12567;
  assign n12576 = n12575 ^ n12568;
  assign n12595 = n12594 ^ n12576;
  assign n12614 = n12613 ^ n12595;
  assign n12644 = ~n12518 & ~n12549;
  assign n12645 = n12565 & ~n12644;
  assign n12646 = n12518 & n12549;
  assign n12647 = ~n12521 & ~n12534;
  assign n12648 = ~n12595 & ~n12647;
  assign n12649 = ~n12646 & ~n12648;
  assign n12650 = ~n12645 & n12649;
  assign n12651 = n12646 & ~n12647;
  assign n12652 = n12595 & ~n12651;
  assign n12653 = n12565 & ~n12652;
  assign n12654 = ~n12595 & ~n12644;
  assign n12655 = n12521 & n12534;
  assign n12656 = ~n12654 & ~n12655;
  assign n12657 = ~n12653 & n12656;
  assign n12658 = ~n12650 & ~n12657;
  assign n12637 = x56 & x59;
  assign n12636 = x55 & x60;
  assign n12638 = n12637 ^ n12636;
  assign n12635 = x54 & x61;
  assign n12639 = n12638 ^ n12635;
  assign n12632 = n12571 ^ n12568;
  assign n12633 = ~n12575 & ~n12632;
  assign n12634 = n12633 ^ n12574;
  assign n12640 = n12639 ^ n12634;
  assign n12630 = ~x57 & x58;
  assign n12631 = n12630 ^ n12163;
  assign n12641 = n12640 ^ n12631;
  assign n12624 = n12589 ^ n12588;
  assign n12625 = n12590 & ~n12624;
  assign n12626 = n12625 ^ n11972;
  assign n12627 = n12626 ^ n12036;
  assign n12621 = n12584 ^ n12583;
  assign n12622 = n12586 & ~n12621;
  assign n12623 = n12622 ^ n12585;
  assign n12628 = n12627 ^ n12623;
  assign n12618 = n12591 ^ n12582;
  assign n12619 = ~n12592 & n12618;
  assign n12620 = n12619 ^ n12582;
  assign n12629 = n12628 ^ n12620;
  assign n12642 = n12641 ^ n12629;
  assign n12615 = n12593 ^ n12576;
  assign n12616 = n12594 & n12615;
  assign n12617 = n12616 ^ n12579;
  assign n12643 = n12642 ^ n12617;
  assign n12659 = n12658 ^ n12643;
  assign n12694 = n12620 & n12628;
  assign n12695 = ~n12641 & n12694;
  assign n12696 = ~n12617 & ~n12695;
  assign n12697 = n12641 ^ n12620;
  assign n12698 = ~n12629 & ~n12697;
  assign n12699 = n12698 ^ n12641;
  assign n12700 = ~n12696 & ~n12699;
  assign n12701 = n12658 & n12700;
  assign n12702 = n12617 & n12695;
  assign n12703 = ~n12701 & ~n12702;
  assign n12704 = ~n12620 & ~n12628;
  assign n12705 = n12641 & n12704;
  assign n12706 = n12617 & ~n12705;
  assign n12707 = n12699 & ~n12706;
  assign n12708 = ~n12658 & n12707;
  assign n12709 = ~n12617 & n12705;
  assign n12710 = ~n12708 & ~n12709;
  assign n12711 = n12703 & n12710;
  assign n12674 = x53 & ~n11965;
  assign n12675 = x57 & x58;
  assign n12676 = ~n12674 & ~n12675;
  assign n12677 = x54 & x62;
  assign n12678 = ~x53 & ~n12677;
  assign n12679 = n12676 & ~n12678;
  assign n12680 = x63 ^ x54;
  assign n12681 = n12163 & ~n12680;
  assign n12682 = x58 & n12681;
  assign n12683 = ~n12679 & ~n12682;
  assign n12684 = ~n11977 & ~n12678;
  assign n12685 = ~x58 & n12680;
  assign n12686 = n12685 ^ n12675;
  assign n12687 = n12684 & n12686;
  assign n12688 = n12687 ^ n12675;
  assign n12689 = n12683 & ~n12688;
  assign n12671 = n12636 ^ n12635;
  assign n12672 = n12638 & ~n12671;
  assign n12673 = n12672 ^ n12637;
  assign n12690 = n12689 ^ n12673;
  assign n12668 = x57 & x59;
  assign n12667 = x56 & x60;
  assign n12669 = n12668 ^ n12667;
  assign n12666 = x55 & x61;
  assign n12670 = n12669 ^ n12666;
  assign n12691 = n12690 ^ n12670;
  assign n12663 = n12626 ^ n12623;
  assign n12664 = n12627 & ~n12663;
  assign n12665 = n12664 ^ n12036;
  assign n12692 = n12691 ^ n12665;
  assign n12660 = n12639 ^ n12631;
  assign n12661 = ~n12640 & ~n12660;
  assign n12662 = n12661 ^ n12634;
  assign n12693 = n12692 ^ n12662;
  assign n12712 = n12711 ^ n12693;
  assign n12713 = n12662 & ~n12711;
  assign n12714 = ~n12665 & n12691;
  assign n12715 = ~n12713 & ~n12714;
  assign n12739 = ~x58 & x59;
  assign n12740 = n12739 ^ n12354;
  assign n12736 = n12673 ^ n12670;
  assign n12737 = ~n12690 & ~n12736;
  assign n12738 = n12737 ^ n12689;
  assign n12741 = n12740 ^ n12738;
  assign n12731 = x57 & x60;
  assign n12730 = x56 & x61;
  assign n12732 = n12731 ^ n12730;
  assign n12723 = x54 & x63;
  assign n12733 = n12732 ^ n12723;
  assign n12727 = n12667 ^ n12666;
  assign n12728 = n12669 & ~n12727;
  assign n12729 = n12728 ^ n12668;
  assign n12734 = n12733 ^ n12729;
  assign n12716 = ~x53 & ~n12418;
  assign n12717 = ~x54 & ~x63;
  assign n12718 = x58 & x62;
  assign n12719 = ~n12717 & n12718;
  assign n12720 = ~n12716 & n12719;
  assign n12721 = x58 & x63;
  assign n12722 = n12339 & n12721;
  assign n12724 = n12163 & n12723;
  assign n12725 = ~n12722 & ~n12724;
  assign n12726 = ~n12720 & n12725;
  assign n12735 = n12734 ^ n12726;
  assign n12742 = n12741 ^ n12735;
  assign n12743 = ~n12662 & n12710;
  assign n12744 = n12743 ^ n12703;
  assign n12745 = ~n12742 & n12744;
  assign n12746 = n12745 ^ n12703;
  assign n12747 = n12715 & ~n12746;
  assign n12748 = n12662 & n12703;
  assign n12749 = n12714 & n12742;
  assign n12750 = n12748 & n12749;
  assign n12751 = n12742 ^ n12691;
  assign n12752 = n12692 & n12751;
  assign n12753 = ~n12703 & n12752;
  assign n12754 = ~n12750 & ~n12753;
  assign n12755 = ~n12747 & n12754;
  assign n12756 = n12665 & ~n12691;
  assign n12757 = n12703 & ~n12742;
  assign n12758 = ~n12709 & n12742;
  assign n12759 = ~n12708 & n12758;
  assign n12760 = n12662 & ~n12759;
  assign n12761 = ~n12757 & ~n12760;
  assign n12762 = ~n12756 & ~n12761;
  assign n12763 = ~n12743 & n12757;
  assign n12764 = n12762 & ~n12763;
  assign n12765 = n12742 & n12756;
  assign n12766 = n12743 & n12765;
  assign n12767 = n12742 ^ n12665;
  assign n12768 = n12692 & n12767;
  assign n12769 = ~n12710 & n12768;
  assign n12770 = ~n12766 & ~n12769;
  assign n12771 = ~n12764 & n12770;
  assign n12772 = n12755 & n12771;
  assign n12802 = n12742 ^ n12714;
  assign n12803 = n12710 & ~n12748;
  assign n12804 = n12803 ^ n12742;
  assign n12805 = ~n12802 & ~n12804;
  assign n12806 = n12805 ^ n12714;
  assign n12807 = ~n12762 & ~n12806;
  assign n12797 = n12740 ^ n12735;
  assign n12798 = ~n12741 & n12797;
  assign n12799 = n12798 ^ n12738;
  assign n12794 = n12733 ^ n12726;
  assign n12795 = n12734 & n12794;
  assign n12796 = n12795 ^ n12729;
  assign n12800 = n12799 ^ n12796;
  assign n12781 = x59 & n12354;
  assign n12782 = x58 & x59;
  assign n12783 = x55 & x63;
  assign n12784 = ~n12782 & ~n12783;
  assign n12785 = ~n12781 & n12784;
  assign n12786 = x59 & x63;
  assign n12787 = n12530 & n12786;
  assign n12788 = x59 & x62;
  assign n12789 = n12783 & n12788;
  assign n12790 = ~n12787 & ~n12789;
  assign n12791 = ~n12785 & n12790;
  assign n12778 = n12730 ^ n12723;
  assign n12779 = n12732 & ~n12778;
  assign n12780 = n12779 ^ n12731;
  assign n12792 = n12791 ^ n12780;
  assign n12775 = x57 & x61;
  assign n12774 = x58 & x60;
  assign n12776 = n12775 ^ n12774;
  assign n12773 = x56 & x62;
  assign n12777 = n12776 ^ n12773;
  assign n12793 = n12792 ^ n12777;
  assign n12801 = n12800 ^ n12793;
  assign n12808 = n12807 ^ n12801;
  assign n12826 = n12796 ^ n12792;
  assign n12827 = ~n12793 & n12826;
  assign n12828 = n12827 ^ n12796;
  assign n12829 = ~n12799 & n12828;
  assign n12830 = n12777 & n12792;
  assign n12831 = n12796 & n12830;
  assign n12832 = ~n12829 & ~n12831;
  assign n12833 = n12807 & ~n12832;
  assign n12834 = ~n12777 & ~n12792;
  assign n12835 = ~n12796 & n12834;
  assign n12836 = ~n12831 & ~n12835;
  assign n12837 = n12800 & ~n12836;
  assign n12838 = ~n12833 & ~n12837;
  assign n12839 = ~n12799 & ~n12835;
  assign n12840 = ~n12828 & ~n12839;
  assign n12841 = ~n12807 & n12840;
  assign n12842 = n12838 & ~n12841;
  assign n12819 = ~x63 & ~n12780;
  assign n12820 = n12781 & ~n12819;
  assign n12821 = ~n12780 & ~n12787;
  assign n12822 = ~n12784 & ~n12821;
  assign n12823 = ~n12820 & ~n12822;
  assign n12815 = n12773 & n12776;
  assign n12816 = n7409 & n12675;
  assign n12817 = ~n12815 & ~n12816;
  assign n12813 = x56 & x63;
  assign n12812 = x58 & x61;
  assign n12814 = n12813 ^ n12812;
  assign n12818 = n12817 ^ n12814;
  assign n12824 = n12823 ^ n12818;
  assign n12810 = x57 & x62;
  assign n12809 = ~x59 & x60;
  assign n12811 = n12810 ^ n12809;
  assign n12825 = n12824 ^ n12811;
  assign n12843 = n12842 ^ n12825;
  assign n12859 = ~n12796 & n12799;
  assign n12860 = n12825 & ~n12859;
  assign n12861 = ~n12830 & ~n12860;
  assign n12862 = n12796 & ~n12799;
  assign n12863 = n12825 & ~n12834;
  assign n12864 = ~n12862 & ~n12863;
  assign n12865 = ~n12861 & ~n12864;
  assign n12866 = ~n12807 & ~n12865;
  assign n12867 = n12834 & ~n12860;
  assign n12868 = ~n12825 & n12832;
  assign n12869 = ~n12867 & ~n12868;
  assign n12870 = ~n12866 & n12869;
  assign n12853 = n12814 & ~n12817;
  assign n12854 = n12721 & n12730;
  assign n12855 = ~n12853 & ~n12854;
  assign n12850 = x59 & x61;
  assign n12851 = n12850 ^ n12718;
  assign n12849 = x57 & x63;
  assign n12852 = n12851 ^ n12849;
  assign n12856 = n12855 ^ n12852;
  assign n12847 = ~x59 & ~n12810;
  assign n12848 = x60 & ~n12847;
  assign n12857 = n12856 ^ n12848;
  assign n12844 = n12818 ^ n12811;
  assign n12845 = n12824 & n12844;
  assign n12846 = n12845 ^ n12823;
  assign n12858 = n12857 ^ n12846;
  assign n12871 = n12870 ^ n12858;
  assign n12881 = ~x60 & x61;
  assign n12882 = n12881 ^ n12788;
  assign n12883 = n12882 ^ n12721;
  assign n12878 = n12850 ^ n12849;
  assign n12879 = n12851 & ~n12878;
  assign n12880 = n12879 ^ n12718;
  assign n12884 = n12883 ^ n12880;
  assign n12875 = n12852 ^ n12848;
  assign n12876 = ~n12856 & ~n12875;
  assign n12877 = n12876 ^ n12855;
  assign n12885 = n12884 ^ n12877;
  assign n12872 = n12870 ^ n12857;
  assign n12873 = ~n12858 & ~n12872;
  assign n12874 = n12873 ^ n12870;
  assign n12886 = n12885 ^ n12874;
  assign n12894 = ~n12721 & n12877;
  assign n12895 = ~n12874 & n12877;
  assign n12896 = ~n12894 & ~n12895;
  assign n12897 = ~n12880 & ~n12882;
  assign n12898 = ~n12896 & n12897;
  assign n12901 = n12882 ^ n12880;
  assign n12902 = n12880 ^ n12877;
  assign n12903 = ~n12901 & ~n12902;
  assign n12904 = n12903 ^ n12877;
  assign n12905 = ~n12721 & n12904;
  assign n12899 = n12880 & n12882;
  assign n12900 = ~n12877 & n12899;
  assign n12906 = n12905 ^ n12900;
  assign n12907 = n12874 & n12906;
  assign n12908 = n12907 ^ n12905;
  assign n12909 = ~n12898 & ~n12908;
  assign n12910 = ~n12874 & ~n12900;
  assign n12911 = n12721 & ~n12904;
  assign n12912 = ~n12910 & n12911;
  assign n12913 = n12909 & ~n12912;
  assign n12887 = n12786 ^ n8432;
  assign n12888 = ~x61 & ~x62;
  assign n12889 = x60 & ~n12888;
  assign n12890 = n12889 ^ n12887;
  assign n12891 = n12887 & n12890;
  assign n12892 = ~x59 & n12891;
  assign n12893 = n12892 ^ n12890;
  assign n12914 = n12913 ^ n12893;
  assign n12923 = n12721 & ~n12895;
  assign n12924 = n12893 & ~n12897;
  assign n12925 = ~n12923 & ~n12924;
  assign n12926 = n12893 & ~n12894;
  assign n12927 = ~n12899 & ~n12926;
  assign n12928 = ~n12874 & n12927;
  assign n12929 = ~n12893 & n12904;
  assign n12930 = ~n12928 & ~n12929;
  assign n12931 = ~n12925 & n12930;
  assign n12915 = x59 & n7409;
  assign n12916 = x62 & ~n12786;
  assign n12917 = ~n12915 & ~n12916;
  assign n12918 = x60 & x63;
  assign n12919 = ~n12881 & ~n12918;
  assign n12920 = ~n12917 & ~n12919;
  assign n12921 = ~x62 & ~n12918;
  assign n12922 = ~n12920 & ~n12921;
  assign n12932 = n12931 ^ n12922;
  assign n12933 = ~x59 & x61;
  assign n12934 = n12931 & ~n12933;
  assign n12935 = n10350 & ~n12934;
  assign n12936 = ~n12888 & ~n12935;
  assign n12937 = ~x60 & ~n12936;
  assign n12938 = ~x61 & ~n10350;
  assign n12939 = ~n12931 & n12938;
  assign n12940 = x63 & ~n12915;
  assign n12941 = ~x62 & ~n12940;
  assign n12942 = ~n12939 & ~n12941;
  assign n12943 = x60 & ~n12938;
  assign n12944 = x59 & ~x61;
  assign n12945 = n10350 & ~n12944;
  assign n12946 = n12943 & ~n12945;
  assign n12947 = n12931 & n12946;
  assign n12948 = n12942 & ~n12947;
  assign n12949 = ~n12937 & n12948;
  assign n12950 = n8976 & n12931;
  assign n12951 = ~x61 & ~n12950;
  assign n12952 = n10350 & ~n12951;
  assign n12953 = n7409 & n12931;
  assign n12954 = ~x62 & ~n12915;
  assign n12955 = ~n12953 & n12954;
  assign n12956 = x63 & n12955;
  assign n12957 = ~n12952 & ~n12956;
  assign n12958 = x63 & ~n12955;
  assign y0 = x0;
  assign y1 = 1'b0;
  assign y2 = n65;
  assign y3 = n67;
  assign y4 = n72;
  assign y5 = ~n83;
  assign y6 = ~n96;
  assign y7 = ~n115;
  assign y8 = ~n146;
  assign y9 = n164;
  assign y10 = n197;
  assign y11 = ~n219;
  assign y12 = n255;
  assign y13 = n299;
  assign y14 = ~n335;
  assign y15 = n382;
  assign y16 = n427;
  assign y17 = n480;
  assign y18 = n538;
  assign y19 = n598;
  assign y20 = n664;
  assign y21 = n724;
  assign y22 = n795;
  assign y23 = ~n865;
  assign y24 = n937;
  assign y25 = ~n1014;
  assign y26 = ~n1094;
  assign y27 = n1186;
  assign y28 = ~n1271;
  assign y29 = n1355;
  assign y30 = ~n1452;
  assign y31 = n1551;
  assign y32 = ~n1649;
  assign y33 = n1747;
  assign y34 = n1845;
  assign y35 = n1964;
  assign y36 = ~n2083;
  assign y37 = ~n2193;
  assign y38 = ~n2313;
  assign y39 = n2432;
  assign y40 = ~n2557;
  assign y41 = ~n2678;
  assign y42 = ~n2816;
  assign y43 = ~n2947;
  assign y44 = n3087;
  assign y45 = ~n3225;
  assign y46 = n3371;
  assign y47 = ~n3514;
  assign y48 = n3668;
  assign y49 = ~n3812;
  assign y50 = n3956;
  assign y51 = n4121;
  assign y52 = ~n4277;
  assign y53 = n4435;
  assign y54 = ~n4608;
  assign y55 = n4777;
  assign y56 = n4939;
  assign y57 = ~n5111;
  assign y58 = ~n5280;
  assign y59 = n5468;
  assign y60 = n5654;
  assign y61 = ~n5832;
  assign y62 = ~n6022;
  assign y63 = n6215;
  assign y64 = n6403;
  assign y65 = ~n6605;
  assign y66 = n6794;
  assign y67 = n6989;
  assign y68 = ~n7174;
  assign y69 = ~n7352;
  assign y70 = ~n7537;
  assign y71 = n7709;
  assign y72 = ~n7877;
  assign y73 = ~n8049;
  assign y74 = ~n8216;
  assign y75 = ~n8386;
  assign y76 = n8548;
  assign y77 = ~n8708;
  assign y78 = n8863;
  assign y79 = ~n9017;
  assign y80 = n9167;
  assign y81 = n9310;
  assign y82 = n9458;
  assign y83 = n9599;
  assign y84 = ~n9741;
  assign y85 = n9879;
  assign y86 = ~n10004;
  assign y87 = n10134;
  assign y88 = ~n10280;
  assign y89 = n10403;
  assign y90 = n10517;
  assign y91 = n10626;
  assign y92 = n10731;
  assign y93 = ~n10844;
  assign y94 = ~n10958;
  assign y95 = n11078;
  assign y96 = ~n11196;
  assign y97 = ~n11290;
  assign y98 = ~n11389;
  assign y99 = ~n11486;
  assign y100 = n11575;
  assign y101 = ~n11672;
  assign y102 = n11756;
  assign y103 = n11841;
  assign y104 = n11918;
  assign y105 = n12002;
  assign y106 = n12082;
  assign y107 = n12147;
  assign y108 = n12212;
  assign y109 = n12276;
  assign y110 = n12334;
  assign y111 = ~n12403;
  assign y112 = n12462;
  assign y113 = n12515;
  assign y114 = n12566;
  assign y115 = ~n12614;
  assign y116 = ~n12659;
  assign y117 = n12712;
  assign y118 = ~n12772;
  assign y119 = ~n12808;
  assign y120 = n12843;
  assign y121 = n12871;
  assign y122 = ~n12886;
  assign y123 = n12914;
  assign y124 = n12932;
  assign y125 = n12949;
  assign y126 = ~n12957;
  assign y127 = n12958;
endmodule
