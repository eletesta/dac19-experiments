module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129;
  wire n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370;
  assign n514 = x127 & x255;
  assign n513 = x383 & x511;
  assign n515 = n514 ^ n513;
  assign n516 = ~x378 & x506;
  assign n517 = ~x377 & x505;
  assign n518 = ~n516 & ~n517;
  assign n519 = x377 & ~x505;
  assign n520 = x504 ^ x376;
  assign n521 = x503 ^ x375;
  assign n522 = ~x374 & x502;
  assign n523 = n522 ^ x503;
  assign n524 = n523 ^ x503;
  assign n525 = x374 & ~x502;
  assign n526 = x501 ^ x373;
  assign n527 = x500 ^ x372;
  assign n528 = ~x371 & x499;
  assign n529 = n528 ^ x500;
  assign n530 = n529 ^ x500;
  assign n531 = x369 & ~x497;
  assign n532 = x368 & ~x496;
  assign n533 = ~n531 & ~n532;
  assign n534 = ~x368 & x496;
  assign n535 = x495 ^ x367;
  assign n536 = x494 ^ x366;
  assign n537 = x365 & ~x493;
  assign n538 = n537 ^ x494;
  assign n539 = n538 ^ x494;
  assign n540 = ~x365 & x493;
  assign n541 = x492 ^ x364;
  assign n542 = x491 ^ x363;
  assign n543 = x362 & ~x490;
  assign n544 = n543 ^ x491;
  assign n545 = n544 ^ x491;
  assign n546 = ~x362 & x490;
  assign n547 = x489 ^ x361;
  assign n548 = ~x360 & x488;
  assign n549 = n548 ^ x489;
  assign n550 = n549 ^ x489;
  assign n551 = x360 & ~x488;
  assign n552 = x487 ^ x359;
  assign n553 = x358 & ~x486;
  assign n554 = n553 ^ x487;
  assign n555 = n554 ^ x487;
  assign n556 = x357 & ~x485;
  assign n557 = x356 & ~x484;
  assign n558 = ~n556 & ~n557;
  assign n559 = ~x356 & x484;
  assign n560 = x483 ^ x355;
  assign n561 = x482 ^ x354;
  assign n562 = x353 & ~x481;
  assign n563 = n562 ^ x482;
  assign n564 = n563 ^ x482;
  assign n565 = ~x351 & x479;
  assign n566 = ~x350 & x478;
  assign n567 = ~n565 & ~n566;
  assign n568 = x350 & ~x478;
  assign n569 = x477 ^ x349;
  assign n570 = x476 ^ x348;
  assign n571 = ~x347 & x475;
  assign n572 = n571 ^ x476;
  assign n573 = n572 ^ x476;
  assign n574 = x347 & ~x475;
  assign n575 = x474 ^ x346;
  assign n576 = x473 ^ x345;
  assign n577 = ~x344 & x472;
  assign n578 = n577 ^ x473;
  assign n579 = n578 ^ x473;
  assign n580 = x344 & ~x472;
  assign n581 = x471 ^ x343;
  assign n582 = x342 & ~x470;
  assign n583 = n582 ^ x471;
  assign n584 = n583 ^ x471;
  assign n585 = x341 & ~x469;
  assign n586 = x340 & ~x468;
  assign n587 = ~n585 & ~n586;
  assign n588 = ~x340 & x468;
  assign n589 = x467 ^ x339;
  assign n590 = x466 ^ x338;
  assign n591 = x337 & ~x465;
  assign n592 = n591 ^ x466;
  assign n593 = n592 ^ x466;
  assign n594 = ~x337 & x465;
  assign n595 = ~x336 & x464;
  assign n596 = ~n594 & ~n595;
  assign n597 = x336 & ~x464;
  assign n598 = x463 ^ x335;
  assign n599 = x462 ^ x334;
  assign n600 = ~x333 & x461;
  assign n601 = n600 ^ x462;
  assign n602 = n601 ^ x462;
  assign n603 = x333 & ~x461;
  assign n604 = x460 ^ x332;
  assign n605 = x459 ^ x331;
  assign n606 = ~x330 & x458;
  assign n607 = n606 ^ x459;
  assign n608 = n607 ^ x459;
  assign n609 = x330 & ~x458;
  assign n610 = x457 ^ x329;
  assign n611 = x456 ^ x328;
  assign n612 = ~x327 & x455;
  assign n613 = n612 ^ x456;
  assign n614 = n613 ^ x456;
  assign n615 = ~x325 & x453;
  assign n616 = ~x326 & x454;
  assign n617 = ~n615 & ~n616;
  assign n618 = ~x323 & x451;
  assign n619 = ~x324 & x452;
  assign n620 = ~n618 & ~n619;
  assign n621 = n617 & n620;
  assign n622 = x323 & ~x451;
  assign n623 = x450 ^ x322;
  assign n624 = x449 ^ x321;
  assign n625 = ~x320 & x448;
  assign n626 = n625 ^ x449;
  assign n627 = n626 ^ x449;
  assign n628 = x315 & ~x443;
  assign n629 = x442 ^ x314;
  assign n630 = x313 & ~x441;
  assign n631 = n630 ^ x442;
  assign n632 = n631 ^ x442;
  assign n633 = ~x311 & x439;
  assign n634 = ~x310 & x438;
  assign n635 = ~n633 & ~n634;
  assign n636 = x310 & ~x438;
  assign n637 = x437 ^ x309;
  assign n638 = x436 ^ x308;
  assign n639 = ~x307 & x435;
  assign n640 = n639 ^ x436;
  assign n641 = n640 ^ x436;
  assign n642 = ~x297 & x425;
  assign n643 = ~x298 & x426;
  assign n644 = ~n642 & ~n643;
  assign n645 = ~x295 & x423;
  assign n646 = ~x296 & x424;
  assign n647 = ~n645 & ~n646;
  assign n648 = n644 & n647;
  assign n649 = x295 & ~x423;
  assign n650 = x422 ^ x294;
  assign n651 = x421 ^ x293;
  assign n652 = ~x292 & x420;
  assign n653 = n652 ^ x421;
  assign n654 = n653 ^ x421;
  assign n655 = x292 & ~x420;
  assign n656 = x419 ^ x291;
  assign n657 = x290 & ~x418;
  assign n658 = n657 ^ x419;
  assign n659 = n658 ^ x419;
  assign n660 = x289 & ~x417;
  assign n661 = x288 & ~x416;
  assign n662 = ~n660 & ~n661;
  assign n663 = ~x288 & x416;
  assign n664 = x415 ^ x287;
  assign n665 = x414 ^ x286;
  assign n666 = x285 & ~x413;
  assign n667 = n666 ^ x414;
  assign n668 = n667 ^ x414;
  assign n669 = ~x285 & x413;
  assign n670 = ~x284 & x412;
  assign n671 = ~n669 & ~n670;
  assign n672 = x284 & ~x412;
  assign n673 = x411 ^ x283;
  assign n674 = x410 ^ x282;
  assign n675 = ~x281 & x409;
  assign n676 = n675 ^ x410;
  assign n677 = n676 ^ x410;
  assign n678 = x279 & ~x407;
  assign n679 = x278 & ~x406;
  assign n680 = ~n678 & ~n679;
  assign n681 = ~x278 & x406;
  assign n682 = x405 ^ x277;
  assign n683 = x404 ^ x276;
  assign n684 = x275 & ~x403;
  assign n685 = n684 ^ x404;
  assign n686 = n685 ^ x404;
  assign n687 = ~x275 & x403;
  assign n688 = x402 ^ x274;
  assign n689 = x401 ^ x273;
  assign n690 = x272 & ~x400;
  assign n691 = n690 ^ x401;
  assign n692 = n691 ^ x401;
  assign n693 = ~x272 & x400;
  assign n694 = x399 ^ x271;
  assign n695 = ~x270 & x398;
  assign n696 = n695 ^ x399;
  assign n697 = n696 ^ x399;
  assign n698 = x270 & ~x398;
  assign n699 = x397 ^ x269;
  assign n700 = x268 & ~x396;
  assign n701 = n700 ^ x397;
  assign n702 = n701 ^ x397;
  assign n703 = ~x268 & x396;
  assign n704 = x395 ^ x267;
  assign n705 = ~x266 & x394;
  assign n706 = n705 ^ x395;
  assign n707 = n706 ^ x395;
  assign n708 = ~x263 & x391;
  assign n709 = ~x262 & x390;
  assign n710 = ~n708 & ~n709;
  assign n711 = x262 & ~x390;
  assign n712 = x389 ^ x261;
  assign n713 = x388 ^ x260;
  assign n714 = ~x259 & x387;
  assign n715 = n714 ^ x388;
  assign n716 = n715 ^ x388;
  assign n717 = x259 & ~x387;
  assign n718 = x258 & ~x386;
  assign n719 = ~n717 & ~n718;
  assign n720 = ~x258 & x386;
  assign n721 = x385 ^ x257;
  assign n722 = x256 & ~x384;
  assign n723 = n722 ^ x385;
  assign n724 = ~n721 & ~n723;
  assign n725 = n724 ^ x385;
  assign n726 = ~n720 & ~n725;
  assign n727 = n719 & ~n726;
  assign n728 = n727 ^ x388;
  assign n729 = n728 ^ x388;
  assign n730 = ~n716 & ~n729;
  assign n731 = n730 ^ x388;
  assign n732 = ~n713 & n731;
  assign n733 = n732 ^ x260;
  assign n734 = n733 ^ x389;
  assign n735 = ~n712 & ~n734;
  assign n736 = n735 ^ x389;
  assign n737 = ~n711 & n736;
  assign n738 = n710 & ~n737;
  assign n739 = x264 & ~x392;
  assign n740 = x263 & ~x391;
  assign n741 = ~n739 & ~n740;
  assign n742 = ~n738 & n741;
  assign n743 = ~x265 & x393;
  assign n744 = ~x264 & x392;
  assign n745 = ~n743 & ~n744;
  assign n746 = ~n742 & n745;
  assign n747 = x266 & ~x394;
  assign n748 = x265 & ~x393;
  assign n749 = ~n747 & ~n748;
  assign n750 = ~n746 & n749;
  assign n751 = n750 ^ x395;
  assign n752 = n751 ^ x395;
  assign n753 = ~n707 & ~n752;
  assign n754 = n753 ^ x395;
  assign n755 = ~n704 & n754;
  assign n756 = n755 ^ x267;
  assign n757 = ~n703 & n756;
  assign n758 = n757 ^ x397;
  assign n759 = n758 ^ x397;
  assign n760 = ~n702 & ~n759;
  assign n761 = n760 ^ x397;
  assign n762 = ~n699 & ~n761;
  assign n763 = n762 ^ x269;
  assign n764 = ~n698 & ~n763;
  assign n765 = n764 ^ x399;
  assign n766 = n765 ^ x399;
  assign n767 = ~n697 & ~n766;
  assign n768 = n767 ^ x399;
  assign n769 = ~n694 & n768;
  assign n770 = n769 ^ x271;
  assign n771 = ~n693 & n770;
  assign n772 = n771 ^ x401;
  assign n773 = n772 ^ x401;
  assign n774 = ~n692 & ~n773;
  assign n775 = n774 ^ x401;
  assign n776 = ~n689 & ~n775;
  assign n777 = n776 ^ x273;
  assign n778 = n777 ^ x402;
  assign n779 = ~n688 & ~n778;
  assign n780 = n779 ^ x402;
  assign n781 = ~n687 & ~n780;
  assign n782 = n781 ^ x404;
  assign n783 = n782 ^ x404;
  assign n784 = ~n686 & ~n783;
  assign n785 = n784 ^ x404;
  assign n786 = ~n683 & ~n785;
  assign n787 = n786 ^ x276;
  assign n788 = n787 ^ x405;
  assign n789 = ~n682 & ~n788;
  assign n790 = n789 ^ x405;
  assign n791 = ~n681 & ~n790;
  assign n792 = n680 & ~n791;
  assign n793 = ~x280 & x408;
  assign n794 = ~x279 & x407;
  assign n795 = ~n793 & ~n794;
  assign n796 = ~n792 & n795;
  assign n797 = x281 & ~x409;
  assign n798 = x280 & ~x408;
  assign n799 = ~n797 & ~n798;
  assign n800 = ~n796 & n799;
  assign n801 = n800 ^ x410;
  assign n802 = n801 ^ x410;
  assign n803 = ~n677 & ~n802;
  assign n804 = n803 ^ x410;
  assign n805 = ~n674 & n804;
  assign n806 = n805 ^ x282;
  assign n807 = n806 ^ x411;
  assign n808 = ~n673 & ~n807;
  assign n809 = n808 ^ x411;
  assign n810 = ~n672 & n809;
  assign n811 = n671 & ~n810;
  assign n812 = n811 ^ x414;
  assign n813 = n812 ^ x414;
  assign n814 = ~n668 & ~n813;
  assign n815 = n814 ^ x414;
  assign n816 = ~n665 & ~n815;
  assign n817 = n816 ^ x286;
  assign n818 = n817 ^ x415;
  assign n819 = ~n664 & ~n818;
  assign n820 = n819 ^ x415;
  assign n821 = ~n663 & ~n820;
  assign n822 = n662 & ~n821;
  assign n823 = ~x290 & x418;
  assign n824 = ~x289 & x417;
  assign n825 = ~n823 & ~n824;
  assign n826 = ~n822 & n825;
  assign n827 = n826 ^ x419;
  assign n828 = n827 ^ x419;
  assign n829 = ~n659 & ~n828;
  assign n830 = n829 ^ x419;
  assign n831 = ~n656 & ~n830;
  assign n832 = n831 ^ x291;
  assign n833 = ~n655 & ~n832;
  assign n834 = n833 ^ x421;
  assign n835 = n834 ^ x421;
  assign n836 = ~n654 & ~n835;
  assign n837 = n836 ^ x421;
  assign n838 = ~n651 & n837;
  assign n839 = n838 ^ x293;
  assign n840 = n839 ^ x422;
  assign n841 = ~n650 & ~n840;
  assign n842 = n841 ^ x422;
  assign n843 = ~n649 & n842;
  assign n844 = n648 & ~n843;
  assign n845 = x299 & ~x427;
  assign n846 = x298 & ~x426;
  assign n847 = ~n845 & ~n846;
  assign n848 = x425 ^ x297;
  assign n849 = x296 & ~x424;
  assign n850 = n849 ^ x425;
  assign n851 = ~n848 & ~n850;
  assign n852 = n851 ^ x425;
  assign n853 = ~n643 & ~n852;
  assign n854 = n847 & ~n853;
  assign n855 = ~n844 & n854;
  assign n856 = ~x302 & x430;
  assign n857 = ~x301 & x429;
  assign n858 = ~n856 & ~n857;
  assign n859 = ~x299 & x427;
  assign n860 = ~x300 & x428;
  assign n861 = ~n859 & ~n860;
  assign n862 = n858 & n861;
  assign n863 = ~n855 & n862;
  assign n864 = x302 & ~x430;
  assign n865 = x303 & ~x431;
  assign n866 = ~n864 & ~n865;
  assign n867 = x429 ^ x301;
  assign n868 = x300 & ~x428;
  assign n869 = n868 ^ x429;
  assign n870 = ~n867 & ~n869;
  assign n871 = n870 ^ x429;
  assign n872 = ~n856 & ~n871;
  assign n873 = n866 & ~n872;
  assign n874 = ~n863 & n873;
  assign n875 = ~x304 & x432;
  assign n876 = ~x303 & x431;
  assign n877 = ~n875 & ~n876;
  assign n878 = ~n874 & n877;
  assign n879 = x305 & ~x433;
  assign n880 = x304 & ~x432;
  assign n881 = ~n879 & ~n880;
  assign n882 = ~n878 & n881;
  assign n883 = ~x306 & x434;
  assign n884 = ~x305 & x433;
  assign n885 = ~n883 & ~n884;
  assign n886 = ~n882 & n885;
  assign n887 = x307 & ~x435;
  assign n888 = x306 & ~x434;
  assign n889 = ~n887 & ~n888;
  assign n890 = ~n886 & n889;
  assign n891 = n890 ^ x436;
  assign n892 = n891 ^ x436;
  assign n893 = ~n641 & ~n892;
  assign n894 = n893 ^ x436;
  assign n895 = ~n638 & n894;
  assign n896 = n895 ^ x308;
  assign n897 = n896 ^ x437;
  assign n898 = ~n637 & ~n897;
  assign n899 = n898 ^ x437;
  assign n900 = ~n636 & n899;
  assign n901 = n635 & ~n900;
  assign n902 = x312 & ~x440;
  assign n903 = x311 & ~x439;
  assign n904 = ~n902 & ~n903;
  assign n905 = ~n901 & n904;
  assign n906 = ~x313 & x441;
  assign n907 = ~x312 & x440;
  assign n908 = ~n906 & ~n907;
  assign n909 = ~n905 & n908;
  assign n910 = n909 ^ x442;
  assign n911 = n910 ^ x442;
  assign n912 = ~n632 & ~n911;
  assign n913 = n912 ^ x442;
  assign n914 = ~n629 & ~n913;
  assign n915 = n914 ^ x314;
  assign n916 = ~n628 & ~n915;
  assign n917 = ~x315 & x443;
  assign n918 = ~x316 & x444;
  assign n919 = ~n917 & ~n918;
  assign n920 = ~x318 & x446;
  assign n921 = ~x317 & x445;
  assign n922 = ~n920 & ~n921;
  assign n923 = ~x319 & x447;
  assign n924 = n922 & ~n923;
  assign n925 = n919 & n924;
  assign n926 = ~n916 & n925;
  assign n927 = x317 & ~x445;
  assign n928 = x316 & ~x444;
  assign n929 = ~n927 & ~n928;
  assign n930 = n924 & ~n929;
  assign n931 = x320 & ~x448;
  assign n932 = x447 ^ x319;
  assign n933 = x318 & ~x446;
  assign n934 = n933 ^ x447;
  assign n935 = ~n932 & n934;
  assign n936 = n935 ^ x319;
  assign n937 = ~n931 & ~n936;
  assign n938 = ~n930 & n937;
  assign n939 = ~n926 & n938;
  assign n940 = n939 ^ x449;
  assign n941 = n940 ^ x449;
  assign n942 = ~n627 & ~n941;
  assign n943 = n942 ^ x449;
  assign n944 = ~n624 & n943;
  assign n945 = n944 ^ x321;
  assign n946 = n945 ^ x450;
  assign n947 = ~n623 & ~n946;
  assign n948 = n947 ^ x450;
  assign n949 = ~n622 & n948;
  assign n950 = n621 & ~n949;
  assign n951 = x327 & ~x455;
  assign n952 = x326 & ~x454;
  assign n953 = ~n951 & ~n952;
  assign n954 = x453 ^ x325;
  assign n955 = x324 & ~x452;
  assign n956 = n955 ^ x453;
  assign n957 = ~n954 & ~n956;
  assign n958 = n957 ^ x453;
  assign n959 = ~n616 & ~n958;
  assign n960 = n953 & ~n959;
  assign n961 = ~n950 & n960;
  assign n962 = n961 ^ x456;
  assign n963 = n962 ^ x456;
  assign n964 = ~n614 & ~n963;
  assign n965 = n964 ^ x456;
  assign n966 = ~n611 & n965;
  assign n967 = n966 ^ x328;
  assign n968 = n967 ^ x457;
  assign n969 = ~n610 & ~n968;
  assign n970 = n969 ^ x457;
  assign n971 = ~n609 & n970;
  assign n972 = n971 ^ x459;
  assign n973 = n972 ^ x459;
  assign n974 = ~n608 & ~n973;
  assign n975 = n974 ^ x459;
  assign n976 = ~n605 & n975;
  assign n977 = n976 ^ x331;
  assign n978 = n977 ^ x460;
  assign n979 = ~n604 & ~n978;
  assign n980 = n979 ^ x460;
  assign n981 = ~n603 & n980;
  assign n982 = n981 ^ x462;
  assign n983 = n982 ^ x462;
  assign n984 = ~n602 & ~n983;
  assign n985 = n984 ^ x462;
  assign n986 = ~n599 & n985;
  assign n987 = n986 ^ x334;
  assign n988 = n987 ^ x463;
  assign n989 = ~n598 & ~n988;
  assign n990 = n989 ^ x463;
  assign n991 = ~n597 & n990;
  assign n992 = n596 & ~n991;
  assign n993 = n992 ^ x466;
  assign n994 = n993 ^ x466;
  assign n995 = ~n593 & ~n994;
  assign n996 = n995 ^ x466;
  assign n997 = ~n590 & ~n996;
  assign n998 = n997 ^ x338;
  assign n999 = n998 ^ x467;
  assign n1000 = ~n589 & ~n999;
  assign n1001 = n1000 ^ x467;
  assign n1002 = ~n588 & ~n1001;
  assign n1003 = n587 & ~n1002;
  assign n1004 = ~x342 & x470;
  assign n1005 = ~x341 & x469;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = ~n1003 & n1006;
  assign n1008 = n1007 ^ x471;
  assign n1009 = n1008 ^ x471;
  assign n1010 = ~n584 & ~n1009;
  assign n1011 = n1010 ^ x471;
  assign n1012 = ~n581 & ~n1011;
  assign n1013 = n1012 ^ x343;
  assign n1014 = ~n580 & ~n1013;
  assign n1015 = n1014 ^ x473;
  assign n1016 = n1015 ^ x473;
  assign n1017 = ~n579 & ~n1016;
  assign n1018 = n1017 ^ x473;
  assign n1019 = ~n576 & n1018;
  assign n1020 = n1019 ^ x345;
  assign n1021 = n1020 ^ x474;
  assign n1022 = ~n575 & ~n1021;
  assign n1023 = n1022 ^ x474;
  assign n1024 = ~n574 & n1023;
  assign n1025 = n1024 ^ x476;
  assign n1026 = n1025 ^ x476;
  assign n1027 = ~n573 & ~n1026;
  assign n1028 = n1027 ^ x476;
  assign n1029 = ~n570 & n1028;
  assign n1030 = n1029 ^ x348;
  assign n1031 = n1030 ^ x477;
  assign n1032 = ~n569 & ~n1031;
  assign n1033 = n1032 ^ x477;
  assign n1034 = ~n568 & n1033;
  assign n1035 = n567 & ~n1034;
  assign n1036 = x352 & ~x480;
  assign n1037 = x351 & ~x479;
  assign n1038 = ~n1036 & ~n1037;
  assign n1039 = ~n1035 & n1038;
  assign n1040 = ~x353 & x481;
  assign n1041 = ~x352 & x480;
  assign n1042 = ~n1040 & ~n1041;
  assign n1043 = ~n1039 & n1042;
  assign n1044 = n1043 ^ x482;
  assign n1045 = n1044 ^ x482;
  assign n1046 = ~n564 & ~n1045;
  assign n1047 = n1046 ^ x482;
  assign n1048 = ~n561 & ~n1047;
  assign n1049 = n1048 ^ x354;
  assign n1050 = n1049 ^ x483;
  assign n1051 = ~n560 & ~n1050;
  assign n1052 = n1051 ^ x483;
  assign n1053 = ~n559 & ~n1052;
  assign n1054 = n558 & ~n1053;
  assign n1055 = ~x358 & x486;
  assign n1056 = ~x357 & x485;
  assign n1057 = ~n1055 & ~n1056;
  assign n1058 = ~n1054 & n1057;
  assign n1059 = n1058 ^ x487;
  assign n1060 = n1059 ^ x487;
  assign n1061 = ~n555 & ~n1060;
  assign n1062 = n1061 ^ x487;
  assign n1063 = ~n552 & ~n1062;
  assign n1064 = n1063 ^ x359;
  assign n1065 = ~n551 & ~n1064;
  assign n1066 = n1065 ^ x489;
  assign n1067 = n1066 ^ x489;
  assign n1068 = ~n550 & ~n1067;
  assign n1069 = n1068 ^ x489;
  assign n1070 = ~n547 & n1069;
  assign n1071 = n1070 ^ x361;
  assign n1072 = ~n546 & n1071;
  assign n1073 = n1072 ^ x491;
  assign n1074 = n1073 ^ x491;
  assign n1075 = ~n545 & ~n1074;
  assign n1076 = n1075 ^ x491;
  assign n1077 = ~n542 & ~n1076;
  assign n1078 = n1077 ^ x363;
  assign n1079 = n1078 ^ x492;
  assign n1080 = ~n541 & ~n1079;
  assign n1081 = n1080 ^ x492;
  assign n1082 = ~n540 & ~n1081;
  assign n1083 = n1082 ^ x494;
  assign n1084 = n1083 ^ x494;
  assign n1085 = ~n539 & ~n1084;
  assign n1086 = n1085 ^ x494;
  assign n1087 = ~n536 & ~n1086;
  assign n1088 = n1087 ^ x366;
  assign n1089 = n1088 ^ x495;
  assign n1090 = ~n535 & ~n1089;
  assign n1091 = n1090 ^ x495;
  assign n1092 = ~n534 & ~n1091;
  assign n1093 = n533 & ~n1092;
  assign n1094 = ~x370 & x498;
  assign n1095 = ~x369 & x497;
  assign n1096 = ~n1094 & ~n1095;
  assign n1097 = ~n1093 & n1096;
  assign n1098 = x371 & ~x499;
  assign n1099 = x370 & ~x498;
  assign n1100 = ~n1098 & ~n1099;
  assign n1101 = ~n1097 & n1100;
  assign n1102 = n1101 ^ x500;
  assign n1103 = n1102 ^ x500;
  assign n1104 = ~n530 & ~n1103;
  assign n1105 = n1104 ^ x500;
  assign n1106 = ~n527 & n1105;
  assign n1107 = n1106 ^ x372;
  assign n1108 = n1107 ^ x501;
  assign n1109 = ~n526 & ~n1108;
  assign n1110 = n1109 ^ x501;
  assign n1111 = ~n525 & n1110;
  assign n1112 = n1111 ^ x503;
  assign n1113 = n1112 ^ x503;
  assign n1114 = ~n524 & ~n1113;
  assign n1115 = n1114 ^ x503;
  assign n1116 = ~n521 & n1115;
  assign n1117 = n1116 ^ x375;
  assign n1118 = n1117 ^ x504;
  assign n1119 = ~n520 & ~n1118;
  assign n1120 = n1119 ^ x504;
  assign n1121 = ~n519 & n1120;
  assign n1122 = n518 & ~n1121;
  assign n1123 = x379 & ~x507;
  assign n1124 = x378 & ~x506;
  assign n1125 = ~n1123 & ~n1124;
  assign n1126 = ~n1122 & n1125;
  assign n1127 = ~x381 & x509;
  assign n1128 = ~x382 & x510;
  assign n1129 = ~n1127 & ~n1128;
  assign n1130 = ~x379 & x507;
  assign n1131 = ~x380 & x508;
  assign n1132 = ~n1130 & ~n1131;
  assign n1133 = n1129 & n1132;
  assign n1134 = ~n1126 & n1133;
  assign n1135 = ~x383 & x511;
  assign n1136 = x382 & ~x510;
  assign n1137 = ~n1135 & ~n1136;
  assign n1138 = x509 ^ x381;
  assign n1139 = x380 & ~x508;
  assign n1140 = n1139 ^ x509;
  assign n1141 = ~n1138 & ~n1140;
  assign n1142 = n1141 ^ x509;
  assign n1143 = ~n1128 & ~n1142;
  assign n1144 = n1137 & ~n1143;
  assign n1145 = ~n1134 & n1144;
  assign n1146 = x383 & ~x511;
  assign n1147 = ~n1145 & ~n1146;
  assign n1148 = x510 ^ x382;
  assign n1149 = ~n1147 & n1148;
  assign n1150 = n1149 ^ x382;
  assign n1151 = ~x125 & x253;
  assign n1152 = ~x126 & x254;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = ~x123 & x251;
  assign n1155 = ~x124 & x252;
  assign n1156 = ~n1154 & ~n1155;
  assign n1157 = n1153 & n1156;
  assign n1158 = x123 & ~x251;
  assign n1159 = x250 ^ x122;
  assign n1160 = x249 ^ x121;
  assign n1161 = ~x120 & x248;
  assign n1162 = n1161 ^ x249;
  assign n1163 = n1162 ^ x249;
  assign n1164 = x120 & ~x248;
  assign n1165 = x247 ^ x119;
  assign n1166 = x118 & ~x246;
  assign n1167 = n1166 ^ x247;
  assign n1168 = n1167 ^ x247;
  assign n1169 = ~x118 & x246;
  assign n1170 = x245 ^ x117;
  assign n1171 = x244 ^ x116;
  assign n1172 = x115 & ~x243;
  assign n1173 = n1172 ^ x244;
  assign n1174 = n1173 ^ x244;
  assign n1175 = ~x115 & x243;
  assign n1176 = x242 ^ x114;
  assign n1177 = x241 ^ x113;
  assign n1178 = x112 & ~x240;
  assign n1179 = n1178 ^ x241;
  assign n1180 = n1179 ^ x241;
  assign n1181 = ~x112 & x240;
  assign n1182 = ~x111 & x239;
  assign n1183 = ~n1181 & ~n1182;
  assign n1184 = x111 & ~x239;
  assign n1185 = x238 ^ x110;
  assign n1186 = x237 ^ x109;
  assign n1187 = ~x108 & x236;
  assign n1188 = n1187 ^ x237;
  assign n1189 = n1188 ^ x237;
  assign n1190 = x108 & ~x236;
  assign n1191 = x107 & ~x235;
  assign n1192 = ~n1190 & ~n1191;
  assign n1193 = ~x107 & x235;
  assign n1194 = x234 ^ x106;
  assign n1195 = x233 ^ x105;
  assign n1196 = x104 & ~x232;
  assign n1197 = n1196 ^ x233;
  assign n1198 = n1197 ^ x233;
  assign n1199 = ~x104 & x232;
  assign n1200 = ~x103 & x231;
  assign n1201 = ~n1199 & ~n1200;
  assign n1202 = x103 & ~x231;
  assign n1203 = x230 ^ x102;
  assign n1204 = x229 ^ x101;
  assign n1205 = ~x100 & x228;
  assign n1206 = n1205 ^ x229;
  assign n1207 = n1206 ^ x229;
  assign n1208 = x100 & ~x228;
  assign n1209 = x99 & ~x227;
  assign n1210 = ~n1208 & ~n1209;
  assign n1211 = ~x99 & x227;
  assign n1212 = x226 ^ x98;
  assign n1213 = x225 ^ x97;
  assign n1214 = x96 & ~x224;
  assign n1215 = n1214 ^ x225;
  assign n1216 = n1215 ^ x225;
  assign n1217 = ~x96 & x224;
  assign n1218 = x223 ^ x95;
  assign n1219 = x222 ^ x94;
  assign n1220 = x93 & ~x221;
  assign n1221 = n1220 ^ x222;
  assign n1222 = n1221 ^ x222;
  assign n1223 = ~x93 & x221;
  assign n1224 = x220 ^ x92;
  assign n1225 = ~x91 & x219;
  assign n1226 = n1225 ^ x220;
  assign n1227 = n1226 ^ x220;
  assign n1228 = x91 & ~x219;
  assign n1229 = x218 ^ x90;
  assign n1230 = x89 & ~x217;
  assign n1231 = n1230 ^ x218;
  assign n1232 = n1231 ^ x218;
  assign n1233 = x84 & ~x212;
  assign n1234 = x83 & ~x211;
  assign n1235 = ~n1233 & ~n1234;
  assign n1236 = ~x83 & x211;
  assign n1237 = x210 ^ x82;
  assign n1238 = x209 ^ x81;
  assign n1239 = x80 & ~x208;
  assign n1240 = n1239 ^ x209;
  assign n1241 = n1240 ^ x209;
  assign n1242 = ~x70 & x198;
  assign n1243 = ~x69 & x197;
  assign n1244 = ~n1242 & ~n1243;
  assign n1245 = ~x68 & x196;
  assign n1246 = n1244 & ~n1245;
  assign n1247 = x195 ^ x67;
  assign n1248 = ~x66 & x194;
  assign n1249 = n1248 ^ x195;
  assign n1250 = n1249 ^ x195;
  assign n1251 = x66 & ~x194;
  assign n1252 = x193 ^ x65;
  assign n1253 = x192 ^ x64;
  assign n1254 = ~x63 & x191;
  assign n1255 = n1254 ^ x192;
  assign n1256 = n1255 ^ x192;
  assign n1257 = x59 & ~x187;
  assign n1258 = x58 & ~x186;
  assign n1259 = ~n1257 & ~n1258;
  assign n1260 = ~x58 & x186;
  assign n1261 = x185 ^ x57;
  assign n1262 = x184 ^ x56;
  assign n1263 = x55 & ~x183;
  assign n1264 = n1263 ^ x184;
  assign n1265 = n1264 ^ x184;
  assign n1266 = x52 & ~x180;
  assign n1267 = x51 & ~x179;
  assign n1268 = ~n1266 & ~n1267;
  assign n1269 = ~x51 & x179;
  assign n1270 = x178 ^ x50;
  assign n1271 = x177 ^ x49;
  assign n1272 = x48 & ~x176;
  assign n1273 = n1272 ^ x177;
  assign n1274 = n1273 ^ x177;
  assign n1275 = x39 & ~x167;
  assign n1276 = x166 ^ x38;
  assign n1277 = x37 & ~x165;
  assign n1278 = n1277 ^ x166;
  assign n1279 = n1278 ^ x166;
  assign n1280 = ~x35 & x163;
  assign n1281 = ~x34 & x162;
  assign n1282 = ~n1280 & ~n1281;
  assign n1283 = x34 & ~x162;
  assign n1284 = x161 ^ x33;
  assign n1285 = x160 ^ x32;
  assign n1286 = ~x31 & x159;
  assign n1287 = n1286 ^ x160;
  assign n1288 = n1287 ^ x160;
  assign n1289 = x31 & ~x159;
  assign n1290 = x158 ^ x30;
  assign n1291 = x157 ^ x29;
  assign n1292 = ~x28 & x156;
  assign n1293 = n1292 ^ x157;
  assign n1294 = n1293 ^ x157;
  assign n1295 = x28 & ~x156;
  assign n1296 = x155 ^ x27;
  assign n1297 = x154 ^ x26;
  assign n1298 = ~x25 & x153;
  assign n1299 = n1298 ^ x154;
  assign n1300 = n1299 ^ x154;
  assign n1301 = x21 & ~x149;
  assign n1302 = x20 & ~x148;
  assign n1303 = ~n1301 & ~n1302;
  assign n1304 = ~x20 & x148;
  assign n1305 = x147 ^ x19;
  assign n1306 = x146 ^ x18;
  assign n1307 = x17 & ~x145;
  assign n1308 = n1307 ^ x146;
  assign n1309 = n1308 ^ x146;
  assign n1310 = ~x17 & x145;
  assign n1311 = x144 ^ x16;
  assign n1312 = x143 ^ x15;
  assign n1313 = x14 & ~x142;
  assign n1314 = n1313 ^ x143;
  assign n1315 = n1314 ^ x143;
  assign n1316 = ~x14 & x142;
  assign n1317 = x141 ^ x13;
  assign n1318 = ~x12 & x140;
  assign n1319 = n1318 ^ x141;
  assign n1320 = n1319 ^ x141;
  assign n1321 = x12 & ~x140;
  assign n1322 = x139 ^ x11;
  assign n1323 = x10 & ~x138;
  assign n1324 = n1323 ^ x139;
  assign n1325 = n1324 ^ x139;
  assign n1326 = ~x10 & x138;
  assign n1327 = x137 ^ x9;
  assign n1328 = x136 ^ x8;
  assign n1329 = x7 & ~x135;
  assign n1330 = n1329 ^ x136;
  assign n1331 = n1330 ^ x136;
  assign n1332 = ~x7 & x135;
  assign n1333 = x134 ^ x6;
  assign n1334 = x133 ^ x5;
  assign n1335 = x4 & ~x132;
  assign n1336 = n1335 ^ x133;
  assign n1337 = n1336 ^ x133;
  assign n1338 = x3 & ~x131;
  assign n1339 = x2 & ~x130;
  assign n1340 = ~n1338 & ~n1339;
  assign n1341 = ~x2 & x130;
  assign n1342 = x129 ^ x1;
  assign n1343 = x0 & ~x128;
  assign n1344 = n1343 ^ x129;
  assign n1345 = ~n1342 & ~n1344;
  assign n1346 = n1345 ^ x129;
  assign n1347 = ~n1341 & ~n1346;
  assign n1348 = n1340 & ~n1347;
  assign n1349 = ~x4 & x132;
  assign n1350 = ~x3 & x131;
  assign n1351 = ~n1349 & ~n1350;
  assign n1352 = ~n1348 & n1351;
  assign n1353 = n1352 ^ x133;
  assign n1354 = n1353 ^ x133;
  assign n1355 = ~n1337 & ~n1354;
  assign n1356 = n1355 ^ x133;
  assign n1357 = ~n1334 & ~n1356;
  assign n1358 = n1357 ^ x5;
  assign n1359 = n1358 ^ x134;
  assign n1360 = ~n1333 & ~n1359;
  assign n1361 = n1360 ^ x134;
  assign n1362 = ~n1332 & ~n1361;
  assign n1363 = n1362 ^ x136;
  assign n1364 = n1363 ^ x136;
  assign n1365 = ~n1331 & ~n1364;
  assign n1366 = n1365 ^ x136;
  assign n1367 = ~n1328 & ~n1366;
  assign n1368 = n1367 ^ x8;
  assign n1369 = n1368 ^ x137;
  assign n1370 = ~n1327 & ~n1369;
  assign n1371 = n1370 ^ x137;
  assign n1372 = ~n1326 & ~n1371;
  assign n1373 = n1372 ^ x139;
  assign n1374 = n1373 ^ x139;
  assign n1375 = ~n1325 & ~n1374;
  assign n1376 = n1375 ^ x139;
  assign n1377 = ~n1322 & ~n1376;
  assign n1378 = n1377 ^ x11;
  assign n1379 = ~n1321 & ~n1378;
  assign n1380 = n1379 ^ x141;
  assign n1381 = n1380 ^ x141;
  assign n1382 = ~n1320 & ~n1381;
  assign n1383 = n1382 ^ x141;
  assign n1384 = ~n1317 & n1383;
  assign n1385 = n1384 ^ x13;
  assign n1386 = ~n1316 & n1385;
  assign n1387 = n1386 ^ x143;
  assign n1388 = n1387 ^ x143;
  assign n1389 = ~n1315 & ~n1388;
  assign n1390 = n1389 ^ x143;
  assign n1391 = ~n1312 & ~n1390;
  assign n1392 = n1391 ^ x15;
  assign n1393 = n1392 ^ x144;
  assign n1394 = ~n1311 & ~n1393;
  assign n1395 = n1394 ^ x144;
  assign n1396 = ~n1310 & ~n1395;
  assign n1397 = n1396 ^ x146;
  assign n1398 = n1397 ^ x146;
  assign n1399 = ~n1309 & ~n1398;
  assign n1400 = n1399 ^ x146;
  assign n1401 = ~n1306 & ~n1400;
  assign n1402 = n1401 ^ x18;
  assign n1403 = n1402 ^ x147;
  assign n1404 = ~n1305 & ~n1403;
  assign n1405 = n1404 ^ x147;
  assign n1406 = ~n1304 & ~n1405;
  assign n1407 = n1303 & ~n1406;
  assign n1408 = ~x22 & x150;
  assign n1409 = ~x21 & x149;
  assign n1410 = ~n1408 & ~n1409;
  assign n1411 = ~n1407 & n1410;
  assign n1412 = x23 & ~x151;
  assign n1413 = x22 & ~x150;
  assign n1414 = ~n1412 & ~n1413;
  assign n1415 = ~n1411 & n1414;
  assign n1416 = ~x24 & x152;
  assign n1417 = ~x23 & x151;
  assign n1418 = ~n1416 & ~n1417;
  assign n1419 = ~n1415 & n1418;
  assign n1420 = x25 & ~x153;
  assign n1421 = x24 & ~x152;
  assign n1422 = ~n1420 & ~n1421;
  assign n1423 = ~n1419 & n1422;
  assign n1424 = n1423 ^ x154;
  assign n1425 = n1424 ^ x154;
  assign n1426 = ~n1300 & ~n1425;
  assign n1427 = n1426 ^ x154;
  assign n1428 = ~n1297 & n1427;
  assign n1429 = n1428 ^ x26;
  assign n1430 = n1429 ^ x155;
  assign n1431 = ~n1296 & ~n1430;
  assign n1432 = n1431 ^ x155;
  assign n1433 = ~n1295 & n1432;
  assign n1434 = n1433 ^ x157;
  assign n1435 = n1434 ^ x157;
  assign n1436 = ~n1294 & ~n1435;
  assign n1437 = n1436 ^ x157;
  assign n1438 = ~n1291 & n1437;
  assign n1439 = n1438 ^ x29;
  assign n1440 = n1439 ^ x158;
  assign n1441 = ~n1290 & ~n1440;
  assign n1442 = n1441 ^ x158;
  assign n1443 = ~n1289 & n1442;
  assign n1444 = n1443 ^ x160;
  assign n1445 = n1444 ^ x160;
  assign n1446 = ~n1288 & ~n1445;
  assign n1447 = n1446 ^ x160;
  assign n1448 = ~n1285 & n1447;
  assign n1449 = n1448 ^ x32;
  assign n1450 = n1449 ^ x161;
  assign n1451 = ~n1284 & ~n1450;
  assign n1452 = n1451 ^ x161;
  assign n1453 = ~n1283 & n1452;
  assign n1454 = n1282 & ~n1453;
  assign n1455 = x36 & ~x164;
  assign n1456 = x35 & ~x163;
  assign n1457 = ~n1455 & ~n1456;
  assign n1458 = ~n1454 & n1457;
  assign n1459 = ~x37 & x165;
  assign n1460 = ~x36 & x164;
  assign n1461 = ~n1459 & ~n1460;
  assign n1462 = ~n1458 & n1461;
  assign n1463 = n1462 ^ x166;
  assign n1464 = n1463 ^ x166;
  assign n1465 = ~n1279 & ~n1464;
  assign n1466 = n1465 ^ x166;
  assign n1467 = ~n1276 & ~n1466;
  assign n1468 = n1467 ^ x38;
  assign n1469 = ~n1275 & ~n1468;
  assign n1470 = ~x41 & x169;
  assign n1471 = ~x42 & x170;
  assign n1472 = ~n1470 & ~n1471;
  assign n1473 = ~x39 & x167;
  assign n1474 = ~x40 & x168;
  assign n1475 = ~n1473 & ~n1474;
  assign n1476 = n1472 & n1475;
  assign n1477 = ~n1469 & n1476;
  assign n1478 = x43 & ~x171;
  assign n1479 = x42 & ~x170;
  assign n1480 = ~n1478 & ~n1479;
  assign n1481 = x169 ^ x41;
  assign n1482 = x40 & ~x168;
  assign n1483 = n1482 ^ x169;
  assign n1484 = ~n1481 & ~n1483;
  assign n1485 = n1484 ^ x169;
  assign n1486 = ~n1471 & ~n1485;
  assign n1487 = n1480 & ~n1486;
  assign n1488 = ~n1477 & n1487;
  assign n1489 = ~x46 & x174;
  assign n1490 = ~x45 & x173;
  assign n1491 = ~n1489 & ~n1490;
  assign n1492 = ~x43 & x171;
  assign n1493 = ~x44 & x172;
  assign n1494 = ~n1492 & ~n1493;
  assign n1495 = n1491 & n1494;
  assign n1496 = ~n1488 & n1495;
  assign n1497 = x46 & ~x174;
  assign n1498 = x47 & ~x175;
  assign n1499 = ~n1497 & ~n1498;
  assign n1500 = x173 ^ x45;
  assign n1501 = x44 & ~x172;
  assign n1502 = n1501 ^ x173;
  assign n1503 = ~n1500 & ~n1502;
  assign n1504 = n1503 ^ x173;
  assign n1505 = ~n1489 & ~n1504;
  assign n1506 = n1499 & ~n1505;
  assign n1507 = ~n1496 & n1506;
  assign n1508 = ~x48 & x176;
  assign n1509 = ~x47 & x175;
  assign n1510 = ~n1508 & ~n1509;
  assign n1511 = ~n1507 & n1510;
  assign n1512 = n1511 ^ x177;
  assign n1513 = n1512 ^ x177;
  assign n1514 = ~n1274 & ~n1513;
  assign n1515 = n1514 ^ x177;
  assign n1516 = ~n1271 & ~n1515;
  assign n1517 = n1516 ^ x49;
  assign n1518 = n1517 ^ x178;
  assign n1519 = ~n1270 & ~n1518;
  assign n1520 = n1519 ^ x178;
  assign n1521 = ~n1269 & ~n1520;
  assign n1522 = n1268 & ~n1521;
  assign n1523 = ~x53 & x181;
  assign n1524 = ~x52 & x180;
  assign n1525 = ~n1523 & ~n1524;
  assign n1526 = ~n1522 & n1525;
  assign n1527 = x54 & ~x182;
  assign n1528 = x53 & ~x181;
  assign n1529 = ~n1527 & ~n1528;
  assign n1530 = ~n1526 & n1529;
  assign n1531 = ~x55 & x183;
  assign n1532 = ~x54 & x182;
  assign n1533 = ~n1531 & ~n1532;
  assign n1534 = ~n1530 & n1533;
  assign n1535 = n1534 ^ x184;
  assign n1536 = n1535 ^ x184;
  assign n1537 = ~n1265 & ~n1536;
  assign n1538 = n1537 ^ x184;
  assign n1539 = ~n1262 & ~n1538;
  assign n1540 = n1539 ^ x56;
  assign n1541 = n1540 ^ x185;
  assign n1542 = ~n1261 & ~n1541;
  assign n1543 = n1542 ^ x185;
  assign n1544 = ~n1260 & ~n1543;
  assign n1545 = n1259 & ~n1544;
  assign n1546 = ~x62 & x190;
  assign n1547 = ~x61 & x189;
  assign n1548 = ~n1546 & ~n1547;
  assign n1549 = ~x59 & x187;
  assign n1550 = ~x60 & x188;
  assign n1551 = ~n1549 & ~n1550;
  assign n1552 = n1548 & n1551;
  assign n1553 = ~n1545 & n1552;
  assign n1554 = x63 & ~x191;
  assign n1555 = x62 & ~x190;
  assign n1556 = ~n1554 & ~n1555;
  assign n1557 = x189 ^ x61;
  assign n1558 = x60 & ~x188;
  assign n1559 = n1558 ^ x189;
  assign n1560 = ~n1557 & ~n1559;
  assign n1561 = n1560 ^ x189;
  assign n1562 = ~n1546 & ~n1561;
  assign n1563 = n1556 & ~n1562;
  assign n1564 = ~n1553 & n1563;
  assign n1565 = n1564 ^ x192;
  assign n1566 = n1565 ^ x192;
  assign n1567 = ~n1256 & ~n1566;
  assign n1568 = n1567 ^ x192;
  assign n1569 = ~n1253 & n1568;
  assign n1570 = n1569 ^ x64;
  assign n1571 = n1570 ^ x193;
  assign n1572 = ~n1252 & ~n1571;
  assign n1573 = n1572 ^ x193;
  assign n1574 = ~n1251 & n1573;
  assign n1575 = n1574 ^ x195;
  assign n1576 = n1575 ^ x195;
  assign n1577 = ~n1250 & ~n1576;
  assign n1578 = n1577 ^ x195;
  assign n1579 = ~n1247 & n1578;
  assign n1580 = n1579 ^ x67;
  assign n1581 = n1246 & n1580;
  assign n1582 = x70 & ~x198;
  assign n1583 = x71 & ~x199;
  assign n1584 = ~n1582 & ~n1583;
  assign n1585 = x197 ^ x69;
  assign n1586 = x68 & ~x196;
  assign n1587 = n1586 ^ x197;
  assign n1588 = ~n1585 & ~n1587;
  assign n1589 = n1588 ^ x197;
  assign n1590 = ~n1242 & ~n1589;
  assign n1591 = n1584 & ~n1590;
  assign n1592 = ~n1581 & n1591;
  assign n1593 = ~x72 & x200;
  assign n1594 = ~x71 & x199;
  assign n1595 = ~n1593 & ~n1594;
  assign n1596 = ~n1592 & n1595;
  assign n1597 = x73 & ~x201;
  assign n1598 = x72 & ~x200;
  assign n1599 = ~n1597 & ~n1598;
  assign n1600 = ~n1596 & n1599;
  assign n1601 = ~x74 & x202;
  assign n1602 = ~x73 & x201;
  assign n1603 = ~n1601 & ~n1602;
  assign n1604 = ~n1600 & n1603;
  assign n1605 = x75 & ~x203;
  assign n1606 = x74 & ~x202;
  assign n1607 = ~n1605 & ~n1606;
  assign n1608 = ~n1604 & n1607;
  assign n1609 = ~x76 & x204;
  assign n1610 = ~x75 & x203;
  assign n1611 = ~n1609 & ~n1610;
  assign n1612 = ~n1608 & n1611;
  assign n1613 = x77 & ~x205;
  assign n1614 = x76 & ~x204;
  assign n1615 = ~n1613 & ~n1614;
  assign n1616 = ~n1612 & n1615;
  assign n1617 = ~x78 & x206;
  assign n1618 = ~x77 & x205;
  assign n1619 = ~n1617 & ~n1618;
  assign n1620 = ~n1616 & n1619;
  assign n1621 = x79 & ~x207;
  assign n1622 = x78 & ~x206;
  assign n1623 = ~n1621 & ~n1622;
  assign n1624 = ~n1620 & n1623;
  assign n1625 = ~x80 & x208;
  assign n1626 = ~x79 & x207;
  assign n1627 = ~n1625 & ~n1626;
  assign n1628 = ~n1624 & n1627;
  assign n1629 = n1628 ^ x209;
  assign n1630 = n1629 ^ x209;
  assign n1631 = ~n1241 & ~n1630;
  assign n1632 = n1631 ^ x209;
  assign n1633 = ~n1238 & ~n1632;
  assign n1634 = n1633 ^ x81;
  assign n1635 = n1634 ^ x210;
  assign n1636 = ~n1237 & ~n1635;
  assign n1637 = n1636 ^ x210;
  assign n1638 = ~n1236 & ~n1637;
  assign n1639 = n1235 & ~n1638;
  assign n1640 = ~x85 & x213;
  assign n1641 = ~x84 & x212;
  assign n1642 = ~n1640 & ~n1641;
  assign n1643 = ~n1639 & n1642;
  assign n1644 = x86 & ~x214;
  assign n1645 = x85 & ~x213;
  assign n1646 = ~n1644 & ~n1645;
  assign n1647 = ~n1643 & n1646;
  assign n1648 = ~x87 & x215;
  assign n1649 = ~x86 & x214;
  assign n1650 = ~n1648 & ~n1649;
  assign n1651 = ~n1647 & n1650;
  assign n1652 = x88 & ~x216;
  assign n1653 = x87 & ~x215;
  assign n1654 = ~n1652 & ~n1653;
  assign n1655 = ~n1651 & n1654;
  assign n1656 = ~x89 & x217;
  assign n1657 = ~x88 & x216;
  assign n1658 = ~n1656 & ~n1657;
  assign n1659 = ~n1655 & n1658;
  assign n1660 = n1659 ^ x218;
  assign n1661 = n1660 ^ x218;
  assign n1662 = ~n1232 & ~n1661;
  assign n1663 = n1662 ^ x218;
  assign n1664 = ~n1229 & ~n1663;
  assign n1665 = n1664 ^ x90;
  assign n1666 = ~n1228 & ~n1665;
  assign n1667 = n1666 ^ x220;
  assign n1668 = n1667 ^ x220;
  assign n1669 = ~n1227 & ~n1668;
  assign n1670 = n1669 ^ x220;
  assign n1671 = ~n1224 & n1670;
  assign n1672 = n1671 ^ x92;
  assign n1673 = ~n1223 & n1672;
  assign n1674 = n1673 ^ x222;
  assign n1675 = n1674 ^ x222;
  assign n1676 = ~n1222 & ~n1675;
  assign n1677 = n1676 ^ x222;
  assign n1678 = ~n1219 & ~n1677;
  assign n1679 = n1678 ^ x94;
  assign n1680 = n1679 ^ x223;
  assign n1681 = ~n1218 & ~n1680;
  assign n1682 = n1681 ^ x223;
  assign n1683 = ~n1217 & ~n1682;
  assign n1684 = n1683 ^ x225;
  assign n1685 = n1684 ^ x225;
  assign n1686 = ~n1216 & ~n1685;
  assign n1687 = n1686 ^ x225;
  assign n1688 = ~n1213 & ~n1687;
  assign n1689 = n1688 ^ x97;
  assign n1690 = n1689 ^ x226;
  assign n1691 = ~n1212 & ~n1690;
  assign n1692 = n1691 ^ x226;
  assign n1693 = ~n1211 & ~n1692;
  assign n1694 = n1210 & ~n1693;
  assign n1695 = n1694 ^ x229;
  assign n1696 = n1695 ^ x229;
  assign n1697 = ~n1207 & ~n1696;
  assign n1698 = n1697 ^ x229;
  assign n1699 = ~n1204 & n1698;
  assign n1700 = n1699 ^ x101;
  assign n1701 = n1700 ^ x230;
  assign n1702 = ~n1203 & ~n1701;
  assign n1703 = n1702 ^ x230;
  assign n1704 = ~n1202 & n1703;
  assign n1705 = n1201 & ~n1704;
  assign n1706 = n1705 ^ x233;
  assign n1707 = n1706 ^ x233;
  assign n1708 = ~n1198 & ~n1707;
  assign n1709 = n1708 ^ x233;
  assign n1710 = ~n1195 & ~n1709;
  assign n1711 = n1710 ^ x105;
  assign n1712 = n1711 ^ x234;
  assign n1713 = ~n1194 & ~n1712;
  assign n1714 = n1713 ^ x234;
  assign n1715 = ~n1193 & ~n1714;
  assign n1716 = n1192 & ~n1715;
  assign n1717 = n1716 ^ x237;
  assign n1718 = n1717 ^ x237;
  assign n1719 = ~n1189 & ~n1718;
  assign n1720 = n1719 ^ x237;
  assign n1721 = ~n1186 & n1720;
  assign n1722 = n1721 ^ x109;
  assign n1723 = n1722 ^ x238;
  assign n1724 = ~n1185 & ~n1723;
  assign n1725 = n1724 ^ x238;
  assign n1726 = ~n1184 & n1725;
  assign n1727 = n1183 & ~n1726;
  assign n1728 = n1727 ^ x241;
  assign n1729 = n1728 ^ x241;
  assign n1730 = ~n1180 & ~n1729;
  assign n1731 = n1730 ^ x241;
  assign n1732 = ~n1177 & ~n1731;
  assign n1733 = n1732 ^ x113;
  assign n1734 = n1733 ^ x242;
  assign n1735 = ~n1176 & ~n1734;
  assign n1736 = n1735 ^ x242;
  assign n1737 = ~n1175 & ~n1736;
  assign n1738 = n1737 ^ x244;
  assign n1739 = n1738 ^ x244;
  assign n1740 = ~n1174 & ~n1739;
  assign n1741 = n1740 ^ x244;
  assign n1742 = ~n1171 & ~n1741;
  assign n1743 = n1742 ^ x116;
  assign n1744 = n1743 ^ x245;
  assign n1745 = ~n1170 & ~n1744;
  assign n1746 = n1745 ^ x245;
  assign n1747 = ~n1169 & ~n1746;
  assign n1748 = n1747 ^ x247;
  assign n1749 = n1748 ^ x247;
  assign n1750 = ~n1168 & ~n1749;
  assign n1751 = n1750 ^ x247;
  assign n1752 = ~n1165 & ~n1751;
  assign n1753 = n1752 ^ x119;
  assign n1754 = ~n1164 & ~n1753;
  assign n1755 = n1754 ^ x249;
  assign n1756 = n1755 ^ x249;
  assign n1757 = ~n1163 & ~n1756;
  assign n1758 = n1757 ^ x249;
  assign n1759 = ~n1160 & n1758;
  assign n1760 = n1759 ^ x121;
  assign n1761 = n1760 ^ x250;
  assign n1762 = ~n1159 & ~n1761;
  assign n1763 = n1762 ^ x250;
  assign n1764 = ~n1158 & n1763;
  assign n1765 = n1157 & ~n1764;
  assign n1766 = ~x127 & x255;
  assign n1767 = x126 & ~x254;
  assign n1768 = ~n1766 & ~n1767;
  assign n1769 = x253 ^ x125;
  assign n1770 = x124 & ~x252;
  assign n1771 = n1770 ^ x253;
  assign n1772 = ~n1769 & ~n1771;
  assign n1773 = n1772 ^ x253;
  assign n1774 = ~n1152 & ~n1773;
  assign n1775 = n1768 & ~n1774;
  assign n1776 = ~n1765 & n1775;
  assign n1777 = x127 & ~x255;
  assign n1778 = ~n1776 & ~n1777;
  assign n1779 = x254 ^ x126;
  assign n1780 = ~n1778 & n1779;
  assign n1781 = n1780 ^ x126;
  assign n1782 = ~n1150 & n1781;
  assign n1783 = n1782 ^ n513;
  assign n1784 = n1783 ^ n513;
  assign n1785 = n1769 & ~n1778;
  assign n1786 = n1785 ^ x125;
  assign n1787 = n1138 & ~n1147;
  assign n1788 = n1787 ^ x381;
  assign n1789 = n1786 & ~n1788;
  assign n1790 = x508 ^ x380;
  assign n1791 = ~n1147 & n1790;
  assign n1792 = n1791 ^ x380;
  assign n1793 = x252 ^ x124;
  assign n1794 = ~n1778 & n1793;
  assign n1795 = n1794 ^ x124;
  assign n1796 = ~n1792 & n1795;
  assign n1797 = ~n1789 & ~n1796;
  assign n1798 = n1792 & ~n1795;
  assign n1802 = x507 ^ x379;
  assign n1803 = ~n1147 & n1802;
  assign n1804 = n1803 ^ x379;
  assign n1799 = x251 ^ x123;
  assign n1800 = ~n1778 & n1799;
  assign n1801 = n1800 ^ x123;
  assign n1805 = n1804 ^ n1801;
  assign n1808 = x506 ^ x378;
  assign n1809 = ~n1147 & n1808;
  assign n1810 = n1809 ^ x378;
  assign n1806 = n1159 & ~n1778;
  assign n1807 = n1806 ^ x122;
  assign n1811 = n1810 ^ n1807;
  assign n1812 = n1160 & ~n1778;
  assign n1813 = n1812 ^ x121;
  assign n1814 = x505 ^ x377;
  assign n1815 = ~n1147 & n1814;
  assign n1816 = n1815 ^ x377;
  assign n1817 = n1813 & ~n1816;
  assign n1818 = n1817 ^ n1807;
  assign n1819 = n1818 ^ n1807;
  assign n1820 = ~n1813 & n1816;
  assign n1823 = x248 ^ x120;
  assign n1824 = ~n1778 & n1823;
  assign n1825 = n1824 ^ x120;
  assign n1821 = n520 & ~n1147;
  assign n1822 = n1821 ^ x376;
  assign n1826 = n1825 ^ n1822;
  assign n1829 = n521 & ~n1147;
  assign n1830 = n1829 ^ x375;
  assign n1827 = n1165 & ~n1778;
  assign n1828 = n1827 ^ x119;
  assign n1831 = n1830 ^ n1828;
  assign n1832 = x502 ^ x374;
  assign n1833 = ~n1147 & n1832;
  assign n1834 = n1833 ^ x374;
  assign n1835 = x246 ^ x118;
  assign n1836 = ~n1778 & n1835;
  assign n1837 = n1836 ^ x118;
  assign n1838 = ~n1834 & n1837;
  assign n1839 = n1838 ^ n1828;
  assign n1840 = n1839 ^ n1828;
  assign n1841 = n1177 & ~n1778;
  assign n1842 = n1841 ^ x113;
  assign n1843 = x497 ^ x369;
  assign n1844 = ~n1147 & n1843;
  assign n1845 = n1844 ^ x369;
  assign n1846 = n1842 & ~n1845;
  assign n1847 = x496 ^ x368;
  assign n1848 = ~n1147 & n1847;
  assign n1849 = n1848 ^ x368;
  assign n1850 = x240 ^ x112;
  assign n1851 = ~n1778 & n1850;
  assign n1852 = n1851 ^ x112;
  assign n1853 = ~n1849 & n1852;
  assign n1854 = ~n1846 & ~n1853;
  assign n1855 = n1849 & ~n1852;
  assign n1859 = n535 & ~n1147;
  assign n1860 = n1859 ^ x367;
  assign n1856 = x239 ^ x111;
  assign n1857 = ~n1778 & n1856;
  assign n1858 = n1857 ^ x111;
  assign n1861 = n1860 ^ n1858;
  assign n1864 = n1185 & ~n1778;
  assign n1865 = n1864 ^ x110;
  assign n1862 = n536 & ~n1147;
  assign n1863 = n1862 ^ x366;
  assign n1866 = n1865 ^ n1863;
  assign n1867 = n1186 & ~n1778;
  assign n1868 = n1867 ^ x109;
  assign n1869 = x493 ^ x365;
  assign n1870 = ~n1147 & n1869;
  assign n1871 = n1870 ^ x365;
  assign n1872 = n1868 & ~n1871;
  assign n1873 = n1872 ^ n1863;
  assign n1874 = n1873 ^ n1863;
  assign n1875 = ~n1868 & n1871;
  assign n1878 = x236 ^ x108;
  assign n1879 = ~n1778 & n1878;
  assign n1880 = n1879 ^ x108;
  assign n1876 = n541 & ~n1147;
  assign n1877 = n1876 ^ x364;
  assign n1881 = n1880 ^ n1877;
  assign n1885 = n542 & ~n1147;
  assign n1886 = n1885 ^ x363;
  assign n1882 = x235 ^ x107;
  assign n1883 = ~n1778 & n1882;
  assign n1884 = n1883 ^ x107;
  assign n1887 = n1886 ^ n1884;
  assign n1888 = x490 ^ x362;
  assign n1889 = ~n1147 & n1888;
  assign n1890 = n1889 ^ x362;
  assign n1891 = n1194 & ~n1778;
  assign n1892 = n1891 ^ x106;
  assign n1893 = ~n1890 & n1892;
  assign n1894 = n1893 ^ n1884;
  assign n1895 = n1894 ^ n1884;
  assign n1896 = n1890 & ~n1892;
  assign n1899 = n547 & ~n1147;
  assign n1900 = n1899 ^ x361;
  assign n1897 = n1195 & ~n1778;
  assign n1898 = n1897 ^ x105;
  assign n1901 = n1900 ^ n1898;
  assign n1905 = x232 ^ x104;
  assign n1906 = ~n1778 & n1905;
  assign n1907 = n1906 ^ x104;
  assign n1902 = x488 ^ x360;
  assign n1903 = ~n1147 & n1902;
  assign n1904 = n1903 ^ x360;
  assign n1908 = n1907 ^ n1904;
  assign n1909 = n552 & ~n1147;
  assign n1910 = n1909 ^ x359;
  assign n1911 = x231 ^ x103;
  assign n1912 = ~n1778 & n1911;
  assign n1913 = n1912 ^ x103;
  assign n1914 = ~n1910 & n1913;
  assign n1915 = n1914 ^ n1904;
  assign n1916 = n1915 ^ n1904;
  assign n1917 = n1910 & ~n1913;
  assign n1920 = x486 ^ x358;
  assign n1921 = ~n1147 & n1920;
  assign n1922 = n1921 ^ x358;
  assign n1918 = n1203 & ~n1778;
  assign n1919 = n1918 ^ x102;
  assign n1923 = n1922 ^ n1919;
  assign n1927 = n1204 & ~n1778;
  assign n1928 = n1927 ^ x101;
  assign n1924 = x485 ^ x357;
  assign n1925 = ~n1147 & n1924;
  assign n1926 = n1925 ^ x357;
  assign n1929 = n1928 ^ n1926;
  assign n1930 = x228 ^ x100;
  assign n1931 = ~n1778 & n1930;
  assign n1932 = n1931 ^ x100;
  assign n1933 = x484 ^ x356;
  assign n1934 = ~n1147 & n1933;
  assign n1935 = n1934 ^ x356;
  assign n1936 = n1932 & ~n1935;
  assign n1937 = n1936 ^ n1926;
  assign n1938 = n1937 ^ n1926;
  assign n1939 = ~n1932 & n1935;
  assign n1940 = n560 & ~n1147;
  assign n1941 = n1940 ^ x355;
  assign n1942 = x227 ^ x99;
  assign n1943 = ~n1778 & n1942;
  assign n1944 = n1943 ^ x99;
  assign n1945 = n1941 & ~n1944;
  assign n1946 = ~n1939 & ~n1945;
  assign n1947 = ~n1941 & n1944;
  assign n1950 = n561 & ~n1147;
  assign n1951 = n1950 ^ x354;
  assign n1948 = n1212 & ~n1778;
  assign n1949 = n1948 ^ x98;
  assign n1952 = n1951 ^ n1949;
  assign n1956 = n1213 & ~n1778;
  assign n1957 = n1956 ^ x97;
  assign n1953 = x481 ^ x353;
  assign n1954 = ~n1147 & n1953;
  assign n1955 = n1954 ^ x353;
  assign n1958 = n1957 ^ n1955;
  assign n1959 = x224 ^ x96;
  assign n1960 = ~n1778 & n1959;
  assign n1961 = n1960 ^ x96;
  assign n1962 = x480 ^ x352;
  assign n1963 = ~n1147 & n1962;
  assign n1964 = n1963 ^ x352;
  assign n1965 = ~n1961 & n1964;
  assign n1966 = n1965 ^ n1955;
  assign n1967 = n1966 ^ n1955;
  assign n1968 = n1961 & ~n1964;
  assign n1969 = x479 ^ x351;
  assign n1970 = ~n1147 & n1969;
  assign n1971 = n1970 ^ x351;
  assign n1972 = n1218 & ~n1778;
  assign n1973 = n1972 ^ x95;
  assign n1974 = ~n1971 & n1973;
  assign n1975 = ~n1968 & ~n1974;
  assign n1976 = n1971 & ~n1973;
  assign n1979 = x478 ^ x350;
  assign n1980 = ~n1147 & n1979;
  assign n1981 = n1980 ^ x350;
  assign n1977 = n1219 & ~n1778;
  assign n1978 = n1977 ^ x94;
  assign n1982 = n1981 ^ n1978;
  assign n1986 = n569 & ~n1147;
  assign n1987 = n1986 ^ x349;
  assign n1983 = x221 ^ x93;
  assign n1984 = ~n1778 & n1983;
  assign n1985 = n1984 ^ x93;
  assign n1988 = n1987 ^ n1985;
  assign n1989 = n570 & ~n1147;
  assign n1990 = n1989 ^ x348;
  assign n1991 = n1224 & ~n1778;
  assign n1992 = n1991 ^ x92;
  assign n1993 = ~n1990 & n1992;
  assign n1994 = n1993 ^ n1985;
  assign n1995 = n1994 ^ n1985;
  assign n1996 = x212 ^ x84;
  assign n1997 = ~n1778 & n1996;
  assign n1998 = n1997 ^ x84;
  assign n1999 = x468 ^ x340;
  assign n2000 = ~n1147 & n1999;
  assign n2001 = n2000 ^ x340;
  assign n2002 = ~n1998 & n2001;
  assign n2003 = x211 ^ x83;
  assign n2004 = ~n1778 & n2003;
  assign n2005 = n2004 ^ x83;
  assign n2006 = n589 & ~n1147;
  assign n2007 = n2006 ^ x339;
  assign n2008 = ~n2005 & n2007;
  assign n2009 = ~n2002 & ~n2008;
  assign n2010 = n2005 & ~n2007;
  assign n2013 = n590 & ~n1147;
  assign n2014 = n2013 ^ x338;
  assign n2011 = n1237 & ~n1778;
  assign n2012 = n2011 ^ x82;
  assign n2015 = n2014 ^ n2012;
  assign n2019 = n1238 & ~n1778;
  assign n2020 = n2019 ^ x81;
  assign n2016 = x465 ^ x337;
  assign n2017 = ~n1147 & n2016;
  assign n2018 = n2017 ^ x337;
  assign n2021 = n2020 ^ n2018;
  assign n2022 = x208 ^ x80;
  assign n2023 = ~n1778 & n2022;
  assign n2024 = n2023 ^ x80;
  assign n2025 = x464 ^ x336;
  assign n2026 = ~n1147 & n2025;
  assign n2027 = n2026 ^ x336;
  assign n2028 = ~n2024 & n2027;
  assign n2029 = n2028 ^ n2018;
  assign n2030 = n2029 ^ n2018;
  assign n2031 = n2024 & ~n2027;
  assign n2034 = x207 ^ x79;
  assign n2035 = ~n1778 & n2034;
  assign n2036 = n2035 ^ x79;
  assign n2032 = n598 & ~n1147;
  assign n2033 = n2032 ^ x335;
  assign n2037 = n2036 ^ n2033;
  assign n2041 = n599 & ~n1147;
  assign n2042 = n2041 ^ x334;
  assign n2038 = x206 ^ x78;
  assign n2039 = ~n1778 & n2038;
  assign n2040 = n2039 ^ x78;
  assign n2043 = n2042 ^ n2040;
  assign n2044 = x461 ^ x333;
  assign n2045 = ~n1147 & n2044;
  assign n2046 = n2045 ^ x333;
  assign n2047 = x205 ^ x77;
  assign n2048 = ~n1778 & n2047;
  assign n2049 = n2048 ^ x77;
  assign n2050 = n2046 & ~n2049;
  assign n2051 = n2050 ^ n2040;
  assign n2052 = n2051 ^ n2040;
  assign n2053 = n610 & ~n1147;
  assign n2054 = n2053 ^ x329;
  assign n2055 = x201 ^ x73;
  assign n2056 = ~n1778 & n2055;
  assign n2057 = n2056 ^ x73;
  assign n2058 = n2054 & ~n2057;
  assign n2059 = x202 ^ x74;
  assign n2060 = ~n1778 & n2059;
  assign n2061 = n2060 ^ x74;
  assign n2062 = x458 ^ x330;
  assign n2063 = ~n1147 & n2062;
  assign n2064 = n2063 ^ x330;
  assign n2065 = ~n2061 & n2064;
  assign n2066 = ~n2058 & ~n2065;
  assign n2067 = ~n2054 & n2057;
  assign n2070 = x200 ^ x72;
  assign n2071 = ~n1778 & n2070;
  assign n2072 = n2071 ^ x72;
  assign n2068 = n611 & ~n1147;
  assign n2069 = n2068 ^ x328;
  assign n2073 = n2072 ^ n2069;
  assign n2077 = x199 ^ x71;
  assign n2078 = ~n1778 & n2077;
  assign n2079 = n2078 ^ x71;
  assign n2074 = x455 ^ x327;
  assign n2075 = ~n1147 & n2074;
  assign n2076 = n2075 ^ x327;
  assign n2080 = n2079 ^ n2076;
  assign n2081 = x198 ^ x70;
  assign n2082 = ~n1778 & n2081;
  assign n2083 = n2082 ^ x70;
  assign n2084 = x454 ^ x326;
  assign n2085 = ~n1147 & n2084;
  assign n2086 = n2085 ^ x326;
  assign n2087 = ~n2083 & n2086;
  assign n2088 = n2087 ^ n2076;
  assign n2089 = n2088 ^ n2076;
  assign n2090 = n1585 & ~n1778;
  assign n2091 = n2090 ^ x69;
  assign n2092 = n954 & ~n1147;
  assign n2093 = n2092 ^ x325;
  assign n2094 = n2091 & ~n2093;
  assign n2095 = n2083 & ~n2086;
  assign n2096 = ~n2094 & ~n2095;
  assign n2097 = ~n2091 & n2093;
  assign n2101 = x452 ^ x324;
  assign n2102 = ~n1147 & n2101;
  assign n2103 = n2102 ^ x324;
  assign n2098 = x196 ^ x68;
  assign n2099 = ~n1778 & n2098;
  assign n2100 = n2099 ^ x68;
  assign n2104 = n2103 ^ n2100;
  assign n2108 = n1247 & ~n1778;
  assign n2109 = n2108 ^ x67;
  assign n2105 = x451 ^ x323;
  assign n2106 = ~n1147 & n2105;
  assign n2107 = n2106 ^ x323;
  assign n2110 = n2109 ^ n2107;
  assign n2111 = x194 ^ x66;
  assign n2112 = ~n1778 & n2111;
  assign n2113 = n2112 ^ x66;
  assign n2114 = n623 & ~n1147;
  assign n2115 = n2114 ^ x322;
  assign n2116 = n2113 & ~n2115;
  assign n2117 = n2116 ^ n2107;
  assign n2118 = n2117 ^ n2107;
  assign n2119 = n629 & ~n1147;
  assign n2120 = n2119 ^ x314;
  assign n2121 = x186 ^ x58;
  assign n2122 = ~n1778 & n2121;
  assign n2123 = n2122 ^ x58;
  assign n2124 = ~n2120 & n2123;
  assign n2125 = x443 ^ x315;
  assign n2126 = ~n1147 & n2125;
  assign n2127 = n2126 ^ x315;
  assign n2128 = x187 ^ x59;
  assign n2129 = ~n1778 & n2128;
  assign n2130 = n2129 ^ x59;
  assign n2131 = ~n2127 & n2130;
  assign n2132 = ~n2124 & ~n2131;
  assign n2133 = n2120 & ~n2123;
  assign n2136 = x441 ^ x313;
  assign n2137 = ~n1147 & n2136;
  assign n2138 = n2137 ^ x313;
  assign n2134 = n1261 & ~n1778;
  assign n2135 = n2134 ^ x57;
  assign n2139 = n2138 ^ n2135;
  assign n2143 = n1262 & ~n1778;
  assign n2144 = n2143 ^ x56;
  assign n2140 = x440 ^ x312;
  assign n2141 = ~n1147 & n2140;
  assign n2142 = n2141 ^ x312;
  assign n2145 = n2144 ^ n2142;
  assign n2146 = x439 ^ x311;
  assign n2147 = ~n1147 & n2146;
  assign n2148 = n2147 ^ x311;
  assign n2149 = x183 ^ x55;
  assign n2150 = ~n1778 & n2149;
  assign n2151 = n2150 ^ x55;
  assign n2152 = ~n2148 & n2151;
  assign n2153 = n2152 ^ n2142;
  assign n2154 = n2153 ^ n2142;
  assign n2155 = x182 ^ x54;
  assign n2156 = ~n1778 & n2155;
  assign n2157 = n2156 ^ x54;
  assign n2158 = x438 ^ x310;
  assign n2159 = ~n1147 & n2158;
  assign n2160 = n2159 ^ x310;
  assign n2161 = ~n2157 & n2160;
  assign n2162 = n2148 & ~n2151;
  assign n2163 = ~n2161 & ~n2162;
  assign n2164 = n2157 & ~n2160;
  assign n2168 = n637 & ~n1147;
  assign n2169 = n2168 ^ x309;
  assign n2165 = x181 ^ x53;
  assign n2166 = ~n1778 & n2165;
  assign n2167 = n2166 ^ x53;
  assign n2170 = n2169 ^ n2167;
  assign n2173 = x180 ^ x52;
  assign n2174 = ~n1778 & n2173;
  assign n2175 = n2174 ^ x52;
  assign n2171 = n638 & ~n1147;
  assign n2172 = n2171 ^ x308;
  assign n2176 = n2175 ^ n2172;
  assign n2177 = x435 ^ x307;
  assign n2178 = ~n1147 & n2177;
  assign n2179 = n2178 ^ x307;
  assign n2180 = x179 ^ x51;
  assign n2181 = ~n1778 & n2180;
  assign n2182 = n2181 ^ x51;
  assign n2183 = n2179 & ~n2182;
  assign n2184 = n2183 ^ n2172;
  assign n2185 = n2184 ^ n2172;
  assign n2186 = n1271 & ~n1778;
  assign n2187 = n2186 ^ x49;
  assign n2188 = x433 ^ x305;
  assign n2189 = ~n1147 & n2188;
  assign n2190 = n2189 ^ x305;
  assign n2191 = ~n2187 & n2190;
  assign n2192 = x434 ^ x306;
  assign n2193 = ~n1147 & n2192;
  assign n2194 = n2193 ^ x306;
  assign n2195 = n1270 & ~n1778;
  assign n2196 = n2195 ^ x50;
  assign n2197 = n2194 & ~n2196;
  assign n2198 = ~n2191 & ~n2197;
  assign n2199 = n2187 & ~n2190;
  assign n2203 = x432 ^ x304;
  assign n2204 = ~n1147 & n2203;
  assign n2205 = n2204 ^ x304;
  assign n2200 = x176 ^ x48;
  assign n2201 = ~n1778 & n2200;
  assign n2202 = n2201 ^ x48;
  assign n2206 = n2205 ^ n2202;
  assign n2207 = x175 ^ x47;
  assign n2208 = ~n1778 & n2207;
  assign n2209 = n2208 ^ x47;
  assign n2210 = x431 ^ x303;
  assign n2211 = ~n1147 & n2210;
  assign n2212 = n2211 ^ x303;
  assign n2213 = n2209 & ~n2212;
  assign n2214 = ~n2209 & n2212;
  assign n2218 = x174 ^ x46;
  assign n2219 = ~n1778 & n2218;
  assign n2220 = n2219 ^ x46;
  assign n2215 = x430 ^ x302;
  assign n2216 = ~n1147 & n2215;
  assign n2217 = n2216 ^ x302;
  assign n2221 = n2220 ^ n2217;
  assign n2224 = n1500 & ~n1778;
  assign n2225 = n2224 ^ x45;
  assign n2222 = n867 & ~n1147;
  assign n2223 = n2222 ^ x301;
  assign n2226 = n2225 ^ n2223;
  assign n2227 = x428 ^ x300;
  assign n2228 = ~n1147 & n2227;
  assign n2229 = n2228 ^ x300;
  assign n2230 = x172 ^ x44;
  assign n2231 = ~n1778 & n2230;
  assign n2232 = n2231 ^ x44;
  assign n2233 = ~n2229 & n2232;
  assign n2234 = n2233 ^ n2223;
  assign n2235 = n2234 ^ n2223;
  assign n2236 = x427 ^ x299;
  assign n2237 = ~n1147 & n2236;
  assign n2238 = n2237 ^ x299;
  assign n2239 = x171 ^ x43;
  assign n2240 = ~n1778 & n2239;
  assign n2241 = n2240 ^ x43;
  assign n2242 = n2238 & ~n2241;
  assign n2243 = n2229 & ~n2232;
  assign n2244 = ~n2242 & ~n2243;
  assign n2245 = ~n2238 & n2241;
  assign n2249 = x170 ^ x42;
  assign n2250 = ~n1778 & n2249;
  assign n2251 = n2250 ^ x42;
  assign n2246 = x426 ^ x298;
  assign n2247 = ~n1147 & n2246;
  assign n2248 = n2247 ^ x298;
  assign n2252 = n2251 ^ n2248;
  assign n2255 = n1481 & ~n1778;
  assign n2256 = n2255 ^ x41;
  assign n2253 = n848 & ~n1147;
  assign n2254 = n2253 ^ x297;
  assign n2257 = n2256 ^ n2254;
  assign n2258 = x168 ^ x40;
  assign n2259 = ~n1778 & n2258;
  assign n2260 = n2259 ^ x40;
  assign n2261 = x424 ^ x296;
  assign n2262 = ~n1147 & n2261;
  assign n2263 = n2262 ^ x296;
  assign n2264 = ~n2260 & n2263;
  assign n2265 = n2264 ^ n2254;
  assign n2266 = n2265 ^ n2254;
  assign n2267 = n2260 & ~n2263;
  assign n2271 = x167 ^ x39;
  assign n2272 = ~n1778 & n2271;
  assign n2273 = n2272 ^ x39;
  assign n2268 = x423 ^ x295;
  assign n2269 = ~n1147 & n2268;
  assign n2270 = n2269 ^ x295;
  assign n2274 = n2273 ^ n2270;
  assign n2275 = n1276 & ~n1778;
  assign n2276 = n2275 ^ x38;
  assign n2277 = n650 & ~n1147;
  assign n2278 = n2277 ^ x294;
  assign n2279 = n2276 & ~n2278;
  assign n2280 = ~n2276 & n2278;
  assign n2284 = n651 & ~n1147;
  assign n2285 = n2284 ^ x293;
  assign n2281 = x165 ^ x37;
  assign n2282 = ~n1778 & n2281;
  assign n2283 = n2282 ^ x37;
  assign n2286 = n2285 ^ n2283;
  assign n2290 = x164 ^ x36;
  assign n2291 = ~n1778 & n2290;
  assign n2292 = n2291 ^ x36;
  assign n2287 = x420 ^ x292;
  assign n2288 = ~n1147 & n2287;
  assign n2289 = n2288 ^ x292;
  assign n2293 = n2292 ^ n2289;
  assign n2294 = x163 ^ x35;
  assign n2295 = ~n1778 & n2294;
  assign n2296 = n2295 ^ x35;
  assign n2297 = n656 & ~n1147;
  assign n2298 = n2297 ^ x291;
  assign n2299 = n2296 & ~n2298;
  assign n2300 = n2299 ^ n2289;
  assign n2301 = n2300 ^ n2289;
  assign n2302 = ~n2296 & n2298;
  assign n2306 = x418 ^ x290;
  assign n2307 = ~n1147 & n2306;
  assign n2308 = n2307 ^ x290;
  assign n2303 = x162 ^ x34;
  assign n2304 = ~n1778 & n2303;
  assign n2305 = n2304 ^ x34;
  assign n2309 = n2308 ^ n2305;
  assign n2310 = n1284 & ~n1778;
  assign n2311 = n2310 ^ x33;
  assign n2312 = x417 ^ x289;
  assign n2313 = ~n1147 & n2312;
  assign n2314 = n2313 ^ x289;
  assign n2315 = ~n2311 & n2314;
  assign n2316 = n2311 & ~n2314;
  assign n2320 = n1285 & ~n1778;
  assign n2321 = n2320 ^ x32;
  assign n2317 = x416 ^ x288;
  assign n2318 = ~n1147 & n2317;
  assign n2319 = n2318 ^ x288;
  assign n2322 = n2321 ^ n2319;
  assign n2323 = x159 ^ x31;
  assign n2324 = ~n1778 & n2323;
  assign n2325 = n2324 ^ x31;
  assign n2326 = n664 & ~n1147;
  assign n2327 = n2326 ^ x287;
  assign n2328 = n2325 & ~n2327;
  assign n2329 = ~n2325 & n2327;
  assign n2332 = n665 & ~n1147;
  assign n2333 = n2332 ^ x286;
  assign n2330 = n1290 & ~n1778;
  assign n2331 = n2330 ^ x30;
  assign n2334 = n2333 ^ n2331;
  assign n2338 = n1291 & ~n1778;
  assign n2339 = n2338 ^ x29;
  assign n2335 = x413 ^ x285;
  assign n2336 = ~n1147 & n2335;
  assign n2337 = n2336 ^ x285;
  assign n2340 = n2339 ^ n2337;
  assign n2341 = x156 ^ x28;
  assign n2342 = ~n1778 & n2341;
  assign n2343 = n2342 ^ x28;
  assign n2344 = x412 ^ x284;
  assign n2345 = ~n1147 & n2344;
  assign n2346 = n2345 ^ x284;
  assign n2347 = n2343 & ~n2346;
  assign n2348 = n2347 ^ n2337;
  assign n2349 = n2348 ^ n2337;
  assign n2350 = ~n2343 & n2346;
  assign n2353 = n673 & ~n1147;
  assign n2354 = n2353 ^ x283;
  assign n2351 = n1296 & ~n1778;
  assign n2352 = n2351 ^ x27;
  assign n2355 = n2354 ^ n2352;
  assign n2356 = n1297 & ~n1778;
  assign n2357 = n2356 ^ x26;
  assign n2358 = n674 & ~n1147;
  assign n2359 = n2358 ^ x282;
  assign n2360 = ~n2357 & n2359;
  assign n2361 = n2357 & ~n2359;
  assign n2365 = x153 ^ x25;
  assign n2366 = ~n1778 & n2365;
  assign n2367 = n2366 ^ x25;
  assign n2362 = x409 ^ x281;
  assign n2363 = ~n1147 & n2362;
  assign n2364 = n2363 ^ x281;
  assign n2368 = n2367 ^ n2364;
  assign n2372 = x152 ^ x24;
  assign n2373 = ~n1778 & n2372;
  assign n2374 = n2373 ^ x24;
  assign n2369 = x408 ^ x280;
  assign n2370 = ~n1147 & n2369;
  assign n2371 = n2370 ^ x280;
  assign n2375 = n2374 ^ n2371;
  assign n2376 = x407 ^ x279;
  assign n2377 = ~n1147 & n2376;
  assign n2378 = n2377 ^ x279;
  assign n2379 = x151 ^ x23;
  assign n2380 = ~n1778 & n2379;
  assign n2381 = n2380 ^ x23;
  assign n2382 = n2378 & ~n2381;
  assign n2383 = n2382 ^ n2371;
  assign n2384 = n2383 ^ n2371;
  assign n2385 = x406 ^ x278;
  assign n2386 = ~n1147 & n2385;
  assign n2387 = n2386 ^ x278;
  assign n2388 = x150 ^ x22;
  assign n2389 = ~n1778 & n2388;
  assign n2390 = n2389 ^ x22;
  assign n2391 = ~n2387 & n2390;
  assign n2392 = ~n2378 & n2381;
  assign n2393 = ~n2391 & ~n2392;
  assign n2394 = n2387 & ~n2390;
  assign n2398 = n682 & ~n1147;
  assign n2399 = n2398 ^ x277;
  assign n2395 = x149 ^ x21;
  assign n2396 = ~n1778 & n2395;
  assign n2397 = n2396 ^ x21;
  assign n2400 = n2399 ^ n2397;
  assign n2403 = x148 ^ x20;
  assign n2404 = ~n1778 & n2403;
  assign n2405 = n2404 ^ x20;
  assign n2401 = n683 & ~n1147;
  assign n2402 = n2401 ^ x276;
  assign n2406 = n2405 ^ n2402;
  assign n2407 = x403 ^ x275;
  assign n2408 = ~n1147 & n2407;
  assign n2409 = n2408 ^ x275;
  assign n2410 = n1305 & ~n1778;
  assign n2411 = n2410 ^ x19;
  assign n2412 = ~n2409 & n2411;
  assign n2413 = n2412 ^ n2402;
  assign n2414 = n2413 ^ n2402;
  assign n2415 = n2409 & ~n2411;
  assign n2418 = n1306 & ~n1778;
  assign n2419 = n2418 ^ x18;
  assign n2416 = n688 & ~n1147;
  assign n2417 = n2416 ^ x274;
  assign n2420 = n2419 ^ n2417;
  assign n2421 = x145 ^ x17;
  assign n2422 = ~n1778 & n2421;
  assign n2423 = n2422 ^ x17;
  assign n2424 = n689 & ~n1147;
  assign n2425 = n2424 ^ x273;
  assign n2426 = ~n2423 & n2425;
  assign n2427 = n2423 & ~n2425;
  assign n2430 = x400 ^ x272;
  assign n2431 = ~n1147 & n2430;
  assign n2432 = n2431 ^ x272;
  assign n2428 = n1311 & ~n1778;
  assign n2429 = n2428 ^ x16;
  assign n2433 = n2432 ^ n2429;
  assign n2436 = n1312 & ~n1778;
  assign n2437 = n2436 ^ x15;
  assign n2434 = n694 & ~n1147;
  assign n2435 = n2434 ^ x271;
  assign n2438 = n2437 ^ n2435;
  assign n2439 = x398 ^ x270;
  assign n2440 = ~n1147 & n2439;
  assign n2441 = n2440 ^ x270;
  assign n2442 = x142 ^ x14;
  assign n2443 = ~n1778 & n2442;
  assign n2444 = n2443 ^ x14;
  assign n2445 = n2441 & ~n2444;
  assign n2446 = n2445 ^ n2435;
  assign n2447 = n2446 ^ n2435;
  assign n2448 = x393 ^ x265;
  assign n2449 = ~n1147 & n2448;
  assign n2450 = n2449 ^ x265;
  assign n2451 = n1327 & ~n1778;
  assign n2452 = n2451 ^ x9;
  assign n2453 = ~n2450 & n2452;
  assign n2454 = x138 ^ x10;
  assign n2455 = ~n1778 & n2454;
  assign n2456 = n2455 ^ x10;
  assign n2457 = x394 ^ x266;
  assign n2458 = ~n1147 & n2457;
  assign n2459 = n2458 ^ x266;
  assign n2460 = n2456 & ~n2459;
  assign n2461 = ~n2453 & ~n2460;
  assign n2462 = n2450 & ~n2452;
  assign n2465 = x392 ^ x264;
  assign n2466 = ~n1147 & n2465;
  assign n2467 = n2466 ^ x264;
  assign n2463 = n1328 & ~n1778;
  assign n2464 = n2463 ^ x8;
  assign n2468 = n2467 ^ n2464;
  assign n2472 = x135 ^ x7;
  assign n2473 = ~n1778 & n2472;
  assign n2474 = n2473 ^ x7;
  assign n2469 = x391 ^ x263;
  assign n2470 = ~n1147 & n2469;
  assign n2471 = n2470 ^ x263;
  assign n2475 = n2474 ^ n2471;
  assign n2476 = x390 ^ x262;
  assign n2477 = ~n1147 & n2476;
  assign n2478 = n2477 ^ x262;
  assign n2479 = n1333 & ~n1778;
  assign n2480 = n2479 ^ x6;
  assign n2481 = ~n2478 & n2480;
  assign n2482 = n2481 ^ n2471;
  assign n2483 = n2482 ^ n2471;
  assign n2484 = n2478 & ~n2480;
  assign n2487 = n1334 & ~n1778;
  assign n2488 = n2487 ^ x5;
  assign n2485 = n712 & ~n1147;
  assign n2486 = n2485 ^ x261;
  assign n2489 = n2488 ^ n2486;
  assign n2492 = x132 ^ x4;
  assign n2493 = ~n1778 & n2492;
  assign n2494 = n2493 ^ x4;
  assign n2490 = n713 & ~n1147;
  assign n2491 = n2490 ^ x260;
  assign n2495 = n2494 ^ n2491;
  assign n2496 = x387 ^ x259;
  assign n2497 = ~n1147 & n2496;
  assign n2498 = n2497 ^ x259;
  assign n2499 = x131 ^ x3;
  assign n2500 = ~n1778 & n2499;
  assign n2501 = n2500 ^ x3;
  assign n2502 = ~n2498 & n2501;
  assign n2503 = n2502 ^ n2491;
  assign n2504 = n2503 ^ n2491;
  assign n2505 = x386 ^ x258;
  assign n2506 = ~n1147 & n2505;
  assign n2507 = n2506 ^ x258;
  assign n2508 = x130 ^ x2;
  assign n2509 = ~n1778 & n2508;
  assign n2510 = n2509 ^ x2;
  assign n2511 = n2507 & ~n2510;
  assign n2512 = n2498 & ~n2501;
  assign n2513 = ~n2511 & ~n2512;
  assign n2514 = ~n2507 & n2510;
  assign n2517 = n721 & ~n1147;
  assign n2518 = n2517 ^ x257;
  assign n2515 = n1342 & ~n1778;
  assign n2516 = n2515 ^ x1;
  assign n2519 = n2518 ^ n2516;
  assign n2520 = x384 ^ x256;
  assign n2521 = ~n1147 & n2520;
  assign n2522 = n2521 ^ x256;
  assign n2523 = x128 ^ x0;
  assign n2524 = ~n1778 & n2523;
  assign n2525 = n2524 ^ x0;
  assign n2526 = ~n2522 & n2525;
  assign n2527 = n2526 ^ n2516;
  assign n2528 = ~n2519 & n2527;
  assign n2529 = n2528 ^ n2516;
  assign n2530 = ~n2514 & ~n2529;
  assign n2531 = n2513 & ~n2530;
  assign n2532 = n2531 ^ n2491;
  assign n2533 = n2532 ^ n2491;
  assign n2534 = ~n2504 & ~n2533;
  assign n2535 = n2534 ^ n2491;
  assign n2536 = ~n2495 & ~n2535;
  assign n2537 = n2536 ^ n2494;
  assign n2538 = n2537 ^ n2486;
  assign n2539 = ~n2489 & ~n2538;
  assign n2540 = n2539 ^ n2486;
  assign n2541 = ~n2484 & ~n2540;
  assign n2542 = n2541 ^ n2471;
  assign n2543 = n2542 ^ n2471;
  assign n2544 = ~n2483 & ~n2543;
  assign n2545 = n2544 ^ n2471;
  assign n2546 = ~n2475 & ~n2545;
  assign n2547 = n2546 ^ n2474;
  assign n2548 = n2547 ^ n2464;
  assign n2549 = ~n2468 & n2548;
  assign n2550 = n2549 ^ n2464;
  assign n2551 = ~n2462 & n2550;
  assign n2552 = n2461 & ~n2551;
  assign n2553 = ~n2456 & n2459;
  assign n2554 = n1322 & ~n1778;
  assign n2555 = n2554 ^ x11;
  assign n2556 = n704 & ~n1147;
  assign n2557 = n2556 ^ x267;
  assign n2558 = ~n2555 & n2557;
  assign n2559 = ~n2553 & ~n2558;
  assign n2560 = ~n2552 & n2559;
  assign n2561 = n2555 & ~n2557;
  assign n2562 = x140 ^ x12;
  assign n2563 = ~n1778 & n2562;
  assign n2564 = n2563 ^ x12;
  assign n2565 = x396 ^ x268;
  assign n2566 = ~n1147 & n2565;
  assign n2567 = n2566 ^ x268;
  assign n2568 = n2564 & ~n2567;
  assign n2569 = ~n2561 & ~n2568;
  assign n2570 = ~n2560 & n2569;
  assign n2571 = ~n2564 & n2567;
  assign n2572 = n699 & ~n1147;
  assign n2573 = n2572 ^ x269;
  assign n2574 = n1317 & ~n1778;
  assign n2575 = n2574 ^ x13;
  assign n2576 = n2573 & ~n2575;
  assign n2577 = ~n2571 & ~n2576;
  assign n2578 = ~n2570 & n2577;
  assign n2579 = ~n2573 & n2575;
  assign n2580 = ~n2441 & n2444;
  assign n2581 = ~n2579 & ~n2580;
  assign n2582 = ~n2578 & n2581;
  assign n2583 = n2582 ^ n2435;
  assign n2584 = n2583 ^ n2435;
  assign n2585 = ~n2447 & ~n2584;
  assign n2586 = n2585 ^ n2435;
  assign n2587 = ~n2438 & n2586;
  assign n2588 = n2587 ^ n2437;
  assign n2589 = n2588 ^ n2429;
  assign n2590 = ~n2433 & n2589;
  assign n2591 = n2590 ^ n2429;
  assign n2592 = ~n2427 & ~n2591;
  assign n2593 = ~n2426 & ~n2592;
  assign n2594 = n2593 ^ n2417;
  assign n2595 = ~n2420 & ~n2594;
  assign n2596 = n2595 ^ n2417;
  assign n2597 = ~n2415 & ~n2596;
  assign n2598 = n2597 ^ n2402;
  assign n2599 = n2598 ^ n2402;
  assign n2600 = ~n2414 & ~n2599;
  assign n2601 = n2600 ^ n2402;
  assign n2602 = ~n2406 & ~n2601;
  assign n2603 = n2602 ^ n2405;
  assign n2604 = n2603 ^ n2397;
  assign n2605 = ~n2400 & n2604;
  assign n2606 = n2605 ^ n2397;
  assign n2607 = ~n2394 & n2606;
  assign n2608 = n2393 & ~n2607;
  assign n2609 = n2608 ^ n2371;
  assign n2610 = n2609 ^ n2371;
  assign n2611 = ~n2384 & ~n2610;
  assign n2612 = n2611 ^ n2371;
  assign n2613 = ~n2375 & n2612;
  assign n2614 = n2613 ^ n2374;
  assign n2615 = n2614 ^ n2364;
  assign n2616 = ~n2368 & ~n2615;
  assign n2617 = n2616 ^ n2364;
  assign n2618 = ~n2361 & n2617;
  assign n2619 = ~n2360 & ~n2618;
  assign n2620 = n2619 ^ n2352;
  assign n2621 = ~n2355 & n2620;
  assign n2622 = n2621 ^ n2352;
  assign n2623 = ~n2350 & n2622;
  assign n2624 = n2623 ^ n2337;
  assign n2625 = n2624 ^ n2337;
  assign n2626 = ~n2349 & ~n2625;
  assign n2627 = n2626 ^ n2337;
  assign n2628 = ~n2340 & ~n2627;
  assign n2629 = n2628 ^ n2339;
  assign n2630 = n2629 ^ n2331;
  assign n2631 = ~n2334 & n2630;
  assign n2632 = n2631 ^ n2331;
  assign n2633 = ~n2329 & n2632;
  assign n2634 = ~n2328 & ~n2633;
  assign n2635 = n2634 ^ n2319;
  assign n2636 = ~n2322 & n2635;
  assign n2637 = n2636 ^ n2319;
  assign n2638 = ~n2316 & n2637;
  assign n2639 = ~n2315 & ~n2638;
  assign n2640 = n2639 ^ n2305;
  assign n2641 = ~n2309 & n2640;
  assign n2642 = n2641 ^ n2305;
  assign n2643 = ~n2302 & n2642;
  assign n2644 = n2643 ^ n2289;
  assign n2645 = n2644 ^ n2289;
  assign n2646 = ~n2301 & ~n2645;
  assign n2647 = n2646 ^ n2289;
  assign n2648 = ~n2293 & ~n2647;
  assign n2649 = n2648 ^ n2292;
  assign n2650 = n2649 ^ n2283;
  assign n2651 = ~n2286 & n2650;
  assign n2652 = n2651 ^ n2283;
  assign n2653 = ~n2280 & n2652;
  assign n2654 = ~n2279 & ~n2653;
  assign n2655 = n2654 ^ n2270;
  assign n2656 = ~n2274 & n2655;
  assign n2657 = n2656 ^ n2270;
  assign n2658 = ~n2267 & n2657;
  assign n2659 = n2658 ^ n2254;
  assign n2660 = n2659 ^ n2254;
  assign n2661 = ~n2266 & ~n2660;
  assign n2662 = n2661 ^ n2254;
  assign n2663 = ~n2257 & n2662;
  assign n2664 = n2663 ^ n2256;
  assign n2665 = n2664 ^ n2248;
  assign n2666 = ~n2252 & ~n2665;
  assign n2667 = n2666 ^ n2248;
  assign n2668 = ~n2245 & n2667;
  assign n2669 = n2244 & ~n2668;
  assign n2670 = n2669 ^ n2223;
  assign n2671 = n2670 ^ n2223;
  assign n2672 = ~n2235 & ~n2671;
  assign n2673 = n2672 ^ n2223;
  assign n2674 = ~n2226 & ~n2673;
  assign n2675 = n2674 ^ n2225;
  assign n2676 = n2675 ^ n2217;
  assign n2677 = ~n2221 & ~n2676;
  assign n2678 = n2677 ^ n2217;
  assign n2679 = ~n2214 & ~n2678;
  assign n2680 = ~n2213 & ~n2679;
  assign n2681 = n2680 ^ n2202;
  assign n2682 = ~n2206 & ~n2681;
  assign n2683 = n2682 ^ n2202;
  assign n2684 = ~n2199 & ~n2683;
  assign n2685 = n2198 & ~n2684;
  assign n2686 = ~n2194 & n2196;
  assign n2687 = ~n2179 & n2182;
  assign n2688 = ~n2686 & ~n2687;
  assign n2689 = ~n2685 & n2688;
  assign n2690 = n2689 ^ n2172;
  assign n2691 = n2690 ^ n2172;
  assign n2692 = ~n2185 & ~n2691;
  assign n2693 = n2692 ^ n2172;
  assign n2694 = ~n2176 & n2693;
  assign n2695 = n2694 ^ n2175;
  assign n2696 = n2695 ^ n2167;
  assign n2697 = ~n2170 & n2696;
  assign n2698 = n2697 ^ n2167;
  assign n2699 = ~n2164 & ~n2698;
  assign n2700 = n2163 & ~n2699;
  assign n2701 = n2700 ^ n2142;
  assign n2702 = n2701 ^ n2142;
  assign n2703 = ~n2154 & ~n2702;
  assign n2704 = n2703 ^ n2142;
  assign n2705 = ~n2145 & ~n2704;
  assign n2706 = n2705 ^ n2144;
  assign n2707 = n2706 ^ n2135;
  assign n2708 = ~n2139 & n2707;
  assign n2709 = n2708 ^ n2135;
  assign n2710 = ~n2133 & n2709;
  assign n2711 = n2132 & ~n2710;
  assign n2712 = n2127 & ~n2130;
  assign n2713 = x188 ^ x60;
  assign n2714 = ~n1778 & n2713;
  assign n2715 = n2714 ^ x60;
  assign n2716 = x444 ^ x316;
  assign n2717 = ~n1147 & n2716;
  assign n2718 = n2717 ^ x316;
  assign n2719 = ~n2715 & n2718;
  assign n2720 = ~n2712 & ~n2719;
  assign n2721 = ~n2711 & n2720;
  assign n2722 = n2715 & ~n2718;
  assign n2723 = x445 ^ x317;
  assign n2724 = ~n1147 & n2723;
  assign n2725 = n2724 ^ x317;
  assign n2726 = n1557 & ~n1778;
  assign n2727 = n2726 ^ x61;
  assign n2728 = ~n2725 & n2727;
  assign n2729 = ~n2722 & ~n2728;
  assign n2730 = ~n2721 & n2729;
  assign n2731 = n2725 & ~n2727;
  assign n2732 = x190 ^ x62;
  assign n2733 = ~n1778 & n2732;
  assign n2734 = n2733 ^ x62;
  assign n2735 = x446 ^ x318;
  assign n2736 = ~n1147 & n2735;
  assign n2737 = n2736 ^ x318;
  assign n2738 = ~n2734 & n2737;
  assign n2739 = ~n2731 & ~n2738;
  assign n2740 = ~n2730 & n2739;
  assign n2741 = n2734 & ~n2737;
  assign n2742 = x191 ^ x63;
  assign n2743 = ~n1778 & n2742;
  assign n2744 = n2743 ^ x63;
  assign n2745 = n932 & ~n1147;
  assign n2746 = n2745 ^ x319;
  assign n2747 = n2744 & ~n2746;
  assign n2748 = ~n2741 & ~n2747;
  assign n2749 = ~n2740 & n2748;
  assign n2750 = ~n2744 & n2746;
  assign n2751 = n1253 & ~n1778;
  assign n2752 = n2751 ^ x64;
  assign n2753 = x448 ^ x320;
  assign n2754 = ~n1147 & n2753;
  assign n2755 = n2754 ^ x320;
  assign n2756 = ~n2752 & n2755;
  assign n2757 = ~n2750 & ~n2756;
  assign n2758 = ~n2749 & n2757;
  assign n2759 = n2752 & ~n2755;
  assign n2760 = n1252 & ~n1778;
  assign n2761 = n2760 ^ x65;
  assign n2762 = n624 & ~n1147;
  assign n2763 = n2762 ^ x321;
  assign n2764 = n2761 & ~n2763;
  assign n2765 = ~n2759 & ~n2764;
  assign n2766 = ~n2758 & n2765;
  assign n2767 = ~n2761 & n2763;
  assign n2768 = ~n2113 & n2115;
  assign n2769 = ~n2767 & ~n2768;
  assign n2770 = ~n2766 & n2769;
  assign n2771 = n2770 ^ n2107;
  assign n2772 = n2771 ^ n2107;
  assign n2773 = ~n2118 & ~n2772;
  assign n2774 = n2773 ^ n2107;
  assign n2775 = ~n2110 & ~n2774;
  assign n2776 = n2775 ^ n2109;
  assign n2777 = n2776 ^ n2100;
  assign n2778 = ~n2104 & n2777;
  assign n2779 = n2778 ^ n2100;
  assign n2780 = ~n2097 & n2779;
  assign n2781 = n2096 & ~n2780;
  assign n2782 = n2781 ^ n2076;
  assign n2783 = n2782 ^ n2076;
  assign n2784 = ~n2089 & ~n2783;
  assign n2785 = n2784 ^ n2076;
  assign n2786 = ~n2080 & n2785;
  assign n2787 = n2786 ^ n2079;
  assign n2788 = n2787 ^ n2069;
  assign n2789 = ~n2073 & ~n2788;
  assign n2790 = n2789 ^ n2069;
  assign n2791 = ~n2067 & n2790;
  assign n2792 = n2066 & ~n2791;
  assign n2793 = n605 & ~n1147;
  assign n2794 = n2793 ^ x331;
  assign n2795 = x203 ^ x75;
  assign n2796 = ~n1778 & n2795;
  assign n2797 = n2796 ^ x75;
  assign n2798 = ~n2794 & n2797;
  assign n2799 = n2061 & ~n2064;
  assign n2800 = ~n2798 & ~n2799;
  assign n2801 = ~n2792 & n2800;
  assign n2802 = x204 ^ x76;
  assign n2803 = ~n1778 & n2802;
  assign n2804 = n2803 ^ x76;
  assign n2805 = n604 & ~n1147;
  assign n2806 = n2805 ^ x332;
  assign n2807 = ~n2804 & n2806;
  assign n2808 = n2794 & ~n2797;
  assign n2809 = ~n2807 & ~n2808;
  assign n2810 = ~n2801 & n2809;
  assign n2811 = ~n2046 & n2049;
  assign n2812 = n2804 & ~n2806;
  assign n2813 = ~n2811 & ~n2812;
  assign n2814 = ~n2810 & n2813;
  assign n2815 = n2814 ^ n2040;
  assign n2816 = n2815 ^ n2040;
  assign n2817 = ~n2052 & ~n2816;
  assign n2818 = n2817 ^ n2040;
  assign n2819 = ~n2043 & ~n2818;
  assign n2820 = n2819 ^ n2042;
  assign n2821 = n2820 ^ n2036;
  assign n2822 = ~n2037 & ~n2821;
  assign n2823 = n2822 ^ n2036;
  assign n2824 = ~n2031 & ~n2823;
  assign n2825 = n2824 ^ n2018;
  assign n2826 = n2825 ^ n2018;
  assign n2827 = ~n2030 & ~n2826;
  assign n2828 = n2827 ^ n2018;
  assign n2829 = ~n2021 & n2828;
  assign n2830 = n2829 ^ n2020;
  assign n2831 = n2830 ^ n2014;
  assign n2832 = ~n2015 & ~n2831;
  assign n2833 = n2832 ^ n2014;
  assign n2834 = ~n2010 & n2833;
  assign n2835 = n2009 & ~n2834;
  assign n2836 = x213 ^ x85;
  assign n2837 = ~n1778 & n2836;
  assign n2838 = n2837 ^ x85;
  assign n2839 = x469 ^ x341;
  assign n2840 = ~n1147 & n2839;
  assign n2841 = n2840 ^ x341;
  assign n2842 = n2838 & ~n2841;
  assign n2843 = n1998 & ~n2001;
  assign n2844 = ~n2842 & ~n2843;
  assign n2845 = ~n2835 & n2844;
  assign n2846 = x470 ^ x342;
  assign n2847 = ~n1147 & n2846;
  assign n2848 = n2847 ^ x342;
  assign n2849 = x214 ^ x86;
  assign n2850 = ~n1778 & n2849;
  assign n2851 = n2850 ^ x86;
  assign n2852 = n2848 & ~n2851;
  assign n2853 = ~n2838 & n2841;
  assign n2854 = ~n2852 & ~n2853;
  assign n2855 = ~n2845 & n2854;
  assign n2856 = ~n2848 & n2851;
  assign n2857 = x215 ^ x87;
  assign n2858 = ~n1778 & n2857;
  assign n2859 = n2858 ^ x87;
  assign n2860 = n581 & ~n1147;
  assign n2861 = n2860 ^ x343;
  assign n2862 = n2859 & ~n2861;
  assign n2863 = ~n2856 & ~n2862;
  assign n2864 = ~n2855 & n2863;
  assign n2865 = x472 ^ x344;
  assign n2866 = ~n1147 & n2865;
  assign n2867 = n2866 ^ x344;
  assign n2868 = x216 ^ x88;
  assign n2869 = ~n1778 & n2868;
  assign n2870 = n2869 ^ x88;
  assign n2871 = n2867 & ~n2870;
  assign n2872 = ~n2859 & n2861;
  assign n2873 = ~n2871 & ~n2872;
  assign n2874 = ~n2864 & n2873;
  assign n2875 = n576 & ~n1147;
  assign n2876 = n2875 ^ x345;
  assign n2877 = x217 ^ x89;
  assign n2878 = ~n1778 & n2877;
  assign n2879 = n2878 ^ x89;
  assign n2880 = ~n2876 & n2879;
  assign n2881 = ~n2867 & n2870;
  assign n2882 = ~n2880 & ~n2881;
  assign n2883 = ~n2874 & n2882;
  assign n2884 = n575 & ~n1147;
  assign n2885 = n2884 ^ x346;
  assign n2886 = n1229 & ~n1778;
  assign n2887 = n2886 ^ x90;
  assign n2888 = n2885 & ~n2887;
  assign n2889 = n2876 & ~n2879;
  assign n2890 = ~n2888 & ~n2889;
  assign n2891 = ~n2883 & n2890;
  assign n2892 = x219 ^ x91;
  assign n2893 = ~n1778 & n2892;
  assign n2894 = n2893 ^ x91;
  assign n2895 = x475 ^ x347;
  assign n2896 = ~n1147 & n2895;
  assign n2897 = n2896 ^ x347;
  assign n2898 = n2894 & ~n2897;
  assign n2899 = ~n2885 & n2887;
  assign n2900 = ~n2898 & ~n2899;
  assign n2901 = ~n2891 & n2900;
  assign n2902 = n1990 & ~n1992;
  assign n2903 = ~n2894 & n2897;
  assign n2904 = ~n2902 & ~n2903;
  assign n2905 = ~n2901 & n2904;
  assign n2906 = n2905 ^ n1985;
  assign n2907 = n2906 ^ n1985;
  assign n2908 = ~n1995 & ~n2907;
  assign n2909 = n2908 ^ n1985;
  assign n2910 = ~n1988 & n2909;
  assign n2911 = n2910 ^ n1987;
  assign n2912 = n2911 ^ n1981;
  assign n2913 = ~n1982 & n2912;
  assign n2914 = n2913 ^ n1981;
  assign n2915 = ~n1976 & ~n2914;
  assign n2916 = n1975 & ~n2915;
  assign n2917 = n2916 ^ n1955;
  assign n2918 = n2917 ^ n1955;
  assign n2919 = ~n1967 & ~n2918;
  assign n2920 = n2919 ^ n1955;
  assign n2921 = ~n1958 & n2920;
  assign n2922 = n2921 ^ n1957;
  assign n2923 = n2922 ^ n1951;
  assign n2924 = ~n1952 & ~n2923;
  assign n2925 = n2924 ^ n1951;
  assign n2926 = ~n1947 & n2925;
  assign n2927 = n1946 & ~n2926;
  assign n2928 = n2927 ^ n1926;
  assign n2929 = n2928 ^ n1926;
  assign n2930 = ~n1938 & ~n2929;
  assign n2931 = n2930 ^ n1926;
  assign n2932 = ~n1929 & ~n2931;
  assign n2933 = n2932 ^ n1928;
  assign n2934 = n2933 ^ n1922;
  assign n2935 = ~n1923 & ~n2934;
  assign n2936 = n2935 ^ n1922;
  assign n2937 = ~n1917 & ~n2936;
  assign n2938 = n2937 ^ n1904;
  assign n2939 = n2938 ^ n1904;
  assign n2940 = ~n1916 & ~n2939;
  assign n2941 = n2940 ^ n1904;
  assign n2942 = ~n1908 & ~n2941;
  assign n2943 = n2942 ^ n1907;
  assign n2944 = n2943 ^ n1900;
  assign n2945 = ~n1901 & ~n2944;
  assign n2946 = n2945 ^ n1900;
  assign n2947 = ~n1896 & ~n2946;
  assign n2948 = n2947 ^ n1884;
  assign n2949 = n2948 ^ n1884;
  assign n2950 = ~n1895 & ~n2949;
  assign n2951 = n2950 ^ n1884;
  assign n2952 = ~n1887 & n2951;
  assign n2953 = n2952 ^ n1886;
  assign n2954 = n2953 ^ n1877;
  assign n2955 = ~n1881 & n2954;
  assign n2956 = n2955 ^ n1877;
  assign n2957 = ~n1875 & ~n2956;
  assign n2958 = n2957 ^ n1863;
  assign n2959 = n2958 ^ n1863;
  assign n2960 = ~n1874 & ~n2959;
  assign n2961 = n2960 ^ n1863;
  assign n2962 = ~n1866 & ~n2961;
  assign n2963 = n2962 ^ n1865;
  assign n2964 = n2963 ^ n1860;
  assign n2965 = ~n1861 & ~n2964;
  assign n2966 = n2965 ^ n1860;
  assign n2967 = ~n1855 & ~n2966;
  assign n2968 = n1854 & ~n2967;
  assign n2969 = x498 ^ x370;
  assign n2970 = ~n1147 & n2969;
  assign n2971 = n2970 ^ x370;
  assign n2972 = n1176 & ~n1778;
  assign n2973 = n2972 ^ x114;
  assign n2974 = n2971 & ~n2973;
  assign n2975 = ~n1842 & n1845;
  assign n2976 = ~n2974 & ~n2975;
  assign n2977 = ~n2968 & n2976;
  assign n2978 = x499 ^ x371;
  assign n2979 = ~n1147 & n2978;
  assign n2980 = n2979 ^ x371;
  assign n2981 = x243 ^ x115;
  assign n2982 = ~n1778 & n2981;
  assign n2983 = n2982 ^ x115;
  assign n2984 = ~n2980 & n2983;
  assign n2985 = ~n2971 & n2973;
  assign n2986 = ~n2984 & ~n2985;
  assign n2987 = ~n2977 & n2986;
  assign n2988 = n1171 & ~n1778;
  assign n2989 = n2988 ^ x116;
  assign n2990 = n527 & ~n1147;
  assign n2991 = n2990 ^ x372;
  assign n2992 = ~n2989 & n2991;
  assign n2993 = n2980 & ~n2983;
  assign n2994 = ~n2992 & ~n2993;
  assign n2995 = ~n2987 & n2994;
  assign n2996 = n1170 & ~n1778;
  assign n2997 = n2996 ^ x117;
  assign n2998 = n526 & ~n1147;
  assign n2999 = n2998 ^ x373;
  assign n3000 = n2997 & ~n2999;
  assign n3001 = n2989 & ~n2991;
  assign n3002 = ~n3000 & ~n3001;
  assign n3003 = ~n2995 & n3002;
  assign n3004 = n1834 & ~n1837;
  assign n3005 = ~n2997 & n2999;
  assign n3006 = ~n3004 & ~n3005;
  assign n3007 = ~n3003 & n3006;
  assign n3008 = n3007 ^ n1828;
  assign n3009 = n3008 ^ n1828;
  assign n3010 = ~n1840 & ~n3009;
  assign n3011 = n3010 ^ n1828;
  assign n3012 = ~n1831 & n3011;
  assign n3013 = n3012 ^ n1830;
  assign n3014 = n3013 ^ n1822;
  assign n3015 = ~n1826 & n3014;
  assign n3016 = n3015 ^ n1822;
  assign n3017 = ~n1820 & ~n3016;
  assign n3018 = n3017 ^ n1807;
  assign n3019 = n3018 ^ n1807;
  assign n3020 = ~n1819 & ~n3019;
  assign n3021 = n3020 ^ n1807;
  assign n3022 = ~n1811 & n3021;
  assign n3023 = n3022 ^ n1810;
  assign n3024 = n3023 ^ n1804;
  assign n3025 = ~n1805 & n3024;
  assign n3026 = n3025 ^ n1804;
  assign n3027 = ~n1798 & ~n3026;
  assign n3028 = n1797 & ~n3027;
  assign n3029 = n1150 & ~n1781;
  assign n3030 = ~n1786 & n1788;
  assign n3031 = ~n3029 & ~n3030;
  assign n3032 = ~n3028 & n3031;
  assign n3033 = n3032 ^ n513;
  assign n3034 = n3033 ^ n513;
  assign n3035 = ~n1784 & ~n3034;
  assign n3036 = n3035 ^ n513;
  assign n3037 = ~n515 & n3036;
  assign n3038 = n3037 ^ n514;
  assign n3039 = n2525 ^ n2522;
  assign n3040 = ~n3038 & n3039;
  assign n3041 = n3040 ^ n2522;
  assign n3042 = n2519 & ~n3038;
  assign n3043 = n3042 ^ n2518;
  assign n3044 = n2510 ^ n2507;
  assign n3045 = ~n3038 & n3044;
  assign n3046 = n3045 ^ n2507;
  assign n3047 = n2501 ^ n2498;
  assign n3048 = ~n3038 & n3047;
  assign n3049 = n3048 ^ n2498;
  assign n3050 = n2495 & n3038;
  assign n3051 = n3050 ^ n2494;
  assign n3052 = n2489 & n3038;
  assign n3053 = n3052 ^ n2488;
  assign n3054 = n2480 ^ n2478;
  assign n3055 = ~n3038 & n3054;
  assign n3056 = n3055 ^ n2478;
  assign n3057 = n2475 & n3038;
  assign n3058 = n3057 ^ n2474;
  assign n3059 = n2468 & ~n3038;
  assign n3060 = n3059 ^ n2467;
  assign n3061 = n2452 ^ n2450;
  assign n3062 = ~n3038 & n3061;
  assign n3063 = n3062 ^ n2450;
  assign n3064 = n2459 ^ n2456;
  assign n3065 = n3038 & n3064;
  assign n3066 = n3065 ^ n2456;
  assign n3067 = n2557 ^ n2555;
  assign n3068 = n3038 & n3067;
  assign n3069 = n3068 ^ n2555;
  assign n3070 = n2567 ^ n2564;
  assign n3071 = n3038 & n3070;
  assign n3072 = n3071 ^ n2564;
  assign n3073 = n2575 ^ n2573;
  assign n3074 = ~n3038 & n3073;
  assign n3075 = n3074 ^ n2573;
  assign n3076 = n2444 ^ n2441;
  assign n3077 = ~n3038 & n3076;
  assign n3078 = n3077 ^ n2441;
  assign n3079 = n2438 & n3038;
  assign n3080 = n3079 ^ n2437;
  assign n3081 = n2433 & ~n3038;
  assign n3082 = n3081 ^ n2432;
  assign n3083 = n2425 ^ n2423;
  assign n3084 = n3038 & n3083;
  assign n3085 = n3084 ^ n2423;
  assign n3086 = n2420 & n3038;
  assign n3087 = n3086 ^ n2419;
  assign n3088 = n2411 ^ n2409;
  assign n3089 = ~n3038 & n3088;
  assign n3090 = n3089 ^ n2409;
  assign n3091 = n2406 & n3038;
  assign n3092 = n3091 ^ n2405;
  assign n3093 = n2400 & ~n3038;
  assign n3094 = n3093 ^ n2399;
  assign n3095 = n2390 ^ n2387;
  assign n3096 = ~n3038 & n3095;
  assign n3097 = n3096 ^ n2387;
  assign n3098 = n2381 ^ n2378;
  assign n3099 = ~n3038 & n3098;
  assign n3100 = n3099 ^ n2378;
  assign n3101 = n2375 & n3038;
  assign n3102 = n3101 ^ n2374;
  assign n3103 = n2368 & n3038;
  assign n3104 = n3103 ^ n2367;
  assign n3105 = n2359 ^ n2357;
  assign n3106 = n3038 & n3105;
  assign n3107 = n3106 ^ n2357;
  assign n3108 = n2355 & ~n3038;
  assign n3109 = n3108 ^ n2354;
  assign n3110 = n2346 ^ n2343;
  assign n3111 = n3038 & n3110;
  assign n3112 = n3111 ^ n2343;
  assign n3113 = n2340 & n3038;
  assign n3114 = n3113 ^ n2339;
  assign n3115 = n2334 & ~n3038;
  assign n3116 = n3115 ^ n2333;
  assign n3117 = n2327 ^ n2325;
  assign n3118 = n3038 & n3117;
  assign n3119 = n3118 ^ n2325;
  assign n3120 = n2322 & n3038;
  assign n3121 = n3120 ^ n2321;
  assign n3122 = n2314 ^ n2311;
  assign n3123 = n3038 & n3122;
  assign n3124 = n3123 ^ n2311;
  assign n3125 = n2309 & ~n3038;
  assign n3126 = n3125 ^ n2308;
  assign n3127 = n2298 ^ n2296;
  assign n3128 = n3038 & n3127;
  assign n3129 = n3128 ^ n2296;
  assign n3130 = n2293 & n3038;
  assign n3131 = n3130 ^ n2292;
  assign n3132 = n2286 & ~n3038;
  assign n3133 = n3132 ^ n2285;
  assign n3134 = n2278 ^ n2276;
  assign n3135 = n3038 & n3134;
  assign n3136 = n3135 ^ n2276;
  assign n3137 = n2274 & n3038;
  assign n3138 = n3137 ^ n2273;
  assign n3139 = n2263 ^ n2260;
  assign n3140 = n3038 & n3139;
  assign n3141 = n3140 ^ n2260;
  assign n3142 = n2257 & n3038;
  assign n3143 = n3142 ^ n2256;
  assign n3144 = n2252 & n3038;
  assign n3145 = n3144 ^ n2251;
  assign n3146 = n2241 ^ n2238;
  assign n3147 = ~n3038 & n3146;
  assign n3148 = n3147 ^ n2238;
  assign n3149 = n2232 ^ n2229;
  assign n3150 = ~n3038 & n3149;
  assign n3151 = n3150 ^ n2229;
  assign n3152 = n2226 & n3038;
  assign n3153 = n3152 ^ n2225;
  assign n3154 = n2221 & n3038;
  assign n3155 = n3154 ^ n2220;
  assign n3156 = n2212 ^ n2209;
  assign n3157 = n3038 & n3156;
  assign n3158 = n3157 ^ n2209;
  assign n3159 = n2206 & ~n3038;
  assign n3160 = n3159 ^ n2205;
  assign n3161 = n2190 ^ n2187;
  assign n3162 = n3038 & n3161;
  assign n3163 = n3162 ^ n2187;
  assign n3164 = n2196 ^ n2194;
  assign n3165 = ~n3038 & n3164;
  assign n3166 = n3165 ^ n2194;
  assign n3167 = n2182 ^ n2179;
  assign n3168 = ~n3038 & n3167;
  assign n3169 = n3168 ^ n2179;
  assign n3170 = n2176 & n3038;
  assign n3171 = n3170 ^ n2175;
  assign n3172 = n2170 & ~n3038;
  assign n3173 = n3172 ^ n2169;
  assign n3174 = n2160 ^ n2157;
  assign n3175 = n3038 & n3174;
  assign n3176 = n3175 ^ n2157;
  assign n3177 = n2151 ^ n2148;
  assign n3178 = ~n3038 & n3177;
  assign n3179 = n3178 ^ n2148;
  assign n3180 = n2145 & n3038;
  assign n3181 = n3180 ^ n2144;
  assign n3182 = n2139 & ~n3038;
  assign n3183 = n3182 ^ n2138;
  assign n3184 = n2123 ^ n2120;
  assign n3185 = ~n3038 & n3184;
  assign n3186 = n3185 ^ n2120;
  assign n3187 = n2130 ^ n2127;
  assign n3188 = ~n3038 & n3187;
  assign n3189 = n3188 ^ n2127;
  assign n3190 = n2718 ^ n2715;
  assign n3191 = n3038 & n3190;
  assign n3192 = n3191 ^ n2715;
  assign n3193 = n2727 ^ n2725;
  assign n3194 = ~n3038 & n3193;
  assign n3195 = n3194 ^ n2725;
  assign n3196 = n2737 ^ n2734;
  assign n3197 = n3038 & n3196;
  assign n3198 = n3197 ^ n2734;
  assign n3199 = n2746 ^ n2744;
  assign n3200 = n3038 & n3199;
  assign n3201 = n3200 ^ n2744;
  assign n3202 = n2755 ^ n2752;
  assign n3203 = n3038 & n3202;
  assign n3204 = n3203 ^ n2752;
  assign n3205 = n2763 ^ n2761;
  assign n3206 = n3038 & n3205;
  assign n3207 = n3206 ^ n2761;
  assign n3208 = n2115 ^ n2113;
  assign n3209 = n3038 & n3208;
  assign n3210 = n3209 ^ n2113;
  assign n3211 = n2110 & n3038;
  assign n3212 = n3211 ^ n2109;
  assign n3213 = n2104 & ~n3038;
  assign n3214 = n3213 ^ n2103;
  assign n3215 = n2093 ^ n2091;
  assign n3216 = n3038 & n3215;
  assign n3217 = n3216 ^ n2091;
  assign n3218 = n2086 ^ n2083;
  assign n3219 = n3038 & n3218;
  assign n3220 = n3219 ^ n2083;
  assign n3221 = n2080 & n3038;
  assign n3222 = n3221 ^ n2079;
  assign n3223 = n2073 & n3038;
  assign n3224 = n3223 ^ n2072;
  assign n3225 = n2057 ^ n2054;
  assign n3226 = ~n3038 & n3225;
  assign n3227 = n3226 ^ n2054;
  assign n3228 = n2064 ^ n2061;
  assign n3229 = n3038 & n3228;
  assign n3230 = n3229 ^ n2061;
  assign n3231 = n2797 ^ n2794;
  assign n3232 = ~n3038 & n3231;
  assign n3233 = n3232 ^ n2794;
  assign n3234 = n2806 ^ n2804;
  assign n3235 = n3038 & n3234;
  assign n3236 = n3235 ^ n2804;
  assign n3237 = n2049 ^ n2046;
  assign n3238 = ~n3038 & n3237;
  assign n3239 = n3238 ^ n2046;
  assign n3240 = n2043 & ~n3038;
  assign n3241 = n3240 ^ n2042;
  assign n3242 = n2037 & n3038;
  assign n3243 = n3242 ^ n2036;
  assign n3244 = n2027 ^ n2024;
  assign n3245 = n3038 & n3244;
  assign n3246 = n3245 ^ n2024;
  assign n3247 = n2021 & n3038;
  assign n3248 = n3247 ^ n2020;
  assign n3249 = n2015 & ~n3038;
  assign n3250 = n3249 ^ n2014;
  assign n3251 = n2007 ^ n2005;
  assign n3252 = n3038 & n3251;
  assign n3253 = n3252 ^ n2005;
  assign n3254 = n2001 ^ n1998;
  assign n3255 = n3038 & n3254;
  assign n3256 = n3255 ^ n1998;
  assign n3257 = n2841 ^ n2838;
  assign n3258 = n3038 & n3257;
  assign n3259 = n3258 ^ n2838;
  assign n3260 = n2851 ^ n2848;
  assign n3261 = ~n3038 & n3260;
  assign n3262 = n3261 ^ n2848;
  assign n3263 = n2861 ^ n2859;
  assign n3264 = n3038 & n3263;
  assign n3265 = n3264 ^ n2859;
  assign n3266 = n2870 ^ n2867;
  assign n3267 = ~n3038 & n3266;
  assign n3268 = n3267 ^ n2867;
  assign n3269 = n2879 ^ n2876;
  assign n3270 = ~n3038 & n3269;
  assign n3271 = n3270 ^ n2876;
  assign n3272 = n2887 ^ n2885;
  assign n3273 = ~n3038 & n3272;
  assign n3274 = n3273 ^ n2885;
  assign n3275 = n2897 ^ n2894;
  assign n3276 = n3038 & n3275;
  assign n3277 = n3276 ^ n2894;
  assign n3278 = n1992 ^ n1990;
  assign n3279 = ~n3038 & n3278;
  assign n3280 = n3279 ^ n1990;
  assign n3281 = n1988 & ~n3038;
  assign n3282 = n3281 ^ n1987;
  assign n3283 = n1982 & ~n3038;
  assign n3284 = n3283 ^ n1981;
  assign n3285 = n1973 ^ n1971;
  assign n3286 = ~n3038 & n3285;
  assign n3287 = n3286 ^ n1971;
  assign n3288 = n1964 ^ n1961;
  assign n3289 = n3038 & n3288;
  assign n3290 = n3289 ^ n1961;
  assign n3291 = n1958 & n3038;
  assign n3292 = n3291 ^ n1957;
  assign n3293 = n1952 & ~n3038;
  assign n3294 = n3293 ^ n1951;
  assign n3295 = n1944 ^ n1941;
  assign n3296 = ~n3038 & n3295;
  assign n3297 = n3296 ^ n1941;
  assign n3298 = n1935 ^ n1932;
  assign n3299 = n3038 & n3298;
  assign n3300 = n3299 ^ n1932;
  assign n3301 = n1929 & n3038;
  assign n3302 = n3301 ^ n1928;
  assign n3303 = n1923 & ~n3038;
  assign n3304 = n3303 ^ n1922;
  assign n3305 = n1913 ^ n1910;
  assign n3306 = ~n3038 & n3305;
  assign n3307 = n3306 ^ n1910;
  assign n3308 = n1908 & n3038;
  assign n3309 = n3308 ^ n1907;
  assign n3310 = n1901 & ~n3038;
  assign n3311 = n3310 ^ n1900;
  assign n3312 = n1892 ^ n1890;
  assign n3313 = ~n3038 & n3312;
  assign n3314 = n3313 ^ n1890;
  assign n3315 = n1887 & ~n3038;
  assign n3316 = n3315 ^ n1886;
  assign n3317 = n1881 & n3038;
  assign n3318 = n3317 ^ n1880;
  assign n3319 = n1871 ^ n1868;
  assign n3320 = n3038 & n3319;
  assign n3321 = n3320 ^ n1868;
  assign n3322 = n1866 & n3038;
  assign n3323 = n3322 ^ n1865;
  assign n3324 = n1861 & ~n3038;
  assign n3325 = n3324 ^ n1860;
  assign n3326 = n1852 ^ n1849;
  assign n3327 = ~n3038 & n3326;
  assign n3328 = n3327 ^ n1849;
  assign n3329 = n1845 ^ n1842;
  assign n3330 = n3038 & n3329;
  assign n3331 = n3330 ^ n1842;
  assign n3332 = n2973 ^ n2971;
  assign n3333 = ~n3038 & n3332;
  assign n3334 = n3333 ^ n2971;
  assign n3335 = n2983 ^ n2980;
  assign n3336 = ~n3038 & n3335;
  assign n3337 = n3336 ^ n2980;
  assign n3338 = n2991 ^ n2989;
  assign n3339 = n3038 & n3338;
  assign n3340 = n3339 ^ n2989;
  assign n3341 = n2999 ^ n2997;
  assign n3342 = n3038 & n3341;
  assign n3343 = n3342 ^ n2997;
  assign n3344 = n1837 ^ n1834;
  assign n3345 = ~n3038 & n3344;
  assign n3346 = n3345 ^ n1834;
  assign n3347 = n1831 & ~n3038;
  assign n3348 = n3347 ^ n1830;
  assign n3349 = n1826 & n3038;
  assign n3350 = n3349 ^ n1825;
  assign n3351 = n1816 ^ n1813;
  assign n3352 = n3038 & n3351;
  assign n3353 = n3352 ^ n1813;
  assign n3354 = n1811 & ~n3038;
  assign n3355 = n3354 ^ n1810;
  assign n3356 = n1805 & ~n3038;
  assign n3357 = n3356 ^ n1804;
  assign n3358 = n1795 ^ n1792;
  assign n3359 = ~n3038 & n3358;
  assign n3360 = n3359 ^ n1792;
  assign n3361 = n1788 ^ n1786;
  assign n3362 = n3038 & n3361;
  assign n3363 = n3362 ^ n1786;
  assign n3364 = n1781 ^ n1150;
  assign n3365 = ~n3038 & n3364;
  assign n3366 = n3365 ^ n1150;
  assign n3367 = n513 & n514;
  assign n3368 = n1778 ^ n1147;
  assign n3369 = ~n3038 & n3368;
  assign n3370 = n3369 ^ n1147;
  assign y0 = n3041;
  assign y1 = n3043;
  assign y2 = n3046;
  assign y3 = n3049;
  assign y4 = n3051;
  assign y5 = n3053;
  assign y6 = n3056;
  assign y7 = n3058;
  assign y8 = n3060;
  assign y9 = n3063;
  assign y10 = n3066;
  assign y11 = n3069;
  assign y12 = n3072;
  assign y13 = n3075;
  assign y14 = n3078;
  assign y15 = n3080;
  assign y16 = n3082;
  assign y17 = n3085;
  assign y18 = n3087;
  assign y19 = n3090;
  assign y20 = n3092;
  assign y21 = n3094;
  assign y22 = n3097;
  assign y23 = n3100;
  assign y24 = n3102;
  assign y25 = n3104;
  assign y26 = n3107;
  assign y27 = n3109;
  assign y28 = n3112;
  assign y29 = n3114;
  assign y30 = n3116;
  assign y31 = n3119;
  assign y32 = n3121;
  assign y33 = n3124;
  assign y34 = n3126;
  assign y35 = n3129;
  assign y36 = n3131;
  assign y37 = n3133;
  assign y38 = n3136;
  assign y39 = n3138;
  assign y40 = n3141;
  assign y41 = n3143;
  assign y42 = n3145;
  assign y43 = n3148;
  assign y44 = n3151;
  assign y45 = n3153;
  assign y46 = n3155;
  assign y47 = n3158;
  assign y48 = n3160;
  assign y49 = n3163;
  assign y50 = n3166;
  assign y51 = n3169;
  assign y52 = n3171;
  assign y53 = n3173;
  assign y54 = n3176;
  assign y55 = n3179;
  assign y56 = n3181;
  assign y57 = n3183;
  assign y58 = n3186;
  assign y59 = n3189;
  assign y60 = n3192;
  assign y61 = n3195;
  assign y62 = n3198;
  assign y63 = n3201;
  assign y64 = n3204;
  assign y65 = n3207;
  assign y66 = n3210;
  assign y67 = n3212;
  assign y68 = n3214;
  assign y69 = n3217;
  assign y70 = n3220;
  assign y71 = n3222;
  assign y72 = n3224;
  assign y73 = n3227;
  assign y74 = n3230;
  assign y75 = n3233;
  assign y76 = n3236;
  assign y77 = n3239;
  assign y78 = n3241;
  assign y79 = n3243;
  assign y80 = n3246;
  assign y81 = n3248;
  assign y82 = n3250;
  assign y83 = n3253;
  assign y84 = n3256;
  assign y85 = n3259;
  assign y86 = n3262;
  assign y87 = n3265;
  assign y88 = n3268;
  assign y89 = n3271;
  assign y90 = n3274;
  assign y91 = n3277;
  assign y92 = n3280;
  assign y93 = n3282;
  assign y94 = n3284;
  assign y95 = n3287;
  assign y96 = n3290;
  assign y97 = n3292;
  assign y98 = n3294;
  assign y99 = n3297;
  assign y100 = n3300;
  assign y101 = n3302;
  assign y102 = n3304;
  assign y103 = n3307;
  assign y104 = n3309;
  assign y105 = n3311;
  assign y106 = n3314;
  assign y107 = n3316;
  assign y108 = n3318;
  assign y109 = n3321;
  assign y110 = n3323;
  assign y111 = n3325;
  assign y112 = n3328;
  assign y113 = n3331;
  assign y114 = n3334;
  assign y115 = n3337;
  assign y116 = n3340;
  assign y117 = n3343;
  assign y118 = n3346;
  assign y119 = n3348;
  assign y120 = n3350;
  assign y121 = n3353;
  assign y122 = n3355;
  assign y123 = n3357;
  assign y124 = n3360;
  assign y125 = n3363;
  assign y126 = n3366;
  assign y127 = n3367;
  assign y128 = ~n3370;
  assign y129 = n3038;
endmodule
