module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141;
  wire n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148;
  assign n148 = ~x8 & ~x10;
  assign n149 = ~x14 & ~x21;
  assign n150 = n148 & n149;
  assign n151 = ~x13 & n150;
  assign n152 = ~x4 & ~x9;
  assign n153 = ~x12 & n152;
  assign n154 = ~x7 & n153;
  assign n155 = n151 & n154;
  assign n156 = ~x12 & ~x13;
  assign n157 = n156 ^ x9;
  assign n159 = ~x6 & ~x7;
  assign n160 = x12 & x13;
  assign n161 = n159 & ~n160;
  assign n158 = x7 ^ x6;
  assign n162 = n161 ^ n158;
  assign n163 = n162 ^ n161;
  assign n164 = n161 ^ n156;
  assign n165 = n164 ^ n161;
  assign n166 = n163 & n165;
  assign n167 = n166 ^ n161;
  assign n168 = n157 & n167;
  assign n169 = n168 ^ n161;
  assign n170 = n155 & ~n169;
  assign n171 = ~x5 & ~x22;
  assign n172 = ~x11 & n171;
  assign n173 = ~x18 & ~x19;
  assign n174 = ~x16 & n173;
  assign n175 = n172 & n174;
  assign n176 = n170 & n175;
  assign n177 = ~x17 & n176;
  assign n178 = x54 & ~n177;
  assign n179 = ~x0 & ~n178;
  assign n180 = x7 & ~n151;
  assign n186 = x10 ^ x8;
  assign n181 = x21 ^ x14;
  assign n182 = x14 ^ x13;
  assign n183 = n181 & n182;
  assign n184 = n183 ^ x14;
  assign n185 = n148 & ~n184;
  assign n187 = n186 ^ n185;
  assign n188 = n186 ^ x7;
  assign n189 = ~x13 & n149;
  assign n190 = n189 ^ n186;
  assign n191 = ~n186 & ~n190;
  assign n192 = n191 ^ n186;
  assign n193 = ~n188 & ~n192;
  assign n194 = n193 ^ n191;
  assign n195 = n194 ^ n186;
  assign n196 = n195 ^ n189;
  assign n197 = n187 & ~n196;
  assign n198 = n197 ^ n185;
  assign n199 = ~n180 & n198;
  assign n200 = ~x6 & n174;
  assign n201 = n153 & n200;
  assign n202 = n199 & n201;
  assign n203 = ~x17 & x54;
  assign n204 = n172 & n203;
  assign n205 = n202 & n204;
  assign n206 = ~x9 & ~x11;
  assign n207 = n206 ^ n171;
  assign n208 = x54 & ~x56;
  assign n209 = n207 & n208;
  assign n210 = ~n205 & ~n209;
  assign n211 = ~n179 & n210;
  assign n212 = ~x3 & ~x129;
  assign n213 = ~n211 & n212;
  assign n214 = ~n176 & n203;
  assign n215 = ~x1 & n212;
  assign n216 = ~n214 & n215;
  assign n217 = ~x5 & ~n169;
  assign n218 = n203 & n212;
  assign n219 = n174 & n218;
  assign n220 = ~x11 & ~x22;
  assign n221 = ~x4 & n220;
  assign n222 = n150 & n221;
  assign n223 = n219 & n222;
  assign n224 = ~n217 & n223;
  assign n225 = x5 & ~n170;
  assign n226 = n224 & ~n225;
  assign n227 = ~n216 & ~n226;
  assign n228 = ~x42 & ~x44;
  assign n229 = ~x40 & n228;
  assign n230 = ~x38 & ~x50;
  assign n231 = n229 & n230;
  assign n232 = ~x41 & ~x46;
  assign n233 = ~x47 & ~x48;
  assign n234 = n232 & n233;
  assign n235 = ~x43 & n234;
  assign n236 = n231 & n235;
  assign n237 = ~x24 & ~x49;
  assign n238 = ~x45 & n237;
  assign n239 = n236 & n238;
  assign n240 = x82 & ~n239;
  assign n241 = x122 & x127;
  assign n242 = ~x82 & n241;
  assign n243 = ~n240 & ~n242;
  assign n244 = ~x15 & ~x20;
  assign n245 = x82 & ~n244;
  assign n246 = n243 & ~n245;
  assign n247 = x2 & ~n246;
  assign n248 = ~x2 & n244;
  assign n249 = n238 & n248;
  assign n250 = n235 & n249;
  assign n251 = x82 & ~n250;
  assign n252 = x82 & ~n230;
  assign n253 = ~n251 & ~n252;
  assign n254 = x82 & ~n229;
  assign n255 = n253 & ~n254;
  assign n256 = ~n241 & n255;
  assign n257 = ~x65 & n256;
  assign n258 = ~n247 & ~n257;
  assign n259 = ~x129 & ~n258;
  assign n260 = ~x61 & ~x118;
  assign n261 = ~x129 & n260;
  assign n262 = ~n177 & n261;
  assign n263 = ~x123 & ~x129;
  assign n264 = x0 & ~x113;
  assign n265 = n263 & n264;
  assign n266 = ~n262 & ~n265;
  assign n267 = n172 & n218;
  assign n268 = n202 & n267;
  assign n269 = x10 & n268;
  assign n270 = ~x54 & n212;
  assign n271 = x4 & n270;
  assign n272 = ~n269 & ~n271;
  assign n273 = ~x16 & n267;
  assign n274 = n170 & n273;
  assign n275 = ~x29 & ~x59;
  assign n276 = n173 & n275;
  assign n277 = n274 & n276;
  assign n278 = ~x25 & x28;
  assign n279 = n277 & n278;
  assign n280 = x5 & n270;
  assign n281 = ~n279 & ~n280;
  assign n282 = x25 & ~x28;
  assign n283 = n277 & n282;
  assign n284 = x6 & n270;
  assign n285 = ~n283 & ~n284;
  assign n286 = x8 & n268;
  assign n287 = x7 & n270;
  assign n288 = ~n286 & ~n287;
  assign n289 = x21 & n268;
  assign n290 = x8 & n270;
  assign n291 = ~n289 & ~n290;
  assign n292 = ~x5 & n219;
  assign n293 = n170 & n292;
  assign n294 = x11 & ~x22;
  assign n295 = n293 & n294;
  assign n296 = x9 & n270;
  assign n297 = ~n295 & ~n296;
  assign n298 = x14 & n268;
  assign n299 = x10 & n270;
  assign n300 = ~n298 & ~n299;
  assign n301 = n293 ^ n270;
  assign n302 = n301 ^ n270;
  assign n303 = n270 ^ x22;
  assign n304 = n303 ^ n270;
  assign n305 = n302 & n304;
  assign n306 = n305 ^ n270;
  assign n307 = ~x11 & n306;
  assign n308 = n307 ^ n270;
  assign n309 = x18 & ~x19;
  assign n310 = n274 & n309;
  assign n311 = x12 & n270;
  assign n312 = ~n310 & ~n311;
  assign n313 = x29 & x54;
  assign n314 = ~x59 & n313;
  assign n315 = ~x25 & ~x28;
  assign n316 = n314 & n315;
  assign n317 = n212 & n316;
  assign n318 = n177 & n317;
  assign n319 = x13 & n270;
  assign n320 = ~n318 & ~n319;
  assign n321 = x13 & n268;
  assign n322 = x14 & n270;
  assign n323 = ~n321 & ~n322;
  assign n324 = x15 & ~n243;
  assign n325 = ~x15 & n239;
  assign n326 = n325 ^ x70;
  assign n327 = n326 ^ n325;
  assign n328 = n325 ^ n241;
  assign n329 = n328 ^ n325;
  assign n330 = ~n327 & ~n329;
  assign n331 = n330 ^ n325;
  assign n332 = ~x82 & n331;
  assign n333 = n332 ^ n325;
  assign n334 = ~n324 & ~n333;
  assign n335 = ~x70 & ~n241;
  assign n336 = n248 & ~n335;
  assign n337 = ~x129 & ~n336;
  assign n338 = ~n334 & n337;
  assign n339 = x6 & n226;
  assign n340 = x16 & n270;
  assign n341 = ~n339 & ~n340;
  assign n342 = ~x29 & x59;
  assign n343 = n315 & n342;
  assign n344 = n218 & n343;
  assign n345 = n176 & n344;
  assign n346 = x17 & n270;
  assign n347 = ~n345 & ~n346;
  assign n348 = x16 & n173;
  assign n349 = n267 & n348;
  assign n350 = n170 & n349;
  assign n351 = x18 & n270;
  assign n352 = ~n350 & ~n351;
  assign n353 = x54 & n212;
  assign n354 = x17 & n353;
  assign n355 = n176 & n354;
  assign n356 = x19 & n270;
  assign n357 = ~n355 & ~n356;
  assign n358 = n325 ^ x20;
  assign n359 = x82 & ~n358;
  assign n360 = ~x82 & ~n241;
  assign n361 = x20 & ~n360;
  assign n362 = ~x71 & ~n241;
  assign n363 = x2 & x82;
  assign n364 = ~n362 & ~n363;
  assign n365 = ~n361 & n364;
  assign n366 = ~x129 & ~n365;
  assign n367 = ~n359 & n366;
  assign n368 = ~x18 & x19;
  assign n369 = n274 & n368;
  assign n370 = x21 & n270;
  assign n371 = ~n369 & ~n370;
  assign n372 = n170 & n224;
  assign n373 = x22 & n270;
  assign n374 = ~n372 & ~n373;
  assign n375 = ~x23 & x55;
  assign n376 = x61 & ~x129;
  assign n377 = ~n375 & n376;
  assign n378 = x63 & n256;
  assign n381 = x82 & n236;
  assign n382 = ~x45 & n381;
  assign n379 = x82 & ~n249;
  assign n380 = n241 & ~n379;
  assign n383 = n382 ^ n380;
  assign n384 = n383 ^ n382;
  assign n385 = x82 & ~n382;
  assign n386 = n385 ^ n382;
  assign n387 = n386 ^ n382;
  assign n388 = ~n384 & ~n387;
  assign n389 = n388 ^ n382;
  assign n390 = ~x24 & ~n389;
  assign n391 = n390 ^ n382;
  assign n392 = ~x129 & ~n391;
  assign n393 = ~n378 & n392;
  assign n394 = ~x26 & ~x27;
  assign n395 = ~x53 & ~x58;
  assign n396 = ~x85 & n395;
  assign n397 = x26 & x27;
  assign n398 = n396 & ~n397;
  assign n399 = ~n394 & n398;
  assign n400 = x53 & x58;
  assign n401 = ~x85 & ~n400;
  assign n402 = n401 ^ n395;
  assign n403 = n402 ^ n401;
  assign n404 = n401 ^ x85;
  assign n405 = n403 & n404;
  assign n406 = n405 ^ n401;
  assign n407 = n394 & n406;
  assign n408 = ~n399 & ~n407;
  assign n409 = ~x116 & ~n408;
  assign n410 = ~x95 & ~x100;
  assign n411 = ~x97 & n410;
  assign n412 = ~x110 & ~n411;
  assign n413 = n394 & n396;
  assign n414 = n412 & n413;
  assign n415 = ~x39 & ~x52;
  assign n416 = ~x51 & n415;
  assign n417 = x26 & x116;
  assign n418 = n416 & n417;
  assign n419 = n398 & ~n418;
  assign n420 = ~n414 & n419;
  assign n421 = ~n409 & ~n420;
  assign n422 = x27 & x116;
  assign n423 = ~n416 & n422;
  assign n424 = n212 & ~n423;
  assign n425 = x116 & ~n394;
  assign n426 = ~x25 & ~n425;
  assign n427 = n424 & ~n426;
  assign n428 = ~n421 & n427;
  assign n429 = ~x96 & ~x110;
  assign n430 = n429 ^ x116;
  assign n431 = ~x85 & n430;
  assign n432 = n431 ^ x116;
  assign n433 = x100 & n432;
  assign n434 = n212 & n394;
  assign n435 = n395 & n434;
  assign n436 = n433 & n435;
  assign n437 = ~n428 & ~n436;
  assign n438 = x116 & n416;
  assign n439 = n396 & ~n438;
  assign n440 = x26 & ~x27;
  assign n441 = n212 & n440;
  assign n442 = n439 & n441;
  assign n443 = ~n436 & ~n442;
  assign n444 = ~x26 & x27;
  assign n445 = n439 & n444;
  assign n446 = x85 & x116;
  assign n447 = ~x95 & ~n446;
  assign n448 = n394 & n395;
  assign n449 = ~n447 & n448;
  assign n450 = ~x100 & n449;
  assign n451 = n432 & n450;
  assign n452 = ~n445 & ~n451;
  assign n453 = n212 & ~n452;
  assign n454 = ~x26 & x28;
  assign n455 = ~n412 & n454;
  assign n456 = ~n418 & ~n455;
  assign n457 = ~x27 & n396;
  assign n458 = ~n456 & n457;
  assign n459 = n453 ^ n409;
  assign n460 = n459 ^ n453;
  assign n461 = n453 ^ x28;
  assign n462 = n460 & n461;
  assign n463 = n462 ^ n453;
  assign n464 = ~n458 & ~n463;
  assign n465 = n212 & ~n464;
  assign n466 = ~n412 & n413;
  assign n467 = ~n409 & ~n466;
  assign n468 = x29 & ~n467;
  assign n469 = x53 & x116;
  assign n470 = n401 & ~n469;
  assign n471 = n434 & n470;
  assign n472 = ~x53 & x97;
  assign n473 = n410 & n429;
  assign n474 = n473 ^ x116;
  assign n475 = x116 ^ x58;
  assign n476 = n475 ^ x116;
  assign n477 = n476 ^ n472;
  assign n478 = n474 & ~n477;
  assign n479 = n478 ^ n473;
  assign n480 = n472 & n479;
  assign n481 = n480 ^ x53;
  assign n482 = n471 & n481;
  assign n483 = ~n409 & n482;
  assign n484 = ~n468 & ~n483;
  assign n485 = n212 & ~n484;
  assign n486 = x106 ^ x88;
  assign n487 = n486 ^ x88;
  assign n488 = x60 ^ x30;
  assign n489 = x109 & n488;
  assign n490 = n489 ^ x30;
  assign n491 = n490 ^ x88;
  assign n492 = ~n487 & n491;
  assign n493 = n492 ^ x88;
  assign n494 = ~x129 & n493;
  assign n495 = x106 ^ x89;
  assign n496 = n495 ^ x89;
  assign n497 = x31 ^ x30;
  assign n498 = ~x109 & n497;
  assign n499 = n498 ^ x30;
  assign n500 = n499 ^ x89;
  assign n501 = ~n496 & n500;
  assign n502 = n501 ^ x89;
  assign n503 = ~x129 & n502;
  assign n504 = x106 ^ x99;
  assign n505 = n504 ^ x99;
  assign n506 = x32 ^ x31;
  assign n507 = ~x109 & n506;
  assign n508 = n507 ^ x31;
  assign n509 = n508 ^ x99;
  assign n510 = ~n505 & n509;
  assign n511 = n510 ^ x99;
  assign n512 = ~x129 & n511;
  assign n513 = x106 ^ x90;
  assign n514 = n513 ^ x90;
  assign n515 = x33 ^ x32;
  assign n516 = ~x109 & n515;
  assign n517 = n516 ^ x32;
  assign n518 = n517 ^ x90;
  assign n519 = ~n514 & n518;
  assign n520 = n519 ^ x90;
  assign n521 = ~x129 & n520;
  assign n522 = x106 ^ x91;
  assign n523 = n522 ^ x91;
  assign n524 = x34 ^ x33;
  assign n525 = ~x109 & n524;
  assign n526 = n525 ^ x33;
  assign n527 = n526 ^ x91;
  assign n528 = ~n523 & n527;
  assign n529 = n528 ^ x91;
  assign n530 = ~x129 & n529;
  assign n531 = x106 ^ x92;
  assign n532 = n531 ^ x92;
  assign n533 = x35 ^ x34;
  assign n534 = ~x109 & n533;
  assign n535 = n534 ^ x34;
  assign n536 = n535 ^ x92;
  assign n537 = ~n532 & n536;
  assign n538 = n537 ^ x92;
  assign n539 = ~x129 & n538;
  assign n540 = x106 ^ x98;
  assign n541 = n540 ^ x98;
  assign n542 = x36 ^ x35;
  assign n543 = ~x109 & n542;
  assign n544 = n543 ^ x35;
  assign n545 = n544 ^ x98;
  assign n546 = ~n541 & n545;
  assign n547 = n546 ^ x98;
  assign n548 = ~x129 & n547;
  assign n549 = x106 ^ x93;
  assign n550 = n549 ^ x93;
  assign n551 = x37 ^ x36;
  assign n552 = ~x109 & n551;
  assign n553 = n552 ^ x36;
  assign n554 = n553 ^ x93;
  assign n555 = ~n550 & n554;
  assign n556 = n555 ^ x93;
  assign n557 = ~x129 & n556;
  assign n558 = x74 ^ x38;
  assign n559 = ~n241 & ~n558;
  assign n560 = n559 ^ x38;
  assign n561 = n253 & ~n560;
  assign n562 = n229 ^ x38;
  assign n563 = x82 & ~n562;
  assign n564 = ~x129 & ~n563;
  assign n565 = ~n561 & n564;
  assign n566 = ~x51 & x109;
  assign n567 = ~x52 & n566;
  assign n568 = n567 ^ x39;
  assign n569 = ~x106 & ~n568;
  assign n570 = ~x129 & ~n569;
  assign n571 = ~x73 & ~n241;
  assign n572 = n253 & ~n571;
  assign n573 = ~n254 & ~n572;
  assign n574 = x82 & ~n228;
  assign n575 = ~n242 & ~n574;
  assign n576 = x40 & ~n575;
  assign n577 = ~n573 & ~n576;
  assign n578 = ~x129 & ~n577;
  assign n579 = ~x46 & n231;
  assign n580 = n579 ^ x41;
  assign n581 = x82 & ~n580;
  assign n582 = ~x129 & ~n581;
  assign n583 = x76 ^ x41;
  assign n584 = ~n241 & ~n583;
  assign n585 = n584 ^ x41;
  assign n586 = ~n251 & ~n585;
  assign n587 = n582 & ~n586;
  assign n588 = n228 & ~n255;
  assign n589 = x44 & x82;
  assign n590 = ~n242 & ~n589;
  assign n591 = x42 & ~n590;
  assign n592 = ~x72 & ~n241;
  assign n593 = ~n574 & n592;
  assign n594 = ~n591 & ~n593;
  assign n595 = ~n588 & n594;
  assign n596 = ~x129 & ~n595;
  assign n597 = n231 & n232;
  assign n598 = n597 ^ x43;
  assign n599 = x82 & ~n598;
  assign n600 = ~x129 & ~n599;
  assign n601 = x77 ^ x43;
  assign n602 = ~n241 & ~n601;
  assign n603 = n602 ^ x43;
  assign n604 = ~n251 & ~n603;
  assign n605 = n600 & ~n604;
  assign n606 = x67 ^ x44;
  assign n607 = ~n241 & ~n606;
  assign n608 = n607 ^ x44;
  assign n609 = n255 & ~n608;
  assign n610 = ~x129 & ~n589;
  assign n611 = ~n609 & n610;
  assign n612 = ~x68 & ~n241;
  assign n613 = ~n379 & ~n612;
  assign n614 = ~n385 & ~n613;
  assign n615 = x45 & ~n360;
  assign n616 = ~n381 & n615;
  assign n617 = ~n614 & ~n616;
  assign n618 = ~x129 & ~n617;
  assign n619 = x75 ^ x46;
  assign n620 = ~n241 & ~n619;
  assign n621 = n620 ^ x46;
  assign n622 = n255 & ~n621;
  assign n623 = n231 ^ x46;
  assign n624 = x82 & ~n623;
  assign n625 = ~x129 & ~n624;
  assign n626 = ~n622 & n625;
  assign n627 = ~x43 & n597;
  assign n628 = n627 ^ x47;
  assign n629 = x82 & ~n628;
  assign n630 = x64 ^ x47;
  assign n631 = ~n241 & ~n630;
  assign n632 = n631 ^ x47;
  assign n633 = ~n251 & ~n632;
  assign n634 = ~x129 & ~n633;
  assign n635 = ~n629 & n634;
  assign n636 = ~x47 & n627;
  assign n637 = n636 ^ x48;
  assign n638 = x82 & ~n637;
  assign n639 = x48 & ~n360;
  assign n640 = ~x62 & ~n241;
  assign n641 = ~n639 & ~n640;
  assign n642 = ~n379 & n641;
  assign n643 = ~x129 & ~n642;
  assign n644 = ~n638 & n643;
  assign n645 = ~x24 & n382;
  assign n646 = x49 & ~n360;
  assign n647 = ~n645 & n646;
  assign n648 = x82 & ~n248;
  assign n649 = ~x69 & ~n241;
  assign n650 = ~n648 & ~n649;
  assign n651 = ~n240 & ~n650;
  assign n652 = ~n647 & ~n651;
  assign n653 = ~x129 & ~n652;
  assign n654 = ~x66 & ~n241;
  assign n655 = n250 & ~n654;
  assign n656 = ~n242 & ~n252;
  assign n657 = ~n254 & n656;
  assign n658 = ~n655 & n657;
  assign n659 = ~x50 & ~n658;
  assign n660 = ~x38 & n229;
  assign n661 = n252 & n660;
  assign n662 = x66 & n360;
  assign n663 = ~x129 & ~n662;
  assign n664 = ~n661 & n663;
  assign n665 = ~n659 & n664;
  assign n666 = x109 ^ x51;
  assign n667 = ~x106 & ~n666;
  assign n668 = ~x129 & ~n667;
  assign n669 = n566 ^ x52;
  assign n670 = ~x106 & ~n669;
  assign n671 = ~x129 & ~n670;
  assign n672 = ~x129 & ~n256;
  assign n673 = x114 & ~x122;
  assign n674 = n263 & n673;
  assign n675 = ~n398 & ~n407;
  assign n676 = n212 & ~n675;
  assign n677 = ~x37 & ~x58;
  assign n678 = n677 ^ x94;
  assign n679 = x58 & ~x116;
  assign n680 = n679 ^ n677;
  assign n681 = n677 ^ n417;
  assign n682 = ~n677 & n681;
  assign n683 = n682 ^ n677;
  assign n684 = ~n680 & ~n683;
  assign n685 = n684 ^ n682;
  assign n686 = n685 ^ n677;
  assign n687 = n686 ^ n417;
  assign n688 = ~n678 & n687;
  assign n689 = n688 ^ x94;
  assign n690 = n676 & n689;
  assign n691 = x58 & x116;
  assign n692 = x60 ^ x57;
  assign n693 = n691 & n692;
  assign n694 = n693 ^ x57;
  assign n695 = n676 & n694;
  assign n696 = n416 & n425;
  assign n697 = ~n679 & ~n696;
  assign n698 = n676 & ~n697;
  assign n699 = x59 & ~n467;
  assign n700 = x96 & n414;
  assign n701 = ~n699 & ~n700;
  assign n702 = n212 & ~n701;
  assign n703 = ~x117 & ~x122;
  assign n704 = x123 ^ x60;
  assign n705 = n703 & n704;
  assign n706 = n705 ^ x60;
  assign n707 = ~x114 & ~x122;
  assign n708 = x123 & ~x129;
  assign n709 = n707 & n708;
  assign n710 = x132 & x133;
  assign n711 = x131 & n710;
  assign n712 = ~x138 & n711;
  assign n713 = x136 & ~x137;
  assign n714 = n712 & n713;
  assign n715 = n714 ^ x62;
  assign n716 = n715 ^ x62;
  assign n717 = x140 ^ x62;
  assign n718 = n716 & ~n717;
  assign n719 = n718 ^ x62;
  assign n720 = ~x129 & n719;
  assign n721 = n714 ^ x63;
  assign n722 = n721 ^ x63;
  assign n723 = x142 ^ x63;
  assign n724 = n722 & ~n723;
  assign n725 = n724 ^ x63;
  assign n726 = ~x129 & n725;
  assign n727 = n714 ^ x64;
  assign n728 = n727 ^ x64;
  assign n729 = x139 ^ x64;
  assign n730 = n728 & ~n729;
  assign n731 = n730 ^ x64;
  assign n732 = ~x129 & n731;
  assign n733 = n714 ^ x65;
  assign n734 = n733 ^ x65;
  assign n735 = x146 ^ x65;
  assign n736 = n734 & ~n735;
  assign n737 = n736 ^ x65;
  assign n738 = ~x129 & n737;
  assign n739 = ~x136 & ~x137;
  assign n740 = n712 & n739;
  assign n741 = n740 ^ x66;
  assign n742 = n741 ^ x66;
  assign n743 = x143 ^ x66;
  assign n744 = n742 & ~n743;
  assign n745 = n744 ^ x66;
  assign n746 = ~x129 & n745;
  assign n747 = n740 ^ x67;
  assign n748 = n747 ^ x67;
  assign n749 = x139 ^ x67;
  assign n750 = n748 & ~n749;
  assign n751 = n750 ^ x67;
  assign n752 = ~x129 & n751;
  assign n753 = n714 ^ x68;
  assign n754 = n753 ^ x68;
  assign n755 = x141 ^ x68;
  assign n756 = n754 & ~n755;
  assign n757 = n756 ^ x68;
  assign n758 = ~x129 & n757;
  assign n759 = n714 ^ x69;
  assign n760 = n759 ^ x69;
  assign n761 = x143 ^ x69;
  assign n762 = n760 & ~n761;
  assign n763 = n762 ^ x69;
  assign n764 = ~x129 & n763;
  assign n765 = n714 ^ x70;
  assign n766 = n765 ^ x70;
  assign n767 = x144 ^ x70;
  assign n768 = n766 & ~n767;
  assign n769 = n768 ^ x70;
  assign n770 = ~x129 & n769;
  assign n771 = n714 ^ x71;
  assign n772 = n771 ^ x71;
  assign n773 = x145 ^ x71;
  assign n774 = n772 & ~n773;
  assign n775 = n774 ^ x71;
  assign n776 = ~x129 & n775;
  assign n777 = n740 ^ x72;
  assign n778 = n777 ^ x72;
  assign n779 = x140 ^ x72;
  assign n780 = n778 & ~n779;
  assign n781 = n780 ^ x72;
  assign n782 = ~x129 & n781;
  assign n783 = n740 ^ x73;
  assign n784 = n783 ^ x73;
  assign n785 = x141 ^ x73;
  assign n786 = n784 & ~n785;
  assign n787 = n786 ^ x73;
  assign n788 = ~x129 & n787;
  assign n789 = n740 ^ x74;
  assign n790 = n789 ^ x74;
  assign n791 = x142 ^ x74;
  assign n792 = n790 & ~n791;
  assign n793 = n792 ^ x74;
  assign n794 = ~x129 & n793;
  assign n795 = n740 ^ x75;
  assign n796 = n795 ^ x75;
  assign n797 = x144 ^ x75;
  assign n798 = n796 & ~n797;
  assign n799 = n798 ^ x75;
  assign n800 = ~x129 & n799;
  assign n801 = n740 ^ x76;
  assign n802 = n801 ^ x76;
  assign n803 = x145 ^ x76;
  assign n804 = n802 & ~n803;
  assign n805 = n804 ^ x76;
  assign n806 = ~x129 & n805;
  assign n807 = n740 ^ x77;
  assign n808 = n807 ^ x77;
  assign n809 = x146 ^ x77;
  assign n810 = n808 & ~n809;
  assign n811 = n810 ^ x77;
  assign n812 = ~x129 & n811;
  assign n813 = ~x136 & x137;
  assign n814 = n712 & n813;
  assign n815 = n814 ^ x78;
  assign n816 = n815 ^ x78;
  assign n817 = x142 ^ x78;
  assign n818 = n816 & n817;
  assign n819 = n818 ^ x78;
  assign n820 = ~x129 & n819;
  assign n821 = n814 ^ x79;
  assign n822 = n821 ^ x79;
  assign n823 = x143 ^ x79;
  assign n824 = n822 & n823;
  assign n825 = n824 ^ x79;
  assign n826 = ~x129 & n825;
  assign n827 = n814 ^ x80;
  assign n828 = n827 ^ x80;
  assign n829 = x144 ^ x80;
  assign n830 = n828 & n829;
  assign n831 = n830 ^ x80;
  assign n832 = ~x129 & n831;
  assign n833 = n814 ^ x81;
  assign n834 = n833 ^ x81;
  assign n835 = x145 ^ x81;
  assign n836 = n834 & n835;
  assign n837 = n836 ^ x81;
  assign n838 = ~x129 & n837;
  assign n839 = n814 ^ x82;
  assign n840 = n839 ^ x82;
  assign n841 = x146 ^ x82;
  assign n842 = n840 & n841;
  assign n843 = n842 ^ x82;
  assign n844 = ~x129 & n843;
  assign n845 = x62 ^ x31;
  assign n846 = ~x137 & ~n845;
  assign n847 = n846 ^ x31;
  assign n848 = ~x138 & n847;
  assign n849 = ~x137 & x138;
  assign n850 = x89 & n849;
  assign n851 = x136 & ~n850;
  assign n852 = ~n848 & n851;
  assign n853 = x138 ^ x115;
  assign n854 = n853 ^ x115;
  assign n855 = x115 ^ x87;
  assign n856 = ~n854 & ~n855;
  assign n857 = n856 ^ x115;
  assign n858 = n813 & n857;
  assign n859 = x138 ^ x119;
  assign n860 = n859 ^ x119;
  assign n861 = x119 ^ x72;
  assign n862 = ~n860 & ~n861;
  assign n863 = n862 ^ x119;
  assign n864 = n739 & ~n863;
  assign n865 = ~n858 & ~n864;
  assign n866 = ~n852 & n865;
  assign n867 = n814 ^ x84;
  assign n868 = n867 ^ x84;
  assign n869 = x141 ^ x84;
  assign n870 = n868 & n869;
  assign n871 = n870 ^ x84;
  assign n872 = ~x129 & n871;
  assign n873 = x96 & n412;
  assign n874 = ~x85 & ~n873;
  assign n875 = n435 & ~n446;
  assign n876 = ~n874 & n875;
  assign n877 = n814 ^ x86;
  assign n878 = n877 ^ x86;
  assign n879 = x139 ^ x86;
  assign n880 = n878 & n879;
  assign n881 = n880 ^ x86;
  assign n882 = ~x129 & n881;
  assign n883 = n814 ^ x87;
  assign n884 = n883 ^ x87;
  assign n885 = x140 ^ x87;
  assign n886 = n884 & n885;
  assign n887 = n886 ^ x87;
  assign n888 = ~x129 & n887;
  assign n889 = x136 & x137;
  assign n890 = n712 & n889;
  assign n891 = n890 ^ x88;
  assign n892 = n891 ^ x88;
  assign n893 = x139 ^ x88;
  assign n894 = n892 & n893;
  assign n895 = n894 ^ x88;
  assign n896 = ~x129 & n895;
  assign n897 = n890 ^ x89;
  assign n898 = n897 ^ x89;
  assign n899 = x140 ^ x89;
  assign n900 = n898 & n899;
  assign n901 = n900 ^ x89;
  assign n902 = ~x129 & n901;
  assign n903 = n890 ^ x90;
  assign n904 = n903 ^ x90;
  assign n905 = x142 ^ x90;
  assign n906 = n904 & n905;
  assign n907 = n906 ^ x90;
  assign n908 = ~x129 & n907;
  assign n909 = n890 ^ x91;
  assign n910 = n909 ^ x91;
  assign n911 = x143 ^ x91;
  assign n912 = n910 & n911;
  assign n913 = n912 ^ x91;
  assign n914 = ~x129 & n913;
  assign n915 = n890 ^ x92;
  assign n916 = n915 ^ x92;
  assign n917 = x144 ^ x92;
  assign n918 = n916 & n917;
  assign n919 = n918 ^ x92;
  assign n920 = ~x129 & n919;
  assign n921 = n890 ^ x93;
  assign n922 = n921 ^ x93;
  assign n923 = x146 ^ x93;
  assign n924 = n922 & n923;
  assign n925 = n924 ^ x93;
  assign n926 = ~x129 & n925;
  assign n927 = x82 & x138;
  assign n928 = n739 & n927;
  assign n929 = n711 & n928;
  assign n930 = n929 ^ x94;
  assign n931 = n930 ^ x94;
  assign n932 = x142 ^ x94;
  assign n933 = n931 & n932;
  assign n934 = n933 ^ x94;
  assign n935 = ~x129 & n934;
  assign n936 = ~x3 & ~x110;
  assign n937 = ~n711 & ~n936;
  assign n938 = n937 ^ x143;
  assign n939 = n938 ^ x143;
  assign n940 = x143 ^ x95;
  assign n941 = n940 ^ x143;
  assign n942 = ~n939 & n941;
  assign n943 = n942 ^ x143;
  assign n944 = ~n929 & n943;
  assign n945 = n944 ^ x143;
  assign n946 = ~x129 & n945;
  assign n947 = ~n929 & ~n937;
  assign n948 = x96 & n947;
  assign n949 = x146 & n929;
  assign n950 = ~n948 & ~n949;
  assign n951 = ~x129 & ~n950;
  assign n952 = x97 & n947;
  assign n953 = x145 & n929;
  assign n954 = ~n952 & ~n953;
  assign n955 = ~x129 & ~n954;
  assign n956 = n890 ^ x98;
  assign n957 = n956 ^ x98;
  assign n958 = x145 ^ x98;
  assign n959 = n957 & n958;
  assign n960 = n959 ^ x98;
  assign n961 = ~x129 & n960;
  assign n962 = n890 ^ x99;
  assign n963 = n962 ^ x99;
  assign n964 = x141 ^ x99;
  assign n965 = n963 & n964;
  assign n966 = n965 ^ x99;
  assign n967 = ~x129 & n966;
  assign n968 = x100 & n947;
  assign n969 = x144 & n929;
  assign n970 = ~n968 & ~n969;
  assign n971 = ~x129 & ~n970;
  assign n972 = x37 & n889;
  assign n973 = x82 & n813;
  assign n974 = ~n972 & ~n973;
  assign n975 = ~x65 & n713;
  assign n976 = ~x138 & ~n975;
  assign n977 = n974 & n976;
  assign n978 = x93 & n713;
  assign n979 = x138 & ~n978;
  assign n980 = x96 & n813;
  assign n981 = n979 & ~n980;
  assign n982 = ~n977 & ~n981;
  assign n983 = x138 ^ x124;
  assign n984 = n983 ^ x124;
  assign n985 = x124 ^ x77;
  assign n986 = ~n984 & ~n985;
  assign n987 = n986 ^ x124;
  assign n988 = n739 & n987;
  assign n989 = ~n982 & ~n988;
  assign n990 = x34 & n889;
  assign n991 = ~x138 & ~n990;
  assign n992 = x79 & n813;
  assign n993 = n991 & ~n992;
  assign n994 = ~x69 & n713;
  assign n995 = ~x66 & n739;
  assign n996 = ~n994 & ~n995;
  assign n997 = n993 & n996;
  assign n998 = x95 & n813;
  assign n999 = x138 & ~n998;
  assign n1000 = x91 & n713;
  assign n1001 = n999 & ~n1000;
  assign n1002 = ~n997 & ~n1001;
  assign n1003 = ~x74 & n739;
  assign n1004 = x137 ^ x63;
  assign n1005 = n1004 ^ x63;
  assign n1006 = x63 ^ x33;
  assign n1007 = n1005 & ~n1006;
  assign n1008 = n1007 ^ x63;
  assign n1009 = x136 & ~n1008;
  assign n1010 = ~n1003 & ~n1009;
  assign n1011 = x78 & n813;
  assign n1012 = ~x138 & ~n1011;
  assign n1013 = n1010 & n1012;
  assign n1014 = x94 & n813;
  assign n1015 = x138 & ~n1014;
  assign n1016 = x90 & n713;
  assign n1017 = n1015 & ~n1016;
  assign n1018 = ~n1013 & ~n1017;
  assign n1019 = ~x73 & n739;
  assign n1020 = ~x138 & ~n1019;
  assign n1021 = ~x68 & n713;
  assign n1022 = n1020 & ~n1021;
  assign n1023 = x32 & n889;
  assign n1024 = x84 & n813;
  assign n1025 = ~n1023 & ~n1024;
  assign n1026 = n1022 & n1025;
  assign n1027 = ~x112 & n813;
  assign n1028 = x138 & ~n1027;
  assign n1029 = x99 & n713;
  assign n1030 = n1028 & ~n1029;
  assign n1031 = ~n1026 & ~n1030;
  assign n1037 = x70 & n713;
  assign n1038 = ~x35 & n889;
  assign n1039 = ~n1037 & ~n1038;
  assign n1040 = x137 ^ x80;
  assign n1041 = n1040 ^ x80;
  assign n1042 = x80 ^ x75;
  assign n1043 = ~n1041 & ~n1042;
  assign n1044 = n1043 ^ x80;
  assign n1045 = ~x136 & ~n1044;
  assign n1046 = n1039 & ~n1045;
  assign n1032 = x125 & n739;
  assign n1033 = x100 & n813;
  assign n1034 = ~n1032 & ~n1033;
  assign n1035 = x92 & n713;
  assign n1036 = n1034 & ~n1035;
  assign n1047 = n1046 ^ n1036;
  assign n1048 = x138 & ~n1047;
  assign n1049 = n1048 ^ n1046;
  assign n1050 = ~n414 & ~n446;
  assign n1051 = n212 & ~n1050;
  assign n1052 = x71 ^ x36;
  assign n1053 = ~x137 & ~n1052;
  assign n1054 = n1053 ^ x36;
  assign n1055 = n1054 ^ x137;
  assign n1056 = n1055 ^ n1054;
  assign n1057 = n1054 ^ x98;
  assign n1058 = n1057 ^ n1054;
  assign n1059 = ~n1056 & n1058;
  assign n1060 = n1059 ^ n1054;
  assign n1061 = x138 & n1060;
  assign n1062 = n1061 ^ n1054;
  assign n1063 = x136 & n1062;
  assign n1064 = x138 ^ x76;
  assign n1065 = n1064 ^ x76;
  assign n1066 = x76 ^ x23;
  assign n1067 = n1065 & ~n1066;
  assign n1068 = n1067 ^ x76;
  assign n1069 = n739 & ~n1068;
  assign n1070 = x138 ^ x97;
  assign n1071 = n1070 ^ x97;
  assign n1072 = x97 ^ x81;
  assign n1073 = ~n1071 & n1072;
  assign n1074 = n1073 ^ x97;
  assign n1075 = n813 & n1074;
  assign n1076 = ~n1069 & ~n1075;
  assign n1077 = ~n1063 & n1076;
  assign n1078 = x64 ^ x30;
  assign n1079 = ~x137 & ~n1078;
  assign n1080 = n1079 ^ x30;
  assign n1081 = ~x138 & n1080;
  assign n1082 = x88 & n849;
  assign n1083 = x136 & ~n1082;
  assign n1084 = ~n1081 & n1083;
  assign n1085 = x138 ^ x120;
  assign n1086 = n1085 ^ x120;
  assign n1087 = x120 ^ x67;
  assign n1088 = ~n1086 & ~n1087;
  assign n1089 = n1088 ^ x120;
  assign n1090 = n739 & ~n1089;
  assign n1091 = x138 ^ x111;
  assign n1092 = n1091 ^ x111;
  assign n1093 = x111 ^ x86;
  assign n1094 = ~n1092 & n1093;
  assign n1095 = n1094 ^ x111;
  assign n1096 = n813 & ~n1095;
  assign n1097 = ~n1090 & ~n1096;
  assign n1098 = ~n1084 & n1097;
  assign n1099 = ~n416 & n444;
  assign n1100 = ~n440 & ~n1099;
  assign n1101 = x116 & n212;
  assign n1102 = ~n1100 & n1101;
  assign n1103 = x58 ^ x53;
  assign n1104 = ~n472 & n1103;
  assign n1105 = n1101 & n1104;
  assign n1106 = ~x129 & n711;
  assign n1107 = n928 ^ x139;
  assign n1108 = n1107 ^ x139;
  assign n1109 = x139 ^ x111;
  assign n1110 = ~n1108 & n1109;
  assign n1111 = n1110 ^ x139;
  assign n1112 = n1106 & n1111;
  assign n1113 = n928 ^ x141;
  assign n1114 = n1113 ^ x141;
  assign n1115 = x141 ^ x112;
  assign n1116 = ~n1114 & ~n1115;
  assign n1117 = n1116 ^ x141;
  assign n1118 = n1106 & n1117;
  assign n1119 = x113 ^ x54;
  assign n1120 = n1119 ^ x113;
  assign n1121 = n220 ^ x113;
  assign n1122 = n1120 & n1121;
  assign n1123 = n1122 ^ x113;
  assign n1124 = n212 & ~n1123;
  assign n1125 = n928 ^ x140;
  assign n1126 = n1125 ^ x140;
  assign n1127 = x140 ^ x115;
  assign n1128 = ~n1126 & ~n1127;
  assign n1129 = n1128 ^ x140;
  assign n1130 = n1106 & n1129;
  assign n1131 = ~n154 & n353;
  assign n1132 = x122 & ~x129;
  assign n1133 = ~x54 & x118;
  assign n1134 = ~n316 & ~n1133;
  assign n1135 = ~x129 & ~n1134;
  assign n1136 = ~x129 & ~n410;
  assign n1137 = ~x120 & n936;
  assign n1138 = ~x111 & ~x129;
  assign n1139 = ~n1137 & n1138;
  assign n1140 = x81 & x120;
  assign n1141 = ~x129 & n1140;
  assign n1142 = ~x129 & ~x134;
  assign n1143 = ~x129 & ~x135;
  assign n1144 = x57 & ~x129;
  assign n1145 = ~x96 & x125;
  assign n1146 = ~x3 & ~n1145;
  assign n1147 = ~x129 & ~n1146;
  assign n1148 = ~x126 & n710;
  assign y0 = x108;
  assign y1 = x83;
  assign y2 = x104;
  assign y3 = x103;
  assign y4 = x102;
  assign y5 = x105;
  assign y6 = x107;
  assign y7 = x101;
  assign y8 = x126;
  assign y9 = x121;
  assign y10 = x1;
  assign y11 = x0;
  assign y12 = ~1'b0;
  assign y13 = x130;
  assign y14 = x128;
  assign y15 = ~n213;
  assign y16 = n227;
  assign y17 = n259;
  assign y18 = ~n266;
  assign y19 = ~n272;
  assign y20 = ~n281;
  assign y21 = ~n285;
  assign y22 = ~n288;
  assign y23 = ~n291;
  assign y24 = ~n297;
  assign y25 = ~n300;
  assign y26 = n308;
  assign y27 = ~n312;
  assign y28 = ~n320;
  assign y29 = ~n323;
  assign y30 = n338;
  assign y31 = ~n341;
  assign y32 = ~n347;
  assign y33 = ~n352;
  assign y34 = ~n357;
  assign y35 = n367;
  assign y36 = ~n371;
  assign y37 = ~n374;
  assign y38 = n377;
  assign y39 = n393;
  assign y40 = ~n437;
  assign y41 = ~n443;
  assign y42 = n453;
  assign y43 = n465;
  assign y44 = n485;
  assign y45 = n494;
  assign y46 = n503;
  assign y47 = n512;
  assign y48 = n521;
  assign y49 = n530;
  assign y50 = n539;
  assign y51 = n548;
  assign y52 = n557;
  assign y53 = n565;
  assign y54 = n570;
  assign y55 = n578;
  assign y56 = n587;
  assign y57 = n596;
  assign y58 = n605;
  assign y59 = n611;
  assign y60 = n618;
  assign y61 = n626;
  assign y62 = n635;
  assign y63 = n644;
  assign y64 = n653;
  assign y65 = n665;
  assign y66 = n668;
  assign y67 = n671;
  assign y68 = n482;
  assign y69 = ~n672;
  assign y70 = n674;
  assign y71 = n690;
  assign y72 = n695;
  assign y73 = n698;
  assign y74 = n702;
  assign y75 = n706;
  assign y76 = n709;
  assign y77 = ~n720;
  assign y78 = ~n726;
  assign y79 = ~n732;
  assign y80 = ~n738;
  assign y81 = ~n746;
  assign y82 = ~n752;
  assign y83 = ~n758;
  assign y84 = ~n764;
  assign y85 = ~n770;
  assign y86 = ~n776;
  assign y87 = ~n782;
  assign y88 = ~n788;
  assign y89 = ~n794;
  assign y90 = ~n800;
  assign y91 = ~n806;
  assign y92 = ~n812;
  assign y93 = n820;
  assign y94 = n826;
  assign y95 = n832;
  assign y96 = n838;
  assign y97 = n844;
  assign y98 = n866;
  assign y99 = n872;
  assign y100 = n876;
  assign y101 = n882;
  assign y102 = n888;
  assign y103 = n896;
  assign y104 = n902;
  assign y105 = n908;
  assign y106 = n914;
  assign y107 = n920;
  assign y108 = n926;
  assign y109 = n935;
  assign y110 = n946;
  assign y111 = n951;
  assign y112 = n955;
  assign y113 = n961;
  assign y114 = n967;
  assign y115 = n971;
  assign y116 = ~n989;
  assign y117 = n1002;
  assign y118 = n1018;
  assign y119 = n1031;
  assign y120 = n1049;
  assign y121 = n1051;
  assign y122 = ~n1077;
  assign y123 = n1098;
  assign y124 = n1102;
  assign y125 = n1105;
  assign y126 = n1112;
  assign y127 = n1118;
  assign y128 = n1124;
  assign y129 = ~n263;
  assign y130 = n1130;
  assign y131 = n1131;
  assign y132 = ~n1132;
  assign y133 = n1135;
  assign y134 = n1136;
  assign y135 = n1139;
  assign y136 = n1141;
  assign y137 = ~n1142;
  assign y138 = ~n1143;
  assign y139 = n1144;
  assign y140 = n1147;
  assign y141 = n1148;
endmodule
