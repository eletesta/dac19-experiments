module top(n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886);
  input n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127;
  output n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886;
  wire n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821;
  assign n206 = n52 ^ n116;
  assign n195 = n54 ^ n118;
  assign n180 = n56 ^ n120;
  assign n822 = n0 ^ n64;
  assign n217 = n50 ^ n114;
  assign n752 = n11 & n75;
  assign n691 = n23 & n87;
  assign n695 = n42 & n106;
  assign n692 = n48 & n112;
  assign n697 = n39 & n103;
  assign n699 = n15 & n79;
  assign n700 = n20 & n84;
  assign n739 = n9 & n73;
  assign n702 = n16 & n80;
  assign n703 = n27 & n91;
  assign n704 = n58 & n122;
  assign n736 = n38 & n102;
  assign n705 = n5 & n69;
  assign n776 = n40 & n104;
  assign n709 = n52 & n116;
  assign n710 = n59 & n123;
  assign n711 = n62 & n126;
  assign n714 = n57 & n121;
  assign n715 = n13 & n77;
  assign n716 = n21 & n85;
  assign n719 = n31 & n95;
  assign n717 = n29 & n93;
  assign n734 = n49 & n113;
  assign n720 = n10 & n74;
  assign n721 = n37 & n101;
  assign n723 = n56 & n120;
  assign n724 = n33 & n97;
  assign n725 = n8 & n72;
  assign n726 = n60 & n124;
  assign n730 = n46 & n110;
  assign n728 = n12 & n76;
  assign n729 = n43 & n107;
  assign n722 = n6 & n70;
  assign n733 = n41 & n105;
  assign n735 = n47 & n111;
  assign n727 = n25 & n89;
  assign n737 = n1 & n65;
  assign n738 = n34 & n98;
  assign n741 = n32 & n96;
  assign n558 = n64 & n0;
  assign n685 = n2 & n66;
  assign n718 = n14 & n78;
  assign n742 = n30 & n94;
  assign n743 = n24 & n88;
  assign n744 = n28 & n92;
  assign n664 = n45 & n109;
  assign n746 = n50 & n114;
  assign n775 = n26 & n90;
  assign n749 = n44 & n108;
  assign n753 = n115 & n51;
  assign n803 = n17 & n81;
  assign n708 = n19 & n83;
  assign n754 = n61 & n125;
  assign n755 = n22 & n86;
  assign n701 = n53 & n117;
  assign n698 = n63 & n127;
  assign n740 = n3 & n67;
  assign n696 = n119 & n55;
  assign n745 = n36 & n100;
  assign n751 = n7 & n71;
  assign n645 = n18 & n82;
  assign n767 = n35 & n99;
  assign n774 = n54 & n118;
  assign n750 = n4 & n68;
  assign n757 = ~n52;
  assign n796 = ~n120;
  assign n761 = ~n13;
  assign n689 = ~n86;
  assign n802 = ~n33;
  assign n672 = ~n9;
  assign n679 = ~n76;
  assign n795 = ~n99;
  assign n653 = ~n7;
  assign n818 = ~n119;
  assign n684 = ~n24;
  assign n638 = ~n47;
  assign n649 = ~n126;
  assign n648 = ~n62;
  assign n798 = ~n48;
  assign n758 = ~n81;
  assign n759 = ~n17;
  assign n800 = ~n2;
  assign n780 = ~n42;
  assign n642 = ~n31;
  assign n763 = ~n15;
  assign n683 = ~n88;
  assign n783 = ~n40;
  assign n765 = ~n105;
  assign n820 = ~n94;
  assign n687 = ~n125;
  assign n674 = ~n25;
  assign n772 = ~n59;
  assign n678 = ~n23;
  assign n768 = ~n69;
  assign n655 = ~n46;
  assign n668 = ~n45;
  assign n660 = ~n102;
  assign n809 = ~n3;
  assign n658 = ~n118;
  assign n797 = ~n56;
  assign n731 = ~n70;
  assign n654 = ~n110;
  assign n693 = ~n100;
  assign n815 = ~n8;
  assign n747 = ~n85;
  assign n646 = ~n93;
  assign n792 = ~n107;
  assign n643 = ~n103;
  assign n805 = ~n65;
  assign n611 = ~n113;
  assign n748 = ~n21;
  assign n712 = ~n80;
  assign n686 = ~n61;
  assign n810 = ~n68;
  assign n777 = ~n108;
  assign n676 = ~n10;
  assign n707 = ~n98;
  assign n801 = ~n97;
  assign n659 = ~n54;
  assign n669 = ~n37;
  assign n713 = ~n16;
  assign n650 = ~n121;
  assign n694 = ~n36;
  assign n690 = ~n22;
  assign n675 = ~n74;
  assign n681 = ~n82;
  assign n791 = ~n19;
  assign n673 = ~n89;
  assign n647 = ~n29;
  assign n612 = ~n112;
  assign n665 = ~n90;
  assign n808 = ~n67;
  assign n605 = ~n122;
  assign n786 = ~n92;
  assign n706 = ~n34;
  assign n788 = ~n78;
  assign n793 = ~n43;
  assign n644 = ~n39;
  assign n641 = ~n95;
  assign n807 = ~n96;
  assign n804 = ~n1;
  assign n769 = ~n5;
  assign n770 = ~n115;
  assign n600 = ~n117;
  assign n817 = ~n124;
  assign n766 = ~n41;
  assign n760 = ~n77;
  assign n688 = ~n53;
  assign n756 = ~n116;
  assign n782 = ~n104;
  assign n816 = ~n60;
  assign n662 = ~n75;
  assign n789 = ~n14;
  assign n651 = ~n57;
  assign n799 = ~n66;
  assign n819 = ~n55;
  assign n652 = ~n71;
  assign n640 = ~n127;
  assign n787 = ~n28;
  assign n785 = ~n50;
  assign n677 = ~n87;
  assign n812 = ~n84;
  assign n657 = ~n27;
  assign n811 = ~n4;
  assign n779 = ~n106;
  assign n806 = ~n32;
  assign n773 = ~n123;
  assign n762 = ~n79;
  assign n764 = ~n58;
  assign n814 = ~n72;
  assign n666 = ~n26;
  assign n667 = ~n109;
  assign n771 = ~n51;
  assign n794 = ~n35;
  assign n781 = ~n49;
  assign n682 = ~n18;
  assign n813 = ~n20;
  assign n778 = ~n44;
  assign n661 = ~n38;
  assign n784 = ~n114;
  assign n663 = ~n11;
  assign n821 = ~n30;
  assign n656 = ~n91;
  assign n637 = ~n111;
  assign n790 = ~n83;
  assign n680 = ~n12;
  assign n639 = ~n63;
  assign n671 = ~n73;
  assign n732 = ~n6;
  assign n670 = ~n101;
  assign n200 = n53 ^ n600;
  assign n167 = n58 ^ n605;
  assign n224 = n49 ^ n611;
  assign n232 = n48 ^ n612;
  assign n636 = n637 & n638;
  assign n570 = n639 & n640;
  assign n632 = n641 & n642;
  assign n606 = n643 & n644;
  assign n438 = ~n645;
  assign n574 = n646 & n647;
  assign n575 = n648 & n649;
  assign n576 = n650 & n651;
  assign n577 = n652 & n653;
  assign n578 = n654 & n655;
  assign n579 = n656 & n657;
  assign n604 = n658 & n659;
  assign n581 = n660 & n661;
  assign n582 = n662 & n663;
  assign n249 = ~n664;
  assign n583 = n665 & n666;
  assign n584 = n667 & n668;
  assign n585 = n669 & n670;
  assign n586 = n671 & n672;
  assign n587 = n673 & n674;
  assign n588 = n675 & n676;
  assign n589 = n677 & n678;
  assign n590 = n679 & n680;
  assign n607 = n681 & n682;
  assign n591 = n683 & n684;
  assign n550 = ~n685;
  assign n593 = n686 & n687;
  assign n594 = n600 & n688;
  assign n595 = n689 & n690;
  assign n403 = ~n691;
  assign n227 = ~n692;
  assign n596 = n693 & n694;
  assign n270 = ~n695;
  assign n186 = ~n696;
  assign n291 = ~n697;
  assign n130 = ~n698;
  assign n459 = ~n699;
  assign n424 = ~n700;
  assign n201 = ~n701;
  assign n452 = ~n702;
  assign n375 = ~n703;
  assign n168 = ~n704;
  assign n529 = ~n705;
  assign n571 = n706 & n707;
  assign n431 = ~n708;
  assign n203 = ~n709;
  assign n158 = ~n710;
  assign n137 = ~n711;
  assign n599 = n712 & n713;
  assign n171 = ~n714;
  assign n473 = ~n715;
  assign n417 = ~n716;
  assign n361 = ~n717;
  assign n466 = ~n718;
  assign n347 = ~n719;
  assign n494 = ~n720;
  assign n304 = ~n721;
  assign n522 = ~n722;
  assign n177 = ~n723;
  assign n333 = ~n724;
  assign n508 = ~n725;
  assign n151 = ~n726;
  assign n389 = ~n727;
  assign n480 = ~n728;
  assign n263 = ~n729;
  assign n242 = ~n730;
  assign n573 = n731 & n732;
  assign n277 = ~n733;
  assign n225 = ~n734;
  assign n235 = ~n735;
  assign n298 = ~n736;
  assign n556 = ~n737;
  assign n325 = ~n738;
  assign n501 = ~n739;
  assign n543 = ~n740;
  assign n339 = ~n741;
  assign n354 = ~n742;
  assign n396 = ~n743;
  assign n368 = ~n744;
  assign n312 = ~n745;
  assign n215 = ~n746;
  assign n609 = n747 & n748;
  assign n256 = ~n749;
  assign n536 = ~n750;
  assign n515 = ~n751;
  assign n487 = ~n752;
  assign n213 = ~n753;
  assign n144 = ~n754;
  assign n410 = ~n755;
  assign n598 = n756 & n757;
  assign n580 = n758 & n759;
  assign n592 = n760 & n761;
  assign n603 = n762 & n763;
  assign n608 = n605 & n764;
  assign n597 = n765 & n766;
  assign n318 = ~n767;
  assign n610 = n768 & n769;
  assign n613 = n770 & n771;
  assign n601 = n772 & n773;
  assign n193 = ~n774;
  assign n382 = ~n775;
  assign n284 = ~n776;
  assign n615 = n777 & n778;
  assign n614 = n779 & n780;
  assign n616 = n611 & n781;
  assign n617 = n782 & n783;
  assign n618 = n784 & n785;
  assign n619 = n786 & n787;
  assign n620 = n788 & n789;
  assign n572 = n790 & n791;
  assign n621 = n792 & n793;
  assign n622 = n794 & n795;
  assign n623 = n796 & n797;
  assign n624 = n612 & n798;
  assign n625 = n799 & n800;
  assign n626 = n801 & n802;
  assign n445 = ~n803;
  assign n627 = n804 & n805;
  assign n628 = n806 & n807;
  assign n629 = n808 & n809;
  assign n630 = n810 & n811;
  assign n631 = n812 & n813;
  assign n602 = n814 & n815;
  assign n633 = n816 & n817;
  assign n634 = n818 & n819;
  assign n635 = n820 & n821;
  assign n133 = ~n570;
  assign n328 = ~n571;
  assign n434 = ~n572;
  assign n525 = ~n573;
  assign n364 = ~n574;
  assign n142 = ~n575;
  assign n174 = ~n576;
  assign n518 = ~n577;
  assign n245 = ~n578;
  assign n378 = ~n579;
  assign n448 = ~n580;
  assign n301 = ~n581;
  assign n490 = ~n582;
  assign n385 = ~n583;
  assign n252 = ~n584;
  assign n307 = ~n585;
  assign n504 = ~n586;
  assign n392 = ~n587;
  assign n497 = ~n588;
  assign n406 = ~n589;
  assign n483 = ~n590;
  assign n399 = ~n591;
  assign n476 = ~n592;
  assign n147 = ~n593;
  assign n197 = ~n594;
  assign n413 = ~n595;
  assign n315 = ~n596;
  assign n280 = ~n597;
  assign n207 = ~n598;
  assign n455 = ~n599;
  assign n162 = ~n601;
  assign n511 = ~n602;
  assign n462 = ~n603;
  assign n190 = ~n604;
  assign n294 = ~n606;
  assign n441 = ~n607;
  assign n164 = ~n608;
  assign n420 = ~n609;
  assign n532 = ~n610;
  assign n209 = ~n613;
  assign n273 = ~n614;
  assign n259 = ~n615;
  assign n221 = ~n616;
  assign n287 = ~n617;
  assign n219 = ~n618;
  assign n371 = ~n619;
  assign n469 = ~n620;
  assign n266 = ~n621;
  assign n321 = ~n622;
  assign n181 = ~n623;
  assign n230 = ~n624;
  assign n553 = ~n625;
  assign n336 = ~n626;
  assign n569 = ~n627;
  assign n342 = ~n628;
  assign n546 = ~n629;
  assign n539 = ~n630;
  assign n427 = ~n631;
  assign n350 = ~n632;
  assign n154 = ~n633;
  assign n183 = ~n634;
  assign n357 = ~n635;
  assign n238 = ~n636;
  assign n559 = n307 & n304;
  assign n560 = n321 & n318;
  assign n561 = n328 & n325;
  assign n562 = n342 & n339;
  assign n563 = n133 & n130;
  assign n564 = n142 & n137;
  assign n557 = n569 & n556;
  assign n565 = n147 & n144;
  assign n566 = n154 & n151;
  assign n160 = n162 & n158;
  assign n187 = n183 & n186;
  assign n567 = n209 & n213;
  assign n568 = n569 & n558;
  assign n823 = n557 ^ n558;
  assign n309 = ~n559;
  assign n323 = ~n560;
  assign n330 = ~n561;
  assign n344 = ~n562;
  assign n135 = ~n563;
  assign n140 = ~n564;
  assign n149 = ~n565;
  assign n156 = ~n566;
  assign n211 = ~n567;
  assign n555 = ~n568;
  assign n554 = n555 & n556;
  assign n551 = ~n554;
  assign n548 = n2 ^ n551;
  assign n552 = n551 & n553;
  assign n824 = n66 ^ n548;
  assign n549 = ~n552;
  assign n547 = n549 & n550;
  assign n544 = ~n547;
  assign n541 = n67 ^ n544;
  assign n545 = n544 & n546;
  assign n825 = n3 ^ n541;
  assign n542 = ~n545;
  assign n540 = n542 & n543;
  assign n537 = ~n540;
  assign n533 = n4 ^ n537;
  assign n538 = n537 & n539;
  assign n826 = n68 ^ n533;
  assign n535 = ~n538;
  assign n534 = n535 & n536;
  assign n530 = ~n534;
  assign n527 = n5 ^ n530;
  assign n531 = n530 & n532;
  assign n827 = n69 ^ n527;
  assign n528 = ~n531;
  assign n526 = n528 & n529;
  assign n523 = ~n526;
  assign n520 = n6 ^ n523;
  assign n524 = n523 & n525;
  assign n828 = n70 ^ n520;
  assign n521 = ~n524;
  assign n519 = n521 & n522;
  assign n516 = ~n519;
  assign n513 = n7 ^ n516;
  assign n517 = n516 & n518;
  assign n829 = n71 ^ n513;
  assign n514 = ~n517;
  assign n512 = n514 & n515;
  assign n509 = ~n512;
  assign n506 = n8 ^ n509;
  assign n510 = n509 & n511;
  assign n830 = n72 ^ n506;
  assign n507 = ~n510;
  assign n505 = n507 & n508;
  assign n502 = ~n505;
  assign n499 = n9 ^ n502;
  assign n503 = n502 & n504;
  assign n831 = n73 ^ n499;
  assign n500 = ~n503;
  assign n498 = n500 & n501;
  assign n495 = ~n498;
  assign n492 = n10 ^ n495;
  assign n496 = n495 & n497;
  assign n832 = n74 ^ n492;
  assign n493 = ~n496;
  assign n491 = n493 & n494;
  assign n488 = ~n491;
  assign n485 = n11 ^ n488;
  assign n489 = n488 & n490;
  assign n833 = n75 ^ n485;
  assign n486 = ~n489;
  assign n484 = n486 & n487;
  assign n481 = ~n484;
  assign n477 = n12 ^ n481;
  assign n482 = n481 & n483;
  assign n834 = n76 ^ n477;
  assign n479 = ~n482;
  assign n478 = n479 & n480;
  assign n474 = ~n478;
  assign n471 = n13 ^ n474;
  assign n475 = n474 & n476;
  assign n835 = n77 ^ n471;
  assign n472 = ~n475;
  assign n470 = n472 & n473;
  assign n467 = ~n470;
  assign n464 = n14 ^ n467;
  assign n468 = n467 & n469;
  assign n836 = n78 ^ n464;
  assign n465 = ~n468;
  assign n463 = n465 & n466;
  assign n460 = ~n463;
  assign n457 = n15 ^ n460;
  assign n461 = n460 & n462;
  assign n837 = n79 ^ n457;
  assign n458 = ~n461;
  assign n456 = n458 & n459;
  assign n453 = ~n456;
  assign n450 = n80 ^ n453;
  assign n454 = n453 & n455;
  assign n838 = n16 ^ n450;
  assign n451 = ~n454;
  assign n449 = n451 & n452;
  assign n446 = ~n449;
  assign n443 = n17 ^ n446;
  assign n447 = n446 & n448;
  assign n839 = n81 ^ n443;
  assign n444 = ~n447;
  assign n442 = n444 & n445;
  assign n439 = ~n442;
  assign n436 = n82 ^ n439;
  assign n440 = n439 & n441;
  assign n840 = n18 ^ n436;
  assign n437 = ~n440;
  assign n435 = n437 & n438;
  assign n432 = ~n435;
  assign n429 = n19 ^ n432;
  assign n433 = n432 & n434;
  assign n841 = n83 ^ n429;
  assign n430 = ~n433;
  assign n428 = n430 & n431;
  assign n425 = ~n428;
  assign n421 = n20 ^ n425;
  assign n426 = n425 & n427;
  assign n842 = n84 ^ n421;
  assign n423 = ~n426;
  assign n422 = n423 & n424;
  assign n418 = ~n422;
  assign n414 = n21 ^ n418;
  assign n419 = n418 & n420;
  assign n843 = n85 ^ n414;
  assign n416 = ~n419;
  assign n415 = n416 & n417;
  assign n411 = ~n415;
  assign n407 = n22 ^ n411;
  assign n412 = n411 & n413;
  assign n844 = n86 ^ n407;
  assign n409 = ~n412;
  assign n408 = n409 & n410;
  assign n404 = ~n408;
  assign n400 = n87 ^ n404;
  assign n405 = n404 & n406;
  assign n845 = n23 ^ n400;
  assign n402 = ~n405;
  assign n401 = n402 & n403;
  assign n397 = ~n401;
  assign n393 = n88 ^ n397;
  assign n398 = n397 & n399;
  assign n846 = n24 ^ n393;
  assign n395 = ~n398;
  assign n394 = n395 & n396;
  assign n390 = ~n394;
  assign n387 = n25 ^ n390;
  assign n391 = n390 & n392;
  assign n847 = n89 ^ n387;
  assign n388 = ~n391;
  assign n386 = n388 & n389;
  assign n383 = ~n386;
  assign n380 = n26 ^ n383;
  assign n384 = n383 & n385;
  assign n848 = n90 ^ n380;
  assign n381 = ~n384;
  assign n379 = n381 & n382;
  assign n376 = ~n379;
  assign n373 = n27 ^ n376;
  assign n377 = n376 & n378;
  assign n849 = n91 ^ n373;
  assign n374 = ~n377;
  assign n372 = n374 & n375;
  assign n369 = ~n372;
  assign n366 = n28 ^ n369;
  assign n370 = n369 & n371;
  assign n850 = n92 ^ n366;
  assign n367 = ~n370;
  assign n365 = n367 & n368;
  assign n362 = ~n365;
  assign n359 = n93 ^ n362;
  assign n363 = n362 & n364;
  assign n851 = n29 ^ n359;
  assign n360 = ~n363;
  assign n358 = n360 & n361;
  assign n355 = ~n358;
  assign n352 = n30 ^ n355;
  assign n356 = n355 & n357;
  assign n852 = n94 ^ n352;
  assign n353 = ~n356;
  assign n351 = n353 & n354;
  assign n348 = ~n351;
  assign n345 = n31 ^ n348;
  assign n349 = n348 & n350;
  assign n853 = n95 ^ n345;
  assign n346 = ~n349;
  assign n343 = n346 & n347;
  assign n854 = n343 ^ n344;
  assign n341 = ~n343;
  assign n340 = n341 & n342;
  assign n338 = ~n340;
  assign n337 = n338 & n339;
  assign n334 = ~n337;
  assign n331 = n97 ^ n334;
  assign n335 = n334 & n336;
  assign n855 = n33 ^ n331;
  assign n332 = ~n335;
  assign n329 = n332 & n333;
  assign n856 = n329 ^ n330;
  assign n327 = ~n329;
  assign n326 = n327 & n328;
  assign n324 = ~n326;
  assign n322 = n324 & n325;
  assign n857 = n322 ^ n323;
  assign n320 = ~n322;
  assign n319 = n320 & n321;
  assign n317 = ~n319;
  assign n316 = n317 & n318;
  assign n313 = ~n316;
  assign n310 = n100 ^ n313;
  assign n314 = n313 & n315;
  assign n858 = n36 ^ n310;
  assign n311 = ~n314;
  assign n308 = n311 & n312;
  assign n859 = n308 ^ n309;
  assign n306 = ~n308;
  assign n305 = n306 & n307;
  assign n303 = ~n305;
  assign n302 = n303 & n304;
  assign n299 = ~n302;
  assign n296 = n38 ^ n299;
  assign n300 = n299 & n301;
  assign n860 = n102 ^ n296;
  assign n297 = ~n300;
  assign n295 = n297 & n298;
  assign n292 = ~n295;
  assign n288 = n39 ^ n292;
  assign n293 = n292 & n294;
  assign n861 = n103 ^ n288;
  assign n290 = ~n293;
  assign n289 = n290 & n291;
  assign n285 = ~n289;
  assign n281 = n104 ^ n285;
  assign n286 = n285 & n287;
  assign n862 = n40 ^ n281;
  assign n283 = ~n286;
  assign n282 = n283 & n284;
  assign n278 = ~n282;
  assign n274 = n41 ^ n278;
  assign n279 = n278 & n280;
  assign n863 = n105 ^ n274;
  assign n276 = ~n279;
  assign n275 = n276 & n277;
  assign n271 = ~n275;
  assign n268 = n106 ^ n271;
  assign n272 = n271 & n273;
  assign n864 = n42 ^ n268;
  assign n269 = ~n272;
  assign n267 = n269 & n270;
  assign n264 = ~n267;
  assign n261 = n43 ^ n264;
  assign n265 = n264 & n266;
  assign n865 = n107 ^ n261;
  assign n262 = ~n265;
  assign n260 = n262 & n263;
  assign n257 = ~n260;
  assign n253 = n108 ^ n257;
  assign n258 = n257 & n259;
  assign n866 = n44 ^ n253;
  assign n255 = ~n258;
  assign n254 = n255 & n256;
  assign n250 = ~n254;
  assign n247 = n109 ^ n250;
  assign n251 = n250 & n252;
  assign n867 = n45 ^ n247;
  assign n248 = ~n251;
  assign n246 = n248 & n249;
  assign n243 = ~n246;
  assign n240 = n46 ^ n243;
  assign n244 = n243 & n245;
  assign n868 = n110 ^ n240;
  assign n241 = ~n244;
  assign n239 = n241 & n242;
  assign n236 = ~n239;
  assign n233 = n47 ^ n236;
  assign n237 = n236 & n238;
  assign n869 = n111 ^ n233;
  assign n234 = ~n237;
  assign n231 = n234 & n235;
  assign n870 = n231 ^ n232;
  assign n229 = ~n231;
  assign n228 = n229 & n230;
  assign n226 = ~n228;
  assign n223 = n226 & n227;
  assign n871 = n223 ^ n224;
  assign n222 = n223 & n225;
  assign n220 = ~n222;
  assign n216 = n220 & n221;
  assign n872 = n216 ^ n217;
  assign n218 = n216 & n219;
  assign n214 = ~n218;
  assign n210 = n214 & n215;
  assign n873 = n210 ^ n211;
  assign n212 = n210 & n213;
  assign n208 = ~n212;
  assign n205 = n208 & n209;
  assign n874 = n205 ^ n206;
  assign n204 = n205 & n207;
  assign n202 = ~n204;
  assign n199 = n202 & n203;
  assign n875 = n199 ^ n200;
  assign n198 = n199 & n201;
  assign n196 = ~n198;
  assign n194 = n196 & n197;
  assign n876 = n194 ^ n195;
  assign n192 = ~n194;
  assign n191 = n192 & n193;
  assign n189 = ~n191;
  assign n188 = n189 & n190;
  assign n877 = n187 ^ n188;
  assign n185 = ~n188;
  assign n184 = n185 & n186;
  assign n182 = ~n184;
  assign n179 = n182 & n183;
  assign n878 = n179 ^ n180;
  assign n178 = n179 & n181;
  assign n176 = ~n178;
  assign n175 = n176 & n177;
  assign n172 = ~n175;
  assign n169 = n57 ^ n172;
  assign n173 = n172 & n174;
  assign n879 = n121 ^ n169;
  assign n170 = ~n173;
  assign n166 = n170 & n171;
  assign n880 = n166 ^ n167;
  assign n165 = n166 & n168;
  assign n163 = ~n165;
  assign n161 = n163 & n164;
  assign n881 = n160 ^ n161;
  assign n159 = n161 & n162;
  assign n157 = ~n159;
  assign n155 = n157 & n158;
  assign n882 = n155 ^ n156;
  assign n153 = ~n155;
  assign n152 = n153 & n154;
  assign n150 = ~n152;
  assign n148 = n150 & n151;
  assign n883 = n148 ^ n149;
  assign n146 = ~n148;
  assign n145 = n146 & n147;
  assign n143 = ~n145;
  assign n139 = n143 & n144;
  assign n884 = n139 ^ n140;
  assign n141 = ~n139;
  assign n138 = n141 & n142;
  assign n136 = ~n138;
  assign n134 = n136 & n137;
  assign n885 = n134 ^ n135;
  assign n132 = ~n134;
  assign n131 = n132 & n133;
  assign n129 = ~n131;
  assign n128 = n129 & n130;
  assign n886 = ~n128;
endmodule
