module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63;
  output y0;
  wire n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214;
  assign n65 = x29 & ~x61;
  assign n66 = x28 & ~x60;
  assign n67 = ~n65 & ~n66;
  assign n68 = x30 & ~x62;
  assign n69 = x31 & ~x63;
  assign n70 = ~n68 & ~n69;
  assign n71 = n67 & n70;
  assign n72 = x27 & ~x59;
  assign n73 = ~x26 & ~n72;
  assign n74 = x58 & n73;
  assign n75 = x26 & ~x58;
  assign n76 = ~n72 & ~n75;
  assign n77 = ~x25 & n76;
  assign n78 = x57 & n77;
  assign n79 = ~n74 & ~n78;
  assign n80 = ~x27 & x59;
  assign n81 = x25 & ~x57;
  assign n82 = n76 & ~n81;
  assign n83 = x56 & n82;
  assign n84 = ~x24 & n83;
  assign n85 = ~n80 & ~n84;
  assign n86 = n79 & n85;
  assign n87 = n71 & ~n86;
  assign n88 = ~x24 & n82;
  assign n89 = ~n83 & ~n88;
  assign n90 = n71 & ~n89;
  assign n91 = ~x21 & x53;
  assign n92 = ~x20 & x52;
  assign n93 = ~n91 & ~n92;
  assign n94 = x22 & ~x54;
  assign n95 = x21 & ~x53;
  assign n96 = x23 & ~x55;
  assign n97 = ~n95 & ~n96;
  assign n98 = ~n94 & n97;
  assign n99 = ~n93 & n98;
  assign n100 = x55 ^ x23;
  assign n101 = ~x22 & x54;
  assign n102 = n101 ^ x55;
  assign n103 = ~n100 & ~n102;
  assign n104 = n103 ^ x23;
  assign n105 = ~n99 & n104;
  assign n106 = x20 & ~x52;
  assign n107 = n98 & ~n106;
  assign n108 = ~x16 & x48;
  assign n109 = ~x17 & x49;
  assign n110 = ~n108 & ~n109;
  assign n111 = x18 & ~x50;
  assign n112 = x17 & ~x49;
  assign n113 = x19 & ~x51;
  assign n114 = ~n112 & ~n113;
  assign n115 = ~n111 & n114;
  assign n116 = ~n110 & n115;
  assign n117 = x51 ^ x19;
  assign n118 = ~x18 & x50;
  assign n119 = n118 ^ x51;
  assign n120 = ~n117 & ~n119;
  assign n121 = n120 ^ x19;
  assign n122 = ~n116 & n121;
  assign n123 = n107 & ~n122;
  assign n124 = n105 & ~n123;
  assign n125 = n90 & ~n124;
  assign n126 = ~n87 & ~n125;
  assign n127 = ~x30 & ~n69;
  assign n128 = x62 & n127;
  assign n129 = ~x31 & x63;
  assign n130 = ~x29 & x61;
  assign n131 = ~x28 & ~n65;
  assign n132 = x60 & n131;
  assign n133 = ~n130 & ~n132;
  assign n134 = n70 & ~n133;
  assign n135 = ~n129 & ~n134;
  assign n136 = ~n128 & n135;
  assign n137 = x16 & ~x48;
  assign n138 = ~x15 & x47;
  assign n139 = x15 & ~x47;
  assign n140 = ~x14 & ~n139;
  assign n141 = x46 & n140;
  assign n142 = ~n138 & ~n141;
  assign n143 = x14 & ~x46;
  assign n144 = ~n139 & ~n143;
  assign n145 = ~x13 & x45;
  assign n146 = x13 & ~x45;
  assign n147 = ~x12 & ~n146;
  assign n148 = x44 & n147;
  assign n149 = ~n145 & ~n148;
  assign n150 = n144 & ~n149;
  assign n151 = x12 & ~x44;
  assign n152 = ~n146 & ~n151;
  assign n153 = n144 & n152;
  assign n154 = ~x9 & x41;
  assign n155 = x11 & ~x43;
  assign n156 = x10 & ~x42;
  assign n157 = ~n155 & ~n156;
  assign n158 = n154 & n157;
  assign n159 = ~x10 & ~n155;
  assign n160 = x42 & n159;
  assign n161 = ~n158 & ~n160;
  assign n162 = ~x11 & x43;
  assign n163 = x9 & ~x41;
  assign n164 = x40 & ~n163;
  assign n165 = n157 & n164;
  assign n166 = ~x8 & n165;
  assign n167 = ~n162 & ~n166;
  assign n168 = n161 & n167;
  assign n169 = ~x8 & ~n163;
  assign n170 = n157 & n169;
  assign n171 = ~n165 & ~n170;
  assign n172 = x7 & ~x39;
  assign n173 = ~x6 & ~n172;
  assign n174 = x38 & n173;
  assign n175 = x6 & ~x38;
  assign n176 = ~n172 & ~n175;
  assign n177 = ~x5 & n176;
  assign n178 = x37 & n177;
  assign n179 = ~n174 & ~n178;
  assign n180 = ~x7 & x39;
  assign n181 = x5 & ~x37;
  assign n182 = n176 & ~n181;
  assign n183 = x36 & n182;
  assign n184 = ~x4 & n183;
  assign n185 = ~n180 & ~n184;
  assign n186 = n179 & n185;
  assign n187 = ~x4 & n182;
  assign n188 = ~n183 & ~n187;
  assign n189 = x35 ^ x3;
  assign n190 = x34 ^ x2;
  assign n191 = x33 ^ x1;
  assign n192 = x0 & ~x32;
  assign n193 = n192 ^ x33;
  assign n194 = ~n191 & n193;
  assign n195 = n194 ^ x1;
  assign n196 = n195 ^ x34;
  assign n197 = ~n190 & n196;
  assign n198 = n197 ^ x2;
  assign n199 = n198 ^ x35;
  assign n200 = ~n189 & n199;
  assign n201 = n200 ^ x3;
  assign n202 = ~n188 & ~n201;
  assign n203 = n186 & ~n202;
  assign n204 = ~n171 & ~n203;
  assign n205 = n168 & ~n204;
  assign n206 = n153 & ~n205;
  assign n207 = ~n150 & ~n206;
  assign n208 = n142 & n207;
  assign n209 = ~n137 & ~n208;
  assign n210 = n115 & n209;
  assign n211 = n107 & n210;
  assign n212 = n90 & n211;
  assign n213 = n136 & ~n212;
  assign n214 = n126 & n213;
  assign y0 = ~n214;
endmodule
