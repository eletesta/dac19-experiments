module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63;
  wire n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705;
  assign n65 = x0 & x32;
  assign n76 = x33 & ~n65;
  assign n66 = ~x32 & x33;
  assign n67 = ~x0 & n66;
  assign n69 = x32 & x33;
  assign n68 = x32 & ~x33;
  assign n70 = n69 ^ n68;
  assign n71 = n69 ^ x1;
  assign n72 = n71 ^ n69;
  assign n73 = n70 & n72;
  assign n74 = n73 ^ n69;
  assign n75 = ~n67 & ~n74;
  assign n77 = n76 ^ n75;
  assign n87 = ~n75 & n76;
  assign n84 = x34 ^ x33;
  assign n85 = x0 & n84;
  assign n78 = ~x1 & n66;
  assign n79 = n69 ^ x2;
  assign n80 = n79 ^ n69;
  assign n81 = n70 & n80;
  assign n82 = n81 ^ n69;
  assign n83 = ~n78 & ~n82;
  assign n86 = n85 ^ n83;
  assign n88 = n87 ^ n86;
  assign n114 = ~n83 & n85;
  assign n115 = n83 & ~n85;
  assign n116 = n87 & ~n115;
  assign n117 = ~n114 & ~n116;
  assign n100 = x35 & n84;
  assign n101 = ~x1 & n100;
  assign n102 = x35 ^ x34;
  assign n103 = ~n84 & n102;
  assign n104 = x35 & n103;
  assign n105 = ~x0 & n104;
  assign n106 = ~n101 & ~n105;
  assign n107 = ~x35 & n84;
  assign n108 = x1 & n107;
  assign n109 = ~x35 & n103;
  assign n110 = x0 & n109;
  assign n111 = ~n108 & ~n110;
  assign n112 = n106 & n111;
  assign n95 = x33 ^ x0;
  assign n96 = ~n84 & n95;
  assign n97 = n96 ^ x0;
  assign n98 = x35 & ~n97;
  assign n89 = ~x2 & n66;
  assign n90 = n69 ^ x3;
  assign n91 = n90 ^ n69;
  assign n92 = n70 & n91;
  assign n93 = n92 ^ n69;
  assign n94 = ~n89 & ~n93;
  assign n99 = n98 ^ n94;
  assign n113 = n112 ^ n99;
  assign n118 = n117 ^ n113;
  assign n138 = ~n99 & ~n112;
  assign n139 = n99 & n112;
  assign n140 = ~n117 & ~n139;
  assign n141 = ~n138 & ~n140;
  assign n136 = ~n94 & n98;
  assign n132 = x36 ^ x35;
  assign n133 = x0 & n132;
  assign n125 = x2 & n107;
  assign n126 = x1 & n109;
  assign n127 = ~n125 & ~n126;
  assign n128 = ~x2 & n100;
  assign n129 = ~x1 & n104;
  assign n130 = ~n128 & ~n129;
  assign n131 = n127 & n130;
  assign n134 = n133 ^ n131;
  assign n119 = ~x3 & n66;
  assign n120 = n69 ^ x4;
  assign n121 = n120 ^ n69;
  assign n122 = n70 & n121;
  assign n123 = n122 ^ n69;
  assign n124 = ~n119 & ~n123;
  assign n135 = n134 ^ n124;
  assign n137 = n136 ^ n135;
  assign n142 = n141 ^ n137;
  assign n181 = n135 & n136;
  assign n182 = ~n135 & ~n136;
  assign n183 = ~n141 & ~n182;
  assign n184 = ~n181 & ~n183;
  assign n174 = x35 ^ x0;
  assign n175 = ~n132 & n174;
  assign n176 = n175 ^ x0;
  assign n177 = x37 & ~n176;
  assign n168 = ~x4 & n66;
  assign n169 = n69 ^ x5;
  assign n170 = n169 ^ n69;
  assign n171 = n70 & n170;
  assign n172 = n171 ^ n69;
  assign n173 = ~n168 & ~n172;
  assign n178 = n177 ^ n173;
  assign n160 = x3 & n107;
  assign n161 = x2 & n109;
  assign n162 = ~n160 & ~n161;
  assign n163 = ~x3 & n100;
  assign n164 = ~x2 & n104;
  assign n165 = ~n163 & ~n164;
  assign n166 = n162 & n165;
  assign n147 = x37 & n132;
  assign n148 = ~x1 & n147;
  assign n149 = x37 ^ x36;
  assign n150 = ~n132 & n149;
  assign n151 = x37 & n150;
  assign n152 = ~x0 & n151;
  assign n153 = ~n148 & ~n152;
  assign n154 = ~x37 & n132;
  assign n155 = x1 & n154;
  assign n156 = ~x37 & n150;
  assign n157 = x0 & n156;
  assign n158 = ~n155 & ~n157;
  assign n159 = n153 & n158;
  assign n167 = n166 ^ n159;
  assign n179 = n178 ^ n167;
  assign n143 = n133 ^ n124;
  assign n144 = n131 ^ n124;
  assign n145 = ~n143 & ~n144;
  assign n146 = n145 ^ n133;
  assign n180 = n179 ^ n146;
  assign n185 = n184 ^ n180;
  assign n217 = n146 & ~n179;
  assign n218 = ~n146 & n179;
  assign n219 = ~n184 & ~n218;
  assign n220 = ~n217 & ~n219;
  assign n211 = x38 ^ x37;
  assign n212 = x0 & n211;
  assign n205 = ~x5 & n66;
  assign n206 = n69 ^ x6;
  assign n207 = n206 ^ n69;
  assign n208 = n70 & n207;
  assign n209 = n208 ^ n69;
  assign n210 = ~n205 & ~n209;
  assign n213 = n212 ^ n210;
  assign n198 = ~x4 & n100;
  assign n199 = ~x3 & n104;
  assign n200 = ~n198 & ~n199;
  assign n201 = x4 & n107;
  assign n202 = x3 & n109;
  assign n203 = ~n201 & ~n202;
  assign n204 = n200 & n203;
  assign n214 = n213 ^ n204;
  assign n190 = ~x2 & n147;
  assign n191 = ~x1 & n151;
  assign n192 = ~n190 & ~n191;
  assign n193 = x2 & n154;
  assign n194 = x1 & n156;
  assign n195 = ~n193 & ~n194;
  assign n196 = n192 & n195;
  assign n189 = ~n173 & n177;
  assign n197 = n196 ^ n189;
  assign n215 = n214 ^ n197;
  assign n186 = n178 ^ n159;
  assign n187 = n167 & ~n186;
  assign n188 = n187 ^ n166;
  assign n216 = n215 ^ n188;
  assign n221 = n220 ^ n216;
  assign n271 = ~n188 & ~n215;
  assign n272 = n188 & n215;
  assign n273 = ~n220 & ~n272;
  assign n274 = ~n271 & ~n273;
  assign n261 = x3 & n154;
  assign n262 = x2 & n156;
  assign n263 = ~n261 & ~n262;
  assign n264 = ~x3 & n147;
  assign n265 = ~x2 & n151;
  assign n266 = ~n264 & ~n265;
  assign n267 = n263 & n266;
  assign n247 = x39 & n211;
  assign n248 = ~x1 & n247;
  assign n249 = x39 ^ x38;
  assign n250 = ~n211 & n249;
  assign n251 = x39 & n250;
  assign n252 = ~x0 & n251;
  assign n253 = ~n248 & ~n252;
  assign n254 = ~x39 & n211;
  assign n255 = x1 & n254;
  assign n256 = ~x39 & n250;
  assign n257 = x0 & n256;
  assign n258 = ~n255 & ~n257;
  assign n259 = n253 & n258;
  assign n240 = x5 & n107;
  assign n241 = x4 & n109;
  assign n242 = ~n240 & ~n241;
  assign n243 = ~x5 & n100;
  assign n244 = ~x4 & n104;
  assign n245 = ~n243 & ~n244;
  assign n246 = n242 & n245;
  assign n260 = n259 ^ n246;
  assign n268 = n267 ^ n260;
  assign n234 = x37 ^ x0;
  assign n235 = ~n211 & n234;
  assign n236 = n235 ^ x0;
  assign n237 = x39 & ~n236;
  assign n228 = ~x6 & n66;
  assign n229 = n69 ^ x7;
  assign n230 = n229 ^ n69;
  assign n231 = n70 & n230;
  assign n232 = n231 ^ n69;
  assign n233 = ~n228 & ~n232;
  assign n238 = n237 ^ n233;
  assign n225 = n210 ^ n204;
  assign n226 = ~n213 & ~n225;
  assign n227 = n226 ^ n212;
  assign n239 = n238 ^ n227;
  assign n269 = n268 ^ n239;
  assign n222 = n214 ^ n189;
  assign n223 = ~n197 & ~n222;
  assign n224 = n223 ^ n196;
  assign n270 = n269 ^ n224;
  assign n275 = n274 ^ n270;
  assign n321 = ~n224 & n269;
  assign n322 = n224 & ~n269;
  assign n323 = ~n274 & ~n322;
  assign n324 = ~n321 & ~n323;
  assign n317 = ~n233 & n237;
  assign n309 = ~x6 & n100;
  assign n310 = ~x5 & n104;
  assign n311 = ~n309 & ~n310;
  assign n312 = x6 & n107;
  assign n313 = x5 & n109;
  assign n314 = ~n312 & ~n313;
  assign n315 = n311 & n314;
  assign n302 = ~x4 & n147;
  assign n303 = ~x3 & n151;
  assign n304 = ~n302 & ~n303;
  assign n305 = x4 & n154;
  assign n306 = x3 & n156;
  assign n307 = ~n305 & ~n306;
  assign n308 = n304 & n307;
  assign n316 = n315 ^ n308;
  assign n318 = n317 ^ n316;
  assign n297 = x40 ^ x39;
  assign n298 = x0 & n297;
  assign n291 = ~x7 & n66;
  assign n292 = n69 ^ x8;
  assign n293 = n292 ^ n69;
  assign n294 = n70 & n293;
  assign n295 = n294 ^ n69;
  assign n296 = ~n291 & ~n295;
  assign n299 = n298 ^ n296;
  assign n284 = ~x2 & n247;
  assign n285 = ~x1 & n251;
  assign n286 = ~n284 & ~n285;
  assign n287 = x2 & n254;
  assign n288 = x1 & n256;
  assign n289 = ~n287 & ~n288;
  assign n290 = n286 & n289;
  assign n300 = n299 ^ n290;
  assign n280 = n267 ^ n259;
  assign n281 = n267 ^ n246;
  assign n282 = n280 & ~n281;
  assign n283 = n282 ^ n259;
  assign n301 = n300 ^ n283;
  assign n319 = n318 ^ n301;
  assign n276 = n268 ^ n238;
  assign n277 = n268 ^ n227;
  assign n278 = n276 & n277;
  assign n279 = n278 ^ n238;
  assign n320 = n319 ^ n279;
  assign n325 = n324 ^ n320;
  assign n388 = ~n279 & ~n319;
  assign n389 = n279 & n319;
  assign n390 = ~n324 & ~n389;
  assign n391 = ~n388 & ~n390;
  assign n377 = x5 & n154;
  assign n378 = x4 & n156;
  assign n379 = ~n377 & ~n378;
  assign n380 = ~x5 & n147;
  assign n381 = ~x4 & n151;
  assign n382 = ~n380 & ~n381;
  assign n383 = n379 & n382;
  assign n372 = x39 ^ x0;
  assign n373 = ~n297 & n372;
  assign n374 = n373 ^ x0;
  assign n375 = x41 & ~n374;
  assign n365 = ~x7 & n100;
  assign n366 = ~x6 & n104;
  assign n367 = ~n365 & ~n366;
  assign n368 = x7 & n107;
  assign n369 = x6 & n109;
  assign n370 = ~n368 & ~n369;
  assign n371 = n367 & n370;
  assign n376 = n375 ^ n371;
  assign n384 = n383 ^ n376;
  assign n362 = n296 ^ n290;
  assign n363 = ~n299 & ~n362;
  assign n364 = n363 ^ n298;
  assign n385 = n384 ^ n364;
  assign n346 = x41 & n297;
  assign n347 = ~x1 & n346;
  assign n348 = x41 ^ x40;
  assign n349 = ~n297 & n348;
  assign n350 = x41 & n349;
  assign n351 = ~x0 & n350;
  assign n352 = ~n347 & ~n351;
  assign n353 = ~x41 & n297;
  assign n354 = x1 & n353;
  assign n355 = ~x41 & n349;
  assign n356 = x0 & n355;
  assign n357 = ~n354 & ~n356;
  assign n358 = n352 & n357;
  assign n339 = ~x3 & n247;
  assign n340 = ~x2 & n251;
  assign n341 = ~n339 & ~n340;
  assign n342 = x3 & n254;
  assign n343 = x2 & n256;
  assign n344 = ~n342 & ~n343;
  assign n345 = n341 & n344;
  assign n359 = n358 ^ n345;
  assign n333 = ~x8 & n66;
  assign n334 = n69 ^ x9;
  assign n335 = n334 ^ n69;
  assign n336 = n70 & n335;
  assign n337 = n336 ^ n69;
  assign n338 = ~n333 & ~n337;
  assign n360 = n359 ^ n338;
  assign n330 = n317 ^ n308;
  assign n331 = n316 & n330;
  assign n332 = n331 ^ n315;
  assign n361 = n360 ^ n332;
  assign n386 = n385 ^ n361;
  assign n326 = n318 ^ n300;
  assign n327 = n318 ^ n283;
  assign n328 = n326 & n327;
  assign n329 = n328 ^ n300;
  assign n387 = n386 ^ n329;
  assign n392 = n391 ^ n387;
  assign n449 = n329 & n386;
  assign n450 = ~n329 & ~n386;
  assign n451 = ~n391 & ~n450;
  assign n452 = ~n449 & ~n451;
  assign n438 = x4 & n254;
  assign n439 = x3 & n256;
  assign n440 = ~n438 & ~n439;
  assign n441 = ~x4 & n247;
  assign n442 = ~x3 & n251;
  assign n443 = ~n441 & ~n442;
  assign n444 = n440 & n443;
  assign n435 = x42 ^ x41;
  assign n436 = x0 & n435;
  assign n428 = ~x8 & n100;
  assign n429 = ~x7 & n104;
  assign n430 = ~n428 & ~n429;
  assign n431 = x8 & n107;
  assign n432 = x7 & n109;
  assign n433 = ~n431 & ~n432;
  assign n434 = n430 & n433;
  assign n437 = n436 ^ n434;
  assign n445 = n444 ^ n437;
  assign n426 = ~n371 & n375;
  assign n423 = n358 ^ n338;
  assign n424 = ~n359 & n423;
  assign n425 = n424 ^ n338;
  assign n427 = n426 ^ n425;
  assign n446 = n445 ^ n427;
  assign n414 = ~x6 & n147;
  assign n415 = ~x5 & n151;
  assign n416 = ~n414 & ~n415;
  assign n417 = x6 & n154;
  assign n418 = x5 & n156;
  assign n419 = ~n417 & ~n418;
  assign n420 = n416 & n419;
  assign n406 = ~x2 & n346;
  assign n407 = ~x1 & n350;
  assign n408 = ~n406 & ~n407;
  assign n409 = x2 & n353;
  assign n410 = x1 & n355;
  assign n411 = ~n409 & ~n410;
  assign n412 = n408 & n411;
  assign n400 = ~x9 & n66;
  assign n401 = n69 ^ x10;
  assign n402 = n401 ^ n69;
  assign n403 = n70 & n402;
  assign n404 = n403 ^ n69;
  assign n405 = ~n400 & ~n404;
  assign n413 = n412 ^ n405;
  assign n421 = n420 ^ n413;
  assign n397 = n376 ^ n364;
  assign n398 = n384 & n397;
  assign n399 = n398 ^ n383;
  assign n422 = n421 ^ n399;
  assign n447 = n446 ^ n422;
  assign n393 = n385 ^ n360;
  assign n394 = n385 ^ n332;
  assign n395 = ~n393 & n394;
  assign n396 = n395 ^ n360;
  assign n448 = n447 ^ n396;
  assign n453 = n452 ^ n448;
  assign n528 = ~n396 & ~n447;
  assign n529 = n396 & n447;
  assign n530 = ~n452 & ~n529;
  assign n531 = ~n528 & ~n530;
  assign n516 = ~x7 & n147;
  assign n517 = ~x6 & n151;
  assign n518 = ~n516 & ~n517;
  assign n519 = x7 & n154;
  assign n520 = x6 & n156;
  assign n521 = ~n519 & ~n520;
  assign n522 = n518 & n521;
  assign n503 = ~x43 & n435;
  assign n504 = x1 & n503;
  assign n505 = x43 ^ x42;
  assign n506 = ~n435 & n505;
  assign n507 = ~x43 & n506;
  assign n508 = x0 & n507;
  assign n509 = ~n504 & ~n508;
  assign n510 = x43 & n435;
  assign n511 = ~x1 & n510;
  assign n512 = x43 & n506;
  assign n513 = ~x0 & n512;
  assign n514 = ~n511 & ~n513;
  assign n515 = n509 & n514;
  assign n523 = n522 ^ n515;
  assign n498 = x41 ^ x0;
  assign n499 = ~n435 & n498;
  assign n500 = n499 ^ x0;
  assign n501 = x43 & ~n500;
  assign n491 = x9 & n107;
  assign n492 = x8 & n109;
  assign n493 = ~n491 & ~n492;
  assign n494 = ~x9 & n100;
  assign n495 = ~x8 & n104;
  assign n496 = ~n494 & ~n495;
  assign n497 = n493 & n496;
  assign n502 = n501 ^ n497;
  assign n524 = n523 ^ n502;
  assign n486 = n420 ^ n412;
  assign n487 = n413 & ~n486;
  assign n488 = n487 ^ n405;
  assign n483 = n444 ^ n434;
  assign n484 = ~n437 & ~n483;
  assign n485 = n484 ^ n436;
  assign n489 = n488 ^ n485;
  assign n474 = ~x5 & n247;
  assign n475 = ~x4 & n251;
  assign n476 = ~n474 & ~n475;
  assign n477 = x5 & n254;
  assign n478 = x4 & n256;
  assign n479 = ~n477 & ~n478;
  assign n480 = n476 & n479;
  assign n467 = ~x3 & n346;
  assign n468 = ~x2 & n350;
  assign n469 = ~n467 & ~n468;
  assign n470 = x3 & n353;
  assign n471 = x2 & n355;
  assign n472 = ~n470 & ~n471;
  assign n473 = n469 & n472;
  assign n481 = n480 ^ n473;
  assign n461 = ~x10 & n66;
  assign n462 = n69 ^ x11;
  assign n463 = n462 ^ n69;
  assign n464 = n70 & n463;
  assign n465 = n464 ^ n69;
  assign n466 = ~n461 & ~n465;
  assign n482 = n481 ^ n466;
  assign n490 = n489 ^ n482;
  assign n525 = n524 ^ n490;
  assign n458 = n445 ^ n426;
  assign n459 = n427 & n458;
  assign n460 = n459 ^ n445;
  assign n526 = n525 ^ n460;
  assign n454 = n446 ^ n421;
  assign n455 = n446 ^ n399;
  assign n456 = n454 & ~n455;
  assign n457 = n456 ^ n421;
  assign n527 = n526 ^ n457;
  assign n532 = n531 ^ n527;
  assign n600 = ~n457 & ~n526;
  assign n601 = n457 & n526;
  assign n602 = ~n531 & ~n601;
  assign n603 = ~n600 & ~n602;
  assign n588 = ~x6 & n247;
  assign n589 = ~x5 & n251;
  assign n590 = ~n588 & ~n589;
  assign n591 = x6 & n254;
  assign n592 = x5 & n256;
  assign n593 = ~n591 & ~n592;
  assign n594 = n590 & n593;
  assign n585 = x44 ^ x43;
  assign n586 = x0 & n585;
  assign n578 = x10 & n107;
  assign n579 = x9 & n109;
  assign n580 = ~n578 & ~n579;
  assign n581 = ~x10 & n100;
  assign n582 = ~x9 & n104;
  assign n583 = ~n581 & ~n582;
  assign n584 = n580 & n583;
  assign n587 = n586 ^ n584;
  assign n595 = n594 ^ n587;
  assign n570 = x2 & n503;
  assign n571 = x1 & n507;
  assign n572 = ~n570 & ~n571;
  assign n573 = ~x2 & n510;
  assign n574 = ~x1 & n512;
  assign n575 = ~n573 & ~n574;
  assign n576 = n572 & n575;
  assign n562 = ~x4 & n346;
  assign n563 = ~x3 & n350;
  assign n564 = ~n562 & ~n563;
  assign n565 = x4 & n353;
  assign n566 = x3 & n355;
  assign n567 = ~n565 & ~n566;
  assign n568 = n564 & n567;
  assign n556 = ~x11 & n66;
  assign n557 = n69 ^ x12;
  assign n558 = n557 ^ n69;
  assign n559 = n70 & n558;
  assign n560 = n559 ^ n69;
  assign n561 = ~n556 & ~n560;
  assign n569 = n568 ^ n561;
  assign n577 = n576 ^ n569;
  assign n596 = n595 ^ n577;
  assign n553 = n515 ^ n502;
  assign n554 = n523 & ~n553;
  assign n555 = n554 ^ n522;
  assign n597 = n596 ^ n555;
  assign n543 = ~x8 & n147;
  assign n544 = ~x7 & n151;
  assign n545 = ~n543 & ~n544;
  assign n546 = x8 & n154;
  assign n547 = x7 & n156;
  assign n548 = ~n546 & ~n547;
  assign n549 = n545 & n548;
  assign n542 = ~n497 & n501;
  assign n550 = n549 ^ n542;
  assign n539 = n480 ^ n466;
  assign n540 = ~n481 & n539;
  assign n541 = n540 ^ n466;
  assign n551 = n550 ^ n541;
  assign n536 = n488 ^ n482;
  assign n537 = n489 & n536;
  assign n538 = n537 ^ n482;
  assign n552 = n551 ^ n538;
  assign n598 = n597 ^ n552;
  assign n533 = n490 ^ n460;
  assign n534 = ~n525 & ~n533;
  assign n535 = n534 ^ n524;
  assign n599 = n598 ^ n535;
  assign n604 = n603 ^ n599;
  assign n691 = ~n535 & ~n598;
  assign n692 = n535 & n598;
  assign n693 = ~n603 & ~n692;
  assign n694 = ~n691 & ~n693;
  assign n679 = x5 & n353;
  assign n680 = x4 & n355;
  assign n681 = ~n679 & ~n680;
  assign n682 = ~x5 & n346;
  assign n683 = ~x4 & n350;
  assign n684 = ~n682 & ~n683;
  assign n685 = n681 & n684;
  assign n671 = x7 & n254;
  assign n672 = x6 & n256;
  assign n673 = ~n671 & ~n672;
  assign n674 = ~x7 & n247;
  assign n675 = ~x6 & n251;
  assign n676 = ~n674 & ~n675;
  assign n677 = n673 & n676;
  assign n664 = ~x11 & n100;
  assign n665 = ~x10 & n104;
  assign n666 = ~n664 & ~n665;
  assign n667 = x11 & n107;
  assign n668 = x10 & n109;
  assign n669 = ~n667 & ~n668;
  assign n670 = n666 & n669;
  assign n678 = n677 ^ n670;
  assign n686 = n685 ^ n678;
  assign n650 = x45 & n585;
  assign n651 = ~x1 & n650;
  assign n652 = x45 ^ x44;
  assign n653 = ~n585 & n652;
  assign n654 = x45 & n653;
  assign n655 = ~x0 & n654;
  assign n656 = ~n651 & ~n655;
  assign n657 = ~x45 & n585;
  assign n658 = x1 & n657;
  assign n659 = ~x45 & n653;
  assign n660 = x0 & n659;
  assign n661 = ~n658 & ~n660;
  assign n662 = n656 & n661;
  assign n642 = ~x9 & n147;
  assign n643 = ~x8 & n151;
  assign n644 = ~n642 & ~n643;
  assign n645 = x9 & n154;
  assign n646 = x8 & n156;
  assign n647 = ~n645 & ~n646;
  assign n648 = n644 & n647;
  assign n635 = x3 & n503;
  assign n636 = x2 & n507;
  assign n637 = ~n635 & ~n636;
  assign n638 = ~x3 & n510;
  assign n639 = ~x2 & n512;
  assign n640 = ~n638 & ~n639;
  assign n641 = n637 & n640;
  assign n649 = n648 ^ n641;
  assign n663 = n662 ^ n649;
  assign n687 = n686 ^ n663;
  assign n632 = n542 ^ n541;
  assign n633 = ~n550 & n632;
  assign n634 = n633 ^ n549;
  assign n688 = n687 ^ n634;
  assign n624 = x43 ^ x0;
  assign n625 = ~n585 & n624;
  assign n626 = n625 ^ x0;
  assign n627 = x45 & ~n626;
  assign n618 = ~x12 & n66;
  assign n619 = n69 ^ x13;
  assign n620 = n619 ^ n69;
  assign n621 = n70 & n620;
  assign n622 = n621 ^ n69;
  assign n623 = ~n618 & ~n622;
  assign n628 = n627 ^ n623;
  assign n614 = n594 ^ n586;
  assign n615 = n594 ^ n584;
  assign n616 = ~n614 & ~n615;
  assign n617 = n616 ^ n586;
  assign n629 = n628 ^ n617;
  assign n611 = n576 ^ n568;
  assign n612 = n569 & ~n611;
  assign n613 = n612 ^ n561;
  assign n630 = n629 ^ n613;
  assign n608 = n577 ^ n555;
  assign n609 = ~n596 & ~n608;
  assign n610 = n609 ^ n595;
  assign n631 = n630 ^ n610;
  assign n689 = n688 ^ n631;
  assign n605 = n597 ^ n551;
  assign n606 = n552 & n605;
  assign n607 = n606 ^ n597;
  assign n690 = n689 ^ n607;
  assign n695 = n694 ^ n690;
  assign n775 = n607 & ~n689;
  assign n776 = ~n607 & n689;
  assign n777 = ~n694 & ~n776;
  assign n778 = ~n775 & ~n777;
  assign n767 = x46 ^ x45;
  assign n768 = x0 & n767;
  assign n761 = ~x13 & n66;
  assign n762 = n69 ^ x14;
  assign n763 = n762 ^ n69;
  assign n764 = n70 & n763;
  assign n765 = n764 ^ n69;
  assign n766 = ~n761 & ~n765;
  assign n769 = n768 ^ n766;
  assign n754 = ~x12 & n100;
  assign n755 = ~x11 & n104;
  assign n756 = ~n754 & ~n755;
  assign n757 = x12 & n107;
  assign n758 = x11 & n109;
  assign n759 = ~n757 & ~n758;
  assign n760 = n756 & n759;
  assign n770 = n769 ^ n760;
  assign n750 = n685 ^ n670;
  assign n751 = n678 & ~n750;
  assign n752 = n751 ^ n677;
  assign n747 = n662 ^ n641;
  assign n748 = n649 & ~n747;
  assign n749 = n748 ^ n648;
  assign n753 = n752 ^ n749;
  assign n771 = n770 ^ n753;
  assign n737 = x10 & n154;
  assign n738 = x9 & n156;
  assign n739 = ~n737 & ~n738;
  assign n740 = ~x10 & n147;
  assign n741 = ~x9 & n151;
  assign n742 = ~n740 & ~n741;
  assign n743 = n739 & n742;
  assign n729 = x8 & n254;
  assign n730 = x7 & n256;
  assign n731 = ~n729 & ~n730;
  assign n732 = ~x8 & n247;
  assign n733 = ~x7 & n251;
  assign n734 = ~n732 & ~n733;
  assign n735 = n731 & n734;
  assign n722 = ~x6 & n346;
  assign n723 = ~x5 & n350;
  assign n724 = ~n722 & ~n723;
  assign n725 = x6 & n353;
  assign n726 = x5 & n355;
  assign n727 = ~n725 & ~n726;
  assign n728 = n724 & n727;
  assign n736 = n735 ^ n728;
  assign n744 = n743 ^ n736;
  assign n720 = ~n623 & n627;
  assign n712 = x4 & n503;
  assign n713 = x3 & n507;
  assign n714 = ~n712 & ~n713;
  assign n715 = ~x4 & n510;
  assign n716 = ~x3 & n512;
  assign n717 = ~n715 & ~n716;
  assign n718 = n714 & n717;
  assign n705 = x2 & n657;
  assign n706 = x1 & n659;
  assign n707 = ~n705 & ~n706;
  assign n708 = ~x2 & n650;
  assign n709 = ~x1 & n654;
  assign n710 = ~n708 & ~n709;
  assign n711 = n707 & n710;
  assign n719 = n718 ^ n711;
  assign n721 = n720 ^ n719;
  assign n745 = n744 ^ n721;
  assign n702 = n617 ^ n613;
  assign n703 = ~n629 & n702;
  assign n704 = n703 ^ n628;
  assign n746 = n745 ^ n704;
  assign n772 = n771 ^ n746;
  assign n699 = n663 ^ n634;
  assign n700 = n687 & ~n699;
  assign n701 = n700 ^ n686;
  assign n773 = n772 ^ n701;
  assign n696 = n688 ^ n610;
  assign n697 = n631 & n696;
  assign n698 = n697 ^ n630;
  assign n774 = n773 ^ n698;
  assign n779 = n778 ^ n774;
  assign n878 = n698 & ~n773;
  assign n879 = ~n698 & n773;
  assign n880 = ~n778 & ~n879;
  assign n881 = ~n878 & ~n880;
  assign n865 = ~x3 & n650;
  assign n866 = ~x2 & n654;
  assign n867 = ~n865 & ~n866;
  assign n868 = x3 & n657;
  assign n869 = x2 & n659;
  assign n870 = ~n868 & ~n869;
  assign n871 = n867 & n870;
  assign n860 = x45 ^ x0;
  assign n861 = ~n767 & n860;
  assign n862 = n861 ^ x0;
  assign n863 = x47 & ~n862;
  assign n854 = ~x14 & n66;
  assign n855 = n69 ^ x15;
  assign n856 = n855 ^ n69;
  assign n857 = n70 & n856;
  assign n858 = n857 ^ n69;
  assign n859 = ~n854 & ~n858;
  assign n864 = n863 ^ n859;
  assign n872 = n871 ^ n864;
  assign n851 = n766 ^ n760;
  assign n852 = ~n769 & ~n851;
  assign n853 = n852 ^ n768;
  assign n873 = n872 ^ n853;
  assign n848 = n720 ^ n711;
  assign n849 = n719 & n848;
  assign n850 = n849 ^ n718;
  assign n874 = n873 ^ n850;
  assign n845 = n770 ^ n752;
  assign n846 = ~n753 & ~n845;
  assign n847 = n846 ^ n770;
  assign n875 = n874 ^ n847;
  assign n835 = x9 & n254;
  assign n836 = x8 & n256;
  assign n837 = ~n835 & ~n836;
  assign n838 = ~x9 & n247;
  assign n839 = ~x8 & n251;
  assign n840 = ~n838 & ~n839;
  assign n841 = n837 & n840;
  assign n827 = ~x13 & n100;
  assign n828 = ~x12 & n104;
  assign n829 = ~n827 & ~n828;
  assign n830 = x13 & n107;
  assign n831 = x12 & n109;
  assign n832 = ~n830 & ~n831;
  assign n833 = n829 & n832;
  assign n814 = ~x47 & n767;
  assign n815 = x1 & n814;
  assign n816 = x47 ^ x46;
  assign n817 = ~n767 & n816;
  assign n818 = ~x47 & n817;
  assign n819 = x0 & n818;
  assign n820 = ~n815 & ~n819;
  assign n821 = x47 & n767;
  assign n822 = ~x1 & n821;
  assign n823 = x47 & n817;
  assign n824 = ~x0 & n823;
  assign n825 = ~n822 & ~n824;
  assign n826 = n820 & n825;
  assign n834 = n833 ^ n826;
  assign n842 = n841 ^ n834;
  assign n805 = x5 & n503;
  assign n806 = x4 & n507;
  assign n807 = ~n805 & ~n806;
  assign n808 = ~x5 & n510;
  assign n809 = ~x4 & n512;
  assign n810 = ~n808 & ~n809;
  assign n811 = n807 & n810;
  assign n797 = ~x7 & n346;
  assign n798 = ~x6 & n350;
  assign n799 = ~n797 & ~n798;
  assign n800 = x7 & n353;
  assign n801 = x6 & n355;
  assign n802 = ~n800 & ~n801;
  assign n803 = n799 & n802;
  assign n790 = ~x11 & n147;
  assign n791 = ~x10 & n151;
  assign n792 = ~n790 & ~n791;
  assign n793 = x11 & n154;
  assign n794 = x10 & n156;
  assign n795 = ~n793 & ~n794;
  assign n796 = n792 & n795;
  assign n804 = n803 ^ n796;
  assign n812 = n811 ^ n804;
  assign n786 = n743 ^ n735;
  assign n787 = n743 ^ n728;
  assign n788 = n786 & ~n787;
  assign n789 = n788 ^ n735;
  assign n813 = n812 ^ n789;
  assign n843 = n842 ^ n813;
  assign n783 = n721 ^ n704;
  assign n784 = ~n745 & n783;
  assign n785 = n784 ^ n744;
  assign n844 = n843 ^ n785;
  assign n876 = n875 ^ n844;
  assign n780 = n746 ^ n701;
  assign n781 = n772 & n780;
  assign n782 = n781 ^ n771;
  assign n877 = n876 ^ n782;
  assign n882 = n881 ^ n877;
  assign n977 = n782 & ~n876;
  assign n978 = ~n782 & n876;
  assign n979 = ~n881 & ~n978;
  assign n980 = ~n977 & ~n979;
  assign n970 = ~n859 & n863;
  assign n967 = n841 ^ n826;
  assign n968 = n834 & ~n967;
  assign n969 = n968 ^ n833;
  assign n971 = n970 ^ n969;
  assign n963 = n811 ^ n803;
  assign n964 = n811 ^ n796;
  assign n965 = n963 & ~n964;
  assign n966 = n965 ^ n803;
  assign n972 = n971 ^ n966;
  assign n960 = n864 ^ n853;
  assign n961 = n872 & n960;
  assign n962 = n961 ^ n871;
  assign n973 = n972 ^ n962;
  assign n956 = n842 ^ n812;
  assign n957 = n842 ^ n789;
  assign n958 = n956 & ~n957;
  assign n959 = n958 ^ n812;
  assign n974 = n973 ^ n959;
  assign n946 = x8 & n353;
  assign n947 = x7 & n355;
  assign n948 = ~n946 & ~n947;
  assign n949 = ~x8 & n346;
  assign n950 = ~x7 & n350;
  assign n951 = ~n949 & ~n950;
  assign n952 = n948 & n951;
  assign n938 = ~x2 & n821;
  assign n939 = ~x1 & n823;
  assign n940 = ~n938 & ~n939;
  assign n941 = x2 & n814;
  assign n942 = x1 & n818;
  assign n943 = ~n941 & ~n942;
  assign n944 = n940 & n943;
  assign n931 = x10 & n254;
  assign n932 = x9 & n256;
  assign n933 = ~n931 & ~n932;
  assign n934 = ~x10 & n247;
  assign n935 = ~x9 & n251;
  assign n936 = ~n934 & ~n935;
  assign n937 = n933 & n936;
  assign n945 = n944 ^ n937;
  assign n953 = n952 ^ n945;
  assign n926 = x48 ^ x47;
  assign n927 = x0 & n926;
  assign n920 = ~x15 & n66;
  assign n921 = n69 ^ x16;
  assign n922 = n921 ^ n69;
  assign n923 = n70 & n922;
  assign n924 = n923 ^ n69;
  assign n925 = ~n920 & ~n924;
  assign n928 = n927 ^ n925;
  assign n913 = ~x14 & n100;
  assign n914 = ~x13 & n104;
  assign n915 = ~n913 & ~n914;
  assign n916 = x14 & n107;
  assign n917 = x13 & n109;
  assign n918 = ~n916 & ~n917;
  assign n919 = n915 & n918;
  assign n929 = n928 ^ n919;
  assign n905 = x4 & n657;
  assign n906 = x3 & n659;
  assign n907 = ~n905 & ~n906;
  assign n908 = ~x4 & n650;
  assign n909 = ~x3 & n654;
  assign n910 = ~n908 & ~n909;
  assign n911 = n907 & n910;
  assign n897 = x12 & n154;
  assign n898 = x11 & n156;
  assign n899 = ~n897 & ~n898;
  assign n900 = ~x12 & n147;
  assign n901 = ~x11 & n151;
  assign n902 = ~n900 & ~n901;
  assign n903 = n899 & n902;
  assign n890 = ~x6 & n510;
  assign n891 = ~x5 & n512;
  assign n892 = ~n890 & ~n891;
  assign n893 = x6 & n503;
  assign n894 = x5 & n507;
  assign n895 = ~n893 & ~n894;
  assign n896 = n892 & n895;
  assign n904 = n903 ^ n896;
  assign n912 = n911 ^ n904;
  assign n930 = n929 ^ n912;
  assign n954 = n953 ^ n930;
  assign n887 = n850 ^ n847;
  assign n888 = ~n874 & n887;
  assign n889 = n888 ^ n873;
  assign n955 = n954 ^ n889;
  assign n975 = n974 ^ n955;
  assign n883 = n875 ^ n843;
  assign n884 = n875 ^ n785;
  assign n885 = n883 & ~n884;
  assign n886 = n885 ^ n843;
  assign n976 = n975 ^ n886;
  assign n981 = n980 ^ n976;
  assign n1092 = ~n886 & n975;
  assign n1093 = n886 & ~n975;
  assign n1094 = ~n980 & ~n1093;
  assign n1095 = ~n1092 & ~n1094;
  assign n1083 = n925 ^ n919;
  assign n1084 = ~n928 & ~n1083;
  assign n1085 = n1084 ^ n927;
  assign n1080 = n911 ^ n903;
  assign n1081 = ~n904 & n1080;
  assign n1082 = n1081 ^ n911;
  assign n1086 = n1085 ^ n1082;
  assign n1077 = n952 ^ n937;
  assign n1078 = n945 & ~n1077;
  assign n1079 = n1078 ^ n944;
  assign n1087 = n1086 ^ n1079;
  assign n1074 = n969 ^ n966;
  assign n1075 = ~n971 & ~n1074;
  assign n1076 = n1075 ^ n970;
  assign n1088 = n1087 ^ n1076;
  assign n1071 = n953 ^ n912;
  assign n1072 = ~n930 & ~n1071;
  assign n1073 = n1072 ^ n929;
  assign n1089 = n1088 ^ n1073;
  assign n1063 = x47 ^ x0;
  assign n1064 = ~n926 & n1063;
  assign n1065 = n1064 ^ x0;
  assign n1066 = x49 & ~n1065;
  assign n1057 = ~x16 & n66;
  assign n1058 = n69 ^ x17;
  assign n1059 = n1058 ^ n69;
  assign n1060 = n70 & n1059;
  assign n1061 = n1060 ^ n69;
  assign n1062 = ~n1057 & ~n1061;
  assign n1067 = n1066 ^ n1062;
  assign n1049 = x5 & n657;
  assign n1050 = x4 & n659;
  assign n1051 = ~n1049 & ~n1050;
  assign n1052 = ~x5 & n650;
  assign n1053 = ~x4 & n654;
  assign n1054 = ~n1052 & ~n1053;
  assign n1055 = n1051 & n1054;
  assign n1042 = ~x7 & n510;
  assign n1043 = ~x6 & n512;
  assign n1044 = ~n1042 & ~n1043;
  assign n1045 = x7 & n503;
  assign n1046 = x6 & n507;
  assign n1047 = ~n1045 & ~n1046;
  assign n1048 = n1044 & n1047;
  assign n1056 = n1055 ^ n1048;
  assign n1068 = n1067 ^ n1056;
  assign n1033 = ~x13 & n147;
  assign n1034 = ~x12 & n151;
  assign n1035 = ~n1033 & ~n1034;
  assign n1036 = x13 & n154;
  assign n1037 = x12 & n156;
  assign n1038 = ~n1036 & ~n1037;
  assign n1039 = n1035 & n1038;
  assign n1025 = x15 & n107;
  assign n1026 = x14 & n109;
  assign n1027 = ~n1025 & ~n1026;
  assign n1028 = ~x15 & n100;
  assign n1029 = ~x14 & n104;
  assign n1030 = ~n1028 & ~n1029;
  assign n1031 = n1027 & n1030;
  assign n1018 = x9 & n353;
  assign n1019 = x8 & n355;
  assign n1020 = ~n1018 & ~n1019;
  assign n1021 = ~x9 & n346;
  assign n1022 = ~x8 & n350;
  assign n1023 = ~n1021 & ~n1022;
  assign n1024 = n1020 & n1023;
  assign n1032 = n1031 ^ n1024;
  assign n1040 = n1039 ^ n1032;
  assign n1004 = x49 & n926;
  assign n1005 = ~x1 & n1004;
  assign n1006 = x49 ^ x48;
  assign n1007 = ~n926 & n1006;
  assign n1008 = x49 & n1007;
  assign n1009 = ~x0 & n1008;
  assign n1010 = ~n1005 & ~n1009;
  assign n1011 = ~x49 & n926;
  assign n1012 = x1 & n1011;
  assign n1013 = ~x49 & n1007;
  assign n1014 = x0 & n1013;
  assign n1015 = ~n1012 & ~n1014;
  assign n1016 = n1010 & n1015;
  assign n996 = ~x3 & n821;
  assign n997 = ~x2 & n823;
  assign n998 = ~n996 & ~n997;
  assign n999 = x3 & n814;
  assign n1000 = x2 & n818;
  assign n1001 = ~n999 & ~n1000;
  assign n1002 = n998 & n1001;
  assign n989 = ~x11 & n247;
  assign n990 = ~x10 & n251;
  assign n991 = ~n989 & ~n990;
  assign n992 = x11 & n254;
  assign n993 = x10 & n256;
  assign n994 = ~n992 & ~n993;
  assign n995 = n991 & n994;
  assign n1003 = n1002 ^ n995;
  assign n1017 = n1016 ^ n1003;
  assign n1041 = n1040 ^ n1017;
  assign n1069 = n1068 ^ n1041;
  assign n986 = n962 ^ n959;
  assign n987 = ~n973 & ~n986;
  assign n988 = n987 ^ n972;
  assign n1070 = n1069 ^ n988;
  assign n1090 = n1089 ^ n1070;
  assign n982 = n974 ^ n954;
  assign n983 = n974 ^ n889;
  assign n984 = n982 & ~n983;
  assign n985 = n984 ^ n954;
  assign n1091 = n1090 ^ n985;
  assign n1096 = n1095 ^ n1091;
  assign n1201 = n985 & ~n1090;
  assign n1202 = ~n985 & n1090;
  assign n1203 = ~n1095 & ~n1202;
  assign n1204 = ~n1201 & ~n1203;
  assign n1193 = x50 ^ x49;
  assign n1194 = x0 & n1193;
  assign n1187 = ~x17 & n66;
  assign n1188 = n69 ^ x18;
  assign n1189 = n1188 ^ n69;
  assign n1190 = n70 & n1189;
  assign n1191 = n1190 ^ n69;
  assign n1192 = ~n1187 & ~n1191;
  assign n1195 = n1194 ^ n1192;
  assign n1180 = ~x12 & n247;
  assign n1181 = ~x11 & n251;
  assign n1182 = ~n1180 & ~n1181;
  assign n1183 = x12 & n254;
  assign n1184 = x11 & n256;
  assign n1185 = ~n1183 & ~n1184;
  assign n1186 = n1182 & n1185;
  assign n1196 = n1195 ^ n1186;
  assign n1171 = ~x8 & n510;
  assign n1172 = ~x7 & n512;
  assign n1173 = ~n1171 & ~n1172;
  assign n1174 = x8 & n503;
  assign n1175 = x7 & n507;
  assign n1176 = ~n1174 & ~n1175;
  assign n1177 = n1173 & n1176;
  assign n1163 = ~x10 & n346;
  assign n1164 = ~x9 & n350;
  assign n1165 = ~n1163 & ~n1164;
  assign n1166 = x10 & n353;
  assign n1167 = x9 & n355;
  assign n1168 = ~n1166 & ~n1167;
  assign n1169 = n1165 & n1168;
  assign n1156 = ~x14 & n147;
  assign n1157 = ~x13 & n151;
  assign n1158 = ~n1156 & ~n1157;
  assign n1159 = x14 & n154;
  assign n1160 = x13 & n156;
  assign n1161 = ~n1159 & ~n1160;
  assign n1162 = n1158 & n1161;
  assign n1170 = n1169 ^ n1162;
  assign n1178 = n1177 ^ n1170;
  assign n1153 = n1039 ^ n1024;
  assign n1154 = n1032 & ~n1153;
  assign n1155 = n1154 ^ n1031;
  assign n1179 = n1178 ^ n1155;
  assign n1197 = n1196 ^ n1179;
  assign n1149 = n1068 ^ n1040;
  assign n1150 = ~n1041 & n1149;
  assign n1151 = n1150 ^ n1068;
  assign n1146 = n1082 ^ n1079;
  assign n1147 = ~n1086 & ~n1146;
  assign n1148 = n1147 ^ n1085;
  assign n1152 = n1151 ^ n1148;
  assign n1198 = n1197 ^ n1152;
  assign n1135 = x6 & n657;
  assign n1136 = x5 & n659;
  assign n1137 = ~n1135 & ~n1136;
  assign n1138 = ~x6 & n650;
  assign n1139 = ~x5 & n654;
  assign n1140 = ~n1138 & ~n1139;
  assign n1141 = n1137 & n1140;
  assign n1134 = ~n1062 & n1066;
  assign n1142 = n1141 ^ n1134;
  assign n1131 = n1016 ^ n1002;
  assign n1132 = ~n1003 & n1131;
  assign n1133 = n1132 ^ n1016;
  assign n1143 = n1142 ^ n1133;
  assign n1122 = ~x16 & n100;
  assign n1123 = ~x15 & n104;
  assign n1124 = ~n1122 & ~n1123;
  assign n1125 = x16 & n107;
  assign n1126 = x15 & n109;
  assign n1127 = ~n1125 & ~n1126;
  assign n1128 = n1124 & n1127;
  assign n1114 = x4 & n814;
  assign n1115 = x3 & n818;
  assign n1116 = ~n1114 & ~n1115;
  assign n1117 = ~x4 & n821;
  assign n1118 = ~x3 & n823;
  assign n1119 = ~n1117 & ~n1118;
  assign n1120 = n1116 & n1119;
  assign n1107 = x2 & n1011;
  assign n1108 = x1 & n1013;
  assign n1109 = ~n1107 & ~n1108;
  assign n1110 = ~x2 & n1004;
  assign n1111 = ~x1 & n1008;
  assign n1112 = ~n1110 & ~n1111;
  assign n1113 = n1109 & n1112;
  assign n1121 = n1120 ^ n1113;
  assign n1129 = n1128 ^ n1121;
  assign n1104 = n1067 ^ n1048;
  assign n1105 = n1056 & ~n1104;
  assign n1106 = n1105 ^ n1055;
  assign n1130 = n1129 ^ n1106;
  assign n1144 = n1143 ^ n1130;
  assign n1101 = n1087 ^ n1073;
  assign n1102 = ~n1088 & n1101;
  assign n1103 = n1102 ^ n1073;
  assign n1145 = n1144 ^ n1103;
  assign n1199 = n1198 ^ n1145;
  assign n1097 = n1089 ^ n1069;
  assign n1098 = n1089 ^ n988;
  assign n1099 = ~n1097 & ~n1098;
  assign n1100 = n1099 ^ n1069;
  assign n1200 = n1199 ^ n1100;
  assign n1205 = n1204 ^ n1200;
  assign n1328 = ~n1100 & ~n1199;
  assign n1329 = n1100 & n1199;
  assign n1330 = ~n1204 & ~n1329;
  assign n1331 = ~n1328 & ~n1330;
  assign n1315 = ~x3 & n1004;
  assign n1316 = ~x2 & n1008;
  assign n1317 = ~n1315 & ~n1316;
  assign n1318 = x3 & n1011;
  assign n1319 = x2 & n1013;
  assign n1320 = ~n1318 & ~n1319;
  assign n1321 = n1317 & n1320;
  assign n1307 = x13 & n254;
  assign n1308 = x12 & n256;
  assign n1309 = ~n1307 & ~n1308;
  assign n1310 = ~x13 & n247;
  assign n1311 = ~x12 & n251;
  assign n1312 = ~n1310 & ~n1311;
  assign n1313 = n1309 & n1312;
  assign n1300 = x5 & n814;
  assign n1301 = x4 & n818;
  assign n1302 = ~n1300 & ~n1301;
  assign n1303 = ~x5 & n821;
  assign n1304 = ~x4 & n823;
  assign n1305 = ~n1303 & ~n1304;
  assign n1306 = n1302 & n1305;
  assign n1314 = n1313 ^ n1306;
  assign n1322 = n1321 ^ n1314;
  assign n1291 = ~x7 & n650;
  assign n1292 = ~x6 & n654;
  assign n1293 = ~n1291 & ~n1292;
  assign n1294 = x7 & n657;
  assign n1295 = x6 & n659;
  assign n1296 = ~n1294 & ~n1295;
  assign n1297 = n1293 & n1296;
  assign n1283 = ~x15 & n147;
  assign n1284 = ~x14 & n151;
  assign n1285 = ~n1283 & ~n1284;
  assign n1286 = x15 & n154;
  assign n1287 = x14 & n156;
  assign n1288 = ~n1286 & ~n1287;
  assign n1289 = n1285 & n1288;
  assign n1276 = ~x9 & n510;
  assign n1277 = ~x8 & n512;
  assign n1278 = ~n1276 & ~n1277;
  assign n1279 = x9 & n503;
  assign n1280 = x8 & n507;
  assign n1281 = ~n1279 & ~n1280;
  assign n1282 = n1278 & n1281;
  assign n1290 = n1289 ^ n1282;
  assign n1298 = n1297 ^ n1290;
  assign n1273 = n1177 ^ n1169;
  assign n1274 = ~n1170 & n1273;
  assign n1275 = n1274 ^ n1177;
  assign n1299 = n1298 ^ n1275;
  assign n1323 = n1322 ^ n1299;
  assign n1270 = n1196 ^ n1178;
  assign n1271 = ~n1179 & ~n1270;
  assign n1272 = n1271 ^ n1196;
  assign n1324 = n1323 ^ n1272;
  assign n1267 = n1143 ^ n1106;
  assign n1268 = n1130 & n1267;
  assign n1269 = n1268 ^ n1129;
  assign n1325 = n1324 ^ n1269;
  assign n1258 = x49 ^ x0;
  assign n1259 = ~n1193 & n1258;
  assign n1260 = n1259 ^ x0;
  assign n1261 = x51 & ~n1260;
  assign n1252 = ~x18 & n66;
  assign n1253 = n69 ^ x19;
  assign n1254 = n1253 ^ n69;
  assign n1255 = n70 & n1254;
  assign n1256 = n1255 ^ n69;
  assign n1257 = ~n1252 & ~n1256;
  assign n1262 = n1261 ^ n1257;
  assign n1249 = n1192 ^ n1186;
  assign n1250 = ~n1195 & ~n1249;
  assign n1251 = n1250 ^ n1194;
  assign n1263 = n1262 ^ n1251;
  assign n1246 = n1128 ^ n1120;
  assign n1247 = ~n1121 & n1246;
  assign n1248 = n1247 ^ n1128;
  assign n1264 = n1263 ^ n1248;
  assign n1237 = x11 & n353;
  assign n1238 = x10 & n355;
  assign n1239 = ~n1237 & ~n1238;
  assign n1240 = ~x11 & n346;
  assign n1241 = ~x10 & n350;
  assign n1242 = ~n1240 & ~n1241;
  assign n1243 = n1239 & n1242;
  assign n1223 = ~x51 & n1193;
  assign n1224 = x1 & n1223;
  assign n1225 = x51 ^ x50;
  assign n1226 = ~n1193 & n1225;
  assign n1227 = ~x51 & n1226;
  assign n1228 = x0 & n1227;
  assign n1229 = ~n1224 & ~n1228;
  assign n1230 = x51 & n1193;
  assign n1231 = ~x1 & n1230;
  assign n1232 = x51 & n1226;
  assign n1233 = ~x0 & n1232;
  assign n1234 = ~n1231 & ~n1233;
  assign n1235 = n1229 & n1234;
  assign n1216 = x17 & n107;
  assign n1217 = x16 & n109;
  assign n1218 = ~n1216 & ~n1217;
  assign n1219 = ~x17 & n100;
  assign n1220 = ~x16 & n104;
  assign n1221 = ~n1219 & ~n1220;
  assign n1222 = n1218 & n1221;
  assign n1236 = n1235 ^ n1222;
  assign n1244 = n1243 ^ n1236;
  assign n1213 = n1134 ^ n1133;
  assign n1214 = ~n1142 & n1213;
  assign n1215 = n1214 ^ n1141;
  assign n1245 = n1244 ^ n1215;
  assign n1265 = n1264 ^ n1245;
  assign n1210 = n1197 ^ n1151;
  assign n1211 = n1152 & ~n1210;
  assign n1212 = n1211 ^ n1197;
  assign n1266 = n1265 ^ n1212;
  assign n1326 = n1325 ^ n1266;
  assign n1206 = n1198 ^ n1144;
  assign n1207 = n1198 ^ n1103;
  assign n1208 = ~n1206 & n1207;
  assign n1209 = n1208 ^ n1144;
  assign n1327 = n1326 ^ n1209;
  assign n1332 = n1331 ^ n1327;
  assign n1452 = n1209 & n1326;
  assign n1453 = ~n1209 & ~n1326;
  assign n1454 = ~n1331 & ~n1453;
  assign n1455 = ~n1452 & ~n1454;
  assign n1439 = x16 & n154;
  assign n1440 = x15 & n156;
  assign n1441 = ~n1439 & ~n1440;
  assign n1442 = ~x16 & n147;
  assign n1443 = ~x15 & n151;
  assign n1444 = ~n1442 & ~n1443;
  assign n1445 = n1441 & n1444;
  assign n1431 = ~x2 & n1230;
  assign n1432 = ~x1 & n1232;
  assign n1433 = ~n1431 & ~n1432;
  assign n1434 = x2 & n1223;
  assign n1435 = x1 & n1227;
  assign n1436 = ~n1434 & ~n1435;
  assign n1437 = n1433 & n1436;
  assign n1424 = ~x12 & n346;
  assign n1425 = ~x11 & n350;
  assign n1426 = ~n1424 & ~n1425;
  assign n1427 = x12 & n353;
  assign n1428 = x11 & n355;
  assign n1429 = ~n1427 & ~n1428;
  assign n1430 = n1426 & n1429;
  assign n1438 = n1437 ^ n1430;
  assign n1446 = n1445 ^ n1438;
  assign n1419 = x52 ^ x51;
  assign n1420 = x0 & n1419;
  assign n1413 = ~x19 & n66;
  assign n1414 = n69 ^ x20;
  assign n1415 = n1414 ^ n69;
  assign n1416 = n70 & n1415;
  assign n1417 = n1416 ^ n69;
  assign n1418 = ~n1413 & ~n1417;
  assign n1421 = n1420 ^ n1418;
  assign n1406 = ~x14 & n247;
  assign n1407 = ~x13 & n251;
  assign n1408 = ~n1406 & ~n1407;
  assign n1409 = x14 & n254;
  assign n1410 = x13 & n256;
  assign n1411 = ~n1409 & ~n1410;
  assign n1412 = n1408 & n1411;
  assign n1422 = n1421 ^ n1412;
  assign n1398 = ~x18 & n100;
  assign n1399 = ~x17 & n104;
  assign n1400 = ~n1398 & ~n1399;
  assign n1401 = x18 & n107;
  assign n1402 = x17 & n109;
  assign n1403 = ~n1401 & ~n1402;
  assign n1404 = n1400 & n1403;
  assign n1390 = ~x4 & n1004;
  assign n1391 = ~x3 & n1008;
  assign n1392 = ~n1390 & ~n1391;
  assign n1393 = x4 & n1011;
  assign n1394 = x3 & n1013;
  assign n1395 = ~n1393 & ~n1394;
  assign n1396 = n1392 & n1395;
  assign n1383 = ~x6 & n821;
  assign n1384 = ~x5 & n823;
  assign n1385 = ~n1383 & ~n1384;
  assign n1386 = x6 & n814;
  assign n1387 = x5 & n818;
  assign n1388 = ~n1386 & ~n1387;
  assign n1389 = n1385 & n1388;
  assign n1397 = n1396 ^ n1389;
  assign n1405 = n1404 ^ n1397;
  assign n1423 = n1422 ^ n1405;
  assign n1447 = n1446 ^ n1423;
  assign n1378 = n1297 ^ n1282;
  assign n1379 = n1290 & ~n1378;
  assign n1380 = n1379 ^ n1289;
  assign n1375 = n1321 ^ n1306;
  assign n1376 = n1314 & ~n1375;
  assign n1377 = n1376 ^ n1313;
  assign n1381 = n1380 ^ n1377;
  assign n1372 = n1243 ^ n1235;
  assign n1373 = ~n1236 & n1372;
  assign n1374 = n1373 ^ n1243;
  assign n1382 = n1381 ^ n1374;
  assign n1448 = n1447 ^ n1382;
  assign n1368 = ~n1257 & n1261;
  assign n1360 = ~x10 & n510;
  assign n1361 = ~x9 & n512;
  assign n1362 = ~n1360 & ~n1361;
  assign n1363 = x10 & n503;
  assign n1364 = x9 & n507;
  assign n1365 = ~n1363 & ~n1364;
  assign n1366 = n1362 & n1365;
  assign n1353 = ~x8 & n650;
  assign n1354 = ~x7 & n654;
  assign n1355 = ~n1353 & ~n1354;
  assign n1356 = x8 & n657;
  assign n1357 = x7 & n659;
  assign n1358 = ~n1356 & ~n1357;
  assign n1359 = n1355 & n1358;
  assign n1367 = n1366 ^ n1359;
  assign n1369 = n1368 ^ n1367;
  assign n1350 = n1251 ^ n1248;
  assign n1351 = ~n1263 & n1350;
  assign n1352 = n1351 ^ n1262;
  assign n1370 = n1369 ^ n1352;
  assign n1346 = n1322 ^ n1298;
  assign n1347 = n1322 ^ n1275;
  assign n1348 = n1346 & ~n1347;
  assign n1349 = n1348 ^ n1298;
  assign n1371 = n1370 ^ n1349;
  assign n1449 = n1448 ^ n1371;
  assign n1341 = n1264 ^ n1244;
  assign n1342 = n1264 ^ n1215;
  assign n1343 = ~n1341 & n1342;
  assign n1344 = n1343 ^ n1244;
  assign n1337 = n1323 ^ n1269;
  assign n1338 = n1272 ^ n1269;
  assign n1339 = n1337 & n1338;
  assign n1340 = n1339 ^ n1323;
  assign n1345 = n1344 ^ n1340;
  assign n1450 = n1449 ^ n1345;
  assign n1333 = n1325 ^ n1265;
  assign n1334 = n1325 ^ n1212;
  assign n1335 = n1333 & ~n1334;
  assign n1336 = n1335 ^ n1265;
  assign n1451 = n1450 ^ n1336;
  assign n1456 = n1455 ^ n1451;
  assign n1592 = n1336 & ~n1450;
  assign n1593 = ~n1336 & n1450;
  assign n1594 = ~n1455 & ~n1593;
  assign n1595 = ~n1592 & ~n1594;
  assign n1571 = x53 & n1419;
  assign n1572 = ~x1 & n1571;
  assign n1573 = x53 ^ x52;
  assign n1574 = ~n1419 & n1573;
  assign n1575 = x53 & n1574;
  assign n1576 = ~x0 & n1575;
  assign n1577 = ~n1572 & ~n1576;
  assign n1578 = ~x53 & n1419;
  assign n1579 = x1 & n1578;
  assign n1580 = ~x53 & n1574;
  assign n1581 = x0 & n1580;
  assign n1582 = ~n1579 & ~n1581;
  assign n1583 = n1577 & n1582;
  assign n1563 = ~x13 & n346;
  assign n1564 = ~x12 & n350;
  assign n1565 = ~n1563 & ~n1564;
  assign n1566 = x13 & n353;
  assign n1567 = x12 & n355;
  assign n1568 = ~n1566 & ~n1567;
  assign n1569 = n1565 & n1568;
  assign n1556 = x3 & n1223;
  assign n1557 = x2 & n1227;
  assign n1558 = ~n1556 & ~n1557;
  assign n1559 = ~x3 & n1230;
  assign n1560 = ~x2 & n1232;
  assign n1561 = ~n1559 & ~n1560;
  assign n1562 = n1558 & n1561;
  assign n1570 = n1569 ^ n1562;
  assign n1584 = n1583 ^ n1570;
  assign n1548 = ~x5 & n1004;
  assign n1549 = ~x4 & n1008;
  assign n1550 = ~n1548 & ~n1549;
  assign n1551 = x5 & n1011;
  assign n1552 = x4 & n1013;
  assign n1553 = ~n1551 & ~n1552;
  assign n1554 = n1550 & n1553;
  assign n1540 = x7 & n814;
  assign n1541 = x6 & n818;
  assign n1542 = ~n1540 & ~n1541;
  assign n1543 = ~x7 & n821;
  assign n1544 = ~x6 & n823;
  assign n1545 = ~n1543 & ~n1544;
  assign n1546 = n1542 & n1545;
  assign n1533 = ~x15 & n247;
  assign n1534 = ~x14 & n251;
  assign n1535 = ~n1533 & ~n1534;
  assign n1536 = x15 & n254;
  assign n1537 = x14 & n256;
  assign n1538 = ~n1536 & ~n1537;
  assign n1539 = n1535 & n1538;
  assign n1547 = n1546 ^ n1539;
  assign n1555 = n1554 ^ n1547;
  assign n1585 = n1584 ^ n1555;
  assign n1530 = n1368 ^ n1359;
  assign n1531 = n1367 & n1530;
  assign n1532 = n1531 ^ n1366;
  assign n1586 = n1585 ^ n1532;
  assign n1527 = n1446 ^ n1405;
  assign n1528 = ~n1423 & ~n1527;
  assign n1529 = n1528 ^ n1422;
  assign n1587 = n1586 ^ n1529;
  assign n1517 = ~x11 & n510;
  assign n1518 = ~x10 & n512;
  assign n1519 = ~n1517 & ~n1518;
  assign n1520 = x11 & n503;
  assign n1521 = x10 & n507;
  assign n1522 = ~n1520 & ~n1521;
  assign n1523 = n1519 & n1522;
  assign n1509 = ~x17 & n147;
  assign n1510 = ~x16 & n151;
  assign n1511 = ~n1509 & ~n1510;
  assign n1512 = x17 & n154;
  assign n1513 = x16 & n156;
  assign n1514 = ~n1512 & ~n1513;
  assign n1515 = n1511 & n1514;
  assign n1503 = ~x20 & n66;
  assign n1504 = n69 ^ x21;
  assign n1505 = n1504 ^ n69;
  assign n1506 = n70 & n1505;
  assign n1507 = n1506 ^ n69;
  assign n1508 = ~n1503 & ~n1507;
  assign n1516 = n1515 ^ n1508;
  assign n1524 = n1523 ^ n1516;
  assign n1499 = n1418 ^ n1412;
  assign n1500 = ~n1421 & ~n1499;
  assign n1501 = n1500 ^ n1420;
  assign n1496 = n1445 ^ n1430;
  assign n1497 = n1438 & ~n1496;
  assign n1498 = n1497 ^ n1437;
  assign n1502 = n1501 ^ n1498;
  assign n1525 = n1524 ^ n1502;
  assign n1486 = x9 & n657;
  assign n1487 = x8 & n659;
  assign n1488 = ~n1486 & ~n1487;
  assign n1489 = ~x9 & n650;
  assign n1490 = ~x8 & n654;
  assign n1491 = ~n1489 & ~n1490;
  assign n1492 = n1488 & n1491;
  assign n1481 = x51 ^ x0;
  assign n1482 = ~n1419 & n1481;
  assign n1483 = n1482 ^ x0;
  assign n1484 = x53 & ~n1483;
  assign n1474 = x19 & n107;
  assign n1475 = x18 & n109;
  assign n1476 = ~n1474 & ~n1475;
  assign n1477 = ~x19 & n100;
  assign n1478 = ~x18 & n104;
  assign n1479 = ~n1477 & ~n1478;
  assign n1480 = n1476 & n1479;
  assign n1485 = n1484 ^ n1480;
  assign n1493 = n1492 ^ n1485;
  assign n1470 = n1404 ^ n1396;
  assign n1471 = n1404 ^ n1389;
  assign n1472 = n1470 & ~n1471;
  assign n1473 = n1472 ^ n1396;
  assign n1494 = n1493 ^ n1473;
  assign n1467 = n1377 ^ n1374;
  assign n1468 = n1381 & ~n1467;
  assign n1469 = n1468 ^ n1380;
  assign n1495 = n1494 ^ n1469;
  assign n1526 = n1525 ^ n1495;
  assign n1588 = n1587 ^ n1526;
  assign n1463 = n1369 ^ n1349;
  assign n1464 = n1352 ^ n1349;
  assign n1465 = ~n1463 & ~n1464;
  assign n1466 = n1465 ^ n1369;
  assign n1589 = n1588 ^ n1466;
  assign n1460 = n1382 ^ n1371;
  assign n1461 = ~n1448 & n1460;
  assign n1462 = n1461 ^ n1447;
  assign n1590 = n1589 ^ n1462;
  assign n1457 = n1449 ^ n1344;
  assign n1458 = ~n1345 & n1457;
  assign n1459 = n1458 ^ n1449;
  assign n1591 = n1590 ^ n1459;
  assign n1596 = n1595 ^ n1591;
  assign n1726 = ~n1459 & ~n1590;
  assign n1727 = n1459 & n1590;
  assign n1728 = ~n1595 & ~n1727;
  assign n1729 = ~n1726 & ~n1728;
  assign n1718 = ~n1480 & n1484;
  assign n1715 = n1523 ^ n1515;
  assign n1716 = n1516 & ~n1715;
  assign n1717 = n1716 ^ n1508;
  assign n1719 = n1718 ^ n1717;
  assign n1712 = n1583 ^ n1569;
  assign n1713 = ~n1570 & n1712;
  assign n1714 = n1713 ^ n1583;
  assign n1720 = n1719 ^ n1714;
  assign n1709 = n1524 ^ n1501;
  assign n1710 = n1502 & ~n1709;
  assign n1711 = n1710 ^ n1524;
  assign n1721 = n1720 ^ n1711;
  assign n1706 = n1555 ^ n1532;
  assign n1707 = n1585 & ~n1706;
  assign n1708 = n1707 ^ n1584;
  assign n1722 = n1721 ^ n1708;
  assign n1695 = x14 & n353;
  assign n1696 = x13 & n355;
  assign n1697 = ~n1695 & ~n1696;
  assign n1698 = ~x14 & n346;
  assign n1699 = ~x13 & n350;
  assign n1700 = ~n1698 & ~n1699;
  assign n1701 = n1697 & n1700;
  assign n1687 = x8 & n814;
  assign n1688 = x7 & n818;
  assign n1689 = ~n1687 & ~n1688;
  assign n1690 = ~x8 & n821;
  assign n1691 = ~x7 & n823;
  assign n1692 = ~n1690 & ~n1691;
  assign n1693 = n1689 & n1692;
  assign n1680 = ~x6 & n1004;
  assign n1681 = ~x5 & n1008;
  assign n1682 = ~n1680 & ~n1681;
  assign n1683 = x6 & n1011;
  assign n1684 = x5 & n1013;
  assign n1685 = ~n1683 & ~n1684;
  assign n1686 = n1682 & n1685;
  assign n1694 = n1693 ^ n1686;
  assign n1702 = n1701 ^ n1694;
  assign n1671 = ~x10 & n650;
  assign n1672 = ~x9 & n654;
  assign n1673 = ~n1671 & ~n1672;
  assign n1674 = x10 & n657;
  assign n1675 = x9 & n659;
  assign n1676 = ~n1674 & ~n1675;
  assign n1677 = n1673 & n1676;
  assign n1663 = ~x18 & n147;
  assign n1664 = ~x17 & n151;
  assign n1665 = ~n1663 & ~n1664;
  assign n1666 = x18 & n154;
  assign n1667 = x17 & n156;
  assign n1668 = ~n1666 & ~n1667;
  assign n1669 = n1665 & n1668;
  assign n1656 = ~x12 & n510;
  assign n1657 = ~x11 & n512;
  assign n1658 = ~n1656 & ~n1657;
  assign n1659 = x12 & n503;
  assign n1660 = x11 & n507;
  assign n1661 = ~n1659 & ~n1660;
  assign n1662 = n1658 & n1661;
  assign n1670 = n1669 ^ n1662;
  assign n1678 = n1677 ^ n1670;
  assign n1653 = n1554 ^ n1539;
  assign n1654 = n1547 & ~n1653;
  assign n1655 = n1654 ^ n1546;
  assign n1679 = n1678 ^ n1655;
  assign n1703 = n1702 ^ n1679;
  assign n1643 = ~x16 & n247;
  assign n1644 = ~x15 & n251;
  assign n1645 = ~n1643 & ~n1644;
  assign n1646 = x16 & n254;
  assign n1647 = x15 & n256;
  assign n1648 = ~n1646 & ~n1647;
  assign n1649 = n1645 & n1648;
  assign n1640 = x54 ^ x53;
  assign n1641 = x0 & n1640;
  assign n1633 = x20 & n107;
  assign n1634 = x19 & n109;
  assign n1635 = ~n1633 & ~n1634;
  assign n1636 = ~x20 & n100;
  assign n1637 = ~x19 & n104;
  assign n1638 = ~n1636 & ~n1637;
  assign n1639 = n1635 & n1638;
  assign n1642 = n1641 ^ n1639;
  assign n1650 = n1649 ^ n1642;
  assign n1624 = x4 & n1223;
  assign n1625 = x3 & n1227;
  assign n1626 = ~n1624 & ~n1625;
  assign n1627 = ~x4 & n1230;
  assign n1628 = ~x3 & n1232;
  assign n1629 = ~n1627 & ~n1628;
  assign n1630 = n1626 & n1629;
  assign n1617 = x2 & n1578;
  assign n1618 = x1 & n1580;
  assign n1619 = ~n1617 & ~n1618;
  assign n1620 = ~x2 & n1571;
  assign n1621 = ~x1 & n1575;
  assign n1622 = ~n1620 & ~n1621;
  assign n1623 = n1619 & n1622;
  assign n1631 = n1630 ^ n1623;
  assign n1611 = ~x21 & n66;
  assign n1612 = n69 ^ x22;
  assign n1613 = n1612 ^ n69;
  assign n1614 = n70 & n1613;
  assign n1615 = n1614 ^ n69;
  assign n1616 = ~n1611 & ~n1615;
  assign n1632 = n1631 ^ n1616;
  assign n1651 = n1650 ^ n1632;
  assign n1608 = n1485 ^ n1473;
  assign n1609 = n1493 & ~n1608;
  assign n1610 = n1609 ^ n1492;
  assign n1652 = n1651 ^ n1610;
  assign n1704 = n1703 ^ n1652;
  assign n1604 = n1525 ^ n1494;
  assign n1605 = n1525 ^ n1469;
  assign n1606 = ~n1604 & n1605;
  assign n1607 = n1606 ^ n1494;
  assign n1705 = n1704 ^ n1607;
  assign n1723 = n1722 ^ n1705;
  assign n1601 = n1586 ^ n1526;
  assign n1602 = ~n1587 & n1601;
  assign n1603 = n1602 ^ n1529;
  assign n1724 = n1723 ^ n1603;
  assign n1597 = n1588 ^ n1462;
  assign n1598 = n1466 ^ n1462;
  assign n1599 = ~n1597 & ~n1598;
  assign n1600 = n1599 ^ n1588;
  assign n1725 = n1724 ^ n1600;
  assign n1730 = n1729 ^ n1725;
  assign n1878 = ~n1600 & n1724;
  assign n1879 = n1600 & ~n1724;
  assign n1880 = ~n1729 & ~n1879;
  assign n1881 = ~n1878 & ~n1880;
  assign n1865 = ~x3 & n1571;
  assign n1866 = ~x2 & n1575;
  assign n1867 = ~n1865 & ~n1866;
  assign n1868 = x3 & n1578;
  assign n1869 = x2 & n1580;
  assign n1870 = ~n1868 & ~n1869;
  assign n1871 = n1867 & n1870;
  assign n1857 = x15 & n353;
  assign n1858 = x14 & n355;
  assign n1859 = ~n1857 & ~n1858;
  assign n1860 = ~x15 & n346;
  assign n1861 = ~x14 & n350;
  assign n1862 = ~n1860 & ~n1861;
  assign n1863 = n1859 & n1862;
  assign n1850 = x5 & n1223;
  assign n1851 = x4 & n1227;
  assign n1852 = ~n1850 & ~n1851;
  assign n1853 = ~x5 & n1230;
  assign n1854 = ~x4 & n1232;
  assign n1855 = ~n1853 & ~n1854;
  assign n1856 = n1852 & n1855;
  assign n1864 = n1863 ^ n1856;
  assign n1872 = n1871 ^ n1864;
  assign n1835 = x55 & n1640;
  assign n1836 = ~x1 & n1835;
  assign n1837 = x55 ^ x54;
  assign n1838 = ~n1640 & n1837;
  assign n1839 = x55 & n1838;
  assign n1840 = ~x0 & n1839;
  assign n1841 = ~n1836 & ~n1840;
  assign n1842 = ~x55 & n1640;
  assign n1843 = x1 & n1842;
  assign n1844 = ~x55 & n1838;
  assign n1845 = x0 & n1844;
  assign n1846 = ~n1843 & ~n1845;
  assign n1847 = n1841 & n1846;
  assign n1827 = x19 & n154;
  assign n1828 = x18 & n156;
  assign n1829 = ~n1827 & ~n1828;
  assign n1830 = ~x19 & n147;
  assign n1831 = ~x18 & n151;
  assign n1832 = ~n1830 & ~n1831;
  assign n1833 = n1829 & n1832;
  assign n1821 = ~x22 & n66;
  assign n1822 = n69 ^ x23;
  assign n1823 = n1822 ^ n69;
  assign n1824 = n70 & n1823;
  assign n1825 = n1824 ^ n69;
  assign n1826 = ~n1821 & ~n1825;
  assign n1834 = n1833 ^ n1826;
  assign n1848 = n1847 ^ n1834;
  assign n1818 = n1701 ^ n1693;
  assign n1819 = ~n1694 & n1818;
  assign n1820 = n1819 ^ n1701;
  assign n1849 = n1848 ^ n1820;
  assign n1873 = n1872 ^ n1849;
  assign n1812 = n1677 ^ n1662;
  assign n1813 = n1670 & ~n1812;
  assign n1814 = n1813 ^ n1669;
  assign n1809 = n1630 ^ n1616;
  assign n1810 = ~n1631 & n1809;
  assign n1811 = n1810 ^ n1616;
  assign n1815 = n1814 ^ n1811;
  assign n1805 = n1649 ^ n1641;
  assign n1806 = n1649 ^ n1639;
  assign n1807 = ~n1805 & ~n1806;
  assign n1808 = n1807 ^ n1641;
  assign n1816 = n1815 ^ n1808;
  assign n1801 = n1702 ^ n1678;
  assign n1802 = n1702 ^ n1655;
  assign n1803 = n1801 & ~n1802;
  assign n1804 = n1803 ^ n1678;
  assign n1817 = n1816 ^ n1804;
  assign n1874 = n1873 ^ n1817;
  assign n1789 = ~x13 & n510;
  assign n1790 = ~x12 & n512;
  assign n1791 = ~n1789 & ~n1790;
  assign n1792 = x13 & n503;
  assign n1793 = x12 & n507;
  assign n1794 = ~n1792 & ~n1793;
  assign n1795 = n1791 & n1794;
  assign n1782 = ~x11 & n650;
  assign n1783 = ~x10 & n654;
  assign n1784 = ~n1782 & ~n1783;
  assign n1785 = x11 & n657;
  assign n1786 = x10 & n659;
  assign n1787 = ~n1785 & ~n1786;
  assign n1788 = n1784 & n1787;
  assign n1796 = n1795 ^ n1788;
  assign n1777 = x53 ^ x0;
  assign n1778 = ~n1640 & n1777;
  assign n1779 = n1778 ^ x0;
  assign n1780 = x55 & ~n1779;
  assign n1770 = ~x21 & n100;
  assign n1771 = ~x20 & n104;
  assign n1772 = ~n1770 & ~n1771;
  assign n1773 = x21 & n107;
  assign n1774 = x20 & n109;
  assign n1775 = ~n1773 & ~n1774;
  assign n1776 = n1772 & n1775;
  assign n1781 = n1780 ^ n1776;
  assign n1797 = n1796 ^ n1781;
  assign n1762 = ~x7 & n1004;
  assign n1763 = ~x6 & n1008;
  assign n1764 = ~n1762 & ~n1763;
  assign n1765 = x7 & n1011;
  assign n1766 = x6 & n1013;
  assign n1767 = ~n1765 & ~n1766;
  assign n1768 = n1764 & n1767;
  assign n1754 = ~x17 & n247;
  assign n1755 = ~x16 & n251;
  assign n1756 = ~n1754 & ~n1755;
  assign n1757 = x17 & n254;
  assign n1758 = x16 & n256;
  assign n1759 = ~n1757 & ~n1758;
  assign n1760 = n1756 & n1759;
  assign n1747 = x9 & n814;
  assign n1748 = x8 & n818;
  assign n1749 = ~n1747 & ~n1748;
  assign n1750 = ~x9 & n821;
  assign n1751 = ~x8 & n823;
  assign n1752 = ~n1750 & ~n1751;
  assign n1753 = n1749 & n1752;
  assign n1761 = n1760 ^ n1753;
  assign n1769 = n1768 ^ n1761;
  assign n1798 = n1797 ^ n1769;
  assign n1744 = n1717 ^ n1714;
  assign n1745 = ~n1719 & ~n1744;
  assign n1746 = n1745 ^ n1718;
  assign n1799 = n1798 ^ n1746;
  assign n1741 = n1632 ^ n1610;
  assign n1742 = ~n1651 & ~n1741;
  assign n1743 = n1742 ^ n1650;
  assign n1800 = n1799 ^ n1743;
  assign n1875 = n1874 ^ n1800;
  assign n1737 = n1711 ^ n1708;
  assign n1738 = ~n1721 & ~n1737;
  assign n1739 = n1738 ^ n1720;
  assign n1734 = n1652 ^ n1607;
  assign n1735 = ~n1704 & n1734;
  assign n1736 = n1735 ^ n1703;
  assign n1740 = n1739 ^ n1736;
  assign n1876 = n1875 ^ n1740;
  assign n1731 = n1705 ^ n1603;
  assign n1732 = n1723 & ~n1731;
  assign n1733 = n1732 ^ n1722;
  assign n1877 = n1876 ^ n1733;
  assign n1882 = n1881 ^ n1877;
  assign n2023 = n1733 & ~n1876;
  assign n2024 = ~n1733 & n1876;
  assign n2025 = ~n1881 & ~n2024;
  assign n2026 = ~n2023 & ~n2025;
  assign n2010 = ~x16 & n346;
  assign n2011 = ~x15 & n350;
  assign n2012 = ~n2010 & ~n2011;
  assign n2013 = x16 & n353;
  assign n2014 = x15 & n355;
  assign n2015 = ~n2013 & ~n2014;
  assign n2016 = n2012 & n2015;
  assign n2002 = x8 & n1011;
  assign n2003 = x7 & n1013;
  assign n2004 = ~n2002 & ~n2003;
  assign n2005 = ~x8 & n1004;
  assign n2006 = ~x7 & n1008;
  assign n2007 = ~n2005 & ~n2006;
  assign n2008 = n2004 & n2007;
  assign n1995 = x10 & n814;
  assign n1996 = x9 & n818;
  assign n1997 = ~n1995 & ~n1996;
  assign n1998 = ~x10 & n821;
  assign n1999 = ~x9 & n823;
  assign n2000 = ~n1998 & ~n1999;
  assign n2001 = n1997 & n2000;
  assign n2009 = n2008 ^ n2001;
  assign n2017 = n2016 ^ n2009;
  assign n1986 = ~x18 & n247;
  assign n1987 = ~x17 & n251;
  assign n1988 = ~n1986 & ~n1987;
  assign n1989 = x18 & n254;
  assign n1990 = x17 & n256;
  assign n1991 = ~n1989 & ~n1990;
  assign n1992 = n1988 & n1991;
  assign n1983 = x56 ^ x55;
  assign n1984 = x0 & n1983;
  assign n1976 = ~x22 & n100;
  assign n1977 = ~x21 & n104;
  assign n1978 = ~n1976 & ~n1977;
  assign n1979 = x22 & n107;
  assign n1980 = x21 & n109;
  assign n1981 = ~n1979 & ~n1980;
  assign n1982 = n1978 & n1981;
  assign n1985 = n1984 ^ n1982;
  assign n1993 = n1992 ^ n1985;
  assign n1967 = ~x6 & n1230;
  assign n1968 = ~x5 & n1232;
  assign n1969 = ~n1967 & ~n1968;
  assign n1970 = x6 & n1223;
  assign n1971 = x5 & n1227;
  assign n1972 = ~n1970 & ~n1971;
  assign n1973 = n1969 & n1972;
  assign n1960 = ~x4 & n1571;
  assign n1961 = ~x3 & n1575;
  assign n1962 = ~n1960 & ~n1961;
  assign n1963 = x4 & n1578;
  assign n1964 = x3 & n1580;
  assign n1965 = ~n1963 & ~n1964;
  assign n1966 = n1962 & n1965;
  assign n1974 = n1973 ^ n1966;
  assign n1954 = ~x23 & n66;
  assign n1955 = n69 ^ x24;
  assign n1956 = n1955 ^ n69;
  assign n1957 = n70 & n1956;
  assign n1958 = n1957 ^ n69;
  assign n1959 = ~n1954 & ~n1958;
  assign n1975 = n1974 ^ n1959;
  assign n1994 = n1993 ^ n1975;
  assign n2018 = n2017 ^ n1994;
  assign n1944 = ~x14 & n510;
  assign n1945 = ~x13 & n512;
  assign n1946 = ~n1944 & ~n1945;
  assign n1947 = x14 & n503;
  assign n1948 = x13 & n507;
  assign n1949 = ~n1947 & ~n1948;
  assign n1950 = n1946 & n1949;
  assign n1936 = ~x2 & n1835;
  assign n1937 = ~x1 & n1839;
  assign n1938 = ~n1936 & ~n1937;
  assign n1939 = x2 & n1842;
  assign n1940 = x1 & n1844;
  assign n1941 = ~n1939 & ~n1940;
  assign n1942 = n1938 & n1941;
  assign n1929 = ~x20 & n147;
  assign n1930 = ~x19 & n151;
  assign n1931 = ~n1929 & ~n1930;
  assign n1932 = x20 & n154;
  assign n1933 = x19 & n156;
  assign n1934 = ~n1932 & ~n1933;
  assign n1935 = n1931 & n1934;
  assign n1943 = n1942 ^ n1935;
  assign n1951 = n1950 ^ n1943;
  assign n1925 = n1847 ^ n1833;
  assign n1926 = n1834 & ~n1925;
  assign n1927 = n1926 ^ n1826;
  assign n1922 = n1768 ^ n1760;
  assign n1923 = ~n1761 & n1922;
  assign n1924 = n1923 ^ n1768;
  assign n1928 = n1927 ^ n1924;
  assign n1952 = n1951 ^ n1928;
  assign n1919 = n1872 ^ n1848;
  assign n1920 = ~n1849 & n1919;
  assign n1921 = n1920 ^ n1872;
  assign n1953 = n1952 ^ n1921;
  assign n2019 = n2018 ^ n1953;
  assign n1907 = ~x12 & n650;
  assign n1908 = ~x11 & n654;
  assign n1909 = ~n1907 & ~n1908;
  assign n1910 = x12 & n657;
  assign n1911 = x11 & n659;
  assign n1912 = ~n1910 & ~n1911;
  assign n1913 = n1909 & n1912;
  assign n1906 = ~n1776 & n1780;
  assign n1914 = n1913 ^ n1906;
  assign n1903 = n1871 ^ n1863;
  assign n1904 = ~n1864 & n1903;
  assign n1905 = n1904 ^ n1871;
  assign n1915 = n1914 ^ n1905;
  assign n1899 = n1788 ^ n1781;
  assign n1900 = n1796 & ~n1899;
  assign n1901 = n1900 ^ n1795;
  assign n1896 = n1814 ^ n1808;
  assign n1897 = ~n1815 & ~n1896;
  assign n1898 = n1897 ^ n1808;
  assign n1902 = n1901 ^ n1898;
  assign n1916 = n1915 ^ n1902;
  assign n1893 = n1769 ^ n1746;
  assign n1894 = n1798 & n1893;
  assign n1895 = n1894 ^ n1797;
  assign n1917 = n1916 ^ n1895;
  assign n1890 = n1873 ^ n1816;
  assign n1891 = n1817 & ~n1890;
  assign n1892 = n1891 ^ n1873;
  assign n1918 = n1917 ^ n1892;
  assign n2020 = n2019 ^ n1918;
  assign n1886 = n1874 ^ n1799;
  assign n1887 = n1874 ^ n1743;
  assign n1888 = n1886 & ~n1887;
  assign n1889 = n1888 ^ n1799;
  assign n2021 = n2020 ^ n1889;
  assign n1883 = n1875 ^ n1739;
  assign n1884 = n1740 & n1883;
  assign n1885 = n1884 ^ n1875;
  assign n2022 = n2021 ^ n1885;
  assign n2027 = n2026 ^ n2022;
  assign n2189 = n1885 & ~n2021;
  assign n2190 = ~n1885 & n2021;
  assign n2191 = ~n2026 & ~n2190;
  assign n2192 = ~n2189 & ~n2191;
  assign n2175 = ~x13 & n650;
  assign n2176 = ~x12 & n654;
  assign n2177 = ~n2175 & ~n2176;
  assign n2178 = x13 & n657;
  assign n2179 = x12 & n659;
  assign n2180 = ~n2178 & ~n2179;
  assign n2181 = n2177 & n2180;
  assign n2161 = x57 & n1983;
  assign n2162 = ~x1 & n2161;
  assign n2163 = x57 ^ x56;
  assign n2164 = ~n1983 & n2163;
  assign n2165 = x57 & n2164;
  assign n2166 = ~x0 & n2165;
  assign n2167 = ~n2162 & ~n2166;
  assign n2168 = ~x57 & n1983;
  assign n2169 = x1 & n2168;
  assign n2170 = ~x57 & n2164;
  assign n2171 = x0 & n2170;
  assign n2172 = ~n2169 & ~n2171;
  assign n2173 = n2167 & n2172;
  assign n2154 = ~x21 & n147;
  assign n2155 = ~x20 & n151;
  assign n2156 = ~n2154 & ~n2155;
  assign n2157 = x21 & n154;
  assign n2158 = x20 & n156;
  assign n2159 = ~n2157 & ~n2158;
  assign n2160 = n2156 & n2159;
  assign n2174 = n2173 ^ n2160;
  assign n2182 = n2181 ^ n2174;
  assign n2150 = n1992 ^ n1982;
  assign n2151 = ~n1985 & ~n2150;
  assign n2152 = n2151 ^ n1984;
  assign n2146 = n1950 ^ n1942;
  assign n2147 = n1950 ^ n1935;
  assign n2148 = n2146 & ~n2147;
  assign n2149 = n2148 ^ n1942;
  assign n2153 = n2152 ^ n2149;
  assign n2183 = n2182 ^ n2153;
  assign n2143 = n1906 ^ n1905;
  assign n2144 = ~n1914 & n2143;
  assign n2145 = n2144 ^ n1913;
  assign n2184 = n2183 ^ n2145;
  assign n2139 = n2017 ^ n1993;
  assign n2140 = n2017 ^ n1975;
  assign n2141 = ~n2139 & ~n2140;
  assign n2142 = n2141 ^ n1993;
  assign n2185 = n2184 ^ n2142;
  assign n2135 = n2018 ^ n1952;
  assign n2136 = ~n1953 & ~n2135;
  assign n2137 = n2136 ^ n2018;
  assign n2131 = n1915 ^ n1901;
  assign n2132 = n1915 ^ n1898;
  assign n2133 = ~n2131 & ~n2132;
  assign n2134 = n2133 ^ n1901;
  assign n2138 = n2137 ^ n2134;
  assign n2186 = n2185 ^ n2138;
  assign n2120 = x3 & n1842;
  assign n2121 = x2 & n1844;
  assign n2122 = ~n2120 & ~n2121;
  assign n2123 = ~x3 & n1835;
  assign n2124 = ~x2 & n1839;
  assign n2125 = ~n2123 & ~n2124;
  assign n2126 = n2122 & n2125;
  assign n2112 = x15 & n503;
  assign n2113 = x14 & n507;
  assign n2114 = ~n2112 & ~n2113;
  assign n2115 = ~x15 & n510;
  assign n2116 = ~x14 & n512;
  assign n2117 = ~n2115 & ~n2116;
  assign n2118 = n2114 & n2117;
  assign n2106 = ~x24 & n66;
  assign n2107 = n69 ^ x25;
  assign n2108 = n2107 ^ n69;
  assign n2109 = n70 & n2108;
  assign n2110 = n2109 ^ n69;
  assign n2111 = ~n2106 & ~n2110;
  assign n2119 = n2118 ^ n2111;
  assign n2127 = n2126 ^ n2119;
  assign n2097 = ~x9 & n1004;
  assign n2098 = ~x8 & n1008;
  assign n2099 = ~n2097 & ~n2098;
  assign n2100 = x9 & n1011;
  assign n2101 = x8 & n1013;
  assign n2102 = ~n2100 & ~n2101;
  assign n2103 = n2099 & n2102;
  assign n2089 = ~x19 & n247;
  assign n2090 = ~x18 & n251;
  assign n2091 = ~n2089 & ~n2090;
  assign n2092 = x19 & n254;
  assign n2093 = x18 & n256;
  assign n2094 = ~n2092 & ~n2093;
  assign n2095 = n2091 & n2094;
  assign n2082 = ~x11 & n821;
  assign n2083 = ~x10 & n823;
  assign n2084 = ~n2082 & ~n2083;
  assign n2085 = x11 & n814;
  assign n2086 = x10 & n818;
  assign n2087 = ~n2085 & ~n2086;
  assign n2088 = n2084 & n2087;
  assign n2096 = n2095 ^ n2088;
  assign n2104 = n2103 ^ n2096;
  assign n2074 = x5 & n1578;
  assign n2075 = x4 & n1580;
  assign n2076 = ~n2074 & ~n2075;
  assign n2077 = ~x5 & n1571;
  assign n2078 = ~x4 & n1575;
  assign n2079 = ~n2077 & ~n2078;
  assign n2080 = n2076 & n2079;
  assign n2066 = ~x17 & n346;
  assign n2067 = ~x16 & n350;
  assign n2068 = ~n2066 & ~n2067;
  assign n2069 = x17 & n353;
  assign n2070 = x16 & n355;
  assign n2071 = ~n2069 & ~n2070;
  assign n2072 = n2068 & n2071;
  assign n2059 = x7 & n1223;
  assign n2060 = x6 & n1227;
  assign n2061 = ~n2059 & ~n2060;
  assign n2062 = ~x7 & n1230;
  assign n2063 = ~x6 & n1232;
  assign n2064 = ~n2062 & ~n2063;
  assign n2065 = n2061 & n2064;
  assign n2073 = n2072 ^ n2065;
  assign n2081 = n2080 ^ n2073;
  assign n2105 = n2104 ^ n2081;
  assign n2128 = n2127 ^ n2105;
  assign n2051 = x55 ^ x0;
  assign n2052 = ~n1983 & n2051;
  assign n2053 = n2052 ^ x0;
  assign n2054 = x57 & ~n2053;
  assign n2044 = x23 & n107;
  assign n2045 = x22 & n109;
  assign n2046 = ~n2044 & ~n2045;
  assign n2047 = ~x23 & n100;
  assign n2048 = ~x22 & n104;
  assign n2049 = ~n2047 & ~n2048;
  assign n2050 = n2046 & n2049;
  assign n2055 = n2054 ^ n2050;
  assign n2040 = n2016 ^ n2008;
  assign n2041 = n2016 ^ n2001;
  assign n2042 = n2040 & ~n2041;
  assign n2043 = n2042 ^ n2008;
  assign n2056 = n2055 ^ n2043;
  assign n2037 = n1973 ^ n1959;
  assign n2038 = ~n1974 & n2037;
  assign n2039 = n2038 ^ n1959;
  assign n2057 = n2056 ^ n2039;
  assign n2034 = n1951 ^ n1927;
  assign n2035 = ~n1928 & n2034;
  assign n2036 = n2035 ^ n1951;
  assign n2058 = n2057 ^ n2036;
  assign n2129 = n2128 ^ n2058;
  assign n2031 = n1895 ^ n1892;
  assign n2032 = n1917 & ~n2031;
  assign n2033 = n2032 ^ n1916;
  assign n2130 = n2129 ^ n2033;
  assign n2187 = n2186 ^ n2130;
  assign n2028 = n1918 ^ n1889;
  assign n2029 = ~n2020 & n2028;
  assign n2030 = n2029 ^ n2019;
  assign n2188 = n2187 ^ n2030;
  assign n2193 = n2192 ^ n2188;
  assign n2349 = n2030 & n2187;
  assign n2350 = ~n2030 & ~n2187;
  assign n2351 = ~n2192 & ~n2350;
  assign n2352 = ~n2349 & ~n2351;
  assign n2340 = n2043 ^ n2039;
  assign n2341 = n2056 & ~n2340;
  assign n2342 = n2341 ^ n2055;
  assign n2337 = n2182 ^ n2152;
  assign n2338 = n2153 & ~n2337;
  assign n2339 = n2338 ^ n2182;
  assign n2343 = n2342 ^ n2339;
  assign n2334 = n2127 ^ n2081;
  assign n2335 = n2105 & ~n2334;
  assign n2336 = n2335 ^ n2104;
  assign n2344 = n2343 ^ n2336;
  assign n2330 = n2183 ^ n2142;
  assign n2331 = n2145 ^ n2142;
  assign n2332 = n2330 & n2331;
  assign n2333 = n2332 ^ n2183;
  assign n2345 = n2344 ^ n2333;
  assign n2327 = n2128 ^ n2057;
  assign n2328 = ~n2058 & n2327;
  assign n2329 = n2328 ^ n2128;
  assign n2346 = n2345 ^ n2329;
  assign n2315 = ~x20 & n247;
  assign n2316 = ~x19 & n251;
  assign n2317 = ~n2315 & ~n2316;
  assign n2318 = x20 & n254;
  assign n2319 = x19 & n256;
  assign n2320 = ~n2318 & ~n2319;
  assign n2321 = n2317 & n2320;
  assign n2312 = x58 ^ x57;
  assign n2313 = x0 & n2312;
  assign n2305 = ~x24 & n100;
  assign n2306 = ~x23 & n104;
  assign n2307 = ~n2305 & ~n2306;
  assign n2308 = x24 & n107;
  assign n2309 = x23 & n109;
  assign n2310 = ~n2308 & ~n2309;
  assign n2311 = n2307 & n2310;
  assign n2314 = n2313 ^ n2311;
  assign n2322 = n2321 ^ n2314;
  assign n2302 = n2181 ^ n2160;
  assign n2303 = n2174 & ~n2302;
  assign n2304 = n2303 ^ n2173;
  assign n2323 = n2322 ^ n2304;
  assign n2293 = ~x6 & n1571;
  assign n2294 = ~x5 & n1575;
  assign n2295 = ~n2293 & ~n2294;
  assign n2296 = x6 & n1578;
  assign n2297 = x5 & n1580;
  assign n2298 = ~n2296 & ~n2297;
  assign n2299 = n2295 & n2298;
  assign n2286 = ~x8 & n1230;
  assign n2287 = ~x7 & n1232;
  assign n2288 = ~n2286 & ~n2287;
  assign n2289 = x8 & n1223;
  assign n2290 = x7 & n1227;
  assign n2291 = ~n2289 & ~n2290;
  assign n2292 = n2288 & n2291;
  assign n2300 = n2299 ^ n2292;
  assign n2280 = ~x25 & n66;
  assign n2281 = n69 ^ x26;
  assign n2282 = n2281 ^ n69;
  assign n2283 = n70 & n2282;
  assign n2284 = n2283 ^ n69;
  assign n2285 = ~n2280 & ~n2284;
  assign n2301 = n2300 ^ n2285;
  assign n2324 = n2323 ^ n2301;
  assign n2269 = ~x18 & n346;
  assign n2270 = ~x17 & n350;
  assign n2271 = ~n2269 & ~n2270;
  assign n2272 = x18 & n353;
  assign n2273 = x17 & n355;
  assign n2274 = ~n2272 & ~n2273;
  assign n2275 = n2271 & n2274;
  assign n2261 = x10 & n1011;
  assign n2262 = x9 & n1013;
  assign n2263 = ~n2261 & ~n2262;
  assign n2264 = ~x10 & n1004;
  assign n2265 = ~x9 & n1008;
  assign n2266 = ~n2264 & ~n2265;
  assign n2267 = n2263 & n2266;
  assign n2254 = x12 & n814;
  assign n2255 = x11 & n818;
  assign n2256 = ~n2254 & ~n2255;
  assign n2257 = ~x12 & n821;
  assign n2258 = ~x11 & n823;
  assign n2259 = ~n2257 & ~n2258;
  assign n2260 = n2256 & n2259;
  assign n2268 = n2267 ^ n2260;
  assign n2276 = n2275 ^ n2268;
  assign n2246 = ~x2 & n2161;
  assign n2247 = ~x1 & n2165;
  assign n2248 = ~n2246 & ~n2247;
  assign n2249 = x2 & n2168;
  assign n2250 = x1 & n2170;
  assign n2251 = ~n2249 & ~n2250;
  assign n2252 = n2248 & n2251;
  assign n2238 = ~x4 & n1835;
  assign n2239 = ~x3 & n1839;
  assign n2240 = ~n2238 & ~n2239;
  assign n2241 = x4 & n1842;
  assign n2242 = x3 & n1844;
  assign n2243 = ~n2241 & ~n2242;
  assign n2244 = n2240 & n2243;
  assign n2231 = ~x16 & n510;
  assign n2232 = ~x15 & n512;
  assign n2233 = ~n2231 & ~n2232;
  assign n2234 = x16 & n503;
  assign n2235 = x15 & n507;
  assign n2236 = ~n2234 & ~n2235;
  assign n2237 = n2233 & n2236;
  assign n2245 = n2244 ^ n2237;
  assign n2253 = n2252 ^ n2245;
  assign n2277 = n2276 ^ n2253;
  assign n2222 = x22 & n154;
  assign n2223 = x21 & n156;
  assign n2224 = ~n2222 & ~n2223;
  assign n2225 = ~x22 & n147;
  assign n2226 = ~x21 & n151;
  assign n2227 = ~n2225 & ~n2226;
  assign n2228 = n2224 & n2227;
  assign n2215 = ~x14 & n650;
  assign n2216 = ~x13 & n654;
  assign n2217 = ~n2215 & ~n2216;
  assign n2218 = x14 & n657;
  assign n2219 = x13 & n659;
  assign n2220 = ~n2218 & ~n2219;
  assign n2221 = n2217 & n2220;
  assign n2229 = n2228 ^ n2221;
  assign n2214 = ~n2050 & n2054;
  assign n2230 = n2229 ^ n2214;
  assign n2278 = n2277 ^ n2230;
  assign n2209 = n2103 ^ n2088;
  assign n2210 = n2096 & ~n2209;
  assign n2211 = n2210 ^ n2095;
  assign n2205 = n2080 ^ n2072;
  assign n2206 = n2080 ^ n2065;
  assign n2207 = n2205 & ~n2206;
  assign n2208 = n2207 ^ n2072;
  assign n2212 = n2211 ^ n2208;
  assign n2201 = n2126 ^ n2111;
  assign n2202 = n2126 ^ n2118;
  assign n2203 = n2201 & ~n2202;
  assign n2204 = n2203 ^ n2111;
  assign n2213 = n2212 ^ n2204;
  assign n2279 = n2278 ^ n2213;
  assign n2325 = n2324 ^ n2279;
  assign n2198 = n2185 ^ n2137;
  assign n2199 = n2138 & ~n2198;
  assign n2200 = n2199 ^ n2185;
  assign n2326 = n2325 ^ n2200;
  assign n2347 = n2346 ^ n2326;
  assign n2194 = n2186 ^ n2129;
  assign n2195 = n2186 ^ n2033;
  assign n2196 = ~n2194 & n2195;
  assign n2197 = n2196 ^ n2129;
  assign n2348 = n2347 ^ n2197;
  assign n2353 = n2352 ^ n2348;
  assign n2526 = ~n2197 & n2347;
  assign n2527 = n2197 & ~n2347;
  assign n2528 = ~n2352 & ~n2527;
  assign n2529 = ~n2526 & ~n2528;
  assign n2516 = n2275 ^ n2267;
  assign n2517 = n2275 ^ n2260;
  assign n2518 = n2516 & ~n2517;
  assign n2519 = n2518 ^ n2267;
  assign n2513 = n2299 ^ n2285;
  assign n2514 = ~n2300 & n2513;
  assign n2515 = n2514 ^ n2285;
  assign n2520 = n2519 ^ n2515;
  assign n2510 = n2252 ^ n2237;
  assign n2511 = n2245 & ~n2510;
  assign n2512 = n2511 ^ n2244;
  assign n2521 = n2520 ^ n2512;
  assign n2506 = n2322 ^ n2301;
  assign n2507 = n2323 & ~n2506;
  assign n2508 = n2507 ^ n2301;
  assign n2503 = n2208 ^ n2204;
  assign n2504 = n2212 & ~n2503;
  assign n2505 = n2504 ^ n2211;
  assign n2509 = n2508 ^ n2505;
  assign n2522 = n2521 ^ n2509;
  assign n2498 = n2324 ^ n2278;
  assign n2499 = n2324 ^ n2213;
  assign n2500 = n2498 & n2499;
  assign n2501 = n2500 ^ n2278;
  assign n2495 = n2342 ^ n2336;
  assign n2496 = ~n2343 & n2495;
  assign n2497 = n2496 ^ n2336;
  assign n2502 = n2501 ^ n2497;
  assign n2523 = n2522 ^ n2502;
  assign n2483 = x15 & n657;
  assign n2484 = x14 & n659;
  assign n2485 = ~n2483 & ~n2484;
  assign n2486 = ~x15 & n650;
  assign n2487 = ~x14 & n654;
  assign n2488 = ~n2486 & ~n2487;
  assign n2489 = n2485 & n2488;
  assign n2478 = x57 ^ x0;
  assign n2479 = ~n2312 & n2478;
  assign n2480 = n2479 ^ x0;
  assign n2481 = x59 & ~n2480;
  assign n2471 = ~x25 & n100;
  assign n2472 = ~x24 & n104;
  assign n2473 = ~n2471 & ~n2472;
  assign n2474 = x25 & n107;
  assign n2475 = x24 & n109;
  assign n2476 = ~n2474 & ~n2475;
  assign n2477 = n2473 & n2476;
  assign n2482 = n2481 ^ n2477;
  assign n2490 = n2489 ^ n2482;
  assign n2468 = n2321 ^ n2311;
  assign n2469 = ~n2314 & ~n2468;
  assign n2470 = n2469 ^ n2313;
  assign n2491 = n2490 ^ n2470;
  assign n2459 = ~x7 & n1571;
  assign n2460 = ~x6 & n1575;
  assign n2461 = ~n2459 & ~n2460;
  assign n2462 = x7 & n1578;
  assign n2463 = x6 & n1580;
  assign n2464 = ~n2462 & ~n2463;
  assign n2465 = n2461 & n2464;
  assign n2451 = x19 & n353;
  assign n2452 = x18 & n355;
  assign n2453 = ~n2451 & ~n2452;
  assign n2454 = ~x19 & n346;
  assign n2455 = ~x18 & n350;
  assign n2456 = ~n2454 & ~n2455;
  assign n2457 = n2453 & n2456;
  assign n2444 = ~x9 & n1230;
  assign n2445 = ~x8 & n1232;
  assign n2446 = ~n2444 & ~n2445;
  assign n2447 = x9 & n1223;
  assign n2448 = x8 & n1227;
  assign n2449 = ~n2447 & ~n2448;
  assign n2450 = n2446 & n2449;
  assign n2458 = n2457 ^ n2450;
  assign n2466 = n2465 ^ n2458;
  assign n2441 = n2221 ^ n2214;
  assign n2442 = n2229 & n2441;
  assign n2443 = n2442 ^ n2228;
  assign n2467 = n2466 ^ n2443;
  assign n2492 = n2491 ^ n2467;
  assign n2431 = ~x5 & n1835;
  assign n2432 = ~x4 & n1839;
  assign n2433 = ~n2431 & ~n2432;
  assign n2434 = x5 & n1842;
  assign n2435 = x4 & n1844;
  assign n2436 = ~n2434 & ~n2435;
  assign n2437 = n2433 & n2436;
  assign n2423 = ~x17 & n510;
  assign n2424 = ~x16 & n512;
  assign n2425 = ~n2423 & ~n2424;
  assign n2426 = x17 & n503;
  assign n2427 = x16 & n507;
  assign n2428 = ~n2426 & ~n2427;
  assign n2429 = n2425 & n2428;
  assign n2417 = ~x26 & n66;
  assign n2418 = n69 ^ x27;
  assign n2419 = n2418 ^ n69;
  assign n2420 = n70 & n2419;
  assign n2421 = n2420 ^ n69;
  assign n2422 = ~n2417 & ~n2421;
  assign n2430 = n2429 ^ n2422;
  assign n2438 = n2437 ^ n2430;
  assign n2408 = ~x11 & n1004;
  assign n2409 = ~x10 & n1008;
  assign n2410 = ~n2408 & ~n2409;
  assign n2411 = x11 & n1011;
  assign n2412 = x10 & n1013;
  assign n2413 = ~n2411 & ~n2412;
  assign n2414 = n2410 & n2413;
  assign n2400 = x21 & n254;
  assign n2401 = x20 & n256;
  assign n2402 = ~n2400 & ~n2401;
  assign n2403 = ~x21 & n247;
  assign n2404 = ~x20 & n251;
  assign n2405 = ~n2403 & ~n2404;
  assign n2406 = n2402 & n2405;
  assign n2393 = ~x13 & n821;
  assign n2394 = ~x12 & n823;
  assign n2395 = ~n2393 & ~n2394;
  assign n2396 = x13 & n814;
  assign n2397 = x12 & n818;
  assign n2398 = ~n2396 & ~n2397;
  assign n2399 = n2395 & n2398;
  assign n2407 = n2406 ^ n2399;
  assign n2415 = n2414 ^ n2407;
  assign n2379 = ~x59 & n2312;
  assign n2380 = x1 & n2379;
  assign n2381 = x59 ^ x58;
  assign n2382 = ~n2312 & n2381;
  assign n2383 = ~x59 & n2382;
  assign n2384 = x0 & n2383;
  assign n2385 = ~n2380 & ~n2384;
  assign n2386 = x59 & n2312;
  assign n2387 = ~x1 & n2386;
  assign n2388 = x59 & n2382;
  assign n2389 = ~x0 & n2388;
  assign n2390 = ~n2387 & ~n2389;
  assign n2391 = n2385 & n2390;
  assign n2371 = x3 & n2168;
  assign n2372 = x2 & n2170;
  assign n2373 = ~n2371 & ~n2372;
  assign n2374 = ~x3 & n2161;
  assign n2375 = ~x2 & n2165;
  assign n2376 = ~n2374 & ~n2375;
  assign n2377 = n2373 & n2376;
  assign n2364 = x23 & n154;
  assign n2365 = x22 & n156;
  assign n2366 = ~n2364 & ~n2365;
  assign n2367 = ~x23 & n147;
  assign n2368 = ~x22 & n151;
  assign n2369 = ~n2367 & ~n2368;
  assign n2370 = n2366 & n2369;
  assign n2378 = n2377 ^ n2370;
  assign n2392 = n2391 ^ n2378;
  assign n2416 = n2415 ^ n2392;
  assign n2439 = n2438 ^ n2416;
  assign n2361 = n2253 ^ n2230;
  assign n2362 = n2277 & n2361;
  assign n2363 = n2362 ^ n2276;
  assign n2440 = n2439 ^ n2363;
  assign n2493 = n2492 ^ n2440;
  assign n2358 = n2333 ^ n2329;
  assign n2359 = ~n2345 & n2358;
  assign n2360 = n2359 ^ n2344;
  assign n2494 = n2493 ^ n2360;
  assign n2524 = n2523 ^ n2494;
  assign n2354 = n2346 ^ n2325;
  assign n2355 = n2346 ^ n2200;
  assign n2356 = ~n2354 & n2355;
  assign n2357 = n2356 ^ n2325;
  assign n2525 = n2524 ^ n2357;
  assign n2530 = n2529 ^ n2525;
  assign n2697 = ~n2357 & ~n2524;
  assign n2698 = n2357 & n2524;
  assign n2699 = ~n2529 & ~n2698;
  assign n2700 = ~n2697 & ~n2699;
  assign n2682 = ~x20 & n346;
  assign n2683 = ~x19 & n350;
  assign n2684 = ~n2682 & ~n2683;
  assign n2685 = x20 & n353;
  assign n2686 = x19 & n355;
  assign n2687 = ~n2685 & ~n2686;
  assign n2688 = n2684 & n2687;
  assign n2674 = ~x14 & n821;
  assign n2675 = ~x13 & n823;
  assign n2676 = ~n2674 & ~n2675;
  assign n2677 = x14 & n814;
  assign n2678 = x13 & n818;
  assign n2679 = ~n2677 & ~n2678;
  assign n2680 = n2676 & n2679;
  assign n2667 = ~x12 & n1004;
  assign n2668 = ~x11 & n1008;
  assign n2669 = ~n2667 & ~n2668;
  assign n2670 = x12 & n1011;
  assign n2671 = x11 & n1013;
  assign n2672 = ~n2670 & ~n2671;
  assign n2673 = n2669 & n2672;
  assign n2681 = n2680 ^ n2673;
  assign n2689 = n2688 ^ n2681;
  assign n2663 = n2437 ^ n2429;
  assign n2664 = n2430 & ~n2663;
  assign n2665 = n2664 ^ n2422;
  assign n2660 = n2391 ^ n2370;
  assign n2661 = n2378 & ~n2660;
  assign n2662 = n2661 ^ n2377;
  assign n2666 = n2665 ^ n2662;
  assign n2690 = n2689 ^ n2666;
  assign n2657 = ~n2477 & n2481;
  assign n2654 = n2414 ^ n2399;
  assign n2655 = n2407 & ~n2654;
  assign n2656 = n2655 ^ n2406;
  assign n2658 = n2657 ^ n2656;
  assign n2651 = n2465 ^ n2450;
  assign n2652 = n2458 & ~n2651;
  assign n2653 = n2652 ^ n2457;
  assign n2659 = n2658 ^ n2653;
  assign n2691 = n2690 ^ n2659;
  assign n2648 = n2438 ^ n2415;
  assign n2649 = ~n2416 & n2648;
  assign n2650 = n2649 ^ n2438;
  assign n2692 = n2691 ^ n2650;
  assign n2638 = ~x4 & n2161;
  assign n2639 = ~x3 & n2165;
  assign n2640 = ~n2638 & ~n2639;
  assign n2641 = x4 & n2168;
  assign n2642 = x3 & n2170;
  assign n2643 = ~n2641 & ~n2642;
  assign n2644 = n2640 & n2643;
  assign n2630 = x18 & n503;
  assign n2631 = x17 & n507;
  assign n2632 = ~n2630 & ~n2631;
  assign n2633 = ~x18 & n510;
  assign n2634 = ~x17 & n512;
  assign n2635 = ~n2633 & ~n2634;
  assign n2636 = n2632 & n2635;
  assign n2623 = ~x6 & n1835;
  assign n2624 = ~x5 & n1839;
  assign n2625 = ~n2623 & ~n2624;
  assign n2626 = x6 & n1842;
  assign n2627 = x5 & n1844;
  assign n2628 = ~n2626 & ~n2627;
  assign n2629 = n2625 & n2628;
  assign n2637 = n2636 ^ n2629;
  assign n2645 = n2644 ^ n2637;
  assign n2620 = n2519 ^ n2512;
  assign n2621 = ~n2520 & n2620;
  assign n2622 = n2621 ^ n2512;
  assign n2646 = n2645 ^ n2622;
  assign n2617 = n2482 ^ n2470;
  assign n2618 = n2490 & n2617;
  assign n2619 = n2618 ^ n2489;
  assign n2647 = n2646 ^ n2619;
  assign n2693 = n2692 ^ n2647;
  assign n2613 = n2492 ^ n2439;
  assign n2614 = n2492 ^ n2363;
  assign n2615 = ~n2613 & n2614;
  assign n2616 = n2615 ^ n2439;
  assign n2694 = n2693 ^ n2616;
  assign n2600 = x22 & n254;
  assign n2601 = x21 & n256;
  assign n2602 = ~n2600 & ~n2601;
  assign n2603 = ~x22 & n247;
  assign n2604 = ~x21 & n251;
  assign n2605 = ~n2603 & ~n2604;
  assign n2606 = n2602 & n2605;
  assign n2597 = x60 ^ x59;
  assign n2598 = x0 & n2597;
  assign n2590 = ~x26 & n100;
  assign n2591 = ~x25 & n104;
  assign n2592 = ~n2590 & ~n2591;
  assign n2593 = x26 & n107;
  assign n2594 = x25 & n109;
  assign n2595 = ~n2593 & ~n2594;
  assign n2596 = n2592 & n2595;
  assign n2599 = n2598 ^ n2596;
  assign n2607 = n2606 ^ n2599;
  assign n2582 = ~x16 & n650;
  assign n2583 = ~x15 & n654;
  assign n2584 = ~n2582 & ~n2583;
  assign n2585 = x16 & n657;
  assign n2586 = x15 & n659;
  assign n2587 = ~n2585 & ~n2586;
  assign n2588 = n2584 & n2587;
  assign n2574 = x24 & n154;
  assign n2575 = x23 & n156;
  assign n2576 = ~n2574 & ~n2575;
  assign n2577 = ~x24 & n147;
  assign n2578 = ~x23 & n151;
  assign n2579 = ~n2577 & ~n2578;
  assign n2580 = n2576 & n2579;
  assign n2567 = ~x2 & n2386;
  assign n2568 = ~x1 & n2388;
  assign n2569 = ~n2567 & ~n2568;
  assign n2570 = x2 & n2379;
  assign n2571 = x1 & n2383;
  assign n2572 = ~n2570 & ~n2571;
  assign n2573 = n2569 & n2572;
  assign n2581 = n2580 ^ n2573;
  assign n2589 = n2588 ^ n2581;
  assign n2608 = n2607 ^ n2589;
  assign n2558 = x10 & n1223;
  assign n2559 = x9 & n1227;
  assign n2560 = ~n2558 & ~n2559;
  assign n2561 = ~x10 & n1230;
  assign n2562 = ~x9 & n1232;
  assign n2563 = ~n2561 & ~n2562;
  assign n2564 = n2560 & n2563;
  assign n2551 = x8 & n1578;
  assign n2552 = x7 & n1580;
  assign n2553 = ~n2551 & ~n2552;
  assign n2554 = ~x8 & n1571;
  assign n2555 = ~x7 & n1575;
  assign n2556 = ~n2554 & ~n2555;
  assign n2557 = n2553 & n2556;
  assign n2565 = n2564 ^ n2557;
  assign n2545 = ~x27 & n66;
  assign n2546 = n69 ^ x28;
  assign n2547 = n2546 ^ n69;
  assign n2548 = n70 & n2547;
  assign n2549 = n2548 ^ n69;
  assign n2550 = ~n2545 & ~n2549;
  assign n2566 = n2565 ^ n2550;
  assign n2609 = n2608 ^ n2566;
  assign n2542 = n2491 ^ n2443;
  assign n2543 = n2467 & n2542;
  assign n2544 = n2543 ^ n2466;
  assign n2610 = n2609 ^ n2544;
  assign n2539 = n2521 ^ n2508;
  assign n2540 = ~n2509 & n2539;
  assign n2541 = n2540 ^ n2521;
  assign n2611 = n2610 ^ n2541;
  assign n2535 = n2522 ^ n2501;
  assign n2536 = n2522 ^ n2497;
  assign n2537 = ~n2535 & ~n2536;
  assign n2538 = n2537 ^ n2501;
  assign n2612 = n2611 ^ n2538;
  assign n2695 = n2694 ^ n2612;
  assign n2531 = n2523 ^ n2493;
  assign n2532 = n2523 ^ n2360;
  assign n2533 = n2531 & n2532;
  assign n2534 = n2533 ^ n2493;
  assign n2696 = n2695 ^ n2534;
  assign n2701 = n2700 ^ n2696;
  assign n2886 = n2534 & n2695;
  assign n2887 = ~n2534 & ~n2695;
  assign n2888 = ~n2700 & ~n2887;
  assign n2889 = ~n2886 & ~n2888;
  assign n2872 = ~x15 & n821;
  assign n2873 = ~x14 & n823;
  assign n2874 = ~n2872 & ~n2873;
  assign n2875 = x15 & n814;
  assign n2876 = x14 & n818;
  assign n2877 = ~n2875 & ~n2876;
  assign n2878 = n2874 & n2877;
  assign n2864 = x27 & n107;
  assign n2865 = x26 & n109;
  assign n2866 = ~n2864 & ~n2865;
  assign n2867 = ~x27 & n100;
  assign n2868 = ~x26 & n104;
  assign n2869 = ~n2867 & ~n2868;
  assign n2870 = n2866 & n2869;
  assign n2857 = ~x23 & n247;
  assign n2858 = ~x22 & n251;
  assign n2859 = ~n2857 & ~n2858;
  assign n2860 = x23 & n254;
  assign n2861 = x22 & n256;
  assign n2862 = ~n2860 & ~n2861;
  assign n2863 = n2859 & n2862;
  assign n2871 = n2870 ^ n2863;
  assign n2879 = n2878 ^ n2871;
  assign n2853 = n2644 ^ n2636;
  assign n2854 = ~n2637 & n2853;
  assign n2855 = n2854 ^ n2644;
  assign n2850 = n2588 ^ n2580;
  assign n2851 = ~n2581 & n2850;
  assign n2852 = n2851 ^ n2588;
  assign n2856 = n2855 ^ n2852;
  assign n2880 = n2879 ^ n2856;
  assign n2843 = n2606 ^ n2598;
  assign n2844 = n2606 ^ n2596;
  assign n2845 = ~n2843 & ~n2844;
  assign n2846 = n2845 ^ n2598;
  assign n2840 = n2564 ^ n2550;
  assign n2841 = ~n2565 & n2840;
  assign n2842 = n2841 ^ n2550;
  assign n2847 = n2846 ^ n2842;
  assign n2837 = n2688 ^ n2673;
  assign n2838 = n2681 & ~n2837;
  assign n2839 = n2838 ^ n2680;
  assign n2848 = n2847 ^ n2839;
  assign n2834 = n2689 ^ n2665;
  assign n2835 = ~n2666 & n2834;
  assign n2836 = n2835 ^ n2689;
  assign n2849 = n2848 ^ n2836;
  assign n2881 = n2880 ^ n2849;
  assign n2826 = x59 ^ x0;
  assign n2827 = ~n2597 & n2826;
  assign n2828 = n2827 ^ x0;
  assign n2829 = x61 & ~n2828;
  assign n2820 = ~x28 & n66;
  assign n2821 = n69 ^ x29;
  assign n2822 = n2821 ^ n69;
  assign n2823 = n70 & n2822;
  assign n2824 = n2823 ^ n69;
  assign n2825 = ~n2820 & ~n2824;
  assign n2830 = n2829 ^ n2825;
  assign n2812 = x3 & n2379;
  assign n2813 = x2 & n2383;
  assign n2814 = ~n2812 & ~n2813;
  assign n2815 = ~x3 & n2386;
  assign n2816 = ~x2 & n2388;
  assign n2817 = ~n2815 & ~n2816;
  assign n2818 = n2814 & n2817;
  assign n2799 = x61 & n2597;
  assign n2800 = ~x1 & n2799;
  assign n2801 = x61 ^ x60;
  assign n2802 = ~n2597 & n2801;
  assign n2803 = x61 & n2802;
  assign n2804 = ~x0 & n2803;
  assign n2805 = ~n2800 & ~n2804;
  assign n2806 = ~x61 & n2597;
  assign n2807 = x1 & n2806;
  assign n2808 = ~x61 & n2802;
  assign n2809 = x0 & n2808;
  assign n2810 = ~n2807 & ~n2809;
  assign n2811 = n2805 & n2810;
  assign n2819 = n2818 ^ n2811;
  assign n2831 = n2830 ^ n2819;
  assign n2796 = n2656 ^ n2653;
  assign n2797 = ~n2658 & ~n2796;
  assign n2798 = n2797 ^ n2657;
  assign n2832 = n2831 ^ n2798;
  assign n2792 = n2607 ^ n2566;
  assign n2793 = n2589 ^ n2566;
  assign n2794 = ~n2792 & ~n2793;
  assign n2795 = n2794 ^ n2607;
  assign n2833 = n2832 ^ n2795;
  assign n2882 = n2881 ^ n2833;
  assign n2781 = ~x19 & n510;
  assign n2782 = ~x18 & n512;
  assign n2783 = ~n2781 & ~n2782;
  assign n2784 = x19 & n503;
  assign n2785 = x18 & n507;
  assign n2786 = ~n2784 & ~n2785;
  assign n2787 = n2783 & n2786;
  assign n2773 = ~x9 & n1571;
  assign n2774 = ~x8 & n1575;
  assign n2775 = ~n2773 & ~n2774;
  assign n2776 = x9 & n1578;
  assign n2777 = x8 & n1580;
  assign n2778 = ~n2776 & ~n2777;
  assign n2779 = n2775 & n2778;
  assign n2766 = x25 & n154;
  assign n2767 = x24 & n156;
  assign n2768 = ~n2766 & ~n2767;
  assign n2769 = ~x25 & n147;
  assign n2770 = ~x24 & n151;
  assign n2771 = ~n2769 & ~n2770;
  assign n2772 = n2768 & n2771;
  assign n2780 = n2779 ^ n2772;
  assign n2788 = n2787 ^ n2780;
  assign n2757 = ~x17 & n650;
  assign n2758 = ~x16 & n654;
  assign n2759 = ~n2757 & ~n2758;
  assign n2760 = x17 & n657;
  assign n2761 = x16 & n659;
  assign n2762 = ~n2760 & ~n2761;
  assign n2763 = n2759 & n2762;
  assign n2749 = ~x7 & n1835;
  assign n2750 = ~x6 & n1839;
  assign n2751 = ~n2749 & ~n2750;
  assign n2752 = x7 & n1842;
  assign n2753 = x6 & n1844;
  assign n2754 = ~n2752 & ~n2753;
  assign n2755 = n2751 & n2754;
  assign n2742 = ~x5 & n2161;
  assign n2743 = ~x4 & n2165;
  assign n2744 = ~n2742 & ~n2743;
  assign n2745 = x5 & n2168;
  assign n2746 = x4 & n2170;
  assign n2747 = ~n2745 & ~n2746;
  assign n2748 = n2744 & n2747;
  assign n2756 = n2755 ^ n2748;
  assign n2764 = n2763 ^ n2756;
  assign n2734 = x11 & n1223;
  assign n2735 = x10 & n1227;
  assign n2736 = ~n2734 & ~n2735;
  assign n2737 = ~x11 & n1230;
  assign n2738 = ~x10 & n1232;
  assign n2739 = ~n2737 & ~n2738;
  assign n2740 = n2736 & n2739;
  assign n2726 = ~x13 & n1004;
  assign n2727 = ~x12 & n1008;
  assign n2728 = ~n2726 & ~n2727;
  assign n2729 = x13 & n1011;
  assign n2730 = x12 & n1013;
  assign n2731 = ~n2729 & ~n2730;
  assign n2732 = n2728 & n2731;
  assign n2719 = ~x21 & n346;
  assign n2720 = ~x20 & n350;
  assign n2721 = ~n2719 & ~n2720;
  assign n2722 = x21 & n353;
  assign n2723 = x20 & n355;
  assign n2724 = ~n2722 & ~n2723;
  assign n2725 = n2721 & n2724;
  assign n2733 = n2732 ^ n2725;
  assign n2741 = n2740 ^ n2733;
  assign n2765 = n2764 ^ n2741;
  assign n2789 = n2788 ^ n2765;
  assign n2715 = n2645 ^ n2619;
  assign n2716 = n2622 ^ n2619;
  assign n2717 = n2715 & ~n2716;
  assign n2718 = n2717 ^ n2645;
  assign n2790 = n2789 ^ n2718;
  assign n2712 = n2690 ^ n2650;
  assign n2713 = n2691 & n2712;
  assign n2714 = n2713 ^ n2650;
  assign n2791 = n2790 ^ n2714;
  assign n2883 = n2882 ^ n2791;
  assign n2708 = n2647 ^ n2616;
  assign n2709 = ~n2693 & ~n2708;
  assign n2710 = n2709 ^ n2692;
  assign n2705 = n2544 ^ n2541;
  assign n2706 = ~n2610 & ~n2705;
  assign n2707 = n2706 ^ n2609;
  assign n2711 = n2710 ^ n2707;
  assign n2884 = n2883 ^ n2711;
  assign n2702 = n2694 ^ n2611;
  assign n2703 = ~n2612 & n2702;
  assign n2704 = n2703 ^ n2694;
  assign n2885 = n2884 ^ n2704;
  assign n2890 = n2889 ^ n2885;
  assign n3068 = n2704 & n2884;
  assign n3069 = ~n2704 & ~n2884;
  assign n3070 = ~n2889 & ~n3069;
  assign n3071 = ~n3068 & ~n3070;
  assign n3054 = x8 & n1842;
  assign n3055 = x7 & n1844;
  assign n3056 = ~n3054 & ~n3055;
  assign n3057 = ~x8 & n1835;
  assign n3058 = ~x7 & n1839;
  assign n3059 = ~n3057 & ~n3058;
  assign n3060 = n3056 & n3059;
  assign n3046 = ~x26 & n147;
  assign n3047 = ~x25 & n151;
  assign n3048 = ~n3046 & ~n3047;
  assign n3049 = x26 & n154;
  assign n3050 = x25 & n156;
  assign n3051 = ~n3049 & ~n3050;
  assign n3052 = n3048 & n3051;
  assign n3039 = ~x20 & n510;
  assign n3040 = ~x19 & n512;
  assign n3041 = ~n3039 & ~n3040;
  assign n3042 = x20 & n503;
  assign n3043 = x19 & n507;
  assign n3044 = ~n3042 & ~n3043;
  assign n3045 = n3041 & n3044;
  assign n3053 = n3052 ^ n3045;
  assign n3061 = n3060 ^ n3053;
  assign n3034 = x62 ^ x61;
  assign n3035 = x0 & n3034;
  assign n3028 = ~x29 & n66;
  assign n3029 = n69 ^ x30;
  assign n3030 = n3029 ^ n69;
  assign n3031 = n70 & n3030;
  assign n3032 = n3031 ^ n69;
  assign n3033 = ~n3028 & ~n3032;
  assign n3036 = n3035 ^ n3033;
  assign n3021 = ~x28 & n100;
  assign n3022 = ~x27 & n104;
  assign n3023 = ~n3021 & ~n3022;
  assign n3024 = x28 & n107;
  assign n3025 = x27 & n109;
  assign n3026 = ~n3024 & ~n3025;
  assign n3027 = n3023 & n3026;
  assign n3037 = n3036 ^ n3027;
  assign n3013 = x4 & n2379;
  assign n3014 = x3 & n2383;
  assign n3015 = ~n3013 & ~n3014;
  assign n3016 = ~x4 & n2386;
  assign n3017 = ~x3 & n2388;
  assign n3018 = ~n3016 & ~n3017;
  assign n3019 = n3015 & n3018;
  assign n3005 = ~x6 & n2161;
  assign n3006 = ~x5 & n2165;
  assign n3007 = ~n3005 & ~n3006;
  assign n3008 = x6 & n2168;
  assign n3009 = x5 & n2170;
  assign n3010 = ~n3008 & ~n3009;
  assign n3011 = n3007 & n3010;
  assign n2998 = ~x18 & n650;
  assign n2999 = ~x17 & n654;
  assign n3000 = ~n2998 & ~n2999;
  assign n3001 = x18 & n657;
  assign n3002 = x17 & n659;
  assign n3003 = ~n3001 & ~n3002;
  assign n3004 = n3000 & n3003;
  assign n3012 = n3011 ^ n3004;
  assign n3020 = n3019 ^ n3012;
  assign n3038 = n3037 ^ n3020;
  assign n3062 = n3061 ^ n3038;
  assign n2995 = n2880 ^ n2848;
  assign n2996 = n2849 & ~n2995;
  assign n2997 = n2996 ^ n2880;
  assign n3063 = n3062 ^ n2997;
  assign n2991 = n2831 ^ n2795;
  assign n2992 = n2798 ^ n2795;
  assign n2993 = ~n2991 & ~n2992;
  assign n2994 = n2993 ^ n2831;
  assign n3064 = n3063 ^ n2994;
  assign n2978 = ~x14 & n1004;
  assign n2979 = ~x13 & n1008;
  assign n2980 = ~n2978 & ~n2979;
  assign n2981 = x14 & n1011;
  assign n2982 = x13 & n1013;
  assign n2983 = ~n2981 & ~n2982;
  assign n2984 = n2980 & n2983;
  assign n2970 = x24 & n254;
  assign n2971 = x23 & n256;
  assign n2972 = ~n2970 & ~n2971;
  assign n2973 = ~x24 & n247;
  assign n2974 = ~x23 & n251;
  assign n2975 = ~n2973 & ~n2974;
  assign n2976 = n2972 & n2975;
  assign n2963 = ~x16 & n821;
  assign n2964 = ~x15 & n823;
  assign n2965 = ~n2963 & ~n2964;
  assign n2966 = x16 & n814;
  assign n2967 = x15 & n818;
  assign n2968 = ~n2966 & ~n2967;
  assign n2969 = n2965 & n2968;
  assign n2977 = n2976 ^ n2969;
  assign n2985 = n2984 ^ n2977;
  assign n2955 = ~x10 & n1571;
  assign n2956 = ~x9 & n1575;
  assign n2957 = ~n2955 & ~n2956;
  assign n2958 = x10 & n1578;
  assign n2959 = x9 & n1580;
  assign n2960 = ~n2958 & ~n2959;
  assign n2961 = n2957 & n2960;
  assign n2947 = ~x22 & n346;
  assign n2948 = ~x21 & n350;
  assign n2949 = ~n2947 & ~n2948;
  assign n2950 = x22 & n353;
  assign n2951 = x21 & n355;
  assign n2952 = ~n2950 & ~n2951;
  assign n2953 = n2949 & n2952;
  assign n2940 = ~x12 & n1230;
  assign n2941 = ~x11 & n1232;
  assign n2942 = ~n2940 & ~n2941;
  assign n2943 = x12 & n1223;
  assign n2944 = x11 & n1227;
  assign n2945 = ~n2943 & ~n2944;
  assign n2946 = n2942 & n2945;
  assign n2954 = n2953 ^ n2946;
  assign n2962 = n2961 ^ n2954;
  assign n2986 = n2985 ^ n2962;
  assign n2937 = n2830 ^ n2811;
  assign n2938 = n2819 & ~n2937;
  assign n2939 = n2938 ^ n2818;
  assign n2987 = n2986 ^ n2939;
  assign n2931 = n2787 ^ n2772;
  assign n2932 = n2780 & ~n2931;
  assign n2933 = n2932 ^ n2779;
  assign n2928 = n2740 ^ n2725;
  assign n2929 = n2733 & ~n2928;
  assign n2930 = n2929 ^ n2732;
  assign n2934 = n2933 ^ n2930;
  assign n2925 = n2763 ^ n2748;
  assign n2926 = n2756 & ~n2925;
  assign n2927 = n2926 ^ n2755;
  assign n2935 = n2934 ^ n2927;
  assign n2922 = n2879 ^ n2855;
  assign n2923 = ~n2856 & n2922;
  assign n2924 = n2923 ^ n2879;
  assign n2936 = n2935 ^ n2924;
  assign n2988 = n2987 ^ n2936;
  assign n2911 = ~x2 & n2799;
  assign n2912 = ~x1 & n2803;
  assign n2913 = ~n2911 & ~n2912;
  assign n2914 = x2 & n2806;
  assign n2915 = x1 & n2808;
  assign n2916 = ~n2914 & ~n2915;
  assign n2917 = n2913 & n2916;
  assign n2910 = ~n2825 & n2829;
  assign n2918 = n2917 ^ n2910;
  assign n2907 = n2878 ^ n2863;
  assign n2908 = n2871 & ~n2907;
  assign n2909 = n2908 ^ n2870;
  assign n2919 = n2918 ^ n2909;
  assign n2904 = n2846 ^ n2839;
  assign n2905 = n2847 & ~n2904;
  assign n2906 = n2905 ^ n2839;
  assign n2920 = n2919 ^ n2906;
  assign n2901 = n2788 ^ n2764;
  assign n2902 = ~n2765 & n2901;
  assign n2903 = n2902 ^ n2788;
  assign n2921 = n2920 ^ n2903;
  assign n2989 = n2988 ^ n2921;
  assign n2897 = n2789 ^ n2714;
  assign n2898 = n2718 ^ n2714;
  assign n2899 = n2897 & ~n2898;
  assign n2900 = n2899 ^ n2789;
  assign n2990 = n2989 ^ n2900;
  assign n3065 = n3064 ^ n2990;
  assign n2894 = n2833 ^ n2791;
  assign n2895 = ~n2882 & ~n2894;
  assign n2896 = n2895 ^ n2881;
  assign n3066 = n3065 ^ n2896;
  assign n2891 = n2883 ^ n2710;
  assign n2892 = ~n2711 & n2891;
  assign n2893 = n2892 ^ n2883;
  assign n3067 = n3066 ^ n2893;
  assign n3072 = n3071 ^ n3067;
  assign n3269 = n2893 & n3066;
  assign n3270 = ~n2893 & ~n3066;
  assign n3271 = ~n3071 & ~n3270;
  assign n3272 = ~n3269 & ~n3271;
  assign n3254 = x7 & n2168;
  assign n3255 = x6 & n2170;
  assign n3256 = ~n3254 & ~n3255;
  assign n3257 = ~x7 & n2161;
  assign n3258 = ~x6 & n2165;
  assign n3259 = ~n3257 & ~n3258;
  assign n3260 = n3256 & n3259;
  assign n3246 = ~x9 & n1835;
  assign n3247 = ~x8 & n1839;
  assign n3248 = ~n3246 & ~n3247;
  assign n3249 = x9 & n1842;
  assign n3250 = x8 & n1844;
  assign n3251 = ~n3249 & ~n3250;
  assign n3252 = n3248 & n3251;
  assign n3239 = x21 & n503;
  assign n3240 = x20 & n507;
  assign n3241 = ~n3239 & ~n3240;
  assign n3242 = ~x21 & n510;
  assign n3243 = ~x20 & n512;
  assign n3244 = ~n3242 & ~n3243;
  assign n3245 = n3241 & n3244;
  assign n3253 = n3252 ^ n3245;
  assign n3261 = n3260 ^ n3253;
  assign n3231 = ~x27 & n147;
  assign n3232 = ~x26 & n151;
  assign n3233 = ~n3231 & ~n3232;
  assign n3234 = x27 & n154;
  assign n3235 = x26 & n156;
  assign n3236 = ~n3234 & ~n3235;
  assign n3237 = n3233 & n3236;
  assign n3223 = x13 & n1223;
  assign n3224 = x12 & n1227;
  assign n3225 = ~n3223 & ~n3224;
  assign n3226 = ~x13 & n1230;
  assign n3227 = ~x12 & n1232;
  assign n3228 = ~n3226 & ~n3227;
  assign n3229 = n3225 & n3228;
  assign n3216 = ~x11 & n1571;
  assign n3217 = ~x10 & n1575;
  assign n3218 = ~n3216 & ~n3217;
  assign n3219 = x11 & n1578;
  assign n3220 = x10 & n1580;
  assign n3221 = ~n3219 & ~n3220;
  assign n3222 = n3218 & n3221;
  assign n3230 = n3229 ^ n3222;
  assign n3238 = n3237 ^ n3230;
  assign n3262 = n3261 ^ n3238;
  assign n3213 = n2933 ^ n2927;
  assign n3214 = ~n2934 & n3213;
  assign n3215 = n3214 ^ n2927;
  assign n3263 = n3262 ^ n3215;
  assign n3209 = n2919 ^ n2903;
  assign n3210 = n2906 ^ n2903;
  assign n3211 = ~n3209 & ~n3210;
  assign n3212 = n3211 ^ n2919;
  assign n3264 = n3263 ^ n3212;
  assign n3206 = n2987 ^ n2935;
  assign n3207 = ~n2936 & n3206;
  assign n3208 = n3207 ^ n2987;
  assign n3265 = n3264 ^ n3208;
  assign n3196 = x61 ^ x0;
  assign n3197 = ~n3034 & n3196;
  assign n3198 = n3197 ^ x0;
  assign n3199 = x63 & ~n3198;
  assign n3190 = ~x30 & n66;
  assign n3191 = n69 ^ x31;
  assign n3192 = n3191 ^ n69;
  assign n3193 = n70 & n3192;
  assign n3194 = n3193 ^ n69;
  assign n3195 = ~n3190 & ~n3194;
  assign n3200 = n3199 ^ n3195;
  assign n3187 = n3033 ^ n3027;
  assign n3188 = ~n3036 & ~n3187;
  assign n3189 = n3188 ^ n3035;
  assign n3201 = n3200 ^ n3189;
  assign n3184 = n2984 ^ n2969;
  assign n3185 = n2977 & ~n3184;
  assign n3186 = n3185 ^ n2976;
  assign n3202 = n3201 ^ n3186;
  assign n3178 = n2961 ^ n2946;
  assign n3179 = n2954 & ~n3178;
  assign n3180 = n3179 ^ n2953;
  assign n3175 = n3060 ^ n3045;
  assign n3176 = n3053 & ~n3175;
  assign n3177 = n3176 ^ n3052;
  assign n3181 = n3180 ^ n3177;
  assign n3172 = n3019 ^ n3004;
  assign n3173 = n3012 & ~n3172;
  assign n3174 = n3173 ^ n3011;
  assign n3182 = n3181 ^ n3174;
  assign n3169 = n2910 ^ n2909;
  assign n3170 = ~n2918 & n3169;
  assign n3171 = n3170 ^ n2917;
  assign n3183 = n3182 ^ n3171;
  assign n3203 = n3202 ^ n3183;
  assign n3159 = ~x23 & n346;
  assign n3160 = ~x22 & n350;
  assign n3161 = ~n3159 & ~n3160;
  assign n3162 = x23 & n353;
  assign n3163 = x22 & n355;
  assign n3164 = ~n3162 & ~n3163;
  assign n3165 = n3161 & n3164;
  assign n3151 = ~x15 & n1004;
  assign n3152 = ~x14 & n1008;
  assign n3153 = ~n3151 & ~n3152;
  assign n3154 = x15 & n1011;
  assign n3155 = x14 & n1013;
  assign n3156 = ~n3154 & ~n3155;
  assign n3157 = n3153 & n3156;
  assign n3144 = x17 & n814;
  assign n3145 = x16 & n818;
  assign n3146 = ~n3144 & ~n3145;
  assign n3147 = ~x17 & n821;
  assign n3148 = ~x16 & n823;
  assign n3149 = ~n3147 & ~n3148;
  assign n3150 = n3146 & n3149;
  assign n3158 = n3157 ^ n3150;
  assign n3166 = n3165 ^ n3158;
  assign n3129 = x63 & n3034;
  assign n3130 = ~x1 & n3129;
  assign n3131 = x63 ^ x62;
  assign n3132 = ~n3034 & n3131;
  assign n3133 = x63 & n3132;
  assign n3134 = ~x0 & n3133;
  assign n3135 = ~n3130 & ~n3134;
  assign n3136 = ~x63 & n3034;
  assign n3137 = x1 & n3136;
  assign n3138 = ~x63 & n3132;
  assign n3139 = x0 & n3138;
  assign n3140 = ~n3137 & ~n3139;
  assign n3141 = n3135 & n3140;
  assign n3121 = ~x29 & n100;
  assign n3122 = ~x28 & n104;
  assign n3123 = ~n3121 & ~n3122;
  assign n3124 = x29 & n107;
  assign n3125 = x28 & n109;
  assign n3126 = ~n3124 & ~n3125;
  assign n3127 = n3123 & n3126;
  assign n3114 = ~x25 & n247;
  assign n3115 = ~x24 & n251;
  assign n3116 = ~n3114 & ~n3115;
  assign n3117 = x25 & n254;
  assign n3118 = x24 & n256;
  assign n3119 = ~n3117 & ~n3118;
  assign n3120 = n3116 & n3119;
  assign n3128 = n3127 ^ n3120;
  assign n3142 = n3141 ^ n3128;
  assign n3106 = ~x3 & n2799;
  assign n3107 = ~x2 & n2803;
  assign n3108 = ~n3106 & ~n3107;
  assign n3109 = x3 & n2806;
  assign n3110 = x2 & n2808;
  assign n3111 = ~n3109 & ~n3110;
  assign n3112 = n3108 & n3111;
  assign n3098 = ~x5 & n2386;
  assign n3099 = ~x4 & n2388;
  assign n3100 = ~n3098 & ~n3099;
  assign n3101 = x5 & n2379;
  assign n3102 = x4 & n2383;
  assign n3103 = ~n3101 & ~n3102;
  assign n3104 = n3100 & n3103;
  assign n3091 = x19 & n657;
  assign n3092 = x18 & n659;
  assign n3093 = ~n3091 & ~n3092;
  assign n3094 = ~x19 & n650;
  assign n3095 = ~x18 & n654;
  assign n3096 = ~n3094 & ~n3095;
  assign n3097 = n3093 & n3096;
  assign n3105 = n3104 ^ n3097;
  assign n3113 = n3112 ^ n3105;
  assign n3143 = n3142 ^ n3113;
  assign n3167 = n3166 ^ n3143;
  assign n3086 = n3061 ^ n3037;
  assign n3087 = n3061 ^ n3020;
  assign n3088 = ~n3086 & ~n3087;
  assign n3089 = n3088 ^ n3037;
  assign n3083 = n2962 ^ n2939;
  assign n3084 = n2986 & ~n3083;
  assign n3085 = n3084 ^ n2985;
  assign n3090 = n3089 ^ n3085;
  assign n3168 = n3167 ^ n3090;
  assign n3204 = n3203 ^ n3168;
  assign n3080 = n2997 ^ n2994;
  assign n3081 = ~n3063 & ~n3080;
  assign n3082 = n3081 ^ n3062;
  assign n3205 = n3204 ^ n3082;
  assign n3266 = n3265 ^ n3205;
  assign n3077 = n2921 ^ n2900;
  assign n3078 = ~n2989 & n3077;
  assign n3079 = n3078 ^ n2988;
  assign n3267 = n3266 ^ n3079;
  assign n3073 = n3064 ^ n2896;
  assign n3074 = n2990 ^ n2896;
  assign n3075 = n3073 & ~n3074;
  assign n3076 = n3075 ^ n3064;
  assign n3268 = n3267 ^ n3076;
  assign n3273 = n3272 ^ n3268;
  assign n3457 = n3076 & ~n3267;
  assign n3458 = ~n3076 & n3267;
  assign n3459 = ~n3272 & ~n3458;
  assign n3460 = ~n3457 & ~n3459;
  assign n3448 = x0 & x63;
  assign n3446 = x31 & n66;
  assign n3447 = n3446 ^ x33;
  assign n3449 = n3448 ^ n3447;
  assign n3439 = ~x30 & n100;
  assign n3440 = ~x29 & n104;
  assign n3441 = ~n3439 & ~n3440;
  assign n3442 = x30 & n107;
  assign n3443 = x29 & n109;
  assign n3444 = ~n3442 & ~n3443;
  assign n3445 = n3441 & n3444;
  assign n3450 = n3449 ^ n3445;
  assign n3435 = n3260 ^ n3252;
  assign n3436 = ~n3253 & n3435;
  assign n3437 = n3436 ^ n3260;
  assign n3432 = n3112 ^ n3104;
  assign n3433 = ~n3105 & n3432;
  assign n3434 = n3433 ^ n3112;
  assign n3438 = n3437 ^ n3434;
  assign n3451 = n3450 ^ n3438;
  assign n3428 = n3166 ^ n3142;
  assign n3429 = ~n3143 & n3428;
  assign n3430 = n3429 ^ n3166;
  assign n3425 = n3189 ^ n3186;
  assign n3426 = ~n3201 & n3425;
  assign n3427 = n3426 ^ n3200;
  assign n3431 = n3430 ^ n3427;
  assign n3452 = n3451 ^ n3431;
  assign n3414 = x20 & n657;
  assign n3415 = x19 & n659;
  assign n3416 = ~n3414 & ~n3415;
  assign n3417 = ~x20 & n650;
  assign n3418 = ~x19 & n654;
  assign n3419 = ~n3417 & ~n3418;
  assign n3420 = n3416 & n3419;
  assign n3406 = ~x10 & n1835;
  assign n3407 = ~x9 & n1839;
  assign n3408 = ~n3406 & ~n3407;
  assign n3409 = x10 & n1842;
  assign n3410 = x9 & n1844;
  assign n3411 = ~n3409 & ~n3410;
  assign n3412 = n3408 & n3411;
  assign n3399 = x8 & n2168;
  assign n3400 = x7 & n2170;
  assign n3401 = ~n3399 & ~n3400;
  assign n3402 = ~x8 & n2161;
  assign n3403 = ~x7 & n2165;
  assign n3404 = ~n3402 & ~n3403;
  assign n3405 = n3401 & n3404;
  assign n3413 = n3412 ^ n3405;
  assign n3421 = n3420 ^ n3413;
  assign n3390 = ~x14 & n1230;
  assign n3391 = ~x13 & n1232;
  assign n3392 = ~n3390 & ~n3391;
  assign n3393 = x14 & n1223;
  assign n3394 = x13 & n1227;
  assign n3395 = ~n3393 & ~n3394;
  assign n3396 = n3392 & n3395;
  assign n3382 = ~x24 & n346;
  assign n3383 = ~x23 & n350;
  assign n3384 = ~n3382 & ~n3383;
  assign n3385 = x24 & n353;
  assign n3386 = x23 & n355;
  assign n3387 = ~n3385 & ~n3386;
  assign n3388 = n3384 & n3387;
  assign n3375 = ~x16 & n1004;
  assign n3376 = ~x15 & n1008;
  assign n3377 = ~n3375 & ~n3376;
  assign n3378 = x16 & n1011;
  assign n3379 = x15 & n1013;
  assign n3380 = ~n3378 & ~n3379;
  assign n3381 = n3377 & n3380;
  assign n3389 = n3388 ^ n3381;
  assign n3397 = n3396 ^ n3389;
  assign n3367 = x22 & n503;
  assign n3368 = x21 & n507;
  assign n3369 = ~n3367 & ~n3368;
  assign n3370 = ~x22 & n510;
  assign n3371 = ~x21 & n512;
  assign n3372 = ~n3370 & ~n3371;
  assign n3373 = n3369 & n3372;
  assign n3359 = x28 & n154;
  assign n3360 = x27 & n156;
  assign n3361 = ~n3359 & ~n3360;
  assign n3362 = ~x28 & n147;
  assign n3363 = ~x27 & n151;
  assign n3364 = ~n3362 & ~n3363;
  assign n3365 = n3361 & n3364;
  assign n3352 = x12 & n1578;
  assign n3353 = x11 & n1580;
  assign n3354 = ~n3352 & ~n3353;
  assign n3355 = ~x12 & n1571;
  assign n3356 = ~x11 & n1575;
  assign n3357 = ~n3355 & ~n3356;
  assign n3358 = n3354 & n3357;
  assign n3366 = n3365 ^ n3358;
  assign n3374 = n3373 ^ n3366;
  assign n3398 = n3397 ^ n3374;
  assign n3422 = n3421 ^ n3398;
  assign n3347 = n3165 ^ n3157;
  assign n3348 = ~n3158 & n3347;
  assign n3349 = n3348 ^ n3165;
  assign n3344 = n3141 ^ n3120;
  assign n3345 = n3128 & ~n3344;
  assign n3346 = n3345 ^ n3127;
  assign n3350 = n3349 ^ n3346;
  assign n3340 = n3237 ^ n3229;
  assign n3341 = n3237 ^ n3222;
  assign n3342 = n3340 & ~n3341;
  assign n3343 = n3342 ^ n3229;
  assign n3351 = n3350 ^ n3343;
  assign n3423 = n3422 ^ n3351;
  assign n3337 = n3238 ^ n3215;
  assign n3338 = n3262 & ~n3337;
  assign n3339 = n3338 ^ n3261;
  assign n3424 = n3423 ^ n3339;
  assign n3453 = n3452 ^ n3424;
  assign n3331 = ~n3195 & n3199;
  assign n3323 = ~x6 & n2386;
  assign n3324 = ~x5 & n2388;
  assign n3325 = ~n3323 & ~n3324;
  assign n3326 = x6 & n2379;
  assign n3327 = x5 & n2383;
  assign n3328 = ~n3326 & ~n3327;
  assign n3329 = n3325 & n3328;
  assign n3316 = ~x4 & n2799;
  assign n3317 = ~x3 & n2803;
  assign n3318 = ~n3316 & ~n3317;
  assign n3319 = x4 & n2806;
  assign n3320 = x3 & n2808;
  assign n3321 = ~n3319 & ~n3320;
  assign n3322 = n3318 & n3321;
  assign n3330 = n3329 ^ n3322;
  assign n3332 = n3331 ^ n3330;
  assign n3308 = x18 & n814;
  assign n3309 = x17 & n818;
  assign n3310 = ~n3308 & ~n3309;
  assign n3311 = ~x18 & n821;
  assign n3312 = ~x17 & n823;
  assign n3313 = ~n3311 & ~n3312;
  assign n3314 = n3310 & n3313;
  assign n3300 = x2 & n3136;
  assign n3301 = x1 & n3138;
  assign n3302 = ~n3300 & ~n3301;
  assign n3303 = ~x2 & n3129;
  assign n3304 = ~x1 & n3133;
  assign n3305 = ~n3303 & ~n3304;
  assign n3306 = n3302 & n3305;
  assign n3293 = ~x26 & n247;
  assign n3294 = ~x25 & n251;
  assign n3295 = ~n3293 & ~n3294;
  assign n3296 = x26 & n254;
  assign n3297 = x25 & n256;
  assign n3298 = ~n3296 & ~n3297;
  assign n3299 = n3295 & n3298;
  assign n3307 = n3306 ^ n3299;
  assign n3315 = n3314 ^ n3307;
  assign n3333 = n3332 ^ n3315;
  assign n3290 = n3177 ^ n3174;
  assign n3291 = n3181 & ~n3290;
  assign n3292 = n3291 ^ n3180;
  assign n3334 = n3333 ^ n3292;
  assign n3287 = n3202 ^ n3182;
  assign n3288 = ~n3183 & ~n3287;
  assign n3289 = n3288 ^ n3202;
  assign n3335 = n3334 ^ n3289;
  assign n3284 = n3167 ^ n3089;
  assign n3285 = n3090 & ~n3284;
  assign n3286 = n3285 ^ n3167;
  assign n3336 = n3335 ^ n3286;
  assign n3454 = n3453 ^ n3336;
  assign n3280 = n3212 ^ n3208;
  assign n3281 = ~n3264 & n3280;
  assign n3282 = n3281 ^ n3263;
  assign n3277 = n3168 ^ n3082;
  assign n3278 = n3204 & ~n3277;
  assign n3279 = n3278 ^ n3203;
  assign n3283 = n3282 ^ n3279;
  assign n3455 = n3454 ^ n3283;
  assign n3274 = n3205 ^ n3079;
  assign n3275 = n3266 & n3274;
  assign n3276 = n3275 ^ n3265;
  assign n3456 = n3455 ^ n3276;
  assign n3461 = n3460 ^ n3456;
  assign n3648 = n3276 & n3455;
  assign n3649 = ~n3276 & ~n3455;
  assign n3650 = ~n3460 & ~n3649;
  assign n3651 = ~n3648 & ~n3650;
  assign n3633 = ~x5 & n2799;
  assign n3634 = ~x4 & n2803;
  assign n3635 = ~n3633 & ~n3634;
  assign n3636 = x5 & n2806;
  assign n3637 = x4 & n2808;
  assign n3638 = ~n3636 & ~n3637;
  assign n3639 = n3635 & n3638;
  assign n3640 = n3639 ^ x33;
  assign n3630 = n3447 ^ n3445;
  assign n3631 = n3449 & n3630;
  assign n3632 = n3631 ^ n3448;
  assign n3641 = n3640 ^ n3632;
  assign n3624 = n3314 ^ n3306;
  assign n3625 = n3314 ^ n3299;
  assign n3626 = n3624 & ~n3625;
  assign n3627 = n3626 ^ n3306;
  assign n3621 = n3396 ^ n3381;
  assign n3622 = n3389 & ~n3621;
  assign n3623 = n3622 ^ n3388;
  assign n3628 = n3627 ^ n3623;
  assign n3617 = n3420 ^ n3412;
  assign n3618 = n3420 ^ n3405;
  assign n3619 = n3617 & ~n3618;
  assign n3620 = n3619 ^ n3412;
  assign n3629 = n3628 ^ n3620;
  assign n3642 = n3641 ^ n3629;
  assign n3614 = n3421 ^ n3374;
  assign n3615 = n3398 & ~n3614;
  assign n3616 = n3615 ^ n3397;
  assign n3643 = n3642 ^ n3616;
  assign n3608 = n3331 ^ n3322;
  assign n3609 = n3330 & n3608;
  assign n3610 = n3609 ^ n3329;
  assign n3605 = n3346 ^ n3343;
  assign n3606 = n3350 & ~n3605;
  assign n3607 = n3606 ^ n3349;
  assign n3611 = n3610 ^ n3607;
  assign n3602 = n3450 ^ n3437;
  assign n3603 = ~n3438 & n3602;
  assign n3604 = n3603 ^ n3450;
  assign n3612 = n3611 ^ n3604;
  assign n3598 = n3451 ^ n3430;
  assign n3599 = n3451 ^ n3427;
  assign n3600 = n3598 & ~n3599;
  assign n3601 = n3600 ^ n3430;
  assign n3613 = n3612 ^ n3601;
  assign n3644 = n3643 ^ n3613;
  assign n3585 = ~x13 & n1571;
  assign n3586 = ~x12 & n1575;
  assign n3587 = ~n3585 & ~n3586;
  assign n3588 = x13 & n1578;
  assign n3589 = x12 & n1580;
  assign n3590 = ~n3588 & ~n3589;
  assign n3591 = n3587 & n3590;
  assign n3577 = x15 & n1223;
  assign n3578 = x14 & n1227;
  assign n3579 = ~n3577 & ~n3578;
  assign n3580 = ~x15 & n1230;
  assign n3581 = ~x14 & n1232;
  assign n3582 = ~n3580 & ~n3581;
  assign n3583 = n3579 & n3582;
  assign n3570 = ~x25 & n346;
  assign n3571 = ~x24 & n350;
  assign n3572 = ~n3570 & ~n3571;
  assign n3573 = x25 & n353;
  assign n3574 = x24 & n355;
  assign n3575 = ~n3573 & ~n3574;
  assign n3576 = n3572 & n3575;
  assign n3584 = n3583 ^ n3576;
  assign n3592 = n3591 ^ n3584;
  assign n3561 = ~x11 & n1835;
  assign n3562 = ~x10 & n1839;
  assign n3563 = ~n3561 & ~n3562;
  assign n3564 = x11 & n1842;
  assign n3565 = x10 & n1844;
  assign n3566 = ~n3564 & ~n3565;
  assign n3567 = n3563 & n3566;
  assign n3553 = ~x29 & n147;
  assign n3554 = ~x28 & n151;
  assign n3555 = ~n3553 & ~n3554;
  assign n3556 = x29 & n154;
  assign n3557 = x28 & n156;
  assign n3558 = ~n3556 & ~n3557;
  assign n3559 = n3555 & n3558;
  assign n3546 = x23 & n503;
  assign n3547 = x22 & n507;
  assign n3548 = ~n3546 & ~n3547;
  assign n3549 = ~x23 & n510;
  assign n3550 = ~x22 & n512;
  assign n3551 = ~n3549 & ~n3550;
  assign n3552 = n3548 & n3551;
  assign n3560 = n3559 ^ n3552;
  assign n3568 = n3567 ^ n3560;
  assign n3538 = x27 & n254;
  assign n3539 = x26 & n256;
  assign n3540 = ~n3538 & ~n3539;
  assign n3541 = ~x27 & n247;
  assign n3542 = ~x26 & n251;
  assign n3543 = ~n3541 & ~n3542;
  assign n3544 = n3540 & n3543;
  assign n3530 = ~x31 & n100;
  assign n3531 = ~x30 & n104;
  assign n3532 = ~n3530 & ~n3531;
  assign n3533 = x31 & n107;
  assign n3534 = x30 & n109;
  assign n3535 = ~n3533 & ~n3534;
  assign n3536 = n3532 & n3535;
  assign n3523 = ~x17 & n1004;
  assign n3524 = ~x16 & n1008;
  assign n3525 = ~n3523 & ~n3524;
  assign n3526 = x17 & n1011;
  assign n3527 = x16 & n1013;
  assign n3528 = ~n3526 & ~n3527;
  assign n3529 = n3525 & n3528;
  assign n3537 = n3536 ^ n3529;
  assign n3545 = n3544 ^ n3537;
  assign n3569 = n3568 ^ n3545;
  assign n3593 = n3592 ^ n3569;
  assign n3514 = x7 & n2379;
  assign n3515 = x6 & n2383;
  assign n3516 = ~n3514 & ~n3515;
  assign n3517 = ~x7 & n2386;
  assign n3518 = ~x6 & n2388;
  assign n3519 = ~n3517 & ~n3518;
  assign n3520 = n3516 & n3519;
  assign n3506 = ~x21 & n650;
  assign n3507 = ~x20 & n654;
  assign n3508 = ~n3506 & ~n3507;
  assign n3509 = x21 & n657;
  assign n3510 = x20 & n659;
  assign n3511 = ~n3509 & ~n3510;
  assign n3512 = n3508 & n3511;
  assign n3499 = ~x9 & n2161;
  assign n3500 = ~x8 & n2165;
  assign n3501 = ~n3499 & ~n3500;
  assign n3502 = x9 & n2168;
  assign n3503 = x8 & n2170;
  assign n3504 = ~n3502 & ~n3503;
  assign n3505 = n3501 & n3504;
  assign n3513 = n3512 ^ n3505;
  assign n3521 = n3520 ^ n3513;
  assign n3496 = x1 & x63;
  assign n3488 = ~x19 & n821;
  assign n3489 = ~x18 & n823;
  assign n3490 = ~n3488 & ~n3489;
  assign n3491 = x19 & n814;
  assign n3492 = x18 & n818;
  assign n3493 = ~n3491 & ~n3492;
  assign n3494 = n3490 & n3493;
  assign n3481 = ~x3 & n3129;
  assign n3482 = ~x2 & n3133;
  assign n3483 = ~n3481 & ~n3482;
  assign n3484 = x3 & n3136;
  assign n3485 = x2 & n3138;
  assign n3486 = ~n3484 & ~n3485;
  assign n3487 = n3483 & n3486;
  assign n3495 = n3494 ^ n3487;
  assign n3497 = n3496 ^ n3495;
  assign n3477 = n3373 ^ n3365;
  assign n3478 = n3373 ^ n3358;
  assign n3479 = n3477 & ~n3478;
  assign n3480 = n3479 ^ n3365;
  assign n3498 = n3497 ^ n3480;
  assign n3522 = n3521 ^ n3498;
  assign n3594 = n3593 ^ n3522;
  assign n3474 = n3315 ^ n3292;
  assign n3475 = ~n3333 & ~n3474;
  assign n3476 = n3475 ^ n3332;
  assign n3595 = n3594 ^ n3476;
  assign n3471 = n3351 ^ n3339;
  assign n3472 = n3423 & ~n3471;
  assign n3473 = n3472 ^ n3422;
  assign n3596 = n3595 ^ n3473;
  assign n3468 = n3289 ^ n3286;
  assign n3469 = n3335 & n3468;
  assign n3470 = n3469 ^ n3334;
  assign n3597 = n3596 ^ n3470;
  assign n3645 = n3644 ^ n3597;
  assign n3465 = n3424 ^ n3336;
  assign n3466 = n3453 & ~n3465;
  assign n3467 = n3466 ^ n3452;
  assign n3646 = n3645 ^ n3467;
  assign n3462 = n3454 ^ n3282;
  assign n3463 = n3283 & n3462;
  assign n3464 = n3463 ^ n3454;
  assign n3647 = n3646 ^ n3464;
  assign n3652 = n3651 ^ n3647;
  assign n3835 = ~n3464 & n3646;
  assign n3836 = n3464 & ~n3646;
  assign n3837 = ~n3651 & ~n3836;
  assign n3838 = ~n3835 & ~n3837;
  assign n3824 = x35 ^ x31;
  assign n3825 = n103 & n3824;
  assign n3826 = ~n100 & ~n3825;
  assign n3827 = n3826 ^ x33;
  assign n3821 = n3496 ^ n3494;
  assign n3822 = ~n3495 & ~n3821;
  assign n3823 = n3822 ^ n3496;
  assign n3828 = n3827 ^ n3823;
  assign n3818 = n3521 ^ n3497;
  assign n3819 = n3498 & ~n3818;
  assign n3820 = n3819 ^ n3521;
  assign n3829 = n3828 ^ n3820;
  assign n3814 = n3592 ^ n3568;
  assign n3815 = n3592 ^ n3545;
  assign n3816 = n3814 & ~n3815;
  assign n3817 = n3816 ^ n3568;
  assign n3830 = n3829 ^ n3817;
  assign n3807 = n3591 ^ n3576;
  assign n3808 = n3584 & ~n3807;
  assign n3809 = n3808 ^ n3583;
  assign n3804 = n3544 ^ n3536;
  assign n3805 = ~n3537 & n3804;
  assign n3806 = n3805 ^ n3544;
  assign n3810 = n3809 ^ n3806;
  assign n3801 = n3567 ^ n3559;
  assign n3802 = ~n3560 & n3801;
  assign n3803 = n3802 ^ n3567;
  assign n3811 = n3810 ^ n3803;
  assign n3797 = n3639 ^ n3632;
  assign n3798 = ~n3640 & n3797;
  assign n3799 = n3798 ^ x33;
  assign n3794 = n3627 ^ n3620;
  assign n3795 = ~n3628 & n3794;
  assign n3796 = n3795 ^ n3620;
  assign n3800 = n3799 ^ n3796;
  assign n3812 = n3811 ^ n3800;
  assign n3790 = n3610 ^ n3604;
  assign n3791 = n3607 ^ n3604;
  assign n3792 = n3790 & ~n3791;
  assign n3793 = n3792 ^ n3610;
  assign n3813 = n3812 ^ n3793;
  assign n3831 = n3830 ^ n3813;
  assign n3777 = ~x8 & n2386;
  assign n3778 = ~x7 & n2388;
  assign n3779 = ~n3777 & ~n3778;
  assign n3780 = x8 & n2379;
  assign n3781 = x7 & n2383;
  assign n3782 = ~n3780 & ~n3781;
  assign n3783 = n3779 & n3782;
  assign n3769 = ~x22 & n650;
  assign n3770 = ~x21 & n654;
  assign n3771 = ~n3769 & ~n3770;
  assign n3772 = x22 & n657;
  assign n3773 = x21 & n659;
  assign n3774 = ~n3772 & ~n3773;
  assign n3775 = n3771 & n3774;
  assign n3762 = ~x10 & n2161;
  assign n3763 = ~x9 & n2165;
  assign n3764 = ~n3762 & ~n3763;
  assign n3765 = x10 & n2168;
  assign n3766 = x9 & n2170;
  assign n3767 = ~n3765 & ~n3766;
  assign n3768 = n3764 & n3767;
  assign n3776 = n3775 ^ n3768;
  assign n3784 = n3783 ^ n3776;
  assign n3759 = x2 & x63;
  assign n3751 = ~x26 & n346;
  assign n3752 = ~x25 & n350;
  assign n3753 = ~n3751 & ~n3752;
  assign n3754 = x26 & n353;
  assign n3755 = x25 & n355;
  assign n3756 = ~n3754 & ~n3755;
  assign n3757 = n3753 & n3756;
  assign n3744 = ~x30 & n147;
  assign n3745 = ~x29 & n151;
  assign n3746 = ~n3744 & ~n3745;
  assign n3747 = x30 & n154;
  assign n3748 = x29 & n156;
  assign n3749 = ~n3747 & ~n3748;
  assign n3750 = n3746 & n3749;
  assign n3758 = n3757 ^ n3750;
  assign n3760 = n3759 ^ n3758;
  assign n3736 = ~x28 & n247;
  assign n3737 = ~x27 & n251;
  assign n3738 = ~n3736 & ~n3737;
  assign n3739 = x28 & n254;
  assign n3740 = x27 & n256;
  assign n3741 = ~n3739 & ~n3740;
  assign n3742 = n3738 & n3741;
  assign n3728 = ~x12 & n1835;
  assign n3729 = ~x11 & n1839;
  assign n3730 = ~n3728 & ~n3729;
  assign n3731 = x12 & n1842;
  assign n3732 = x11 & n1844;
  assign n3733 = ~n3731 & ~n3732;
  assign n3734 = n3730 & n3733;
  assign n3721 = ~x14 & n1571;
  assign n3722 = ~x13 & n1575;
  assign n3723 = ~n3721 & ~n3722;
  assign n3724 = x14 & n1578;
  assign n3725 = x13 & n1580;
  assign n3726 = ~n3724 & ~n3725;
  assign n3727 = n3723 & n3726;
  assign n3735 = n3734 ^ n3727;
  assign n3743 = n3742 ^ n3735;
  assign n3761 = n3760 ^ n3743;
  assign n3785 = n3784 ^ n3761;
  assign n3712 = ~x24 & n510;
  assign n3713 = ~x23 & n512;
  assign n3714 = ~n3712 & ~n3713;
  assign n3715 = x24 & n503;
  assign n3716 = x23 & n507;
  assign n3717 = ~n3715 & ~n3716;
  assign n3718 = n3714 & n3717;
  assign n3704 = ~x18 & n1004;
  assign n3705 = ~x17 & n1008;
  assign n3706 = ~n3704 & ~n3705;
  assign n3707 = x18 & n1011;
  assign n3708 = x17 & n1013;
  assign n3709 = ~n3707 & ~n3708;
  assign n3710 = n3706 & n3709;
  assign n3697 = x16 & n1223;
  assign n3698 = x15 & n1227;
  assign n3699 = ~n3697 & ~n3698;
  assign n3700 = ~x16 & n1230;
  assign n3701 = ~x15 & n1232;
  assign n3702 = ~n3700 & ~n3701;
  assign n3703 = n3699 & n3702;
  assign n3711 = n3710 ^ n3703;
  assign n3719 = n3718 ^ n3711;
  assign n3688 = ~x4 & n3129;
  assign n3689 = ~x3 & n3133;
  assign n3690 = ~n3688 & ~n3689;
  assign n3691 = x4 & n3136;
  assign n3692 = x3 & n3138;
  assign n3693 = ~n3691 & ~n3692;
  assign n3694 = n3690 & n3693;
  assign n3680 = ~x6 & n2799;
  assign n3681 = ~x5 & n2803;
  assign n3682 = ~n3680 & ~n3681;
  assign n3683 = x6 & n2806;
  assign n3684 = x5 & n2808;
  assign n3685 = ~n3683 & ~n3684;
  assign n3686 = n3682 & n3685;
  assign n3673 = x20 & n814;
  assign n3674 = x19 & n818;
  assign n3675 = ~n3673 & ~n3674;
  assign n3676 = ~x20 & n821;
  assign n3677 = ~x19 & n823;
  assign n3678 = ~n3676 & ~n3677;
  assign n3679 = n3675 & n3678;
  assign n3687 = n3686 ^ n3679;
  assign n3695 = n3694 ^ n3687;
  assign n3669 = n3520 ^ n3512;
  assign n3670 = n3520 ^ n3505;
  assign n3671 = n3669 & ~n3670;
  assign n3672 = n3671 ^ n3512;
  assign n3696 = n3695 ^ n3672;
  assign n3720 = n3719 ^ n3696;
  assign n3786 = n3785 ^ n3720;
  assign n3665 = n3641 ^ n3616;
  assign n3666 = n3629 ^ n3616;
  assign n3667 = n3665 & ~n3666;
  assign n3668 = n3667 ^ n3641;
  assign n3787 = n3786 ^ n3668;
  assign n3662 = n3522 ^ n3476;
  assign n3663 = ~n3594 & ~n3662;
  assign n3664 = n3663 ^ n3593;
  assign n3788 = n3787 ^ n3664;
  assign n3659 = n3643 ^ n3612;
  assign n3660 = ~n3613 & n3659;
  assign n3661 = n3660 ^ n3643;
  assign n3789 = n3788 ^ n3661;
  assign n3832 = n3831 ^ n3789;
  assign n3656 = n3473 ^ n3470;
  assign n3657 = n3596 & n3656;
  assign n3658 = n3657 ^ n3595;
  assign n3833 = n3832 ^ n3658;
  assign n3653 = n3597 ^ n3467;
  assign n3654 = ~n3645 & n3653;
  assign n3655 = n3654 ^ n3644;
  assign n3834 = n3833 ^ n3655;
  assign n3839 = n3838 ^ n3834;
  assign n4020 = ~n3655 & ~n3833;
  assign n4021 = n3655 & n3833;
  assign n4022 = ~n3838 & ~n4021;
  assign n4023 = ~n4020 & ~n4022;
  assign n4009 = n3742 ^ n3734;
  assign n4010 = ~n3735 & n4009;
  assign n4011 = n4010 ^ n3742;
  assign n4006 = n3718 ^ n3703;
  assign n4007 = n3711 & ~n4006;
  assign n4008 = n4007 ^ n3710;
  assign n4012 = n4011 ^ n4008;
  assign n4003 = n3783 ^ n3768;
  assign n4004 = n3776 & ~n4003;
  assign n4005 = n4004 ^ n3775;
  assign n4013 = n4012 ^ n4005;
  assign n3999 = n3784 ^ n3760;
  assign n4000 = n3784 ^ n3743;
  assign n4001 = ~n3999 & ~n4000;
  assign n4002 = n4001 ^ n3760;
  assign n4014 = n4013 ^ n4002;
  assign n3995 = n3719 ^ n3695;
  assign n3996 = n3719 ^ n3672;
  assign n3997 = n3995 & ~n3996;
  assign n3998 = n3997 ^ n3695;
  assign n4015 = n4014 ^ n3998;
  assign n3990 = n3828 ^ n3817;
  assign n3991 = n3820 ^ n3817;
  assign n3992 = n3990 & ~n3991;
  assign n3993 = n3992 ^ n3828;
  assign n3987 = n3811 ^ n3799;
  assign n3988 = n3800 & ~n3987;
  assign n3989 = n3988 ^ n3811;
  assign n3994 = n3993 ^ n3989;
  assign n4016 = n4015 ^ n3994;
  assign n3974 = x11 & n2168;
  assign n3975 = x10 & n2170;
  assign n3976 = ~n3974 & ~n3975;
  assign n3977 = ~x11 & n2161;
  assign n3978 = ~x10 & n2165;
  assign n3979 = ~n3977 & ~n3978;
  assign n3980 = n3976 & n3979;
  assign n3966 = ~x29 & n247;
  assign n3967 = ~x28 & n251;
  assign n3968 = ~n3966 & ~n3967;
  assign n3969 = x29 & n254;
  assign n3970 = x28 & n256;
  assign n3971 = ~n3969 & ~n3970;
  assign n3972 = n3968 & n3971;
  assign n3959 = x23 & n657;
  assign n3960 = x22 & n659;
  assign n3961 = ~n3959 & ~n3960;
  assign n3962 = ~x23 & n650;
  assign n3963 = ~x22 & n654;
  assign n3964 = ~n3962 & ~n3963;
  assign n3965 = n3961 & n3964;
  assign n3973 = n3972 ^ n3965;
  assign n3981 = n3980 ^ n3973;
  assign n3950 = ~x7 & n2799;
  assign n3951 = ~x6 & n2803;
  assign n3952 = ~n3950 & ~n3951;
  assign n3953 = x7 & n2806;
  assign n3954 = x6 & n2808;
  assign n3955 = ~n3953 & ~n3954;
  assign n3956 = n3952 & n3955;
  assign n3942 = ~x21 & n821;
  assign n3943 = ~x20 & n823;
  assign n3944 = ~n3942 & ~n3943;
  assign n3945 = x21 & n814;
  assign n3946 = x20 & n818;
  assign n3947 = ~n3945 & ~n3946;
  assign n3948 = n3944 & n3947;
  assign n3935 = x9 & n2379;
  assign n3936 = x8 & n2383;
  assign n3937 = ~n3935 & ~n3936;
  assign n3938 = ~x9 & n2386;
  assign n3939 = ~x8 & n2388;
  assign n3940 = ~n3938 & ~n3939;
  assign n3941 = n3937 & n3940;
  assign n3949 = n3948 ^ n3941;
  assign n3957 = n3956 ^ n3949;
  assign n3927 = ~x13 & n1835;
  assign n3928 = ~x12 & n1839;
  assign n3929 = ~n3927 & ~n3928;
  assign n3930 = x13 & n1842;
  assign n3931 = x12 & n1844;
  assign n3932 = ~n3930 & ~n3931;
  assign n3933 = n3929 & n3932;
  assign n3919 = ~x25 & n510;
  assign n3920 = ~x24 & n512;
  assign n3921 = ~n3919 & ~n3920;
  assign n3922 = x25 & n503;
  assign n3923 = x24 & n507;
  assign n3924 = ~n3922 & ~n3923;
  assign n3925 = n3921 & n3924;
  assign n3912 = ~x15 & n1571;
  assign n3913 = ~x14 & n1575;
  assign n3914 = ~n3912 & ~n3913;
  assign n3915 = x15 & n1578;
  assign n3916 = x14 & n1580;
  assign n3917 = ~n3915 & ~n3916;
  assign n3918 = n3914 & n3917;
  assign n3926 = n3925 ^ n3918;
  assign n3934 = n3933 ^ n3926;
  assign n3958 = n3957 ^ n3934;
  assign n3982 = n3981 ^ n3958;
  assign n3903 = x27 & n353;
  assign n3904 = x26 & n355;
  assign n3905 = ~n3903 & ~n3904;
  assign n3906 = ~x27 & n346;
  assign n3907 = ~x26 & n350;
  assign n3908 = ~n3906 & ~n3907;
  assign n3909 = n3905 & n3908;
  assign n3901 = ~n100 & ~n104;
  assign n3894 = x31 & n154;
  assign n3895 = x30 & n156;
  assign n3896 = ~n3894 & ~n3895;
  assign n3897 = ~x31 & n147;
  assign n3898 = ~x30 & n151;
  assign n3899 = ~n3897 & ~n3898;
  assign n3900 = n3896 & n3899;
  assign n3902 = n3901 ^ n3900;
  assign n3910 = n3909 ^ n3902;
  assign n3885 = ~x17 & n1230;
  assign n3886 = ~x16 & n1232;
  assign n3887 = ~n3885 & ~n3886;
  assign n3888 = x17 & n1223;
  assign n3889 = x16 & n1227;
  assign n3890 = ~n3888 & ~n3889;
  assign n3891 = n3887 & n3890;
  assign n3883 = x3 & x63;
  assign n3876 = ~x19 & n1004;
  assign n3877 = ~x18 & n1008;
  assign n3878 = ~n3876 & ~n3877;
  assign n3879 = x19 & n1011;
  assign n3880 = x18 & n1013;
  assign n3881 = ~n3879 & ~n3880;
  assign n3882 = n3878 & n3881;
  assign n3884 = n3883 ^ n3882;
  assign n3892 = n3891 ^ n3884;
  assign n3873 = n3694 ^ n3686;
  assign n3874 = ~n3687 & n3873;
  assign n3875 = n3874 ^ n3694;
  assign n3893 = n3892 ^ n3875;
  assign n3911 = n3910 ^ n3893;
  assign n3983 = n3982 ^ n3911;
  assign n3862 = x5 & n3136;
  assign n3863 = x4 & n3138;
  assign n3864 = ~n3862 & ~n3863;
  assign n3865 = ~x5 & n3129;
  assign n3866 = ~x4 & n3133;
  assign n3867 = ~n3865 & ~n3866;
  assign n3868 = n3864 & n3867;
  assign n3869 = n3868 ^ n3826;
  assign n3859 = n3759 ^ n3757;
  assign n3860 = ~n3758 & ~n3859;
  assign n3861 = n3860 ^ n3759;
  assign n3870 = n3869 ^ n3861;
  assign n3856 = n3806 ^ n3803;
  assign n3857 = n3810 & ~n3856;
  assign n3858 = n3857 ^ n3809;
  assign n3871 = n3870 ^ n3858;
  assign n3853 = n3826 ^ n3823;
  assign n3854 = ~n3827 & ~n3853;
  assign n3855 = n3854 ^ x33;
  assign n3872 = n3871 ^ n3855;
  assign n3984 = n3983 ^ n3872;
  assign n3850 = n3720 ^ n3668;
  assign n3851 = ~n3786 & ~n3850;
  assign n3852 = n3851 ^ n3785;
  assign n3985 = n3984 ^ n3852;
  assign n3847 = n3830 ^ n3812;
  assign n3848 = n3813 & ~n3847;
  assign n3849 = n3848 ^ n3830;
  assign n3986 = n3985 ^ n3849;
  assign n4017 = n4016 ^ n3986;
  assign n3843 = n3787 ^ n3661;
  assign n3844 = n3664 ^ n3661;
  assign n3845 = ~n3843 & ~n3844;
  assign n3846 = n3845 ^ n3787;
  assign n4018 = n4017 ^ n3846;
  assign n3840 = n3789 ^ n3658;
  assign n3841 = n3832 & n3840;
  assign n3842 = n3841 ^ n3831;
  assign n4019 = n4018 ^ n3842;
  assign n4024 = n4023 ^ n4019;
  assign n4201 = n3842 & ~n4018;
  assign n4202 = ~n3842 & n4018;
  assign n4203 = ~n4023 & ~n4202;
  assign n4204 = ~n4201 & ~n4203;
  assign n4187 = x18 & n1223;
  assign n4188 = x17 & n1227;
  assign n4189 = ~n4187 & ~n4188;
  assign n4190 = ~x18 & n1230;
  assign n4191 = ~x17 & n1232;
  assign n4192 = ~n4190 & ~n4191;
  assign n4193 = n4189 & n4192;
  assign n4179 = ~x26 & n510;
  assign n4180 = ~x25 & n512;
  assign n4181 = ~n4179 & ~n4180;
  assign n4182 = x26 & n503;
  assign n4183 = x25 & n507;
  assign n4184 = ~n4182 & ~n4183;
  assign n4185 = n4181 & n4184;
  assign n4172 = ~x30 & n247;
  assign n4173 = ~x29 & n251;
  assign n4174 = ~n4172 & ~n4173;
  assign n4175 = x30 & n254;
  assign n4176 = x29 & n256;
  assign n4177 = ~n4175 & ~n4176;
  assign n4178 = n4174 & n4177;
  assign n4186 = n4185 ^ n4178;
  assign n4194 = n4193 ^ n4186;
  assign n4168 = n3980 ^ n3965;
  assign n4169 = n3973 & ~n4168;
  assign n4170 = n4169 ^ n3972;
  assign n4164 = n3956 ^ n3948;
  assign n4165 = n3956 ^ n3941;
  assign n4166 = n4164 & ~n4165;
  assign n4167 = n4166 ^ n3948;
  assign n4171 = n4170 ^ n4167;
  assign n4195 = n4194 ^ n4171;
  assign n4157 = n3909 ^ n3901;
  assign n4158 = n3909 ^ n3900;
  assign n4159 = ~n4157 & ~n4158;
  assign n4160 = n4159 ^ n3901;
  assign n4153 = n3891 ^ n3883;
  assign n4154 = n3891 ^ n3882;
  assign n4155 = ~n4153 & ~n4154;
  assign n4156 = n4155 ^ n3883;
  assign n4161 = n4160 ^ n4156;
  assign n4149 = n3933 ^ n3925;
  assign n4150 = n3933 ^ n3918;
  assign n4151 = n4149 & ~n4150;
  assign n4152 = n4151 ^ n3925;
  assign n4162 = n4161 ^ n4152;
  assign n4145 = n3910 ^ n3892;
  assign n4146 = n3910 ^ n3875;
  assign n4147 = n4145 & n4146;
  assign n4148 = n4147 ^ n3892;
  assign n4163 = n4162 ^ n4148;
  assign n4196 = n4195 ^ n4163;
  assign n4138 = x37 ^ x31;
  assign n4139 = n150 & n4138;
  assign n4140 = ~n147 & ~n4139;
  assign n4136 = x4 & x63;
  assign n4129 = x6 & n3136;
  assign n4130 = x5 & n3138;
  assign n4131 = ~n4129 & ~n4130;
  assign n4132 = ~x6 & n3129;
  assign n4133 = ~x5 & n3133;
  assign n4134 = ~n4132 & ~n4133;
  assign n4135 = n4131 & n4134;
  assign n4137 = n4136 ^ n4135;
  assign n4141 = n4140 ^ n4137;
  assign n4125 = n4011 ^ n4005;
  assign n4126 = n4008 ^ n4005;
  assign n4127 = n4125 & ~n4126;
  assign n4128 = n4127 ^ n4011;
  assign n4142 = n4141 ^ n4128;
  assign n4122 = n3868 ^ n3861;
  assign n4123 = n3869 & n4122;
  assign n4124 = n4123 ^ n3826;
  assign n4143 = n4142 ^ n4124;
  assign n4119 = n4002 ^ n3998;
  assign n4120 = ~n4014 & n4119;
  assign n4121 = n4120 ^ n4013;
  assign n4144 = n4143 ^ n4121;
  assign n4197 = n4196 ^ n4144;
  assign n4106 = x22 & n814;
  assign n4107 = x21 & n818;
  assign n4108 = ~n4106 & ~n4107;
  assign n4109 = ~x22 & n821;
  assign n4110 = ~x21 & n823;
  assign n4111 = ~n4109 & ~n4110;
  assign n4112 = n4108 & n4111;
  assign n4098 = ~x28 & n346;
  assign n4099 = ~x27 & n350;
  assign n4100 = ~n4098 & ~n4099;
  assign n4101 = x28 & n353;
  assign n4102 = x27 & n355;
  assign n4103 = ~n4101 & ~n4102;
  assign n4104 = n4100 & n4103;
  assign n4091 = ~x12 & n2161;
  assign n4092 = ~x11 & n2165;
  assign n4093 = ~n4091 & ~n4092;
  assign n4094 = x12 & n2168;
  assign n4095 = x11 & n2170;
  assign n4096 = ~n4094 & ~n4095;
  assign n4097 = n4093 & n4096;
  assign n4105 = n4104 ^ n4097;
  assign n4113 = n4112 ^ n4105;
  assign n4082 = ~x20 & n1004;
  assign n4083 = ~x19 & n1008;
  assign n4084 = ~n4082 & ~n4083;
  assign n4085 = x20 & n1011;
  assign n4086 = x19 & n1013;
  assign n4087 = ~n4085 & ~n4086;
  assign n4088 = n4084 & n4087;
  assign n4074 = x10 & n2379;
  assign n4075 = x9 & n2383;
  assign n4076 = ~n4074 & ~n4075;
  assign n4077 = ~x10 & n2386;
  assign n4078 = ~x9 & n2388;
  assign n4079 = ~n4077 & ~n4078;
  assign n4080 = n4076 & n4079;
  assign n4067 = x8 & n2806;
  assign n4068 = x7 & n2808;
  assign n4069 = ~n4067 & ~n4068;
  assign n4070 = ~x8 & n2799;
  assign n4071 = ~x7 & n2803;
  assign n4072 = ~n4070 & ~n4071;
  assign n4073 = n4069 & n4072;
  assign n4081 = n4080 ^ n4073;
  assign n4089 = n4088 ^ n4081;
  assign n4059 = x14 & n1842;
  assign n4060 = x13 & n1844;
  assign n4061 = ~n4059 & ~n4060;
  assign n4062 = ~x14 & n1835;
  assign n4063 = ~x13 & n1839;
  assign n4064 = ~n4062 & ~n4063;
  assign n4065 = n4061 & n4064;
  assign n4051 = ~x16 & n1571;
  assign n4052 = ~x15 & n1575;
  assign n4053 = ~n4051 & ~n4052;
  assign n4054 = x16 & n1578;
  assign n4055 = x15 & n1580;
  assign n4056 = ~n4054 & ~n4055;
  assign n4057 = n4053 & n4056;
  assign n4044 = ~x24 & n650;
  assign n4045 = ~x23 & n654;
  assign n4046 = ~n4044 & ~n4045;
  assign n4047 = x24 & n657;
  assign n4048 = x23 & n659;
  assign n4049 = ~n4047 & ~n4048;
  assign n4050 = n4046 & n4049;
  assign n4058 = n4057 ^ n4050;
  assign n4066 = n4065 ^ n4058;
  assign n4090 = n4089 ^ n4066;
  assign n4114 = n4113 ^ n4090;
  assign n4041 = n3981 ^ n3957;
  assign n4042 = ~n3958 & n4041;
  assign n4043 = n4042 ^ n3981;
  assign n4115 = n4114 ^ n4043;
  assign n4037 = n3870 ^ n3855;
  assign n4038 = n3858 ^ n3855;
  assign n4039 = ~n4037 & ~n4038;
  assign n4040 = n4039 ^ n3870;
  assign n4116 = n4115 ^ n4040;
  assign n4034 = n3911 ^ n3872;
  assign n4035 = n3983 & n4034;
  assign n4036 = n4035 ^ n3982;
  assign n4117 = n4116 ^ n4036;
  assign n4031 = n4015 ^ n3993;
  assign n4032 = ~n3994 & ~n4031;
  assign n4033 = n4032 ^ n4015;
  assign n4118 = n4117 ^ n4033;
  assign n4198 = n4197 ^ n4118;
  assign n4028 = n3852 ^ n3849;
  assign n4029 = n3985 & n4028;
  assign n4030 = n4029 ^ n3984;
  assign n4199 = n4198 ^ n4030;
  assign n4025 = n3986 ^ n3846;
  assign n4026 = ~n4017 & n4025;
  assign n4027 = n4026 ^ n4016;
  assign n4200 = n4199 ^ n4027;
  assign n4205 = n4204 ^ n4200;
  assign n4376 = n4027 & ~n4199;
  assign n4377 = ~n4027 & n4199;
  assign n4378 = ~n4204 & ~n4377;
  assign n4379 = ~n4376 & ~n4378;
  assign n4361 = ~x25 & n650;
  assign n4362 = ~x24 & n654;
  assign n4363 = ~n4361 & ~n4362;
  assign n4364 = x25 & n657;
  assign n4365 = x24 & n659;
  assign n4366 = ~n4364 & ~n4365;
  assign n4367 = n4363 & n4366;
  assign n4353 = ~x19 & n1230;
  assign n4354 = ~x18 & n1232;
  assign n4355 = ~n4353 & ~n4354;
  assign n4356 = x19 & n1223;
  assign n4357 = x18 & n1227;
  assign n4358 = ~n4356 & ~n4357;
  assign n4359 = n4355 & n4358;
  assign n4346 = x17 & n1578;
  assign n4347 = x16 & n1580;
  assign n4348 = ~n4346 & ~n4347;
  assign n4349 = ~x17 & n1571;
  assign n4350 = ~x16 & n1575;
  assign n4351 = ~n4349 & ~n4350;
  assign n4352 = n4348 & n4351;
  assign n4360 = n4359 ^ n4352;
  assign n4368 = n4367 ^ n4360;
  assign n4342 = n4088 ^ n4080;
  assign n4343 = ~n4081 & n4342;
  assign n4344 = n4343 ^ n4088;
  assign n4338 = n4112 ^ n4104;
  assign n4339 = n4112 ^ n4097;
  assign n4340 = n4338 & ~n4339;
  assign n4341 = n4340 ^ n4104;
  assign n4345 = n4344 ^ n4341;
  assign n4369 = n4368 ^ n4345;
  assign n4333 = n4193 ^ n4178;
  assign n4334 = n4186 & ~n4333;
  assign n4335 = n4334 ^ n4185;
  assign n4336 = n4335 ^ n4140;
  assign n4330 = n4065 ^ n4050;
  assign n4331 = n4058 & ~n4330;
  assign n4332 = n4331 ^ n4057;
  assign n4337 = n4336 ^ n4332;
  assign n4370 = n4369 ^ n4337;
  assign n4327 = n4194 ^ n4170;
  assign n4328 = ~n4171 & n4327;
  assign n4329 = n4328 ^ n4194;
  assign n4371 = n4370 ^ n4329;
  assign n4322 = n4141 ^ n4124;
  assign n4323 = n4128 ^ n4124;
  assign n4324 = n4322 & ~n4323;
  assign n4325 = n4324 ^ n4141;
  assign n4319 = n4195 ^ n4162;
  assign n4320 = n4163 & n4319;
  assign n4321 = n4320 ^ n4195;
  assign n4326 = n4325 ^ n4321;
  assign n4372 = n4371 ^ n4326;
  assign n4306 = ~x9 & n2799;
  assign n4307 = ~x8 & n2803;
  assign n4308 = ~n4306 & ~n4307;
  assign n4309 = x9 & n2806;
  assign n4310 = x8 & n2808;
  assign n4311 = ~n4309 & ~n4310;
  assign n4312 = n4308 & n4311;
  assign n4298 = ~x23 & n821;
  assign n4299 = ~x22 & n823;
  assign n4300 = ~n4298 & ~n4299;
  assign n4301 = x23 & n814;
  assign n4302 = x22 & n818;
  assign n4303 = ~n4301 & ~n4302;
  assign n4304 = n4300 & n4303;
  assign n4291 = ~x11 & n2386;
  assign n4292 = ~x10 & n2388;
  assign n4293 = ~n4291 & ~n4292;
  assign n4294 = x11 & n2379;
  assign n4295 = x10 & n2383;
  assign n4296 = ~n4294 & ~n4295;
  assign n4297 = n4293 & n4296;
  assign n4305 = n4304 ^ n4297;
  assign n4313 = n4312 ^ n4305;
  assign n4282 = ~x27 & n510;
  assign n4283 = ~x26 & n512;
  assign n4284 = ~n4282 & ~n4283;
  assign n4285 = x27 & n503;
  assign n4286 = x26 & n507;
  assign n4287 = ~n4285 & ~n4286;
  assign n4288 = n4284 & n4287;
  assign n4280 = ~n147 & ~n151;
  assign n4273 = ~x31 & n247;
  assign n4274 = ~x30 & n251;
  assign n4275 = ~n4273 & ~n4274;
  assign n4276 = x31 & n254;
  assign n4277 = x30 & n256;
  assign n4278 = ~n4276 & ~n4277;
  assign n4279 = n4275 & n4278;
  assign n4281 = n4280 ^ n4279;
  assign n4289 = n4288 ^ n4281;
  assign n4271 = x5 & x63;
  assign n4263 = ~x21 & n1004;
  assign n4264 = ~x20 & n1008;
  assign n4265 = ~n4263 & ~n4264;
  assign n4266 = x21 & n1011;
  assign n4267 = x20 & n1013;
  assign n4268 = ~n4266 & ~n4267;
  assign n4269 = n4265 & n4268;
  assign n4256 = ~x7 & n3129;
  assign n4257 = ~x6 & n3133;
  assign n4258 = ~n4256 & ~n4257;
  assign n4259 = x7 & n3136;
  assign n4260 = x6 & n3138;
  assign n4261 = ~n4259 & ~n4260;
  assign n4262 = n4258 & n4261;
  assign n4270 = n4269 ^ n4262;
  assign n4272 = n4271 ^ n4270;
  assign n4290 = n4289 ^ n4272;
  assign n4314 = n4313 ^ n4290;
  assign n4252 = n4113 ^ n4089;
  assign n4253 = n4113 ^ n4066;
  assign n4254 = n4252 & ~n4253;
  assign n4255 = n4254 ^ n4089;
  assign n4315 = n4314 ^ n4255;
  assign n4242 = ~x29 & n346;
  assign n4243 = ~x28 & n350;
  assign n4244 = ~n4242 & ~n4243;
  assign n4245 = x29 & n353;
  assign n4246 = x28 & n355;
  assign n4247 = ~n4245 & ~n4246;
  assign n4248 = n4244 & n4247;
  assign n4234 = ~x15 & n1835;
  assign n4235 = ~x14 & n1839;
  assign n4236 = ~n4234 & ~n4235;
  assign n4237 = x15 & n1842;
  assign n4238 = x14 & n1844;
  assign n4239 = ~n4237 & ~n4238;
  assign n4240 = n4236 & n4239;
  assign n4227 = x13 & n2168;
  assign n4228 = x12 & n2170;
  assign n4229 = ~n4227 & ~n4228;
  assign n4230 = ~x13 & n2161;
  assign n4231 = ~x12 & n2165;
  assign n4232 = ~n4230 & ~n4231;
  assign n4233 = n4229 & n4232;
  assign n4241 = n4240 ^ n4233;
  assign n4249 = n4248 ^ n4241;
  assign n4223 = n4140 ^ n4136;
  assign n4224 = n4140 ^ n4135;
  assign n4225 = n4223 & n4224;
  assign n4226 = n4225 ^ n4136;
  assign n4250 = n4249 ^ n4226;
  assign n4219 = n4160 ^ n4152;
  assign n4220 = n4156 ^ n4152;
  assign n4221 = ~n4219 & n4220;
  assign n4222 = n4221 ^ n4160;
  assign n4251 = n4250 ^ n4222;
  assign n4316 = n4315 ^ n4251;
  assign n4216 = n4043 ^ n4040;
  assign n4217 = n4115 & n4216;
  assign n4218 = n4217 ^ n4114;
  assign n4317 = n4316 ^ n4218;
  assign n4212 = n4196 ^ n4143;
  assign n4213 = n4196 ^ n4121;
  assign n4214 = ~n4212 & n4213;
  assign n4215 = n4214 ^ n4143;
  assign n4318 = n4317 ^ n4215;
  assign n4373 = n4372 ^ n4318;
  assign n4209 = n4036 ^ n4033;
  assign n4210 = ~n4117 & n4209;
  assign n4211 = n4210 ^ n4116;
  assign n4374 = n4373 ^ n4211;
  assign n4206 = n4118 ^ n4030;
  assign n4207 = ~n4198 & n4206;
  assign n4208 = n4207 ^ n4197;
  assign n4375 = n4374 ^ n4208;
  assign n4380 = n4379 ^ n4375;
  assign n4540 = n4208 & n4374;
  assign n4541 = ~n4208 & ~n4374;
  assign n4542 = ~n4379 & ~n4541;
  assign n4543 = ~n4540 & ~n4542;
  assign n4527 = n4288 ^ n4280;
  assign n4528 = n4288 ^ n4279;
  assign n4529 = ~n4527 & ~n4528;
  assign n4530 = n4529 ^ n4280;
  assign n4524 = n4367 ^ n4359;
  assign n4525 = ~n4360 & n4524;
  assign n4526 = n4525 ^ n4367;
  assign n4531 = n4530 ^ n4526;
  assign n4521 = n4248 ^ n4233;
  assign n4522 = n4241 & ~n4521;
  assign n4523 = n4522 ^ n4240;
  assign n4532 = n4531 ^ n4523;
  assign n4518 = n4335 ^ n4332;
  assign n4519 = n4336 & ~n4518;
  assign n4520 = n4519 ^ n4140;
  assign n4533 = n4532 ^ n4520;
  assign n4515 = n4368 ^ n4344;
  assign n4516 = ~n4345 & n4515;
  assign n4517 = n4516 ^ n4368;
  assign n4534 = n4533 ^ n4517;
  assign n4504 = ~x10 & n2799;
  assign n4505 = ~x9 & n2803;
  assign n4506 = ~n4504 & ~n4505;
  assign n4507 = x10 & n2806;
  assign n4508 = x9 & n2808;
  assign n4509 = ~n4507 & ~n4508;
  assign n4510 = n4506 & n4509;
  assign n4500 = x39 ^ x31;
  assign n4501 = n250 & n4500;
  assign n4502 = ~n247 & ~n4501;
  assign n4493 = ~x22 & n1004;
  assign n4494 = ~x21 & n1008;
  assign n4495 = ~n4493 & ~n4494;
  assign n4496 = x22 & n1011;
  assign n4497 = x21 & n1013;
  assign n4498 = ~n4496 & ~n4497;
  assign n4499 = n4495 & n4498;
  assign n4503 = n4502 ^ n4499;
  assign n4511 = n4510 ^ n4503;
  assign n4485 = x12 & n2379;
  assign n4486 = x11 & n2383;
  assign n4487 = ~n4485 & ~n4486;
  assign n4488 = ~x12 & n2386;
  assign n4489 = ~x11 & n2388;
  assign n4490 = ~n4488 & ~n4489;
  assign n4491 = n4487 & n4490;
  assign n4477 = ~x24 & n821;
  assign n4478 = ~x23 & n823;
  assign n4479 = ~n4477 & ~n4478;
  assign n4480 = x24 & n814;
  assign n4481 = x23 & n818;
  assign n4482 = ~n4480 & ~n4481;
  assign n4483 = n4479 & n4482;
  assign n4470 = ~x14 & n2161;
  assign n4471 = ~x13 & n2165;
  assign n4472 = ~n4470 & ~n4471;
  assign n4473 = x14 & n2168;
  assign n4474 = x13 & n2170;
  assign n4475 = ~n4473 & ~n4474;
  assign n4476 = n4472 & n4475;
  assign n4484 = n4483 ^ n4476;
  assign n4492 = n4491 ^ n4484;
  assign n4512 = n4511 ^ n4492;
  assign n4461 = ~x30 & n346;
  assign n4462 = ~x29 & n350;
  assign n4463 = ~n4461 & ~n4462;
  assign n4464 = x30 & n353;
  assign n4465 = x29 & n355;
  assign n4466 = ~n4464 & ~n4465;
  assign n4467 = n4463 & n4466;
  assign n4454 = ~x20 & n1230;
  assign n4455 = ~x19 & n1232;
  assign n4456 = ~n4454 & ~n4455;
  assign n4457 = x20 & n1223;
  assign n4458 = x19 & n1227;
  assign n4459 = ~n4457 & ~n4458;
  assign n4460 = n4456 & n4459;
  assign n4468 = n4467 ^ n4460;
  assign n4451 = n4312 ^ n4304;
  assign n4452 = ~n4305 & n4451;
  assign n4453 = n4452 ^ n4312;
  assign n4469 = n4468 ^ n4453;
  assign n4513 = n4512 ^ n4469;
  assign n4448 = n4337 ^ n4329;
  assign n4449 = n4370 & ~n4448;
  assign n4450 = n4449 ^ n4369;
  assign n4514 = n4513 ^ n4450;
  assign n4535 = n4534 ^ n4514;
  assign n4436 = ~x16 & n1835;
  assign n4437 = ~x15 & n1839;
  assign n4438 = ~n4436 & ~n4437;
  assign n4439 = x16 & n1842;
  assign n4440 = x15 & n1844;
  assign n4441 = ~n4439 & ~n4440;
  assign n4442 = n4438 & n4441;
  assign n4428 = ~x26 & n650;
  assign n4429 = ~x25 & n654;
  assign n4430 = ~n4428 & ~n4429;
  assign n4431 = x26 & n657;
  assign n4432 = x25 & n659;
  assign n4433 = ~n4431 & ~n4432;
  assign n4434 = n4430 & n4433;
  assign n4421 = ~x18 & n1571;
  assign n4422 = ~x17 & n1575;
  assign n4423 = ~n4421 & ~n4422;
  assign n4424 = x18 & n1578;
  assign n4425 = x17 & n1580;
  assign n4426 = ~n4424 & ~n4425;
  assign n4427 = n4423 & n4426;
  assign n4435 = n4434 ^ n4427;
  assign n4443 = n4442 ^ n4435;
  assign n4418 = x6 & x63;
  assign n4410 = ~x28 & n510;
  assign n4411 = ~x27 & n512;
  assign n4412 = ~n4410 & ~n4411;
  assign n4413 = x28 & n503;
  assign n4414 = x27 & n507;
  assign n4415 = ~n4413 & ~n4414;
  assign n4416 = n4412 & n4415;
  assign n4403 = ~x8 & n3129;
  assign n4404 = ~x7 & n3133;
  assign n4405 = ~n4403 & ~n4404;
  assign n4406 = x8 & n3136;
  assign n4407 = x7 & n3138;
  assign n4408 = ~n4406 & ~n4407;
  assign n4409 = n4405 & n4408;
  assign n4417 = n4416 ^ n4409;
  assign n4419 = n4418 ^ n4417;
  assign n4400 = n4271 ^ n4269;
  assign n4401 = ~n4270 & ~n4400;
  assign n4402 = n4401 ^ n4271;
  assign n4420 = n4419 ^ n4402;
  assign n4444 = n4443 ^ n4420;
  assign n4396 = n4313 ^ n4289;
  assign n4397 = n4313 ^ n4272;
  assign n4398 = ~n4396 & n4397;
  assign n4399 = n4398 ^ n4289;
  assign n4445 = n4444 ^ n4399;
  assign n4393 = n4226 ^ n4222;
  assign n4394 = ~n4250 & ~n4393;
  assign n4395 = n4394 ^ n4249;
  assign n4446 = n4445 ^ n4395;
  assign n4390 = n4255 ^ n4251;
  assign n4391 = n4315 & ~n4390;
  assign n4392 = n4391 ^ n4314;
  assign n4447 = n4446 ^ n4392;
  assign n4536 = n4535 ^ n4447;
  assign n4387 = n4371 ^ n4325;
  assign n4388 = ~n4326 & n4387;
  assign n4389 = n4388 ^ n4371;
  assign n4537 = n4536 ^ n4389;
  assign n4384 = n4218 ^ n4215;
  assign n4385 = n4317 & ~n4384;
  assign n4386 = n4385 ^ n4316;
  assign n4538 = n4537 ^ n4386;
  assign n4381 = n4318 ^ n4211;
  assign n4382 = n4373 & n4381;
  assign n4383 = n4382 ^ n4372;
  assign n4539 = n4538 ^ n4383;
  assign n4544 = n4543 ^ n4539;
  assign n4700 = ~n4383 & n4538;
  assign n4701 = n4383 & ~n4538;
  assign n4702 = ~n4543 & ~n4701;
  assign n4703 = ~n4700 & ~n4702;
  assign n4688 = n4491 ^ n4483;
  assign n4689 = ~n4484 & n4688;
  assign n4690 = n4689 ^ n4491;
  assign n4685 = n4442 ^ n4434;
  assign n4686 = ~n4435 & n4685;
  assign n4687 = n4686 ^ n4442;
  assign n4691 = n4690 ^ n4687;
  assign n4682 = n4510 ^ n4499;
  assign n4683 = n4503 & ~n4682;
  assign n4684 = n4683 ^ n4502;
  assign n4692 = n4691 ^ n4684;
  assign n4678 = n4460 ^ n4453;
  assign n4679 = ~n4468 & ~n4678;
  assign n4680 = n4679 ^ n4467;
  assign n4675 = n4526 ^ n4523;
  assign n4676 = ~n4531 & ~n4675;
  assign n4677 = n4676 ^ n4530;
  assign n4681 = n4680 ^ n4677;
  assign n4693 = n4692 ^ n4681;
  assign n4672 = n4492 ^ n4469;
  assign n4673 = n4512 & n4672;
  assign n4674 = n4673 ^ n4511;
  assign n4694 = n4693 ^ n4674;
  assign n4668 = n4532 ^ n4517;
  assign n4669 = n4520 ^ n4517;
  assign n4670 = ~n4668 & ~n4669;
  assign n4671 = n4670 ^ n4532;
  assign n4695 = n4694 ^ n4671;
  assign n4662 = x7 & x63;
  assign n4655 = ~x21 & n1230;
  assign n4656 = ~x20 & n1232;
  assign n4657 = ~n4655 & ~n4656;
  assign n4658 = x21 & n1223;
  assign n4659 = x20 & n1227;
  assign n4660 = ~n4658 & ~n4659;
  assign n4661 = n4657 & n4660;
  assign n4663 = n4662 ^ n4661;
  assign n4664 = n4663 ^ n4467;
  assign n4646 = x9 & n3136;
  assign n4647 = x8 & n3138;
  assign n4648 = ~n4646 & ~n4647;
  assign n4649 = ~x9 & n3129;
  assign n4650 = ~x8 & n3133;
  assign n4651 = ~n4649 & ~n4650;
  assign n4652 = n4648 & n4651;
  assign n4638 = x23 & n1011;
  assign n4639 = x22 & n1013;
  assign n4640 = ~n4638 & ~n4639;
  assign n4641 = ~x23 & n1004;
  assign n4642 = ~x22 & n1008;
  assign n4643 = ~n4641 & ~n4642;
  assign n4644 = n4640 & n4643;
  assign n4631 = ~x11 & n2799;
  assign n4632 = ~x10 & n2803;
  assign n4633 = ~n4631 & ~n4632;
  assign n4634 = x11 & n2806;
  assign n4635 = x10 & n2808;
  assign n4636 = ~n4634 & ~n4635;
  assign n4637 = n4633 & n4636;
  assign n4645 = n4644 ^ n4637;
  assign n4653 = n4652 ^ n4645;
  assign n4623 = ~x29 & n510;
  assign n4624 = ~x28 & n512;
  assign n4625 = ~n4623 & ~n4624;
  assign n4626 = x29 & n503;
  assign n4627 = x28 & n507;
  assign n4628 = ~n4626 & ~n4627;
  assign n4629 = n4625 & n4628;
  assign n4615 = x15 & n2168;
  assign n4616 = x14 & n2170;
  assign n4617 = ~n4615 & ~n4616;
  assign n4618 = ~x15 & n2161;
  assign n4619 = ~x14 & n2165;
  assign n4620 = ~n4618 & ~n4619;
  assign n4621 = n4617 & n4620;
  assign n4608 = ~x13 & n2386;
  assign n4609 = ~x12 & n2388;
  assign n4610 = ~n4608 & ~n4609;
  assign n4611 = x13 & n2379;
  assign n4612 = x12 & n2383;
  assign n4613 = ~n4611 & ~n4612;
  assign n4614 = n4610 & n4613;
  assign n4622 = n4621 ^ n4614;
  assign n4630 = n4629 ^ n4622;
  assign n4654 = n4653 ^ n4630;
  assign n4665 = n4664 ^ n4654;
  assign n4598 = x27 & n657;
  assign n4599 = x26 & n659;
  assign n4600 = ~n4598 & ~n4599;
  assign n4601 = ~x27 & n650;
  assign n4602 = ~x26 & n654;
  assign n4603 = ~n4601 & ~n4602;
  assign n4604 = n4600 & n4603;
  assign n4596 = ~n247 & ~n251;
  assign n4589 = ~x31 & n346;
  assign n4590 = ~x30 & n350;
  assign n4591 = ~n4589 & ~n4590;
  assign n4592 = x31 & n353;
  assign n4593 = x30 & n355;
  assign n4594 = ~n4592 & ~n4593;
  assign n4595 = n4591 & n4594;
  assign n4597 = n4596 ^ n4595;
  assign n4605 = n4604 ^ n4597;
  assign n4580 = ~x25 & n821;
  assign n4581 = ~x24 & n823;
  assign n4582 = ~n4580 & ~n4581;
  assign n4583 = x25 & n814;
  assign n4584 = x24 & n818;
  assign n4585 = ~n4583 & ~n4584;
  assign n4586 = n4582 & n4585;
  assign n4572 = ~x19 & n1571;
  assign n4573 = ~x18 & n1575;
  assign n4574 = ~n4572 & ~n4573;
  assign n4575 = x19 & n1578;
  assign n4576 = x18 & n1580;
  assign n4577 = ~n4575 & ~n4576;
  assign n4578 = n4574 & n4577;
  assign n4565 = ~x17 & n1835;
  assign n4566 = ~x16 & n1839;
  assign n4567 = ~n4565 & ~n4566;
  assign n4568 = x17 & n1842;
  assign n4569 = x16 & n1844;
  assign n4570 = ~n4568 & ~n4569;
  assign n4571 = n4567 & n4570;
  assign n4579 = n4578 ^ n4571;
  assign n4587 = n4586 ^ n4579;
  assign n4562 = n4418 ^ n4416;
  assign n4563 = ~n4417 & ~n4562;
  assign n4564 = n4563 ^ n4418;
  assign n4588 = n4587 ^ n4564;
  assign n4606 = n4605 ^ n4588;
  assign n4559 = n4443 ^ n4419;
  assign n4560 = ~n4420 & ~n4559;
  assign n4561 = n4560 ^ n4443;
  assign n4607 = n4606 ^ n4561;
  assign n4666 = n4665 ^ n4607;
  assign n4556 = n4399 ^ n4395;
  assign n4557 = ~n4445 & n4556;
  assign n4558 = n4557 ^ n4444;
  assign n4667 = n4666 ^ n4558;
  assign n4696 = n4695 ^ n4667;
  assign n4552 = n4534 ^ n4513;
  assign n4553 = n4534 ^ n4450;
  assign n4554 = n4552 & n4553;
  assign n4555 = n4554 ^ n4513;
  assign n4697 = n4696 ^ n4555;
  assign n4548 = n4535 ^ n4446;
  assign n4549 = n4535 ^ n4392;
  assign n4550 = ~n4548 & ~n4549;
  assign n4551 = n4550 ^ n4446;
  assign n4698 = n4697 ^ n4551;
  assign n4545 = n4389 ^ n4386;
  assign n4546 = ~n4537 & ~n4545;
  assign n4547 = n4546 ^ n4536;
  assign n4699 = n4698 ^ n4547;
  assign n4704 = n4703 ^ n4699;
  assign n4853 = n4547 & ~n4698;
  assign n4854 = ~n4547 & n4698;
  assign n4855 = ~n4703 & ~n4854;
  assign n4856 = ~n4853 & ~n4855;
  assign n4839 = ~x30 & n510;
  assign n4840 = ~x29 & n512;
  assign n4841 = ~n4839 & ~n4840;
  assign n4842 = x30 & n503;
  assign n4843 = x29 & n507;
  assign n4844 = ~n4842 & ~n4843;
  assign n4845 = n4841 & n4844;
  assign n4836 = n4586 ^ n4578;
  assign n4837 = ~n4579 & n4836;
  assign n4838 = n4837 ^ n4586;
  assign n4846 = n4845 ^ n4838;
  assign n4833 = n4629 ^ n4621;
  assign n4834 = ~n4622 & n4833;
  assign n4835 = n4834 ^ n4629;
  assign n4847 = n4846 ^ n4835;
  assign n4829 = n4661 ^ n4467;
  assign n4830 = ~n4663 & ~n4829;
  assign n4831 = n4830 ^ n4662;
  assign n4826 = n4687 ^ n4684;
  assign n4827 = n4691 & ~n4826;
  assign n4828 = n4827 ^ n4690;
  assign n4832 = n4831 ^ n4828;
  assign n4848 = n4847 ^ n4832;
  assign n4816 = ~x12 & n2799;
  assign n4817 = ~x11 & n2803;
  assign n4818 = ~n4816 & ~n4817;
  assign n4819 = x12 & n2806;
  assign n4820 = x11 & n2808;
  assign n4821 = ~n4819 & ~n4820;
  assign n4822 = n4818 & n4821;
  assign n4808 = ~x24 & n1004;
  assign n4809 = ~x23 & n1008;
  assign n4810 = ~n4808 & ~n4809;
  assign n4811 = x24 & n1011;
  assign n4812 = x23 & n1013;
  assign n4813 = ~n4811 & ~n4812;
  assign n4814 = n4810 & n4813;
  assign n4801 = ~x14 & n2386;
  assign n4802 = ~x13 & n2388;
  assign n4803 = ~n4801 & ~n4802;
  assign n4804 = x14 & n2379;
  assign n4805 = x13 & n2383;
  assign n4806 = ~n4804 & ~n4805;
  assign n4807 = n4803 & n4806;
  assign n4815 = n4814 ^ n4807;
  assign n4823 = n4822 ^ n4815;
  assign n4792 = ~x16 & n2161;
  assign n4793 = ~x15 & n2165;
  assign n4794 = ~n4792 & ~n4793;
  assign n4795 = x16 & n2168;
  assign n4796 = x15 & n2170;
  assign n4797 = ~n4795 & ~n4796;
  assign n4798 = n4794 & n4797;
  assign n4784 = ~x18 & n1835;
  assign n4785 = ~x17 & n1839;
  assign n4786 = ~n4784 & ~n4785;
  assign n4787 = x18 & n1842;
  assign n4788 = x17 & n1844;
  assign n4789 = ~n4787 & ~n4788;
  assign n4790 = n4786 & n4789;
  assign n4777 = x26 & n814;
  assign n4778 = x25 & n818;
  assign n4779 = ~n4777 & ~n4778;
  assign n4780 = ~x26 & n821;
  assign n4781 = ~x25 & n823;
  assign n4782 = ~n4780 & ~n4781;
  assign n4783 = n4779 & n4782;
  assign n4791 = n4790 ^ n4783;
  assign n4799 = n4798 ^ n4791;
  assign n4769 = ~x10 & n3129;
  assign n4770 = ~x9 & n3133;
  assign n4771 = ~n4769 & ~n4770;
  assign n4772 = x10 & n3136;
  assign n4773 = x9 & n3138;
  assign n4774 = ~n4772 & ~n4773;
  assign n4775 = n4771 & n4774;
  assign n4765 = x41 ^ x31;
  assign n4766 = n349 & n4765;
  assign n4767 = ~n346 & ~n4766;
  assign n4758 = x22 & n1223;
  assign n4759 = x21 & n1227;
  assign n4760 = ~n4758 & ~n4759;
  assign n4761 = ~x22 & n1230;
  assign n4762 = ~x21 & n1232;
  assign n4763 = ~n4761 & ~n4762;
  assign n4764 = n4760 & n4763;
  assign n4768 = n4767 ^ n4764;
  assign n4776 = n4775 ^ n4768;
  assign n4800 = n4799 ^ n4776;
  assign n4824 = n4823 ^ n4800;
  assign n4755 = n4692 ^ n4680;
  assign n4756 = ~n4681 & ~n4755;
  assign n4757 = n4756 ^ n4692;
  assign n4825 = n4824 ^ n4757;
  assign n4849 = n4848 ^ n4825;
  assign n4742 = ~x20 & n1571;
  assign n4743 = ~x19 & n1575;
  assign n4744 = ~n4742 & ~n4743;
  assign n4745 = x20 & n1578;
  assign n4746 = x19 & n1580;
  assign n4747 = ~n4745 & ~n4746;
  assign n4748 = n4744 & n4747;
  assign n4740 = x8 & x63;
  assign n4733 = x28 & n657;
  assign n4734 = x27 & n659;
  assign n4735 = ~n4733 & ~n4734;
  assign n4736 = ~x28 & n650;
  assign n4737 = ~x27 & n654;
  assign n4738 = ~n4736 & ~n4737;
  assign n4739 = n4735 & n4738;
  assign n4741 = n4740 ^ n4739;
  assign n4749 = n4748 ^ n4741;
  assign n4728 = n4604 ^ n4596;
  assign n4729 = n4604 ^ n4595;
  assign n4730 = ~n4728 & ~n4729;
  assign n4731 = n4730 ^ n4596;
  assign n4725 = n4652 ^ n4637;
  assign n4726 = n4645 & ~n4725;
  assign n4727 = n4726 ^ n4644;
  assign n4732 = n4731 ^ n4727;
  assign n4750 = n4749 ^ n4732;
  assign n4722 = n4605 ^ n4587;
  assign n4723 = n4588 & ~n4722;
  assign n4724 = n4723 ^ n4605;
  assign n4751 = n4750 ^ n4724;
  assign n4719 = n4664 ^ n4653;
  assign n4720 = ~n4654 & ~n4719;
  assign n4721 = n4720 ^ n4664;
  assign n4752 = n4751 ^ n4721;
  assign n4716 = n4665 ^ n4606;
  assign n4717 = ~n4607 & ~n4716;
  assign n4718 = n4717 ^ n4665;
  assign n4753 = n4752 ^ n4718;
  assign n4713 = n4693 ^ n4671;
  assign n4714 = n4694 & n4713;
  assign n4715 = n4714 ^ n4674;
  assign n4754 = n4753 ^ n4715;
  assign n4850 = n4849 ^ n4754;
  assign n4709 = n4695 ^ n4666;
  assign n4710 = n4695 ^ n4558;
  assign n4711 = n4709 & n4710;
  assign n4712 = n4711 ^ n4666;
  assign n4851 = n4850 ^ n4712;
  assign n4705 = n4555 ^ n4551;
  assign n4706 = n4696 ^ n4551;
  assign n4707 = n4705 & n4706;
  assign n4708 = n4707 ^ n4555;
  assign n4852 = n4851 ^ n4708;
  assign n4857 = n4856 ^ n4852;
  assign n5004 = n4708 & ~n4851;
  assign n5005 = ~n4708 & n4851;
  assign n5006 = ~n4856 & ~n5005;
  assign n5007 = ~n5004 & ~n5006;
  assign n4996 = x9 & x63;
  assign n4988 = ~x23 & n1230;
  assign n4989 = ~x22 & n1232;
  assign n4990 = ~n4988 & ~n4989;
  assign n4991 = x23 & n1223;
  assign n4992 = x22 & n1227;
  assign n4993 = ~n4991 & ~n4992;
  assign n4994 = n4990 & n4993;
  assign n4981 = ~x11 & n3129;
  assign n4982 = ~x10 & n3133;
  assign n4983 = ~n4981 & ~n4982;
  assign n4984 = x11 & n3136;
  assign n4985 = x10 & n3138;
  assign n4986 = ~n4984 & ~n4985;
  assign n4987 = n4983 & n4986;
  assign n4995 = n4994 ^ n4987;
  assign n4997 = n4996 ^ n4995;
  assign n4972 = ~x21 & n1571;
  assign n4973 = ~x20 & n1575;
  assign n4974 = ~n4972 & ~n4973;
  assign n4975 = x21 & n1578;
  assign n4976 = x20 & n1580;
  assign n4977 = ~n4975 & ~n4976;
  assign n4978 = n4974 & n4977;
  assign n4979 = n4978 ^ n4845;
  assign n4969 = n4822 ^ n4814;
  assign n4970 = ~n4815 & n4969;
  assign n4971 = n4970 ^ n4822;
  assign n4980 = n4979 ^ n4971;
  assign n4998 = n4997 ^ n4980;
  assign n4966 = n4838 ^ n4835;
  assign n4967 = ~n4846 & ~n4966;
  assign n4968 = n4967 ^ n4845;
  assign n4999 = n4998 ^ n4968;
  assign n4956 = x25 & n1011;
  assign n4957 = x24 & n1013;
  assign n4958 = ~n4956 & ~n4957;
  assign n4959 = ~x25 & n1004;
  assign n4960 = ~x24 & n1008;
  assign n4961 = ~n4959 & ~n4960;
  assign n4962 = n4958 & n4961;
  assign n4948 = x19 & n1842;
  assign n4949 = x18 & n1844;
  assign n4950 = ~n4948 & ~n4949;
  assign n4951 = ~x19 & n1835;
  assign n4952 = ~x18 & n1839;
  assign n4953 = ~n4951 & ~n4952;
  assign n4954 = n4950 & n4953;
  assign n4941 = ~x17 & n2161;
  assign n4942 = ~x16 & n2165;
  assign n4943 = ~n4941 & ~n4942;
  assign n4944 = x17 & n2168;
  assign n4945 = x16 & n2170;
  assign n4946 = ~n4944 & ~n4945;
  assign n4947 = n4943 & n4946;
  assign n4955 = n4954 ^ n4947;
  assign n4963 = n4962 ^ n4955;
  assign n4932 = x27 & n814;
  assign n4933 = x26 & n818;
  assign n4934 = ~n4932 & ~n4933;
  assign n4935 = ~x27 & n821;
  assign n4936 = ~x26 & n823;
  assign n4937 = ~n4935 & ~n4936;
  assign n4938 = n4934 & n4937;
  assign n4930 = ~n346 & ~n350;
  assign n4923 = ~x31 & n510;
  assign n4924 = ~x30 & n512;
  assign n4925 = ~n4923 & ~n4924;
  assign n4926 = x31 & n503;
  assign n4927 = x30 & n507;
  assign n4928 = ~n4926 & ~n4927;
  assign n4929 = n4925 & n4928;
  assign n4931 = n4930 ^ n4929;
  assign n4939 = n4938 ^ n4931;
  assign n4915 = ~x29 & n650;
  assign n4916 = ~x28 & n654;
  assign n4917 = ~n4915 & ~n4916;
  assign n4918 = x29 & n657;
  assign n4919 = x28 & n659;
  assign n4920 = ~n4918 & ~n4919;
  assign n4921 = n4917 & n4920;
  assign n4907 = ~x15 & n2386;
  assign n4908 = ~x14 & n2388;
  assign n4909 = ~n4907 & ~n4908;
  assign n4910 = x15 & n2379;
  assign n4911 = x14 & n2383;
  assign n4912 = ~n4910 & ~n4911;
  assign n4913 = n4909 & n4912;
  assign n4900 = ~x13 & n2799;
  assign n4901 = ~x12 & n2803;
  assign n4902 = ~n4900 & ~n4901;
  assign n4903 = x13 & n2806;
  assign n4904 = x12 & n2808;
  assign n4905 = ~n4903 & ~n4904;
  assign n4906 = n4902 & n4905;
  assign n4914 = n4913 ^ n4906;
  assign n4922 = n4921 ^ n4914;
  assign n4940 = n4939 ^ n4922;
  assign n4964 = n4963 ^ n4940;
  assign n4896 = n4847 ^ n4831;
  assign n4897 = n4847 ^ n4828;
  assign n4898 = n4896 & n4897;
  assign n4899 = n4898 ^ n4831;
  assign n4965 = n4964 ^ n4899;
  assign n5000 = n4999 ^ n4965;
  assign n4887 = n4748 ^ n4739;
  assign n4888 = ~n4741 & ~n4887;
  assign n4889 = n4888 ^ n4740;
  assign n4883 = n4775 ^ n4767;
  assign n4884 = n4775 ^ n4764;
  assign n4885 = n4883 & ~n4884;
  assign n4886 = n4885 ^ n4767;
  assign n4890 = n4889 ^ n4886;
  assign n4879 = n4798 ^ n4790;
  assign n4880 = n4798 ^ n4783;
  assign n4881 = n4879 & ~n4880;
  assign n4882 = n4881 ^ n4790;
  assign n4891 = n4890 ^ n4882;
  assign n4876 = n4749 ^ n4731;
  assign n4877 = n4732 & n4876;
  assign n4878 = n4877 ^ n4749;
  assign n4892 = n4891 ^ n4878;
  assign n4872 = n4823 ^ n4799;
  assign n4873 = n4823 ^ n4776;
  assign n4874 = n4872 & ~n4873;
  assign n4875 = n4874 ^ n4799;
  assign n4893 = n4892 ^ n4875;
  assign n4868 = n4750 ^ n4721;
  assign n4869 = n4724 ^ n4721;
  assign n4870 = ~n4868 & ~n4869;
  assign n4871 = n4870 ^ n4750;
  assign n4894 = n4893 ^ n4871;
  assign n4864 = n4848 ^ n4824;
  assign n4865 = n4848 ^ n4757;
  assign n4866 = n4864 & ~n4865;
  assign n4867 = n4866 ^ n4824;
  assign n4895 = n4894 ^ n4867;
  assign n5001 = n5000 ^ n4895;
  assign n4861 = n4718 ^ n4715;
  assign n4862 = ~n4753 & n4861;
  assign n4863 = n4862 ^ n4752;
  assign n5002 = n5001 ^ n4863;
  assign n4858 = n4754 ^ n4712;
  assign n4859 = ~n4850 & ~n4858;
  assign n4860 = n4859 ^ n4849;
  assign n5003 = n5002 ^ n4860;
  assign n5008 = n5007 ^ n5003;
  assign n5144 = ~n4860 & ~n5002;
  assign n5145 = n4860 & n5002;
  assign n5146 = ~n5007 & ~n5145;
  assign n5147 = ~n5144 & ~n5146;
  assign n5130 = ~x30 & n650;
  assign n5131 = ~x29 & n654;
  assign n5132 = ~n5130 & ~n5131;
  assign n5133 = x30 & n657;
  assign n5134 = x29 & n659;
  assign n5135 = ~n5133 & ~n5134;
  assign n5136 = n5132 & n5135;
  assign n5122 = ~x20 & n1835;
  assign n5123 = ~x19 & n1839;
  assign n5124 = ~n5122 & ~n5123;
  assign n5125 = x20 & n1842;
  assign n5126 = x19 & n1844;
  assign n5127 = ~n5125 & ~n5126;
  assign n5128 = n5124 & n5127;
  assign n5115 = x22 & n1578;
  assign n5116 = x21 & n1580;
  assign n5117 = ~n5115 & ~n5116;
  assign n5118 = ~x22 & n1571;
  assign n5119 = ~x21 & n1575;
  assign n5120 = ~n5118 & ~n5119;
  assign n5121 = n5117 & n5120;
  assign n5129 = n5128 ^ n5121;
  assign n5137 = n5136 ^ n5129;
  assign n5107 = ~x12 & n3129;
  assign n5108 = ~x11 & n3133;
  assign n5109 = ~n5107 & ~n5108;
  assign n5110 = x12 & n3136;
  assign n5111 = x11 & n3138;
  assign n5112 = ~n5110 & ~n5111;
  assign n5113 = n5109 & n5112;
  assign n5099 = x14 & n2806;
  assign n5100 = x13 & n2808;
  assign n5101 = ~n5099 & ~n5100;
  assign n5102 = ~x14 & n2799;
  assign n5103 = ~x13 & n2803;
  assign n5104 = ~n5102 & ~n5103;
  assign n5105 = n5101 & n5104;
  assign n5092 = x24 & n1223;
  assign n5093 = x23 & n1227;
  assign n5094 = ~n5092 & ~n5093;
  assign n5095 = ~x24 & n1230;
  assign n5096 = ~x23 & n1232;
  assign n5097 = ~n5095 & ~n5096;
  assign n5098 = n5094 & n5097;
  assign n5106 = n5105 ^ n5098;
  assign n5114 = n5113 ^ n5106;
  assign n5138 = n5137 ^ n5114;
  assign n5088 = n4889 ^ n4882;
  assign n5089 = n4886 ^ n4882;
  assign n5090 = ~n5088 & ~n5089;
  assign n5091 = n5090 ^ n4889;
  assign n5139 = n5138 ^ n5091;
  assign n5078 = ~x16 & n2386;
  assign n5079 = ~x15 & n2388;
  assign n5080 = ~n5078 & ~n5079;
  assign n5081 = x16 & n2379;
  assign n5082 = x15 & n2383;
  assign n5083 = ~n5081 & ~n5082;
  assign n5084 = n5080 & n5083;
  assign n5070 = ~x18 & n2161;
  assign n5071 = ~x17 & n2165;
  assign n5072 = ~n5070 & ~n5071;
  assign n5073 = x18 & n2168;
  assign n5074 = x17 & n2170;
  assign n5075 = ~n5073 & ~n5074;
  assign n5076 = n5072 & n5075;
  assign n5063 = ~x26 & n1004;
  assign n5064 = ~x25 & n1008;
  assign n5065 = ~n5063 & ~n5064;
  assign n5066 = x26 & n1011;
  assign n5067 = x25 & n1013;
  assign n5068 = ~n5066 & ~n5067;
  assign n5069 = n5065 & n5068;
  assign n5077 = n5076 ^ n5069;
  assign n5085 = n5084 ^ n5077;
  assign n5060 = x10 & x63;
  assign n5056 = x43 ^ x31;
  assign n5057 = n506 & n5056;
  assign n5058 = ~n510 & ~n5057;
  assign n5049 = ~x28 & n821;
  assign n5050 = ~x27 & n823;
  assign n5051 = ~n5049 & ~n5050;
  assign n5052 = x28 & n814;
  assign n5053 = x27 & n818;
  assign n5054 = ~n5052 & ~n5053;
  assign n5055 = n5051 & n5054;
  assign n5059 = n5058 ^ n5055;
  assign n5061 = n5060 ^ n5059;
  assign n5046 = n4962 ^ n4947;
  assign n5047 = n4955 & ~n5046;
  assign n5048 = n5047 ^ n4954;
  assign n5062 = n5061 ^ n5048;
  assign n5086 = n5085 ^ n5062;
  assign n5043 = n4980 ^ n4968;
  assign n5044 = ~n4998 & n5043;
  assign n5045 = n5044 ^ n4997;
  assign n5087 = n5086 ^ n5045;
  assign n5140 = n5139 ^ n5087;
  assign n5034 = n4921 ^ n4913;
  assign n5035 = ~n4914 & n5034;
  assign n5036 = n5035 ^ n4921;
  assign n5031 = n4996 ^ n4994;
  assign n5032 = ~n4995 & ~n5031;
  assign n5033 = n5032 ^ n4996;
  assign n5037 = n5036 ^ n5033;
  assign n5028 = n4938 ^ n4929;
  assign n5029 = ~n4931 & ~n5028;
  assign n5030 = n5029 ^ n4930;
  assign n5038 = n5037 ^ n5030;
  assign n5025 = n4978 ^ n4971;
  assign n5026 = n4979 & ~n5025;
  assign n5027 = n5026 ^ n4845;
  assign n5039 = n5038 ^ n5027;
  assign n5022 = n4963 ^ n4922;
  assign n5023 = ~n4940 & ~n5022;
  assign n5024 = n5023 ^ n4939;
  assign n5040 = n5039 ^ n5024;
  assign n5019 = n4891 ^ n4875;
  assign n5020 = ~n4892 & ~n5019;
  assign n5021 = n5020 ^ n4875;
  assign n5041 = n5040 ^ n5021;
  assign n5015 = n4999 ^ n4964;
  assign n5016 = n4999 ^ n4899;
  assign n5017 = ~n5015 & n5016;
  assign n5018 = n5017 ^ n4964;
  assign n5042 = n5041 ^ n5018;
  assign n5141 = n5140 ^ n5042;
  assign n5012 = n4871 ^ n4867;
  assign n5013 = n4894 & ~n5012;
  assign n5014 = n5013 ^ n4893;
  assign n5142 = n5141 ^ n5014;
  assign n5009 = n4895 ^ n4863;
  assign n5010 = n5001 & ~n5009;
  assign n5011 = n5010 ^ n5000;
  assign n5143 = n5142 ^ n5011;
  assign n5148 = n5147 ^ n5143;
  assign n5283 = ~n5011 & ~n5142;
  assign n5284 = n5011 & n5142;
  assign n5285 = ~n5147 & ~n5284;
  assign n5286 = ~n5283 & ~n5285;
  assign n5269 = ~x21 & n1835;
  assign n5270 = ~x20 & n1839;
  assign n5271 = ~n5269 & ~n5270;
  assign n5272 = x21 & n1842;
  assign n5273 = x20 & n1844;
  assign n5274 = ~n5272 & ~n5273;
  assign n5275 = n5271 & n5274;
  assign n5267 = x11 & x63;
  assign n5260 = x23 & n1578;
  assign n5261 = x22 & n1580;
  assign n5262 = ~n5260 & ~n5261;
  assign n5263 = ~x23 & n1571;
  assign n5264 = ~x22 & n1575;
  assign n5265 = ~n5263 & ~n5264;
  assign n5266 = n5262 & n5265;
  assign n5268 = n5267 ^ n5266;
  assign n5276 = n5275 ^ n5268;
  assign n5251 = ~x29 & n821;
  assign n5252 = ~x28 & n823;
  assign n5253 = ~n5251 & ~n5252;
  assign n5254 = x29 & n814;
  assign n5255 = x28 & n818;
  assign n5256 = ~n5254 & ~n5255;
  assign n5257 = n5253 & n5256;
  assign n5243 = ~x15 & n2799;
  assign n5244 = ~x14 & n2803;
  assign n5245 = ~n5243 & ~n5244;
  assign n5246 = x15 & n2806;
  assign n5247 = x14 & n2808;
  assign n5248 = ~n5246 & ~n5247;
  assign n5249 = n5245 & n5248;
  assign n5236 = ~x13 & n3129;
  assign n5237 = ~x12 & n3133;
  assign n5238 = ~n5236 & ~n5237;
  assign n5239 = x13 & n3136;
  assign n5240 = x12 & n3138;
  assign n5241 = ~n5239 & ~n5240;
  assign n5242 = n5238 & n5241;
  assign n5250 = n5249 ^ n5242;
  assign n5258 = n5257 ^ n5250;
  assign n5232 = n5113 ^ n5105;
  assign n5233 = n5113 ^ n5098;
  assign n5234 = n5232 & ~n5233;
  assign n5235 = n5234 ^ n5105;
  assign n5259 = n5258 ^ n5235;
  assign n5277 = n5276 ^ n5259;
  assign n5222 = ~x27 & n1004;
  assign n5223 = ~x26 & n1008;
  assign n5224 = ~n5222 & ~n5223;
  assign n5225 = x27 & n1011;
  assign n5226 = x26 & n1013;
  assign n5227 = ~n5225 & ~n5226;
  assign n5228 = n5224 & n5227;
  assign n5220 = ~n510 & ~n512;
  assign n5213 = ~x31 & n650;
  assign n5214 = ~x30 & n654;
  assign n5215 = ~n5213 & ~n5214;
  assign n5216 = x31 & n657;
  assign n5217 = x30 & n659;
  assign n5218 = ~n5216 & ~n5217;
  assign n5219 = n5215 & n5218;
  assign n5221 = n5220 ^ n5219;
  assign n5229 = n5228 ^ n5221;
  assign n5205 = ~x25 & n1230;
  assign n5206 = ~x24 & n1232;
  assign n5207 = ~n5205 & ~n5206;
  assign n5208 = x25 & n1223;
  assign n5209 = x24 & n1227;
  assign n5210 = ~n5208 & ~n5209;
  assign n5211 = n5207 & n5210;
  assign n5197 = x19 & n2168;
  assign n5198 = x18 & n2170;
  assign n5199 = ~n5197 & ~n5198;
  assign n5200 = ~x19 & n2161;
  assign n5201 = ~x18 & n2165;
  assign n5202 = ~n5200 & ~n5201;
  assign n5203 = n5199 & n5202;
  assign n5190 = ~x17 & n2386;
  assign n5191 = ~x16 & n2388;
  assign n5192 = ~n5190 & ~n5191;
  assign n5193 = x17 & n2379;
  assign n5194 = x16 & n2383;
  assign n5195 = ~n5193 & ~n5194;
  assign n5196 = n5192 & n5195;
  assign n5204 = n5203 ^ n5196;
  assign n5212 = n5211 ^ n5204;
  assign n5230 = n5229 ^ n5212;
  assign n5186 = n5136 ^ n5128;
  assign n5187 = n5136 ^ n5121;
  assign n5188 = ~n5186 & n5187;
  assign n5189 = n5188 ^ n5128;
  assign n5231 = n5230 ^ n5189;
  assign n5278 = n5277 ^ n5231;
  assign n5183 = n5114 ^ n5091;
  assign n5184 = ~n5138 & n5183;
  assign n5185 = n5184 ^ n5137;
  assign n5279 = n5278 ^ n5185;
  assign n5175 = n5060 ^ n5058;
  assign n5176 = ~n5059 & ~n5175;
  assign n5177 = n5176 ^ n5060;
  assign n5178 = n5177 ^ n5136;
  assign n5172 = n5084 ^ n5069;
  assign n5173 = n5077 & ~n5172;
  assign n5174 = n5173 ^ n5076;
  assign n5179 = n5178 ^ n5174;
  assign n5167 = n5085 ^ n5061;
  assign n5168 = n5085 ^ n5048;
  assign n5169 = ~n5167 & ~n5168;
  assign n5170 = n5169 ^ n5061;
  assign n5163 = n5036 ^ n5030;
  assign n5164 = n5033 ^ n5030;
  assign n5165 = ~n5163 & ~n5164;
  assign n5166 = n5165 ^ n5036;
  assign n5171 = n5170 ^ n5166;
  assign n5180 = n5179 ^ n5171;
  assign n5159 = n5038 ^ n5024;
  assign n5160 = n5027 ^ n5024;
  assign n5161 = ~n5159 & n5160;
  assign n5162 = n5161 ^ n5038;
  assign n5181 = n5180 ^ n5162;
  assign n5155 = n5139 ^ n5086;
  assign n5156 = n5139 ^ n5045;
  assign n5157 = ~n5155 & n5156;
  assign n5158 = n5157 ^ n5086;
  assign n5182 = n5181 ^ n5158;
  assign n5280 = n5279 ^ n5182;
  assign n5152 = n5021 ^ n5018;
  assign n5153 = ~n5041 & n5152;
  assign n5154 = n5153 ^ n5040;
  assign n5281 = n5280 ^ n5154;
  assign n5149 = n5042 ^ n5014;
  assign n5150 = n5141 & ~n5149;
  assign n5151 = n5150 ^ n5140;
  assign n5282 = n5281 ^ n5151;
  assign n5287 = n5286 ^ n5282;
  assign n5410 = ~n5151 & n5281;
  assign n5411 = n5151 & ~n5281;
  assign n5412 = ~n5286 & ~n5411;
  assign n5413 = ~n5410 & ~n5412;
  assign n5397 = ~x16 & n2799;
  assign n5398 = ~x15 & n2803;
  assign n5399 = ~n5397 & ~n5398;
  assign n5400 = x16 & n2806;
  assign n5401 = x15 & n2808;
  assign n5402 = ~n5400 & ~n5401;
  assign n5403 = n5399 & n5402;
  assign n5389 = x18 & n2379;
  assign n5390 = x17 & n2383;
  assign n5391 = ~n5389 & ~n5390;
  assign n5392 = ~x18 & n2386;
  assign n5393 = ~x17 & n2388;
  assign n5394 = ~n5392 & ~n5393;
  assign n5395 = n5391 & n5394;
  assign n5382 = x26 & n1223;
  assign n5383 = x25 & n1227;
  assign n5384 = ~n5382 & ~n5383;
  assign n5385 = ~x26 & n1230;
  assign n5386 = ~x25 & n1232;
  assign n5387 = ~n5385 & ~n5386;
  assign n5388 = n5384 & n5387;
  assign n5396 = n5395 ^ n5388;
  assign n5404 = n5403 ^ n5396;
  assign n5373 = ~x22 & n1835;
  assign n5374 = ~x21 & n1839;
  assign n5375 = ~n5373 & ~n5374;
  assign n5376 = x22 & n1842;
  assign n5377 = x21 & n1844;
  assign n5378 = ~n5376 & ~n5377;
  assign n5379 = n5375 & n5378;
  assign n5369 = x45 ^ x31;
  assign n5370 = n653 & n5369;
  assign n5371 = ~n650 & ~n5370;
  assign n5362 = ~x28 & n1004;
  assign n5363 = ~x27 & n1008;
  assign n5364 = ~n5362 & ~n5363;
  assign n5365 = x28 & n1011;
  assign n5366 = x27 & n1013;
  assign n5367 = ~n5365 & ~n5366;
  assign n5368 = n5364 & n5367;
  assign n5372 = n5371 ^ n5368;
  assign n5380 = n5379 ^ n5372;
  assign n5360 = x12 & x63;
  assign n5352 = x24 & n1578;
  assign n5353 = x23 & n1580;
  assign n5354 = ~n5352 & ~n5353;
  assign n5355 = ~x24 & n1571;
  assign n5356 = ~x23 & n1575;
  assign n5357 = ~n5355 & ~n5356;
  assign n5358 = n5354 & n5357;
  assign n5345 = x14 & n3136;
  assign n5346 = x13 & n3138;
  assign n5347 = ~n5345 & ~n5346;
  assign n5348 = ~x14 & n3129;
  assign n5349 = ~x13 & n3133;
  assign n5350 = ~n5348 & ~n5349;
  assign n5351 = n5347 & n5350;
  assign n5359 = n5358 ^ n5351;
  assign n5361 = n5360 ^ n5359;
  assign n5381 = n5380 ^ n5361;
  assign n5405 = n5404 ^ n5381;
  assign n5341 = n5276 ^ n5258;
  assign n5342 = ~n5259 & ~n5341;
  assign n5343 = n5342 ^ n5276;
  assign n5338 = n5212 ^ n5189;
  assign n5339 = ~n5230 & ~n5338;
  assign n5340 = n5339 ^ n5229;
  assign n5344 = n5343 ^ n5340;
  assign n5406 = n5405 ^ n5344;
  assign n5330 = n5275 ^ n5266;
  assign n5331 = ~n5268 & ~n5330;
  assign n5332 = n5331 ^ n5267;
  assign n5327 = n5228 ^ n5219;
  assign n5328 = ~n5221 & ~n5327;
  assign n5329 = n5328 ^ n5220;
  assign n5333 = n5332 ^ n5329;
  assign n5324 = n5211 ^ n5196;
  assign n5325 = n5204 & ~n5324;
  assign n5326 = n5325 ^ n5203;
  assign n5334 = n5333 ^ n5326;
  assign n5314 = ~x30 & n821;
  assign n5315 = ~x29 & n823;
  assign n5316 = ~n5314 & ~n5315;
  assign n5317 = x30 & n814;
  assign n5318 = x29 & n818;
  assign n5319 = ~n5317 & ~n5318;
  assign n5320 = n5316 & n5319;
  assign n5307 = ~x20 & n2161;
  assign n5308 = ~x19 & n2165;
  assign n5309 = ~n5307 & ~n5308;
  assign n5310 = x20 & n2168;
  assign n5311 = x19 & n2170;
  assign n5312 = ~n5310 & ~n5311;
  assign n5313 = n5309 & n5312;
  assign n5321 = n5320 ^ n5313;
  assign n5303 = n5257 ^ n5249;
  assign n5304 = n5257 ^ n5242;
  assign n5305 = n5303 & ~n5304;
  assign n5306 = n5305 ^ n5249;
  assign n5322 = n5321 ^ n5306;
  assign n5300 = n5177 ^ n5174;
  assign n5301 = ~n5178 & n5300;
  assign n5302 = n5301 ^ n5136;
  assign n5323 = n5322 ^ n5302;
  assign n5335 = n5334 ^ n5323;
  assign n5297 = n5179 ^ n5170;
  assign n5298 = n5171 & n5297;
  assign n5299 = n5298 ^ n5179;
  assign n5336 = n5335 ^ n5299;
  assign n5294 = n5231 ^ n5185;
  assign n5295 = n5278 & ~n5294;
  assign n5296 = n5295 ^ n5277;
  assign n5337 = n5336 ^ n5296;
  assign n5407 = n5406 ^ n5337;
  assign n5291 = n5162 ^ n5158;
  assign n5292 = n5181 & n5291;
  assign n5293 = n5292 ^ n5180;
  assign n5408 = n5407 ^ n5293;
  assign n5288 = n5182 ^ n5154;
  assign n5289 = n5280 & ~n5288;
  assign n5290 = n5289 ^ n5279;
  assign n5409 = n5408 ^ n5290;
  assign n5414 = n5413 ^ n5409;
  assign n5536 = n5290 & ~n5408;
  assign n5537 = ~n5290 & n5408;
  assign n5538 = ~n5413 & ~n5537;
  assign n5539 = ~n5536 & ~n5538;
  assign n5522 = x27 & n1223;
  assign n5523 = x26 & n1227;
  assign n5524 = ~n5522 & ~n5523;
  assign n5525 = ~x27 & n1230;
  assign n5526 = ~x26 & n1232;
  assign n5527 = ~n5525 & ~n5526;
  assign n5528 = n5524 & n5527;
  assign n5520 = ~n650 & ~n654;
  assign n5513 = ~x31 & n821;
  assign n5514 = ~x30 & n823;
  assign n5515 = ~n5513 & ~n5514;
  assign n5516 = x31 & n814;
  assign n5517 = x30 & n818;
  assign n5518 = ~n5516 & ~n5517;
  assign n5519 = n5515 & n5518;
  assign n5521 = n5520 ^ n5519;
  assign n5529 = n5528 ^ n5521;
  assign n5504 = ~x25 & n1571;
  assign n5505 = ~x24 & n1575;
  assign n5506 = ~n5504 & ~n5505;
  assign n5507 = x25 & n1578;
  assign n5508 = x24 & n1580;
  assign n5509 = ~n5507 & ~n5508;
  assign n5510 = n5506 & n5509;
  assign n5496 = x19 & n2379;
  assign n5497 = x18 & n2383;
  assign n5498 = ~n5496 & ~n5497;
  assign n5499 = ~x19 & n2386;
  assign n5500 = ~x18 & n2388;
  assign n5501 = ~n5499 & ~n5500;
  assign n5502 = n5498 & n5501;
  assign n5489 = ~x17 & n2799;
  assign n5490 = ~x16 & n2803;
  assign n5491 = ~n5489 & ~n5490;
  assign n5492 = x17 & n2806;
  assign n5493 = x16 & n2808;
  assign n5494 = ~n5492 & ~n5493;
  assign n5495 = n5491 & n5494;
  assign n5503 = n5502 ^ n5495;
  assign n5511 = n5510 ^ n5503;
  assign n5481 = ~x29 & n1004;
  assign n5482 = ~x28 & n1008;
  assign n5483 = ~n5481 & ~n5482;
  assign n5484 = x29 & n1011;
  assign n5485 = x28 & n1013;
  assign n5486 = ~n5484 & ~n5485;
  assign n5487 = n5483 & n5486;
  assign n5479 = x13 & x63;
  assign n5472 = x15 & n3136;
  assign n5473 = x14 & n3138;
  assign n5474 = ~n5472 & ~n5473;
  assign n5475 = ~x15 & n3129;
  assign n5476 = ~x14 & n3133;
  assign n5477 = ~n5475 & ~n5476;
  assign n5478 = n5474 & n5477;
  assign n5480 = n5479 ^ n5478;
  assign n5488 = n5487 ^ n5480;
  assign n5512 = n5511 ^ n5488;
  assign n5530 = n5529 ^ n5512;
  assign n5465 = n5379 ^ n5371;
  assign n5466 = n5379 ^ n5368;
  assign n5467 = n5465 & ~n5466;
  assign n5468 = n5467 ^ n5371;
  assign n5461 = n5403 ^ n5395;
  assign n5462 = n5403 ^ n5388;
  assign n5463 = n5461 & ~n5462;
  assign n5464 = n5463 ^ n5395;
  assign n5469 = n5468 ^ n5464;
  assign n5458 = n5360 ^ n5358;
  assign n5459 = ~n5359 & ~n5458;
  assign n5460 = n5459 ^ n5360;
  assign n5470 = n5469 ^ n5460;
  assign n5454 = n5404 ^ n5380;
  assign n5455 = n5404 ^ n5361;
  assign n5456 = n5454 & n5455;
  assign n5457 = n5456 ^ n5380;
  assign n5471 = n5470 ^ n5457;
  assign n5531 = n5530 ^ n5471;
  assign n5442 = ~x21 & n2161;
  assign n5443 = ~x20 & n2165;
  assign n5444 = ~n5442 & ~n5443;
  assign n5445 = x21 & n2168;
  assign n5446 = x20 & n2170;
  assign n5447 = ~n5445 & ~n5446;
  assign n5448 = n5444 & n5447;
  assign n5435 = x23 & n1842;
  assign n5436 = x22 & n1844;
  assign n5437 = ~n5435 & ~n5436;
  assign n5438 = ~x23 & n1835;
  assign n5439 = ~x22 & n1839;
  assign n5440 = ~n5438 & ~n5439;
  assign n5441 = n5437 & n5440;
  assign n5449 = n5448 ^ n5441;
  assign n5450 = n5449 ^ n5320;
  assign n5431 = n5332 ^ n5326;
  assign n5432 = n5329 ^ n5326;
  assign n5433 = ~n5431 & n5432;
  assign n5434 = n5433 ^ n5332;
  assign n5451 = n5450 ^ n5434;
  assign n5428 = n5313 ^ n5306;
  assign n5429 = ~n5321 & ~n5428;
  assign n5430 = n5429 ^ n5320;
  assign n5452 = n5451 ^ n5430;
  assign n5424 = n5334 ^ n5322;
  assign n5425 = n5334 ^ n5302;
  assign n5426 = ~n5424 & ~n5425;
  assign n5427 = n5426 ^ n5322;
  assign n5453 = n5452 ^ n5427;
  assign n5532 = n5531 ^ n5453;
  assign n5421 = n5405 ^ n5343;
  assign n5422 = ~n5344 & n5421;
  assign n5423 = n5422 ^ n5405;
  assign n5533 = n5532 ^ n5423;
  assign n5418 = n5299 ^ n5296;
  assign n5419 = n5336 & ~n5418;
  assign n5420 = n5419 ^ n5335;
  assign n5534 = n5533 ^ n5420;
  assign n5415 = n5337 ^ n5293;
  assign n5416 = n5407 & n5415;
  assign n5417 = n5416 ^ n5406;
  assign n5535 = n5534 ^ n5417;
  assign n5540 = n5539 ^ n5535;
  assign n5653 = n5417 & ~n5534;
  assign n5654 = ~n5417 & n5534;
  assign n5655 = ~n5539 & ~n5654;
  assign n5656 = ~n5653 & ~n5655;
  assign n5640 = ~x24 & n1835;
  assign n5641 = ~x23 & n1839;
  assign n5642 = ~n5640 & ~n5641;
  assign n5643 = x24 & n1842;
  assign n5644 = x23 & n1844;
  assign n5645 = ~n5643 & ~n5644;
  assign n5646 = n5642 & n5645;
  assign n5638 = x14 & x63;
  assign n5631 = ~x30 & n1004;
  assign n5632 = ~x29 & n1008;
  assign n5633 = ~n5631 & ~n5632;
  assign n5634 = x30 & n1011;
  assign n5635 = x29 & n1013;
  assign n5636 = ~n5634 & ~n5635;
  assign n5637 = n5633 & n5636;
  assign n5639 = n5638 ^ n5637;
  assign n5647 = n5646 ^ n5639;
  assign n5622 = ~x16 & n3129;
  assign n5623 = ~x15 & n3133;
  assign n5624 = ~n5622 & ~n5623;
  assign n5625 = x16 & n3136;
  assign n5626 = x15 & n3138;
  assign n5627 = ~n5625 & ~n5626;
  assign n5628 = n5624 & n5627;
  assign n5614 = ~x26 & n1571;
  assign n5615 = ~x25 & n1575;
  assign n5616 = ~n5614 & ~n5615;
  assign n5617 = x26 & n1578;
  assign n5618 = x25 & n1580;
  assign n5619 = ~n5617 & ~n5618;
  assign n5620 = n5616 & n5619;
  assign n5607 = ~x18 & n2799;
  assign n5608 = ~x17 & n2803;
  assign n5609 = ~n5607 & ~n5608;
  assign n5610 = x18 & n2806;
  assign n5611 = x17 & n2808;
  assign n5612 = ~n5610 & ~n5611;
  assign n5613 = n5609 & n5612;
  assign n5621 = n5620 ^ n5613;
  assign n5629 = n5628 ^ n5621;
  assign n5603 = n5487 ^ n5479;
  assign n5604 = n5487 ^ n5478;
  assign n5605 = ~n5603 & ~n5604;
  assign n5606 = n5605 ^ n5479;
  assign n5630 = n5629 ^ n5606;
  assign n5648 = n5647 ^ n5630;
  assign n5597 = x47 ^ x31;
  assign n5598 = n817 & n5597;
  assign n5599 = ~n821 & ~n5598;
  assign n5594 = n5528 ^ n5519;
  assign n5595 = ~n5521 & ~n5594;
  assign n5596 = n5595 ^ n5520;
  assign n5600 = n5599 ^ n5596;
  assign n5591 = n5510 ^ n5502;
  assign n5592 = ~n5503 & n5591;
  assign n5593 = n5592 ^ n5510;
  assign n5601 = n5600 ^ n5593;
  assign n5588 = n5529 ^ n5511;
  assign n5589 = n5512 & ~n5588;
  assign n5590 = n5589 ^ n5529;
  assign n5602 = n5601 ^ n5590;
  assign n5649 = n5648 ^ n5602;
  assign n5576 = x20 & n2379;
  assign n5577 = x19 & n2383;
  assign n5578 = ~n5576 & ~n5577;
  assign n5579 = ~x20 & n2386;
  assign n5580 = ~x19 & n2388;
  assign n5581 = ~n5579 & ~n5580;
  assign n5582 = n5578 & n5581;
  assign n5568 = ~x22 & n2161;
  assign n5569 = ~x21 & n2165;
  assign n5570 = ~n5568 & ~n5569;
  assign n5571 = x22 & n2168;
  assign n5572 = x21 & n2170;
  assign n5573 = ~n5571 & ~n5572;
  assign n5574 = n5570 & n5573;
  assign n5561 = ~x28 & n1230;
  assign n5562 = ~x27 & n1232;
  assign n5563 = ~n5561 & ~n5562;
  assign n5564 = x28 & n1223;
  assign n5565 = x27 & n1227;
  assign n5566 = ~n5564 & ~n5565;
  assign n5567 = n5563 & n5566;
  assign n5575 = n5574 ^ n5567;
  assign n5583 = n5582 ^ n5575;
  assign n5557 = n5448 ^ n5320;
  assign n5558 = n5441 ^ n5320;
  assign n5559 = n5557 & ~n5558;
  assign n5560 = n5559 ^ n5448;
  assign n5584 = n5583 ^ n5560;
  assign n5554 = n5464 ^ n5460;
  assign n5555 = n5469 & n5554;
  assign n5556 = n5555 ^ n5468;
  assign n5585 = n5584 ^ n5556;
  assign n5550 = n5450 ^ n5430;
  assign n5551 = n5434 ^ n5430;
  assign n5552 = ~n5550 & ~n5551;
  assign n5553 = n5552 ^ n5450;
  assign n5586 = n5585 ^ n5553;
  assign n5547 = n5530 ^ n5457;
  assign n5548 = n5471 & n5547;
  assign n5549 = n5548 ^ n5530;
  assign n5587 = n5586 ^ n5549;
  assign n5650 = n5649 ^ n5587;
  assign n5544 = n5531 ^ n5452;
  assign n5545 = n5453 & ~n5544;
  assign n5546 = n5545 ^ n5531;
  assign n5651 = n5650 ^ n5546;
  assign n5541 = n5423 ^ n5420;
  assign n5542 = ~n5533 & ~n5541;
  assign n5543 = n5542 ^ n5532;
  assign n5652 = n5651 ^ n5543;
  assign n5657 = n5656 ^ n5652;
  assign n5765 = ~n5543 & ~n5651;
  assign n5766 = n5543 & n5651;
  assign n5767 = ~n5656 & ~n5766;
  assign n5768 = ~n5765 & ~n5767;
  assign n5752 = ~x23 & n2161;
  assign n5753 = ~x22 & n2165;
  assign n5754 = ~n5752 & ~n5753;
  assign n5755 = x23 & n2168;
  assign n5756 = x22 & n2170;
  assign n5757 = ~n5755 & ~n5756;
  assign n5758 = n5754 & n5757;
  assign n5750 = x15 & x63;
  assign n5743 = x29 & n1223;
  assign n5744 = x28 & n1227;
  assign n5745 = ~n5743 & ~n5744;
  assign n5746 = ~x29 & n1230;
  assign n5747 = ~x28 & n1232;
  assign n5748 = ~n5746 & ~n5747;
  assign n5749 = n5745 & n5748;
  assign n5751 = n5750 ^ n5749;
  assign n5759 = n5758 ^ n5751;
  assign n5739 = n5646 ^ n5637;
  assign n5740 = ~n5639 & ~n5739;
  assign n5741 = n5740 ^ n5638;
  assign n5735 = n5582 ^ n5574;
  assign n5736 = n5582 ^ n5567;
  assign n5737 = n5735 & ~n5736;
  assign n5738 = n5737 ^ n5574;
  assign n5742 = n5741 ^ n5738;
  assign n5760 = n5759 ^ n5742;
  assign n5731 = n5647 ^ n5629;
  assign n5732 = n5630 & ~n5731;
  assign n5733 = n5732 ^ n5647;
  assign n5727 = n5599 ^ n5593;
  assign n5728 = n5596 ^ n5593;
  assign n5729 = ~n5727 & n5728;
  assign n5730 = n5729 ^ n5599;
  assign n5734 = n5733 ^ n5730;
  assign n5761 = n5760 ^ n5734;
  assign n5715 = ~x27 & n1571;
  assign n5716 = ~x26 & n1575;
  assign n5717 = ~n5715 & ~n5716;
  assign n5718 = x27 & n1578;
  assign n5719 = x26 & n1580;
  assign n5720 = ~n5718 & ~n5719;
  assign n5721 = n5717 & n5720;
  assign n5713 = ~n821 & ~n823;
  assign n5706 = ~x31 & n1004;
  assign n5707 = ~x30 & n1008;
  assign n5708 = ~n5706 & ~n5707;
  assign n5709 = x31 & n1011;
  assign n5710 = x30 & n1013;
  assign n5711 = ~n5709 & ~n5710;
  assign n5712 = n5708 & n5711;
  assign n5714 = n5713 ^ n5712;
  assign n5722 = n5721 ^ n5714;
  assign n5698 = x25 & n1842;
  assign n5699 = x24 & n1844;
  assign n5700 = ~n5698 & ~n5699;
  assign n5701 = ~x25 & n1835;
  assign n5702 = ~x24 & n1839;
  assign n5703 = ~n5701 & ~n5702;
  assign n5704 = n5700 & n5703;
  assign n5690 = ~x19 & n2799;
  assign n5691 = ~x18 & n2803;
  assign n5692 = ~n5690 & ~n5691;
  assign n5693 = x19 & n2806;
  assign n5694 = x18 & n2808;
  assign n5695 = ~n5693 & ~n5694;
  assign n5696 = n5692 & n5695;
  assign n5683 = ~x17 & n3129;
  assign n5684 = ~x16 & n3133;
  assign n5685 = ~n5683 & ~n5684;
  assign n5686 = x17 & n3136;
  assign n5687 = x16 & n3138;
  assign n5688 = ~n5686 & ~n5687;
  assign n5689 = n5685 & n5688;
  assign n5697 = n5696 ^ n5689;
  assign n5705 = n5704 ^ n5697;
  assign n5723 = n5722 ^ n5705;
  assign n5674 = x21 & n2379;
  assign n5675 = x20 & n2383;
  assign n5676 = ~n5674 & ~n5675;
  assign n5677 = ~x21 & n2386;
  assign n5678 = ~x20 & n2388;
  assign n5679 = ~n5677 & ~n5678;
  assign n5680 = n5676 & n5679;
  assign n5681 = n5680 ^ n5599;
  assign n5671 = n5628 ^ n5613;
  assign n5672 = n5621 & ~n5671;
  assign n5673 = n5672 ^ n5620;
  assign n5682 = n5681 ^ n5673;
  assign n5724 = n5723 ^ n5682;
  assign n5668 = n5560 ^ n5556;
  assign n5669 = n5584 & ~n5668;
  assign n5670 = n5669 ^ n5583;
  assign n5725 = n5724 ^ n5670;
  assign n5665 = n5648 ^ n5601;
  assign n5666 = n5602 & n5665;
  assign n5667 = n5666 ^ n5648;
  assign n5726 = n5725 ^ n5667;
  assign n5762 = n5761 ^ n5726;
  assign n5661 = n5585 ^ n5549;
  assign n5662 = n5553 ^ n5549;
  assign n5663 = n5661 & ~n5662;
  assign n5664 = n5663 ^ n5585;
  assign n5763 = n5762 ^ n5664;
  assign n5658 = n5587 ^ n5546;
  assign n5659 = ~n5650 & n5658;
  assign n5660 = n5659 ^ n5649;
  assign n5764 = n5763 ^ n5660;
  assign n5769 = n5768 ^ n5764;
  assign n5868 = n5660 & n5763;
  assign n5869 = ~n5660 & ~n5763;
  assign n5870 = ~n5768 & ~n5869;
  assign n5871 = ~n5868 & ~n5870;
  assign n5859 = n5721 ^ n5712;
  assign n5860 = ~n5714 & ~n5859;
  assign n5861 = n5860 ^ n5713;
  assign n5856 = n5704 ^ n5689;
  assign n5857 = n5697 & ~n5856;
  assign n5858 = n5857 ^ n5696;
  assign n5862 = n5861 ^ n5858;
  assign n5853 = n5758 ^ n5749;
  assign n5854 = ~n5751 & ~n5853;
  assign n5855 = n5854 ^ n5750;
  assign n5863 = n5862 ^ n5855;
  assign n5849 = n5680 ^ n5673;
  assign n5850 = n5681 & ~n5849;
  assign n5851 = n5850 ^ n5599;
  assign n5846 = n5759 ^ n5741;
  assign n5847 = n5742 & n5846;
  assign n5848 = n5847 ^ n5759;
  assign n5852 = n5851 ^ n5848;
  assign n5864 = n5863 ^ n5852;
  assign n5839 = x49 ^ x31;
  assign n5840 = n1007 & n5839;
  assign n5841 = ~n1004 & ~n5840;
  assign n5831 = ~x20 & n2799;
  assign n5832 = ~x19 & n2803;
  assign n5833 = ~n5831 & ~n5832;
  assign n5834 = x20 & n2806;
  assign n5835 = x19 & n2808;
  assign n5836 = ~n5834 & ~n5835;
  assign n5837 = n5833 & n5836;
  assign n5824 = ~x22 & n2386;
  assign n5825 = ~x21 & n2388;
  assign n5826 = ~n5824 & ~n5825;
  assign n5827 = x22 & n2379;
  assign n5828 = x21 & n2383;
  assign n5829 = ~n5827 & ~n5828;
  assign n5830 = n5826 & n5829;
  assign n5838 = n5837 ^ n5830;
  assign n5842 = n5841 ^ n5838;
  assign n5815 = x28 & n1578;
  assign n5816 = x27 & n1580;
  assign n5817 = ~n5815 & ~n5816;
  assign n5818 = ~x28 & n1571;
  assign n5819 = ~x27 & n1575;
  assign n5820 = ~n5818 & ~n5819;
  assign n5821 = n5817 & n5820;
  assign n5807 = x24 & n2168;
  assign n5808 = x23 & n2170;
  assign n5809 = ~n5807 & ~n5808;
  assign n5810 = ~x24 & n2161;
  assign n5811 = ~x23 & n2165;
  assign n5812 = ~n5810 & ~n5811;
  assign n5813 = n5809 & n5812;
  assign n5800 = x30 & n1223;
  assign n5801 = x29 & n1227;
  assign n5802 = ~n5800 & ~n5801;
  assign n5803 = ~x30 & n1230;
  assign n5804 = ~x29 & n1232;
  assign n5805 = ~n5803 & ~n5804;
  assign n5806 = n5802 & n5805;
  assign n5814 = n5813 ^ n5806;
  assign n5822 = n5821 ^ n5814;
  assign n5798 = x16 & x63;
  assign n5790 = ~x18 & n3129;
  assign n5791 = ~x17 & n3133;
  assign n5792 = ~n5790 & ~n5791;
  assign n5793 = x18 & n3136;
  assign n5794 = x17 & n3138;
  assign n5795 = ~n5793 & ~n5794;
  assign n5796 = n5792 & n5795;
  assign n5783 = x26 & n1842;
  assign n5784 = x25 & n1844;
  assign n5785 = ~n5783 & ~n5784;
  assign n5786 = ~x26 & n1835;
  assign n5787 = ~x25 & n1839;
  assign n5788 = ~n5786 & ~n5787;
  assign n5789 = n5785 & n5788;
  assign n5797 = n5796 ^ n5789;
  assign n5799 = n5798 ^ n5797;
  assign n5823 = n5822 ^ n5799;
  assign n5843 = n5842 ^ n5823;
  assign n5780 = n5705 ^ n5682;
  assign n5781 = ~n5723 & ~n5780;
  assign n5782 = n5781 ^ n5722;
  assign n5844 = n5843 ^ n5782;
  assign n5777 = n5760 ^ n5733;
  assign n5778 = ~n5734 & ~n5777;
  assign n5779 = n5778 ^ n5760;
  assign n5845 = n5844 ^ n5779;
  assign n5865 = n5864 ^ n5845;
  assign n5773 = n5724 ^ n5667;
  assign n5774 = n5670 ^ n5667;
  assign n5775 = ~n5773 & ~n5774;
  assign n5776 = n5775 ^ n5724;
  assign n5866 = n5865 ^ n5776;
  assign n5770 = n5726 ^ n5664;
  assign n5771 = ~n5762 & n5770;
  assign n5772 = n5771 ^ n5761;
  assign n5867 = n5866 ^ n5772;
  assign n5872 = n5871 ^ n5867;
  assign n5965 = ~n5772 & n5866;
  assign n5966 = n5772 & ~n5866;
  assign n5967 = ~n5871 & ~n5966;
  assign n5968 = ~n5965 & ~n5967;
  assign n5956 = n5798 ^ n5796;
  assign n5957 = ~n5797 & ~n5956;
  assign n5958 = n5957 ^ n5798;
  assign n5959 = n5958 ^ n5841;
  assign n5953 = n5821 ^ n5806;
  assign n5954 = n5814 & ~n5953;
  assign n5955 = n5954 ^ n5813;
  assign n5960 = n5959 ^ n5955;
  assign n5949 = n5841 ^ n5837;
  assign n5950 = ~n5838 & ~n5949;
  assign n5951 = n5950 ^ n5841;
  assign n5946 = n5861 ^ n5855;
  assign n5947 = n5862 & n5946;
  assign n5948 = n5947 ^ n5855;
  assign n5952 = n5951 ^ n5948;
  assign n5961 = n5960 ^ n5952;
  assign n5935 = ~x25 & n2161;
  assign n5936 = ~x24 & n2165;
  assign n5937 = ~n5935 & ~n5936;
  assign n5938 = x25 & n2168;
  assign n5939 = x24 & n2170;
  assign n5940 = ~n5938 & ~n5939;
  assign n5941 = n5937 & n5940;
  assign n5933 = x17 & x63;
  assign n5926 = x19 & n3136;
  assign n5927 = x18 & n3138;
  assign n5928 = ~n5926 & ~n5927;
  assign n5929 = ~x19 & n3129;
  assign n5930 = ~x18 & n3133;
  assign n5931 = ~n5929 & ~n5930;
  assign n5932 = n5928 & n5931;
  assign n5934 = n5933 ^ n5932;
  assign n5942 = n5941 ^ n5934;
  assign n5917 = x21 & n2806;
  assign n5918 = x20 & n2808;
  assign n5919 = ~n5917 & ~n5918;
  assign n5920 = ~x21 & n2799;
  assign n5921 = ~x20 & n2803;
  assign n5922 = ~n5920 & ~n5921;
  assign n5923 = n5919 & n5922;
  assign n5909 = ~x29 & n1571;
  assign n5910 = ~x28 & n1575;
  assign n5911 = ~n5909 & ~n5910;
  assign n5912 = x29 & n1578;
  assign n5913 = x28 & n1580;
  assign n5914 = ~n5912 & ~n5913;
  assign n5915 = n5911 & n5914;
  assign n5902 = ~x23 & n2386;
  assign n5903 = ~x22 & n2388;
  assign n5904 = ~n5902 & ~n5903;
  assign n5905 = x23 & n2379;
  assign n5906 = x22 & n2383;
  assign n5907 = ~n5905 & ~n5906;
  assign n5908 = n5904 & n5907;
  assign n5916 = n5915 ^ n5908;
  assign n5924 = n5923 ^ n5916;
  assign n5894 = ~x27 & n1835;
  assign n5895 = ~x26 & n1839;
  assign n5896 = ~n5894 & ~n5895;
  assign n5897 = x27 & n1842;
  assign n5898 = x26 & n1844;
  assign n5899 = ~n5897 & ~n5898;
  assign n5900 = n5896 & n5899;
  assign n5892 = ~n1004 & ~n1008;
  assign n5885 = ~x31 & n1230;
  assign n5886 = ~x30 & n1232;
  assign n5887 = ~n5885 & ~n5886;
  assign n5888 = x31 & n1223;
  assign n5889 = x30 & n1227;
  assign n5890 = ~n5888 & ~n5889;
  assign n5891 = n5887 & n5890;
  assign n5893 = n5892 ^ n5891;
  assign n5901 = n5900 ^ n5893;
  assign n5925 = n5924 ^ n5901;
  assign n5943 = n5942 ^ n5925;
  assign n5882 = n5842 ^ n5822;
  assign n5883 = n5823 & ~n5882;
  assign n5884 = n5883 ^ n5842;
  assign n5944 = n5943 ^ n5884;
  assign n5879 = n5863 ^ n5851;
  assign n5880 = n5852 & n5879;
  assign n5881 = n5880 ^ n5863;
  assign n5945 = n5944 ^ n5881;
  assign n5962 = n5961 ^ n5945;
  assign n5876 = n5782 ^ n5779;
  assign n5877 = ~n5844 & n5876;
  assign n5878 = n5877 ^ n5843;
  assign n5963 = n5962 ^ n5878;
  assign n5873 = n5845 ^ n5776;
  assign n5874 = n5865 & ~n5873;
  assign n5875 = n5874 ^ n5864;
  assign n5964 = n5963 ^ n5875;
  assign n5969 = n5968 ^ n5964;
  assign n6058 = n5875 & ~n5963;
  assign n6059 = ~n5875 & n5963;
  assign n6060 = ~n5968 & ~n6059;
  assign n6061 = ~n6058 & ~n6060;
  assign n6044 = ~x22 & n2799;
  assign n6045 = ~x21 & n2803;
  assign n6046 = ~n6044 & ~n6045;
  assign n6047 = x22 & n2806;
  assign n6048 = x21 & n2808;
  assign n6049 = ~n6047 & ~n6048;
  assign n6050 = n6046 & n6049;
  assign n6036 = ~x24 & n2386;
  assign n6037 = ~x23 & n2388;
  assign n6038 = ~n6036 & ~n6037;
  assign n6039 = x24 & n2379;
  assign n6040 = x23 & n2383;
  assign n6041 = ~n6039 & ~n6040;
  assign n6042 = n6038 & n6041;
  assign n6029 = x28 & n1842;
  assign n6030 = x27 & n1844;
  assign n6031 = ~n6029 & ~n6030;
  assign n6032 = ~x28 & n1835;
  assign n6033 = ~x27 & n1839;
  assign n6034 = ~n6032 & ~n6033;
  assign n6035 = n6031 & n6034;
  assign n6043 = n6042 ^ n6035;
  assign n6051 = n6050 ^ n6043;
  assign n6024 = n5941 ^ n5933;
  assign n6025 = n5941 ^ n5932;
  assign n6026 = ~n6024 & ~n6025;
  assign n6027 = n6026 ^ n5933;
  assign n6021 = n5923 ^ n5908;
  assign n6022 = n5916 & ~n6021;
  assign n6023 = n6022 ^ n5915;
  assign n6028 = n6027 ^ n6023;
  assign n6052 = n6051 ^ n6028;
  assign n6018 = n5942 ^ n5901;
  assign n6019 = ~n5925 & ~n6018;
  assign n6020 = n6019 ^ n5924;
  assign n6053 = n6052 ^ n6020;
  assign n6008 = x26 & n2168;
  assign n6009 = x25 & n2170;
  assign n6010 = ~n6008 & ~n6009;
  assign n6011 = ~x26 & n2161;
  assign n6012 = ~x25 & n2165;
  assign n6013 = ~n6011 & ~n6012;
  assign n6014 = n6010 & n6013;
  assign n6006 = x18 & x63;
  assign n5999 = ~x30 & n1571;
  assign n6000 = ~x29 & n1575;
  assign n6001 = ~n5999 & ~n6000;
  assign n6002 = x30 & n1578;
  assign n6003 = x29 & n1580;
  assign n6004 = ~n6002 & ~n6003;
  assign n6005 = n6001 & n6004;
  assign n6007 = n6006 ^ n6005;
  assign n6015 = n6014 ^ n6007;
  assign n5994 = x51 ^ x31;
  assign n5995 = n1226 & n5994;
  assign n5996 = ~n1230 & ~n5995;
  assign n5987 = x20 & n3136;
  assign n5988 = x19 & n3138;
  assign n5989 = ~n5987 & ~n5988;
  assign n5990 = ~x20 & n3129;
  assign n5991 = ~x19 & n3133;
  assign n5992 = ~n5990 & ~n5991;
  assign n5993 = n5989 & n5992;
  assign n5997 = n5996 ^ n5993;
  assign n5983 = n5900 ^ n5892;
  assign n5984 = n5900 ^ n5891;
  assign n5985 = ~n5983 & ~n5984;
  assign n5986 = n5985 ^ n5892;
  assign n5998 = n5997 ^ n5986;
  assign n6016 = n6015 ^ n5998;
  assign n5980 = n5958 ^ n5955;
  assign n5981 = ~n5959 & n5980;
  assign n5982 = n5981 ^ n5841;
  assign n6017 = n6016 ^ n5982;
  assign n6054 = n6053 ^ n6017;
  assign n5976 = n5960 ^ n5951;
  assign n5977 = n5960 ^ n5948;
  assign n5978 = n5976 & ~n5977;
  assign n5979 = n5978 ^ n5951;
  assign n6055 = n6054 ^ n5979;
  assign n5973 = n5884 ^ n5881;
  assign n5974 = ~n5944 & n5973;
  assign n5975 = n5974 ^ n5943;
  assign n6056 = n6055 ^ n5975;
  assign n5970 = n5945 ^ n5878;
  assign n5971 = n5962 & n5970;
  assign n5972 = n5971 ^ n5961;
  assign n6057 = n6056 ^ n5972;
  assign n6062 = n6061 ^ n6057;
  assign n6143 = n5972 & n6056;
  assign n6144 = ~n5972 & ~n6056;
  assign n6145 = ~n6061 & ~n6144;
  assign n6146 = ~n6143 & ~n6145;
  assign n6129 = x23 & n2806;
  assign n6130 = x22 & n2808;
  assign n6131 = ~n6129 & ~n6130;
  assign n6132 = ~x23 & n2799;
  assign n6133 = ~x22 & n2803;
  assign n6134 = ~n6132 & ~n6133;
  assign n6135 = n6131 & n6134;
  assign n6122 = ~x21 & n3129;
  assign n6123 = ~x20 & n3133;
  assign n6124 = ~n6122 & ~n6123;
  assign n6125 = x21 & n3136;
  assign n6126 = x20 & n3138;
  assign n6127 = ~n6125 & ~n6126;
  assign n6128 = n6124 & n6127;
  assign n6136 = n6135 ^ n6128;
  assign n6137 = n6136 ^ n5996;
  assign n6114 = ~x29 & n1835;
  assign n6115 = ~x28 & n1839;
  assign n6116 = ~n6114 & ~n6115;
  assign n6117 = x29 & n1842;
  assign n6118 = x28 & n1844;
  assign n6119 = ~n6117 & ~n6118;
  assign n6120 = n6116 & n6119;
  assign n6112 = x19 & x63;
  assign n6105 = ~x25 & n2386;
  assign n6106 = ~x24 & n2388;
  assign n6107 = ~n6105 & ~n6106;
  assign n6108 = x25 & n2379;
  assign n6109 = x24 & n2383;
  assign n6110 = ~n6108 & ~n6109;
  assign n6111 = n6107 & n6110;
  assign n6113 = n6112 ^ n6111;
  assign n6121 = n6120 ^ n6113;
  assign n6138 = n6137 ^ n6121;
  assign n6102 = n5993 ^ n5986;
  assign n6103 = ~n5997 & n6102;
  assign n6104 = n6103 ^ n5996;
  assign n6139 = n6138 ^ n6104;
  assign n6091 = ~x27 & n2161;
  assign n6092 = ~x26 & n2165;
  assign n6093 = ~n6091 & ~n6092;
  assign n6094 = x27 & n2168;
  assign n6095 = x26 & n2170;
  assign n6096 = ~n6094 & ~n6095;
  assign n6097 = n6093 & n6096;
  assign n6089 = ~n1230 & ~n1232;
  assign n6082 = ~x31 & n1571;
  assign n6083 = ~x30 & n1575;
  assign n6084 = ~n6082 & ~n6083;
  assign n6085 = x31 & n1578;
  assign n6086 = x30 & n1580;
  assign n6087 = ~n6085 & ~n6086;
  assign n6088 = n6084 & n6087;
  assign n6090 = n6089 ^ n6088;
  assign n6098 = n6097 ^ n6090;
  assign n6078 = n6014 ^ n6005;
  assign n6079 = ~n6007 & ~n6078;
  assign n6080 = n6079 ^ n6006;
  assign n6075 = n6050 ^ n6042;
  assign n6076 = ~n6043 & n6075;
  assign n6077 = n6076 ^ n6050;
  assign n6081 = n6080 ^ n6077;
  assign n6099 = n6098 ^ n6081;
  assign n6072 = n6051 ^ n6027;
  assign n6073 = n6028 & ~n6072;
  assign n6074 = n6073 ^ n6051;
  assign n6100 = n6099 ^ n6074;
  assign n6069 = n5998 ^ n5982;
  assign n6070 = ~n6016 & ~n6069;
  assign n6071 = n6070 ^ n6015;
  assign n6101 = n6100 ^ n6071;
  assign n6140 = n6139 ^ n6101;
  assign n6066 = n6020 ^ n6017;
  assign n6067 = ~n6053 & n6066;
  assign n6068 = n6067 ^ n6052;
  assign n6141 = n6140 ^ n6068;
  assign n6063 = n5979 ^ n5975;
  assign n6064 = ~n6055 & n6063;
  assign n6065 = n6064 ^ n6054;
  assign n6142 = n6141 ^ n6065;
  assign n6147 = n6146 ^ n6142;
  assign n6222 = ~n6065 & ~n6141;
  assign n6223 = n6065 & n6141;
  assign n6224 = ~n6146 & ~n6223;
  assign n6225 = ~n6222 & ~n6224;
  assign n6214 = x20 & x63;
  assign n6206 = ~x28 & n2161;
  assign n6207 = ~x27 & n2165;
  assign n6208 = ~n6206 & ~n6207;
  assign n6209 = x28 & n2168;
  assign n6210 = x27 & n2170;
  assign n6211 = ~n6209 & ~n6210;
  assign n6212 = n6208 & n6211;
  assign n6199 = ~x22 & n3129;
  assign n6200 = ~x21 & n3133;
  assign n6201 = ~n6199 & ~n6200;
  assign n6202 = x22 & n3136;
  assign n6203 = x21 & n3138;
  assign n6204 = ~n6202 & ~n6203;
  assign n6205 = n6201 & n6204;
  assign n6213 = n6212 ^ n6205;
  assign n6215 = n6214 ^ n6213;
  assign n6191 = ~x24 & n2799;
  assign n6192 = ~x23 & n2803;
  assign n6193 = ~n6191 & ~n6192;
  assign n6194 = x24 & n2806;
  assign n6195 = x23 & n2808;
  assign n6196 = ~n6194 & ~n6195;
  assign n6197 = n6193 & n6196;
  assign n6183 = ~x30 & n1835;
  assign n6184 = ~x29 & n1839;
  assign n6185 = ~n6183 & ~n6184;
  assign n6186 = x30 & n1842;
  assign n6187 = x29 & n1844;
  assign n6188 = ~n6186 & ~n6187;
  assign n6189 = n6185 & n6188;
  assign n6176 = x26 & n2379;
  assign n6177 = x25 & n2383;
  assign n6178 = ~n6176 & ~n6177;
  assign n6179 = ~x26 & n2386;
  assign n6180 = ~x25 & n2388;
  assign n6181 = ~n6179 & ~n6180;
  assign n6182 = n6178 & n6181;
  assign n6190 = n6189 ^ n6182;
  assign n6198 = n6197 ^ n6190;
  assign n6216 = n6215 ^ n6198;
  assign n6173 = n6135 ^ n5996;
  assign n6174 = ~n6136 & n6173;
  assign n6175 = n6174 ^ n5996;
  assign n6217 = n6216 ^ n6175;
  assign n6167 = x53 ^ x31;
  assign n6168 = n1574 & n6167;
  assign n6169 = ~n1571 & ~n6168;
  assign n6164 = n6097 ^ n6088;
  assign n6165 = ~n6090 & ~n6164;
  assign n6166 = n6165 ^ n6089;
  assign n6170 = n6169 ^ n6166;
  assign n6161 = n6120 ^ n6111;
  assign n6162 = ~n6113 & ~n6161;
  assign n6163 = n6162 ^ n6112;
  assign n6171 = n6170 ^ n6163;
  assign n6158 = n6098 ^ n6080;
  assign n6159 = n6081 & n6158;
  assign n6160 = n6159 ^ n6098;
  assign n6172 = n6171 ^ n6160;
  assign n6218 = n6217 ^ n6172;
  assign n6155 = n6121 ^ n6104;
  assign n6156 = ~n6138 & ~n6155;
  assign n6157 = n6156 ^ n6137;
  assign n6219 = n6218 ^ n6157;
  assign n6152 = n6074 ^ n6071;
  assign n6153 = n6100 & n6152;
  assign n6154 = n6153 ^ n6099;
  assign n6220 = n6219 ^ n6154;
  assign n6148 = n6139 ^ n6068;
  assign n6149 = n6101 ^ n6068;
  assign n6150 = ~n6148 & ~n6149;
  assign n6151 = n6150 ^ n6139;
  assign n6221 = n6220 ^ n6151;
  assign n6226 = n6225 ^ n6221;
  assign n6296 = ~n6151 & n6220;
  assign n6297 = n6151 & ~n6220;
  assign n6298 = ~n6225 & ~n6297;
  assign n6299 = ~n6296 & ~n6298;
  assign n6284 = ~x27 & n2386;
  assign n6285 = ~x26 & n2388;
  assign n6286 = ~n6284 & ~n6285;
  assign n6287 = x27 & n2379;
  assign n6288 = x26 & n2383;
  assign n6289 = ~n6287 & ~n6288;
  assign n6290 = n6286 & n6289;
  assign n6282 = ~n1571 & ~n1575;
  assign n6275 = x31 & n1842;
  assign n6276 = x30 & n1844;
  assign n6277 = ~n6275 & ~n6276;
  assign n6278 = ~x31 & n1835;
  assign n6279 = ~x30 & n1839;
  assign n6280 = ~n6278 & ~n6279;
  assign n6281 = n6277 & n6280;
  assign n6283 = n6282 ^ n6281;
  assign n6291 = n6290 ^ n6283;
  assign n6266 = x23 & n3136;
  assign n6267 = x22 & n3138;
  assign n6268 = ~n6266 & ~n6267;
  assign n6269 = ~x23 & n3129;
  assign n6270 = ~x22 & n3133;
  assign n6271 = ~n6269 & ~n6270;
  assign n6272 = n6268 & n6271;
  assign n6258 = ~x25 & n2799;
  assign n6259 = ~x24 & n2803;
  assign n6260 = ~n6258 & ~n6259;
  assign n6261 = x25 & n2806;
  assign n6262 = x24 & n2808;
  assign n6263 = ~n6261 & ~n6262;
  assign n6264 = n6260 & n6263;
  assign n6251 = x29 & n2168;
  assign n6252 = x28 & n2170;
  assign n6253 = ~n6251 & ~n6252;
  assign n6254 = ~x29 & n2161;
  assign n6255 = ~x28 & n2165;
  assign n6256 = ~n6254 & ~n6255;
  assign n6257 = n6253 & n6256;
  assign n6265 = n6264 ^ n6257;
  assign n6273 = n6272 ^ n6265;
  assign n6248 = n6214 ^ n6212;
  assign n6249 = ~n6213 & ~n6248;
  assign n6250 = n6249 ^ n6214;
  assign n6274 = n6273 ^ n6250;
  assign n6292 = n6291 ^ n6274;
  assign n6243 = x21 & x63;
  assign n6244 = n6243 ^ n6169;
  assign n6240 = n6197 ^ n6182;
  assign n6241 = n6190 & ~n6240;
  assign n6242 = n6241 ^ n6189;
  assign n6245 = n6244 ^ n6242;
  assign n6236 = n6169 ^ n6163;
  assign n6237 = n6166 ^ n6163;
  assign n6238 = n6236 & ~n6237;
  assign n6239 = n6238 ^ n6169;
  assign n6246 = n6245 ^ n6239;
  assign n6233 = n6198 ^ n6175;
  assign n6234 = ~n6216 & ~n6233;
  assign n6235 = n6234 ^ n6215;
  assign n6247 = n6246 ^ n6235;
  assign n6293 = n6292 ^ n6247;
  assign n6230 = n6217 ^ n6171;
  assign n6231 = ~n6172 & n6230;
  assign n6232 = n6231 ^ n6217;
  assign n6294 = n6293 ^ n6232;
  assign n6227 = n6157 ^ n6154;
  assign n6228 = ~n6219 & ~n6227;
  assign n6229 = n6228 ^ n6218;
  assign n6295 = n6294 ^ n6229;
  assign n6300 = n6299 ^ n6295;
  assign n6365 = n6229 & ~n6294;
  assign n6366 = ~n6229 & n6294;
  assign n6367 = ~n6299 & ~n6366;
  assign n6368 = ~n6365 & ~n6367;
  assign n6357 = x55 ^ x31;
  assign n6358 = n1838 & n6357;
  assign n6359 = ~n1835 & ~n6358;
  assign n6349 = x24 & n3136;
  assign n6350 = x23 & n3138;
  assign n6351 = ~n6349 & ~n6350;
  assign n6352 = ~x24 & n3129;
  assign n6353 = ~x23 & n3133;
  assign n6354 = ~n6352 & ~n6353;
  assign n6355 = n6351 & n6354;
  assign n6342 = ~x26 & n2799;
  assign n6343 = ~x25 & n2803;
  assign n6344 = ~n6342 & ~n6343;
  assign n6345 = x26 & n2806;
  assign n6346 = x25 & n2808;
  assign n6347 = ~n6345 & ~n6346;
  assign n6348 = n6344 & n6347;
  assign n6356 = n6355 ^ n6348;
  assign n6360 = n6359 ^ n6356;
  assign n6338 = n6290 ^ n6281;
  assign n6339 = ~n6283 & ~n6338;
  assign n6340 = n6339 ^ n6282;
  assign n6334 = n6272 ^ n6264;
  assign n6335 = n6272 ^ n6257;
  assign n6336 = n6334 & ~n6335;
  assign n6337 = n6336 ^ n6264;
  assign n6341 = n6340 ^ n6337;
  assign n6361 = n6360 ^ n6341;
  assign n6324 = x30 & n2168;
  assign n6325 = x29 & n2170;
  assign n6326 = ~n6324 & ~n6325;
  assign n6327 = ~x30 & n2161;
  assign n6328 = ~x29 & n2165;
  assign n6329 = ~n6327 & ~n6328;
  assign n6330 = n6326 & n6329;
  assign n6322 = x22 & x63;
  assign n6315 = ~x28 & n2386;
  assign n6316 = ~x27 & n2388;
  assign n6317 = ~n6315 & ~n6316;
  assign n6318 = x28 & n2379;
  assign n6319 = x27 & n2383;
  assign n6320 = ~n6318 & ~n6319;
  assign n6321 = n6317 & n6320;
  assign n6323 = n6322 ^ n6321;
  assign n6331 = n6330 ^ n6323;
  assign n6312 = n6242 ^ n6169;
  assign n6313 = ~n6244 & ~n6312;
  assign n6314 = n6313 ^ n6243;
  assign n6332 = n6331 ^ n6314;
  assign n6308 = n6291 ^ n6273;
  assign n6309 = n6291 ^ n6250;
  assign n6310 = ~n6308 & ~n6309;
  assign n6311 = n6310 ^ n6273;
  assign n6333 = n6332 ^ n6311;
  assign n6362 = n6361 ^ n6333;
  assign n6304 = n6245 ^ n6235;
  assign n6305 = n6239 ^ n6235;
  assign n6306 = n6304 & ~n6305;
  assign n6307 = n6306 ^ n6245;
  assign n6363 = n6362 ^ n6307;
  assign n6301 = n6247 ^ n6232;
  assign n6302 = ~n6293 & ~n6301;
  assign n6303 = n6302 ^ n6292;
  assign n6364 = n6363 ^ n6303;
  assign n6369 = n6368 ^ n6364;
  assign n6427 = ~n6303 & n6363;
  assign n6428 = n6303 & ~n6363;
  assign n6429 = ~n6368 & ~n6428;
  assign n6430 = ~n6427 & ~n6429;
  assign n6420 = x23 & x63;
  assign n6412 = x29 & n2379;
  assign n6413 = x28 & n2383;
  assign n6414 = ~n6412 & ~n6413;
  assign n6415 = ~x29 & n2386;
  assign n6416 = ~x28 & n2388;
  assign n6417 = ~n6415 & ~n6416;
  assign n6418 = n6414 & n6417;
  assign n6405 = ~x25 & n3129;
  assign n6406 = ~x24 & n3133;
  assign n6407 = ~n6405 & ~n6406;
  assign n6408 = x25 & n3136;
  assign n6409 = x24 & n3138;
  assign n6410 = ~n6408 & ~n6409;
  assign n6411 = n6407 & n6410;
  assign n6419 = n6418 ^ n6411;
  assign n6421 = n6420 ^ n6419;
  assign n6401 = n6359 ^ n6355;
  assign n6402 = ~n6356 & n6401;
  assign n6403 = n6402 ^ n6359;
  assign n6404 = n6403 ^ n6330;
  assign n6422 = n6421 ^ n6404;
  assign n6392 = ~x27 & n2799;
  assign n6393 = ~x26 & n2803;
  assign n6394 = ~n6392 & ~n6393;
  assign n6395 = x27 & n2806;
  assign n6396 = x26 & n2808;
  assign n6397 = ~n6395 & ~n6396;
  assign n6398 = n6394 & n6397;
  assign n6390 = ~n1835 & ~n1839;
  assign n6383 = ~x31 & n2161;
  assign n6384 = ~x30 & n2165;
  assign n6385 = ~n6383 & ~n6384;
  assign n6386 = x31 & n2168;
  assign n6387 = x30 & n2170;
  assign n6388 = ~n6386 & ~n6387;
  assign n6389 = n6385 & n6388;
  assign n6391 = n6390 ^ n6389;
  assign n6399 = n6398 ^ n6391;
  assign n6379 = n6330 ^ n6322;
  assign n6380 = n6330 ^ n6321;
  assign n6381 = n6379 & n6380;
  assign n6382 = n6381 ^ n6322;
  assign n6400 = n6399 ^ n6382;
  assign n6423 = n6422 ^ n6400;
  assign n6376 = n6360 ^ n6340;
  assign n6377 = n6341 & ~n6376;
  assign n6378 = n6377 ^ n6360;
  assign n6424 = n6423 ^ n6378;
  assign n6373 = n6314 ^ n6311;
  assign n6374 = ~n6332 & n6373;
  assign n6375 = n6374 ^ n6331;
  assign n6425 = n6424 ^ n6375;
  assign n6370 = n6333 ^ n6307;
  assign n6371 = n6362 & ~n6370;
  assign n6372 = n6371 ^ n6361;
  assign n6426 = n6425 ^ n6372;
  assign n6431 = n6430 ^ n6426;
  assign n6482 = n6372 & n6425;
  assign n6483 = ~n6372 & ~n6425;
  assign n6484 = ~n6430 & ~n6483;
  assign n6485 = ~n6482 & ~n6484;
  assign n6469 = ~x30 & n2386;
  assign n6470 = ~x29 & n2388;
  assign n6471 = ~n6469 & ~n6470;
  assign n6472 = x30 & n2379;
  assign n6473 = x29 & n2383;
  assign n6474 = ~n6472 & ~n6473;
  assign n6475 = n6471 & n6474;
  assign n6462 = ~x28 & n2799;
  assign n6463 = ~x27 & n2803;
  assign n6464 = ~n6462 & ~n6463;
  assign n6465 = x28 & n2806;
  assign n6466 = x27 & n2808;
  assign n6467 = ~n6465 & ~n6466;
  assign n6468 = n6464 & n6467;
  assign n6476 = n6475 ^ n6468;
  assign n6459 = n6420 ^ n6418;
  assign n6460 = ~n6419 & ~n6459;
  assign n6461 = n6460 ^ n6420;
  assign n6477 = n6476 ^ n6461;
  assign n6454 = x57 ^ x31;
  assign n6455 = n2164 & n6454;
  assign n6456 = ~n2161 & ~n6455;
  assign n6452 = x24 & x63;
  assign n6445 = x26 & n3136;
  assign n6446 = x25 & n3138;
  assign n6447 = ~n6445 & ~n6446;
  assign n6448 = ~x26 & n3129;
  assign n6449 = ~x25 & n3133;
  assign n6450 = ~n6448 & ~n6449;
  assign n6451 = n6447 & n6450;
  assign n6453 = n6452 ^ n6451;
  assign n6457 = n6456 ^ n6453;
  assign n6442 = n6398 ^ n6389;
  assign n6443 = ~n6391 & ~n6442;
  assign n6444 = n6443 ^ n6390;
  assign n6458 = n6457 ^ n6444;
  assign n6478 = n6477 ^ n6458;
  assign n6438 = n6421 ^ n6330;
  assign n6439 = n6421 ^ n6403;
  assign n6440 = ~n6438 & n6439;
  assign n6441 = n6440 ^ n6330;
  assign n6479 = n6478 ^ n6441;
  assign n6435 = n6422 ^ n6382;
  assign n6436 = n6400 & ~n6435;
  assign n6437 = n6436 ^ n6399;
  assign n6480 = n6479 ^ n6437;
  assign n6432 = n6378 ^ n6375;
  assign n6433 = ~n6424 & ~n6432;
  assign n6434 = n6433 ^ n6423;
  assign n6481 = n6480 ^ n6434;
  assign n6486 = n6485 ^ n6481;
  assign n6532 = n6434 & n6480;
  assign n6533 = ~n6434 & ~n6480;
  assign n6534 = ~n6485 & ~n6533;
  assign n6535 = ~n6532 & ~n6534;
  assign n6525 = x25 & x63;
  assign n6518 = ~x29 & n2799;
  assign n6519 = ~x28 & n2803;
  assign n6520 = ~n6518 & ~n6519;
  assign n6521 = x29 & n2806;
  assign n6522 = x28 & n2808;
  assign n6523 = ~n6521 & ~n6522;
  assign n6524 = n6520 & n6523;
  assign n6526 = n6525 ^ n6524;
  assign n6527 = n6526 ^ n6475;
  assign n6509 = x27 & n3136;
  assign n6510 = x26 & n3138;
  assign n6511 = ~n6509 & ~n6510;
  assign n6512 = ~x27 & n3129;
  assign n6513 = ~x26 & n3133;
  assign n6514 = ~n6512 & ~n6513;
  assign n6515 = n6511 & n6514;
  assign n6507 = ~n2161 & ~n2165;
  assign n6500 = ~x31 & n2386;
  assign n6501 = ~x30 & n2388;
  assign n6502 = ~n6500 & ~n6501;
  assign n6503 = x31 & n2379;
  assign n6504 = x30 & n2383;
  assign n6505 = ~n6503 & ~n6504;
  assign n6506 = n6502 & n6505;
  assign n6508 = n6507 ^ n6506;
  assign n6516 = n6515 ^ n6508;
  assign n6496 = n6456 ^ n6452;
  assign n6497 = n6456 ^ n6451;
  assign n6498 = ~n6496 & ~n6497;
  assign n6499 = n6498 ^ n6452;
  assign n6517 = n6516 ^ n6499;
  assign n6528 = n6527 ^ n6517;
  assign n6493 = n6468 ^ n6461;
  assign n6494 = ~n6476 & n6493;
  assign n6495 = n6494 ^ n6475;
  assign n6529 = n6528 ^ n6495;
  assign n6490 = n6477 ^ n6444;
  assign n6491 = n6458 & n6490;
  assign n6492 = n6491 ^ n6457;
  assign n6530 = n6529 ^ n6492;
  assign n6487 = n6441 ^ n6437;
  assign n6488 = n6479 & n6487;
  assign n6489 = n6488 ^ n6478;
  assign n6531 = n6530 ^ n6489;
  assign n6536 = n6535 ^ n6531;
  assign n6576 = ~n6489 & n6530;
  assign n6577 = n6489 & ~n6530;
  assign n6578 = ~n6535 & ~n6577;
  assign n6579 = ~n6576 & ~n6578;
  assign n6564 = x28 & n3136;
  assign n6565 = x27 & n3138;
  assign n6566 = ~n6564 & ~n6565;
  assign n6567 = ~x28 & n3129;
  assign n6568 = ~x27 & n3133;
  assign n6569 = ~n6567 & ~n6568;
  assign n6570 = n6566 & n6569;
  assign n6562 = x26 & x63;
  assign n6555 = ~x30 & n2799;
  assign n6556 = ~x29 & n2803;
  assign n6557 = ~n6555 & ~n6556;
  assign n6558 = x30 & n2806;
  assign n6559 = x29 & n2808;
  assign n6560 = ~n6558 & ~n6559;
  assign n6561 = n6557 & n6560;
  assign n6563 = n6562 ^ n6561;
  assign n6571 = n6570 ^ n6563;
  assign n6551 = x59 ^ x31;
  assign n6552 = n2382 & n6551;
  assign n6553 = ~n2386 & ~n6552;
  assign n6547 = n6515 ^ n6507;
  assign n6548 = n6515 ^ n6506;
  assign n6549 = ~n6547 & ~n6548;
  assign n6550 = n6549 ^ n6507;
  assign n6554 = n6553 ^ n6550;
  assign n6572 = n6571 ^ n6554;
  assign n6543 = n6525 ^ n6475;
  assign n6544 = n6524 ^ n6475;
  assign n6545 = ~n6543 & ~n6544;
  assign n6546 = n6545 ^ n6525;
  assign n6573 = n6572 ^ n6546;
  assign n6540 = n6527 ^ n6516;
  assign n6541 = ~n6517 & n6540;
  assign n6542 = n6541 ^ n6527;
  assign n6574 = n6573 ^ n6542;
  assign n6537 = n6495 ^ n6492;
  assign n6538 = n6529 & ~n6537;
  assign n6539 = n6538 ^ n6528;
  assign n6575 = n6574 ^ n6539;
  assign n6580 = n6579 ^ n6575;
  assign n6614 = n6539 & n6574;
  assign n6615 = ~n6539 & ~n6574;
  assign n6616 = ~n6579 & ~n6615;
  assign n6617 = ~n6614 & ~n6616;
  assign n6609 = x27 & x63;
  assign n6607 = ~n2386 & ~n2388;
  assign n6600 = x31 & n2806;
  assign n6601 = x30 & n2808;
  assign n6602 = ~n6600 & ~n6601;
  assign n6603 = ~x31 & n2799;
  assign n6604 = ~x30 & n2803;
  assign n6605 = ~n6603 & ~n6604;
  assign n6606 = n6602 & n6605;
  assign n6608 = n6607 ^ n6606;
  assign n6610 = n6609 ^ n6608;
  assign n6591 = ~x29 & n3129;
  assign n6592 = ~x28 & n3133;
  assign n6593 = ~n6591 & ~n6592;
  assign n6594 = x29 & n3136;
  assign n6595 = x28 & n3138;
  assign n6596 = ~n6594 & ~n6595;
  assign n6597 = n6593 & n6596;
  assign n6598 = n6597 ^ n6553;
  assign n6588 = n6570 ^ n6561;
  assign n6589 = ~n6563 & ~n6588;
  assign n6590 = n6589 ^ n6562;
  assign n6599 = n6598 ^ n6590;
  assign n6611 = n6610 ^ n6599;
  assign n6584 = n6571 ^ n6553;
  assign n6585 = n6571 ^ n6550;
  assign n6586 = n6584 & ~n6585;
  assign n6587 = n6586 ^ n6553;
  assign n6612 = n6611 ^ n6587;
  assign n6581 = n6572 ^ n6542;
  assign n6582 = n6573 & ~n6581;
  assign n6583 = n6582 ^ n6546;
  assign n6613 = n6612 ^ n6583;
  assign n6618 = n6617 ^ n6613;
  assign n6644 = n6583 & ~n6612;
  assign n6645 = ~n6583 & n6612;
  assign n6646 = ~n6617 & ~n6645;
  assign n6647 = ~n6644 & ~n6646;
  assign n6637 = x61 ^ x31;
  assign n6638 = n2802 & n6637;
  assign n6639 = ~n2799 & ~n6638;
  assign n6635 = x28 & x63;
  assign n6628 = ~x30 & n3129;
  assign n6629 = ~x29 & n3133;
  assign n6630 = ~n6628 & ~n6629;
  assign n6631 = x30 & n3136;
  assign n6632 = x29 & n3138;
  assign n6633 = ~n6631 & ~n6632;
  assign n6634 = n6630 & n6633;
  assign n6636 = n6635 ^ n6634;
  assign n6640 = n6639 ^ n6636;
  assign n6625 = n6609 ^ n6607;
  assign n6626 = n6608 & n6625;
  assign n6627 = n6626 ^ n6609;
  assign n6641 = n6640 ^ n6627;
  assign n6622 = n6597 ^ n6590;
  assign n6623 = n6598 & n6622;
  assign n6624 = n6623 ^ n6553;
  assign n6642 = n6641 ^ n6624;
  assign n6619 = n6599 ^ n6587;
  assign n6620 = ~n6611 & ~n6619;
  assign n6621 = n6620 ^ n6610;
  assign n6643 = n6642 ^ n6621;
  assign n6648 = n6647 ^ n6643;
  assign n6670 = ~n6621 & n6642;
  assign n6671 = n6621 & ~n6642;
  assign n6672 = ~n6647 & ~n6671;
  assign n6673 = ~n6670 & ~n6672;
  assign n6665 = x29 & x63;
  assign n6663 = ~n2799 & ~n2803;
  assign n6656 = x31 & n3136;
  assign n6657 = x30 & n3138;
  assign n6658 = ~n6656 & ~n6657;
  assign n6659 = ~x31 & n3129;
  assign n6660 = ~x30 & n3133;
  assign n6661 = ~n6659 & ~n6660;
  assign n6662 = n6658 & n6661;
  assign n6664 = n6663 ^ n6662;
  assign n6666 = n6665 ^ n6664;
  assign n6667 = n6666 ^ n6639;
  assign n6652 = n6639 ^ n6635;
  assign n6653 = n6639 ^ n6634;
  assign n6654 = n6652 & n6653;
  assign n6655 = n6654 ^ n6635;
  assign n6668 = n6667 ^ n6655;
  assign n6649 = n6627 ^ n6624;
  assign n6650 = ~n6641 & n6649;
  assign n6651 = n6650 ^ n6640;
  assign n6669 = n6668 ^ n6651;
  assign n6674 = n6673 ^ n6669;
  assign n6688 = ~n6651 & n6668;
  assign n6689 = n6651 & ~n6668;
  assign n6690 = ~n6673 & ~n6689;
  assign n6691 = ~n6688 & ~n6690;
  assign n6684 = x30 & x63;
  assign n6681 = x63 ^ x31;
  assign n6682 = n3132 & n6681;
  assign n6683 = ~n3129 & ~n6682;
  assign n6685 = n6684 ^ n6683;
  assign n6678 = n6665 ^ n6663;
  assign n6679 = n6664 & n6678;
  assign n6680 = n6679 ^ n6665;
  assign n6686 = n6685 ^ n6680;
  assign n6675 = n6666 ^ n6655;
  assign n6676 = n6667 & n6675;
  assign n6677 = n6676 ^ n6639;
  assign n6687 = n6686 ^ n6677;
  assign n6692 = n6691 ^ n6687;
  assign n6700 = ~n3034 & ~n3132;
  assign n6701 = n6700 ^ x31;
  assign n6702 = x63 & ~n6701;
  assign n6703 = n6702 ^ n6684;
  assign n6697 = n6683 ^ n6680;
  assign n6698 = n6685 & n6697;
  assign n6699 = n6698 ^ n6684;
  assign n6704 = n6703 ^ n6699;
  assign n6693 = ~n6677 & n6686;
  assign n6694 = n6677 & ~n6686;
  assign n6695 = ~n6691 & ~n6694;
  assign n6696 = ~n6693 & ~n6695;
  assign n6705 = n6704 ^ n6696;
  assign y0 = n65;
  assign y1 = ~n77;
  assign y2 = ~n88;
  assign y3 = ~n118;
  assign y4 = ~n142;
  assign y5 = n185;
  assign y6 = ~n221;
  assign y7 = n275;
  assign y8 = ~n325;
  assign y9 = ~n392;
  assign y10 = ~n453;
  assign y11 = ~n532;
  assign y12 = ~n604;
  assign y13 = n695;
  assign y14 = n779;
  assign y15 = n882;
  assign y16 = n981;
  assign y17 = n1096;
  assign y18 = ~n1205;
  assign y19 = ~n1332;
  assign y20 = n1456;
  assign y21 = ~n1596;
  assign y22 = n1730;
  assign y23 = n1882;
  assign y24 = n2027;
  assign y25 = ~n2193;
  assign y26 = n2353;
  assign y27 = ~n2530;
  assign y28 = ~n2701;
  assign y29 = ~n2890;
  assign y30 = ~n3072;
  assign y31 = n3273;
  assign y32 = ~n3461;
  assign y33 = n3652;
  assign y34 = ~n3839;
  assign y35 = n4024;
  assign y36 = n4205;
  assign y37 = ~n4380;
  assign y38 = n4544;
  assign y39 = n4704;
  assign y40 = n4857;
  assign y41 = ~n5008;
  assign y42 = ~n5148;
  assign y43 = n5287;
  assign y44 = n5414;
  assign y45 = n5540;
  assign y46 = ~n5657;
  assign y47 = ~n5769;
  assign y48 = n5872;
  assign y49 = n5969;
  assign y50 = ~n6062;
  assign y51 = ~n6147;
  assign y52 = n6226;
  assign y53 = n6300;
  assign y54 = n6369;
  assign y55 = ~n6431;
  assign y56 = ~n6486;
  assign y57 = n6536;
  assign y58 = ~n6580;
  assign y59 = n6618;
  assign y60 = n6648;
  assign y61 = n6674;
  assign y62 = n6692;
  assign y63 = ~n6705;
endmodule
