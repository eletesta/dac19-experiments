module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24;
  wire n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350;
  assign n25 = ~x0 & ~x1;
  assign n26 = ~x2 & n25;
  assign n27 = ~x3 & n26;
  assign n28 = ~x4 & n27;
  assign n29 = ~x5 & n28;
  assign n30 = ~x6 & ~x7;
  assign n31 = n29 & n30;
  assign n32 = ~x8 & n31;
  assign n33 = ~x9 & n32;
  assign n34 = ~x10 & n33;
  assign n35 = ~x11 & n34;
  assign n36 = ~x12 & ~x13;
  assign n37 = ~x14 & n36;
  assign n38 = n35 & n37;
  assign n39 = ~x22 & ~n38;
  assign n40 = n39 ^ x15;
  assign n41 = ~x15 & n38;
  assign n42 = ~x22 & ~n41;
  assign n43 = ~x18 & ~x19;
  assign n44 = ~x16 & ~x17;
  assign n45 = n43 & n44;
  assign n46 = ~n42 & n45;
  assign n47 = ~x22 & ~n46;
  assign n48 = n47 ^ x20;
  assign n49 = x22 ^ x21;
  assign n164 = n48 & ~n49;
  assign n165 = ~n40 & n164;
  assign n59 = x18 & ~x19;
  assign n60 = ~x22 & n59;
  assign n102 = x16 & x17;
  assign n103 = ~n41 & n102;
  assign n233 = n60 & n103;
  assign n66 = ~x18 & x19;
  assign n234 = n44 & n66;
  assign n235 = ~n42 & n234;
  assign n236 = ~n233 & ~n235;
  assign n237 = n165 & ~n236;
  assign n52 = x21 ^ x20;
  assign n100 = n49 & ~n52;
  assign n152 = ~n40 & n100;
  assign n70 = n41 ^ x16;
  assign n71 = x17 & ~n70;
  assign n119 = ~x22 & n43;
  assign n156 = n71 & n119;
  assign n75 = x16 & ~x17;
  assign n86 = x18 & x19;
  assign n121 = x22 & n86;
  assign n157 = n75 & n121;
  assign n158 = ~n156 & ~n157;
  assign n238 = n152 & ~n158;
  assign n53 = x21 & x22;
  assign n54 = ~n52 & n53;
  assign n55 = n54 ^ n52;
  assign n56 = ~n48 & n55;
  assign n83 = ~n40 & n56;
  assign n87 = ~x22 & n86;
  assign n136 = n87 & n103;
  assign n137 = ~n46 & ~n136;
  assign n239 = n83 & ~n137;
  assign n240 = ~n238 & ~n239;
  assign n241 = ~n237 & n240;
  assign n61 = x17 ^ x16;
  assign n62 = n41 ^ x17;
  assign n63 = n61 & ~n62;
  assign n64 = n60 & n63;
  assign n65 = ~x16 & x17;
  assign n67 = x22 & n66;
  assign n68 = n65 & n67;
  assign n69 = ~n64 & ~n68;
  assign n287 = ~n69 & n83;
  assign n84 = n40 & ~n49;
  assign n85 = n48 & n84;
  assign n72 = x19 & ~x22;
  assign n73 = ~x18 & n72;
  assign n95 = n63 & n73;
  assign n76 = x22 & n59;
  assign n96 = n65 & n76;
  assign n97 = ~n95 & ~n96;
  assign n288 = n85 & ~n97;
  assign n50 = n48 & n49;
  assign n51 = ~n40 & n50;
  assign n113 = ~x17 & ~n70;
  assign n114 = n87 & n113;
  assign n89 = x22 & n43;
  assign n115 = n89 & n102;
  assign n116 = ~n114 & ~n115;
  assign n289 = n51 & ~n116;
  assign n290 = ~n288 & ~n289;
  assign n291 = ~n287 & n290;
  assign n865 = n241 & n291;
  assign n397 = n40 & n48;
  assign n398 = ~n158 & n397;
  assign n399 = n49 & n398;
  assign n104 = x18 & n44;
  assign n105 = ~n103 & ~n104;
  assign n106 = x18 & n42;
  assign n107 = n106 ^ x22;
  assign n108 = ~n105 & ~n107;
  assign n109 = n44 & n86;
  assign n110 = ~n108 & ~n109;
  assign n111 = ~n72 & ~n110;
  assign n74 = n71 & n73;
  assign n77 = n75 & n76;
  assign n78 = ~n74 & ~n77;
  assign n639 = n78 & n116;
  assign n640 = ~n111 & n639;
  assign n641 = n83 & ~n640;
  assign n642 = ~n399 & ~n641;
  assign n153 = n113 & n119;
  assign n154 = n102 & n121;
  assign n155 = ~n153 & ~n154;
  assign n322 = n152 & ~n155;
  assign n341 = n83 & ~n158;
  assign n130 = n40 & n50;
  assign n519 = ~n116 & n130;
  assign n866 = ~n341 & ~n519;
  assign n867 = ~n322 & n866;
  assign n868 = n642 & n867;
  assign n869 = n865 & n868;
  assign n334 = n83 & ~n236;
  assign n120 = n63 & n119;
  assign n122 = n65 & n121;
  assign n123 = ~n120 & ~n122;
  assign n88 = n71 & n87;
  assign n90 = n75 & n89;
  assign n91 = ~n88 & ~n90;
  assign n101 = n40 & n100;
  assign n200 = ~n91 & n101;
  assign n148 = n91 & n137;
  assign n870 = n85 & ~n148;
  assign n871 = ~n200 & ~n870;
  assign n872 = n123 & n871;
  assign n873 = n84 & ~n872;
  assign n874 = ~n334 & ~n873;
  assign n875 = n869 & n874;
  assign n649 = n51 & ~n236;
  assign n998 = ~n78 & n152;
  assign n1514 = ~n649 & ~n998;
  assign n644 = ~n69 & n101;
  assign n217 = n60 & n71;
  assign n218 = n67 & n75;
  assign n219 = ~n217 & ~n218;
  assign n688 = n130 & ~n219;
  assign n1515 = ~n644 & ~n688;
  assign n1516 = n1514 & n1515;
  assign n144 = x19 & n108;
  assign n145 = n44 & n76;
  assign n146 = ~n144 & ~n145;
  assign n211 = ~n83 & ~n101;
  assign n212 = ~n146 & ~n211;
  assign n410 = n51 & n111;
  assign n138 = n73 & n113;
  assign n139 = n76 & n102;
  assign n140 = ~n138 & ~n139;
  assign n523 = n83 & ~n140;
  assign n1517 = ~n410 & ~n523;
  assign n1518 = ~n212 & n1517;
  assign n1519 = n1516 & n1518;
  assign n485 = ~n97 & n130;
  assign n441 = ~n78 & n101;
  assign n263 = ~n40 & ~n219;
  assign n505 = n164 & n263;
  assign n1520 = ~n441 & ~n505;
  assign n1521 = ~n485 & n1520;
  assign n1522 = n1519 & n1521;
  assign n168 = n60 & n113;
  assign n169 = n67 & n102;
  assign n170 = ~n168 & ~n169;
  assign n330 = n83 & ~n170;
  assign n442 = n130 & ~n155;
  assign n879 = ~n330 & ~n442;
  assign n224 = ~n69 & n152;
  assign n512 = n170 & n219;
  assign n2806 = n85 & ~n512;
  assign n2807 = ~n224 & ~n2806;
  assign n2808 = n879 & n2807;
  assign n266 = ~n111 & n158;
  assign n126 = n63 & n87;
  assign n127 = n65 & n89;
  assign n128 = ~n126 & ~n127;
  assign n149 = n116 & n128;
  assign n2809 = n146 & n149;
  assign n2810 = n266 & n2809;
  assign n2811 = n165 & ~n2810;
  assign n2812 = n2808 & ~n2811;
  assign n2813 = n1522 & n2812;
  assign n366 = ~n128 & n165;
  assign n422 = n83 & ~n128;
  assign n713 = ~n366 & ~n422;
  assign n844 = ~n97 & n101;
  assign n845 = n713 & ~n844;
  assign n188 = n83 & ~n91;
  assign n57 = n40 & n56;
  assign n298 = n57 & ~n155;
  assign n846 = ~n188 & ~n298;
  assign n471 = n101 & ~n155;
  assign n79 = n69 & n78;
  assign n847 = ~n79 & n85;
  assign n848 = ~n471 & ~n847;
  assign n849 = n846 & n848;
  assign n850 = n845 & n849;
  assign n278 = n51 & ~n78;
  assign n372 = ~n123 & n130;
  assign n373 = ~n278 & ~n372;
  assign n456 = n83 & ~n97;
  assign n927 = n50 & ~n91;
  assign n928 = ~n456 & ~n927;
  assign n929 = n373 & n928;
  assign n220 = n101 & ~n219;
  assign n280 = n56 & n263;
  assign n1591 = ~n220 & ~n280;
  assign n2814 = ~n211 & ~n266;
  assign n569 = n51 & ~n170;
  assign n340 = n85 & ~n155;
  assign n394 = ~n140 & n152;
  assign n672 = ~n97 & n152;
  assign n2815 = ~n394 & ~n672;
  assign n2816 = ~n340 & n2815;
  assign n2817 = ~n569 & n2816;
  assign n2818 = ~n2814 & n2817;
  assign n2819 = n1591 & n2818;
  assign n2820 = n929 & n2819;
  assign n2821 = n850 & n2820;
  assign n2822 = n2813 & n2821;
  assign n2823 = n875 & n2822;
  assign n58 = ~n51 & ~n57;
  assign n80 = ~n40 & n69;
  assign n81 = ~n79 & ~n80;
  assign n82 = ~n58 & n81;
  assign n195 = n83 & ~n123;
  assign n331 = n152 & ~n236;
  assign n637 = ~n195 & ~n331;
  assign n638 = ~n82 & n637;
  assign n180 = ~n69 & n165;
  assign n181 = n165 & ~n170;
  assign n182 = ~n180 & ~n181;
  assign n243 = n97 & n219;
  assign n244 = n165 & ~n243;
  assign n374 = n57 & ~n123;
  assign n375 = ~n244 & ~n374;
  assign n376 = n182 & n375;
  assign n377 = n373 & n376;
  assign n1752 = ~n123 & ~n377;
  assign n428 = ~n78 & n130;
  assign n613 = n57 & ~n116;
  assign n836 = ~n428 & ~n613;
  assign n192 = n51 & ~n128;
  assign n402 = n51 & ~n146;
  assign n403 = ~n192 & ~n402;
  assign n141 = n137 & n140;
  assign n1032 = n51 & ~n141;
  assign n1033 = n403 & ~n1032;
  assign n1034 = n836 & n1033;
  assign n225 = ~n69 & n85;
  assign n226 = ~n224 & ~n225;
  assign n1753 = ~n322 & ~n422;
  assign n1754 = n226 & n1753;
  assign n418 = ~n123 & n152;
  assign n419 = n101 & ~n146;
  assign n420 = ~n418 & ~n419;
  assign n421 = ~n220 & n420;
  assign n1755 = ~n330 & n421;
  assign n1756 = n1754 & n1755;
  assign n1757 = n1034 & n1756;
  assign n1758 = ~n1752 & n1757;
  assign n1759 = n638 & n1758;
  assign n378 = ~n85 & n140;
  assign n379 = ~n101 & n123;
  assign n380 = ~n378 & ~n379;
  assign n245 = n51 & ~n155;
  assign n712 = ~n245 & ~n287;
  assign n1760 = ~n380 & n712;
  assign n1761 = n1759 & n1760;
  assign n351 = ~n83 & ~n130;
  assign n352 = ~n155 & ~n351;
  assign n353 = ~n123 & n165;
  assign n354 = ~n128 & n164;
  assign n355 = n40 & n354;
  assign n356 = ~n353 & ~n355;
  assign n357 = ~n352 & n356;
  assign n358 = n57 & ~n140;
  assign n359 = ~n78 & n85;
  assign n360 = ~n358 & ~n359;
  assign n293 = n57 & ~n97;
  assign n361 = n116 & n236;
  assign n362 = n51 & ~n361;
  assign n363 = ~n293 & ~n362;
  assign n364 = n360 & n363;
  assign n365 = n357 & n364;
  assign n367 = n57 & ~n219;
  assign n368 = ~n137 & n152;
  assign n369 = ~n367 & ~n368;
  assign n370 = ~n366 & n369;
  assign n371 = n365 & n370;
  assign n261 = n40 & ~n128;
  assign n262 = n56 & n261;
  assign n721 = ~n262 & ~n441;
  assign n396 = n101 & ~n170;
  assign n730 = ~n280 & ~n396;
  assign n940 = n56 & ~n146;
  assign n941 = n730 & ~n940;
  assign n942 = n721 & n941;
  assign n316 = n130 & ~n236;
  assign n943 = ~n316 & ~n485;
  assign n473 = n84 & ~n140;
  assign n944 = ~n111 & ~n473;
  assign n945 = n48 & ~n944;
  assign n946 = n943 & ~n945;
  assign n947 = n942 & n946;
  assign n2502 = n371 & n947;
  assign n112 = n101 & n111;
  assign n117 = n83 & ~n116;
  assign n118 = ~n112 & ~n117;
  assign n385 = n85 & ~n219;
  assign n1542 = ~n78 & n165;
  assign n1543 = ~n385 & ~n1542;
  assign n2503 = n118 & n1543;
  assign n255 = n97 & n140;
  assign n1765 = n78 & n255;
  assign n1766 = n83 & ~n1765;
  assign n1767 = ~n298 & ~n1766;
  assign n271 = n101 & ~n137;
  assign n2504 = ~n180 & ~n271;
  assign n2505 = n1767 & n2504;
  assign n2506 = n2503 & n2505;
  assign n589 = n85 & n111;
  assign n2507 = n165 & ~n361;
  assign n2508 = ~n589 & ~n2507;
  assign n413 = n51 & ~n91;
  assign n728 = n57 & ~n236;
  assign n2509 = ~n413 & ~n728;
  assign n2510 = n2508 & n2509;
  assign n567 = ~n91 & n152;
  assign n2511 = ~n334 & ~n567;
  assign n693 = n152 & ~n170;
  assign n2512 = ~n693 & ~n998;
  assign n2513 = n2511 & n2512;
  assign n2514 = n2510 & n2513;
  assign n2515 = n2506 & n2514;
  assign n2516 = n2502 & n2515;
  assign n2517 = n1761 & n2516;
  assign n761 = ~n116 & n164;
  assign n762 = ~n225 & ~n761;
  assign n763 = n57 & ~n266;
  assign n764 = n762 & ~n763;
  assign n765 = n182 & n764;
  assign n258 = n83 & ~n155;
  assign n766 = n123 & ~n164;
  assign n767 = ~n258 & n766;
  assign n768 = ~n56 & ~n111;
  assign n769 = n85 & ~n170;
  assign n770 = n768 & ~n769;
  assign n771 = ~n767 & ~n770;
  assign n772 = n83 & ~n266;
  assign n773 = ~n771 & ~n772;
  assign n774 = n765 & n773;
  assign n617 = n140 & n146;
  assign n775 = ~n56 & n617;
  assign n776 = n219 & n236;
  assign n777 = ~n164 & n776;
  assign n778 = ~n775 & ~n777;
  assign n779 = n140 & n170;
  assign n780 = n69 & n779;
  assign n781 = n56 & ~n780;
  assign n782 = ~n293 & ~n781;
  assign n783 = ~n778 & n782;
  assign n557 = ~n288 & ~n298;
  assign n784 = ~n164 & n557;
  assign n785 = n783 & n784;
  assign n786 = n774 & n785;
  assign n787 = n56 & n786;
  assign n381 = n51 & ~n123;
  assign n150 = n148 & n149;
  assign n788 = n83 & ~n150;
  assign n789 = ~n381 & ~n788;
  assign n404 = n69 & n155;
  assign n790 = n130 & ~n404;
  assign n791 = n789 & ~n790;
  assign n792 = ~n410 & n791;
  assign n793 = ~n111 & n123;
  assign n794 = n40 & ~n793;
  assign n795 = n158 & n170;
  assign n796 = ~n794 & n795;
  assign n797 = n50 & ~n796;
  assign n798 = ~n245 & ~n797;
  assign n799 = n792 & n798;
  assign n800 = ~n787 & n799;
  assign n227 = ~n57 & n137;
  assign n317 = n78 & n146;
  assign n502 = ~n130 & n317;
  assign n503 = ~n227 & ~n502;
  assign n159 = n155 & n158;
  assign n160 = n123 & n159;
  assign n801 = n160 & ~n794;
  assign n802 = n100 & ~n801;
  assign n595 = n51 & ~n137;
  assign n803 = n56 & ~n317;
  assign n804 = ~n595 & ~n803;
  assign n805 = ~n802 & n804;
  assign n806 = ~n503 & n805;
  assign n807 = n69 & n512;
  assign n808 = n100 & ~n807;
  assign n423 = n101 & ~n236;
  assign n464 = n111 & n152;
  assign n809 = ~n423 & ~n464;
  assign n810 = ~n808 & n809;
  assign n811 = n806 & n810;
  assign n812 = n800 & n811;
  assign n643 = n638 & n642;
  assign n264 = n50 & n263;
  assign n645 = ~n155 & n164;
  assign n646 = ~n40 & n645;
  assign n647 = ~n644 & ~n646;
  assign n648 = ~n264 & n647;
  assign n563 = n130 & ~n146;
  assign n650 = ~n563 & ~n649;
  assign n651 = n648 & n650;
  assign n652 = n643 & n651;
  assign n171 = n146 & n170;
  assign n653 = n116 & n171;
  assign n654 = n57 & ~n653;
  assign n655 = ~n288 & ~n654;
  assign n656 = ~n442 & ~n464;
  assign n657 = ~n237 & n656;
  assign n658 = n655 & n657;
  assign n659 = n652 & n658;
  assign n382 = ~n158 & n165;
  assign n383 = ~n381 & ~n382;
  assign n384 = ~n380 & n383;
  assign n386 = ~n101 & n140;
  assign n387 = ~n385 & n386;
  assign n388 = n97 & ~n164;
  assign n389 = ~n387 & ~n388;
  assign n390 = n384 & ~n389;
  assign n391 = n377 & n390;
  assign n660 = ~n116 & n152;
  assign n661 = ~n394 & ~n660;
  assign n662 = ~n245 & n661;
  assign n539 = n57 & n111;
  assign n147 = n123 & n146;
  assign n663 = n51 & ~n147;
  assign n664 = ~n539 & ~n663;
  assign n665 = ~n236 & n397;
  assign n666 = ~n595 & ~n665;
  assign n667 = n664 & n666;
  assign n668 = n662 & n667;
  assign n669 = n391 & n668;
  assign n670 = n659 & n669;
  assign n671 = ~n78 & n164;
  assign n129 = n101 & ~n128;
  assign n673 = ~n129 & ~n672;
  assign n674 = ~n671 & n673;
  assign n675 = ~n322 & ~n396;
  assign n676 = n674 & n675;
  assign n286 = n101 & ~n116;
  assign n520 = ~n286 & ~n471;
  assign n521 = ~n519 & n520;
  assign n272 = ~n128 & n152;
  assign n677 = ~n272 & ~n353;
  assign n678 = n170 & n404;
  assign n679 = n85 & ~n678;
  assign n680 = ~n40 & ~n97;
  assign n681 = n158 & ~n680;
  assign n682 = n56 & ~n681;
  assign n683 = ~n679 & ~n682;
  assign n684 = n677 & n683;
  assign n685 = n521 & n684;
  assign n686 = n676 & n685;
  assign n687 = n85 & ~n158;
  assign n689 = n111 & n165;
  assign n690 = ~n688 & ~n689;
  assign n691 = ~n687 & n690;
  assign n577 = n130 & ~n137;
  assign n692 = ~n577 & ~n589;
  assign n694 = ~n83 & ~n693;
  assign n695 = ~n171 & ~n694;
  assign n696 = n692 & ~n695;
  assign n697 = n691 & n696;
  assign n698 = n686 & n697;
  assign n699 = n670 & n698;
  assign n92 = n85 & ~n91;
  assign n93 = ~n83 & ~n92;
  assign n94 = ~n82 & n93;
  assign n98 = n80 & n97;
  assign n99 = ~n94 & ~n98;
  assign n124 = n58 & ~n123;
  assign n125 = n118 & ~n124;
  assign n131 = ~n91 & n130;
  assign n132 = ~n129 & ~n131;
  assign n133 = n125 & n132;
  assign n134 = ~n99 & n133;
  assign n135 = ~n51 & n134;
  assign n142 = ~n85 & n141;
  assign n143 = ~n135 & ~n142;
  assign n151 = n56 & n150;
  assign n161 = n152 & n160;
  assign n162 = ~n151 & ~n161;
  assign n163 = n147 & n162;
  assign n166 = n78 & ~n165;
  assign n167 = ~n163 & ~n166;
  assign n172 = n128 & n171;
  assign n173 = n85 & ~n172;
  assign n174 = n123 & n140;
  assign n175 = ~n83 & n174;
  assign n176 = n78 & ~n101;
  assign n177 = n97 & n176;
  assign n178 = ~n175 & ~n177;
  assign n179 = ~n173 & ~n178;
  assign n183 = ~n116 & n165;
  assign n184 = n182 & ~n183;
  assign n185 = n179 & n184;
  assign n186 = ~n167 & n185;
  assign n187 = ~n143 & n186;
  assign n273 = n130 & ~n140;
  assign n332 = ~n273 & ~n331;
  assign n274 = n51 & ~n69;
  assign n700 = ~n274 & ~n340;
  assign n701 = n332 & n700;
  assign n702 = n187 & n701;
  assign n545 = ~n91 & n165;
  assign n813 = ~n40 & n48;
  assign n814 = ~n236 & n813;
  assign n815 = ~n545 & ~n814;
  assign n299 = n57 & ~n137;
  assign n816 = ~n299 & ~n441;
  assign n817 = n815 & n816;
  assign n221 = ~n146 & n152;
  assign n600 = n57 & ~n146;
  assign n818 = ~n221 & ~n600;
  assign n819 = n118 & n818;
  assign n820 = n817 & n819;
  assign n821 = ~n141 & n164;
  assign n822 = ~n165 & ~n821;
  assign n823 = ~n688 & n822;
  assign n824 = ~n40 & n78;
  assign n825 = ~n823 & ~n824;
  assign n826 = ~n130 & n146;
  assign n445 = ~n101 & n236;
  assign n827 = n137 & n445;
  assign n828 = ~n826 & ~n827;
  assign n829 = n164 & ~n243;
  assign n830 = ~n418 & ~n680;
  assign n831 = ~n829 & n830;
  assign n832 = ~n828 & n831;
  assign n833 = ~n825 & n832;
  assign n834 = n820 & n833;
  assign n835 = n702 & n834;
  assign n343 = n85 & ~n236;
  assign n453 = ~n140 & n165;
  assign n454 = ~n343 & ~n453;
  assign n455 = ~n394 & n454;
  assign n837 = n455 & n836;
  assign n838 = n137 & ~n165;
  assign n839 = ~n768 & ~n838;
  assign n840 = ~n238 & ~n839;
  assign n841 = n837 & n840;
  assign n251 = n155 & n170;
  assign n252 = n165 & ~n251;
  assign n253 = n101 & ~n140;
  assign n254 = ~n252 & ~n253;
  assign n256 = n130 & ~n255;
  assign n257 = n254 & ~n256;
  assign n259 = ~n137 & n165;
  assign n260 = ~n258 & ~n259;
  assign n265 = ~n262 & ~n264;
  assign n267 = n85 & ~n266;
  assign n268 = n265 & ~n267;
  assign n269 = n260 & n268;
  assign n270 = n257 & n269;
  assign n842 = n270 & n805;
  assign n843 = n841 & n842;
  assign n468 = n85 & ~n116;
  assign n216 = n57 & ~n91;
  assign n851 = ~n216 & ~n382;
  assign n852 = ~n468 & n851;
  assign n853 = n850 & n852;
  assign n854 = n843 & n853;
  assign n855 = n835 & n854;
  assign n856 = ~n699 & ~n855;
  assign n857 = ~n812 & ~n856;
  assign n965 = n699 & n855;
  assign n863 = ~x22 & ~n35;
  assign n987 = x12 & ~x22;
  assign n988 = ~n863 & ~n987;
  assign n1077 = x13 & ~x22;
  assign n1078 = n988 & ~n1077;
  assign n1079 = n1078 ^ x14;
  assign n2331 = n965 & ~n1079;
  assign n2332 = n857 & ~n2331;
  assign n964 = n812 & n856;
  assign n2333 = n964 & ~n1079;
  assign n2334 = ~n2332 & ~n2333;
  assign n1068 = ~n50 & n812;
  assign n864 = n863 ^ x12;
  assign n2325 = ~n786 & ~n864;
  assign n2326 = n1068 & ~n2325;
  assign n989 = n988 ^ x13;
  assign n1070 = n786 & n800;
  assign n2327 = n989 & n1070;
  assign n2328 = ~n800 & ~n864;
  assign n2329 = ~n2327 & ~n2328;
  assign n2330 = ~n2326 & n2329;
  assign n2239 = n1079 ^ n989;
  assign n2389 = n800 & n2239;
  assign n2390 = n2389 ^ n989;
  assign n2391 = ~n1068 & ~n2390;
  assign n2392 = ~n786 & n989;
  assign n2393 = ~n2391 & ~n2392;
  assign n2404 = ~n2330 & n2393;
  assign n307 = ~x22 & ~n34;
  assign n308 = n307 ^ x11;
  assign n1734 = n864 ^ n308;
  assign n2387 = ~n786 & n1734;
  assign n2388 = ~n857 & ~n2387;
  assign n2403 = n989 & ~n2388;
  assign n2405 = n2404 ^ n2403;
  assign n2406 = n2334 & n2405;
  assign n2407 = n2406 ^ n2404;
  assign n2408 = ~n786 & n2407;
  assign n2394 = n2393 ^ n2388;
  assign n2395 = ~n2330 & n2334;
  assign n2396 = ~n2394 & n2395;
  assign n2409 = ~n2388 & n2393;
  assign n2468 = ~n2396 & ~n2409;
  assign n2469 = ~n2408 & n2468;
  assign n2464 = ~n800 & ~n1079;
  assign n2230 = ~n308 & ~n864;
  assign n2465 = n2239 ^ n2230;
  assign n2466 = ~n786 & n2465;
  assign n2467 = ~n2464 & ~n2466;
  assign n2470 = n2469 ^ n2467;
  assign n2335 = n2334 ^ n2330;
  assign n314 = ~x22 & ~n33;
  assign n315 = n314 ^ x10;
  assign n311 = ~x22 & ~n32;
  assign n312 = n311 ^ x9;
  assign n1697 = n315 ^ n312;
  assign n439 = ~n334 & ~n381;
  assign n440 = ~n212 & n439;
  assign n443 = ~n441 & ~n442;
  assign n444 = n440 & n443;
  assign n446 = n97 & ~n130;
  assign n447 = ~n445 & ~n446;
  assign n448 = ~n238 & ~n447;
  assign n424 = n152 & ~n219;
  assign n449 = ~n278 & ~n424;
  assign n450 = ~n183 & n449;
  assign n451 = n448 & n450;
  assign n452 = n444 & n451;
  assign n199 = n83 & n111;
  assign n457 = ~n199 & ~n456;
  assign n458 = ~n287 & n457;
  assign n459 = n455 & n458;
  assign n460 = n452 & n459;
  assign n461 = ~n101 & ~n165;
  assign n462 = ~n148 & ~n461;
  assign n463 = n51 & ~n158;
  assign n465 = ~n224 & ~n464;
  assign n466 = ~n463 & n465;
  assign n467 = ~n462 & n466;
  assign n469 = ~n402 & ~n468;
  assign n470 = n467 & n469;
  assign n242 = n130 & ~n170;
  assign n472 = ~n242 & ~n471;
  assign n474 = ~n50 & n170;
  assign n475 = ~n100 & n116;
  assign n476 = ~n40 & ~n475;
  assign n477 = ~n474 & n476;
  assign n478 = ~n473 & ~n477;
  assign n479 = n472 & n478;
  assign n480 = n470 & n479;
  assign n281 = n57 & ~n158;
  assign n481 = ~n188 & ~n281;
  assign n482 = n123 & ~n262;
  assign n483 = n481 & n482;
  assign n484 = n56 & ~n483;
  assign n486 = ~n286 & ~n485;
  assign n344 = n91 & n146;
  assign n345 = n165 & ~n344;
  assign n487 = ~n278 & ~n345;
  assign n336 = n85 & ~n137;
  assign n488 = n85 & ~n146;
  assign n489 = ~n336 & ~n488;
  assign n490 = n487 & n489;
  assign n491 = n486 & n490;
  assign n492 = ~n484 & n491;
  assign n493 = n480 & n492;
  assign n494 = n460 & n493;
  assign n495 = ~n152 & ~n165;
  assign n496 = ~n236 & ~n495;
  assign n497 = n101 & ~n123;
  assign n498 = n51 & ~n243;
  assign n499 = ~n497 & ~n498;
  assign n500 = ~n496 & n499;
  assign n501 = ~n131 & n500;
  assign n504 = ~n129 & ~n503;
  assign n506 = ~n111 & n140;
  assign n507 = n128 & n506;
  assign n508 = n130 & ~n507;
  assign n509 = ~n505 & ~n508;
  assign n510 = n504 & n509;
  assign n511 = n501 & n510;
  assign n513 = n57 & ~n512;
  assign n514 = ~n274 & ~n513;
  assign n515 = ~n200 & ~n418;
  assign n516 = n514 & n515;
  assign n517 = n511 & n516;
  assign n518 = n494 & n517;
  assign n703 = ~n220 & ~n341;
  assign n704 = ~n374 & n703;
  assign n705 = n691 & n704;
  assign n706 = n116 & n219;
  assign n707 = n58 & n706;
  assign n708 = ~n85 & ~n111;
  assign n709 = ~n289 & n708;
  assign n710 = ~n707 & ~n709;
  assign n711 = n705 & ~n710;
  assign n714 = n712 & n713;
  assign n715 = ~n225 & ~n418;
  assign n716 = n656 & n715;
  assign n717 = n714 & n716;
  assign n718 = n711 & n717;
  assign n719 = n373 & ~n567;
  assign n720 = ~n216 & ~n660;
  assign n722 = ~n224 & n721;
  assign n723 = n720 & n722;
  assign n724 = n719 & n723;
  assign n725 = ~n508 & n724;
  assign n726 = ~n192 & ~n200;
  assign n727 = n692 & n726;
  assign n729 = ~n382 & ~n728;
  assign n731 = ~n367 & n730;
  assign n732 = n729 & n731;
  assign n733 = n727 & n732;
  assign n201 = n116 & n158;
  assign n734 = n101 & ~n201;
  assign n735 = ~n195 & ~n734;
  assign n736 = ~n463 & n735;
  assign n737 = ~n563 & ~n645;
  assign n738 = ~n281 & n737;
  assign n739 = n736 & n738;
  assign n740 = n733 & n739;
  assign n741 = n725 & n740;
  assign n742 = n718 & n741;
  assign n743 = n702 & n742;
  assign n744 = ~n518 & ~n743;
  assign n1326 = ~n699 & ~n744;
  assign n2320 = n1326 ^ n315;
  assign n2321 = n1697 & n2320;
  assign n2322 = n2321 ^ n312;
  assign n2323 = n2322 ^ n308;
  assign n2324 = ~n786 & n2323;
  assign n2336 = n2335 ^ n2324;
  assign n966 = ~n812 & n965;
  assign n967 = ~n964 & ~n966;
  assign n1952 = n989 ^ n812;
  assign n2054 = ~n967 & n1952;
  assign n858 = n855 ^ n699;
  assign n2055 = n1079 ^ n812;
  assign n2056 = n858 & n2055;
  assign n2057 = ~n2054 & ~n2056;
  assign n1134 = n800 & ~n1068;
  assign n2050 = n864 & n1134;
  assign n1072 = n800 ^ n786;
  assign n2051 = n308 & n1072;
  assign n2052 = n2051 ^ n786;
  assign n2053 = ~n2050 & n2052;
  assign n2058 = n2057 ^ n2053;
  assign n1907 = n864 ^ n812;
  assign n1951 = ~n967 & ~n1907;
  assign n1953 = n858 & n1952;
  assign n1954 = ~n1951 & ~n1953;
  assign n1950 = n312 & ~n786;
  assign n1955 = n1954 ^ n1950;
  assign n746 = n518 & n743;
  assign n1946 = n746 & ~n1079;
  assign n1947 = n1326 & ~n1946;
  assign n745 = n699 & n744;
  assign n1948 = n745 & ~n1079;
  assign n1949 = ~n1947 & ~n1948;
  assign n2047 = n1950 ^ n1949;
  assign n2048 = n1955 & ~n2047;
  assign n2049 = n2048 ^ n1954;
  assign n2317 = n2057 ^ n2049;
  assign n2318 = ~n2058 & n2317;
  assign n2319 = n2318 ^ n2049;
  assign n2337 = n2336 ^ n2319;
  assign n2414 = n308 & ~n2335;
  assign n2415 = n2337 & n2414;
  assign n2416 = ~n2319 & n2322;
  assign n2417 = ~n2415 & ~n2416;
  assign n2418 = ~n786 & ~n2417;
  assign n2419 = n2322 ^ n2319;
  assign n2420 = n2323 & ~n2419;
  assign n2421 = ~n786 & n2420;
  assign n2422 = n2421 ^ n2319;
  assign n2423 = n2335 & ~n2422;
  assign n2424 = ~n2418 & ~n2423;
  assign n2397 = n786 & n2394;
  assign n2398 = n2388 & ~n2393;
  assign n2399 = ~n308 & n2398;
  assign n2400 = ~n2397 & ~n2399;
  assign n2401 = n2330 & ~n2400;
  assign n2402 = ~n2396 & ~n2401;
  assign n2410 = ~n2397 & ~n2409;
  assign n2411 = ~n2334 & ~n2410;
  assign n2412 = ~n2408 & ~n2411;
  assign n2413 = n2402 & n2412;
  assign n2425 = n2424 ^ n2413;
  assign n749 = ~x22 & ~n29;
  assign n750 = n749 ^ x6;
  assign n1647 = n750 & ~n786;
  assign n906 = ~n50 & ~n99;
  assign n323 = n69 & n146;
  assign n907 = ~n323 & ~n813;
  assign n908 = n170 & ~n907;
  assign n909 = ~n906 & ~n908;
  assign n910 = ~n497 & ~n909;
  assign n911 = n56 & ~n150;
  assign n912 = ~n51 & ~n911;
  assign n913 = ~n128 & ~n912;
  assign n914 = ~n271 & ~n423;
  assign n915 = ~n336 & n914;
  assign n916 = ~n273 & n915;
  assign n917 = ~n687 & n916;
  assign n918 = ~n913 & n917;
  assign n551 = ~n299 & ~n463;
  assign n552 = ~n129 & ~n394;
  assign n553 = n551 & n552;
  assign n919 = n164 & n680;
  assign n920 = ~n220 & ~n261;
  assign n921 = ~n919 & n920;
  assign n922 = ~n199 & n921;
  assign n923 = n676 & n922;
  assign n924 = n553 & n923;
  assign n925 = n918 & n924;
  assign n926 = n910 & n925;
  assign n342 = ~n340 & ~n341;
  assign n346 = ~n343 & ~n345;
  assign n347 = n342 & n346;
  assign n930 = n648 & n929;
  assign n931 = n347 & n930;
  assign n932 = ~n272 & ~n442;
  assign n933 = n116 & n123;
  assign n934 = n83 & ~n933;
  assign n935 = n932 & ~n934;
  assign n609 = ~n299 & ~n523;
  assign n936 = ~n238 & ~n589;
  assign n937 = n609 & n936;
  assign n938 = n935 & n937;
  assign n939 = n931 & n938;
  assign n948 = ~n183 & ~n488;
  assign n949 = n776 & n933;
  assign n950 = n57 & ~n949;
  assign n951 = ~n221 & ~n950;
  assign n952 = n948 & n951;
  assign n953 = n369 & n952;
  assign n954 = n947 & n953;
  assign n955 = n939 & n954;
  assign n956 = n926 & n955;
  assign n189 = n78 & ~n188;
  assign n190 = ~n83 & ~n152;
  assign n191 = ~n189 & ~n190;
  assign n193 = ~n112 & ~n192;
  assign n194 = ~n191 & n193;
  assign n196 = ~n50 & ~n57;
  assign n197 = ~n170 & ~n196;
  assign n198 = ~n195 & ~n197;
  assign n202 = n152 & ~n201;
  assign n203 = ~n200 & ~n202;
  assign n204 = n128 & n155;
  assign n205 = n130 & ~n204;
  assign n206 = n203 & ~n205;
  assign n207 = ~n199 & n206;
  assign n208 = n198 & n207;
  assign n209 = n194 & n208;
  assign n210 = ~n83 & n209;
  assign n213 = ~n101 & ~n111;
  assign n214 = ~n212 & n213;
  assign n215 = ~n210 & ~n214;
  assign n228 = n69 & n123;
  assign n229 = ~n85 & n228;
  assign n230 = ~n227 & ~n229;
  assign n425 = ~n423 & ~n424;
  assign n426 = ~n422 & n425;
  assign n427 = ~n245 & n426;
  assign n522 = n427 & n521;
  assign n524 = n85 & ~n201;
  assign n525 = ~n263 & ~n524;
  assign n526 = ~n278 & n525;
  assign n527 = ~n523 & n526;
  assign n528 = ~n85 & n236;
  assign n529 = n69 & n140;
  assign n530 = ~n56 & n529;
  assign n531 = ~n528 & ~n530;
  assign n532 = ~n274 & ~n531;
  assign n325 = n116 & n155;
  assign n533 = n152 & ~n325;
  assign n534 = n532 & ~n533;
  assign n535 = n527 & n534;
  assign n536 = n522 & n535;
  assign n537 = ~n230 & n536;
  assign n538 = ~n215 & n537;
  assign n540 = ~n396 & ~n410;
  assign n541 = ~n539 & n540;
  assign n542 = n257 & n541;
  assign n543 = ~n330 & ~n464;
  assign n544 = ~n131 & n543;
  assign n546 = ~n287 & ~n545;
  assign n547 = ~n271 & ~n464;
  assign n548 = n546 & n547;
  assign n549 = n544 & n548;
  assign n550 = n542 & n549;
  assign n554 = n383 & n553;
  assign n555 = n365 & n554;
  assign n556 = n550 & n555;
  assign n558 = ~n57 & ~n272;
  assign n559 = ~n172 & ~n558;
  assign n560 = n557 & ~n559;
  assign n561 = n85 & ~n147;
  assign n562 = ~n331 & ~n561;
  assign n564 = ~n413 & ~n563;
  assign n565 = n562 & n564;
  assign n566 = n560 & n565;
  assign n568 = n369 & ~n567;
  assign n570 = ~n340 & ~n497;
  assign n571 = ~n569 & n570;
  assign n572 = n568 & n571;
  assign n573 = n566 & n572;
  assign n574 = n556 & n573;
  assign n575 = n538 & n574;
  assign n993 = n454 & n562;
  assign n411 = n101 & ~n158;
  assign n994 = ~n180 & ~n411;
  assign n995 = n993 & n994;
  assign n996 = ~n353 & ~n645;
  assign n997 = n360 & n996;
  assign n999 = ~n289 & ~n998;
  assign n1000 = ~n239 & ~n688;
  assign n1001 = n999 & n1000;
  assign n1002 = n997 & n1001;
  assign n1003 = n995 & n1002;
  assign n222 = ~n220 & ~n221;
  assign n223 = ~n216 & n222;
  assign n877 = ~n262 & ~n367;
  assign n584 = ~n111 & n155;
  assign n1004 = n97 & n584;
  assign n1005 = n85 & ~n1004;
  assign n1006 = n877 & ~n1005;
  assign n1007 = n223 & n1006;
  assign n1008 = n1003 & n1007;
  assign n1009 = n910 & n1008;
  assign n1010 = n83 & ~n243;
  assign n1011 = n871 & ~n1010;
  assign n1012 = n260 & n1011;
  assign n1013 = n543 & n1012;
  assign n1014 = n141 & n171;
  assign n1015 = ~n57 & n1014;
  assign n1016 = n171 & n176;
  assign n1017 = n40 & ~n48;
  assign n1018 = ~n1016 & n1017;
  assign n1019 = ~n1015 & n1018;
  assign n610 = ~n224 & ~n374;
  assign n1020 = ~n148 & n152;
  assign n1021 = ~n394 & ~n1020;
  assign n1022 = n158 & n236;
  assign n1023 = n56 & ~n1022;
  assign n1024 = n1021 & ~n1023;
  assign n1025 = n610 & n1024;
  assign n1026 = ~n1019 & n1025;
  assign n1027 = n1013 & n1026;
  assign n888 = ~n50 & ~n152;
  assign n1028 = ~n273 & ~n442;
  assign n1029 = n266 & n1028;
  assign n1030 = ~n888 & ~n1029;
  assign n1031 = n1027 & ~n1030;
  assign n1035 = n165 & ~n1016;
  assign n1036 = ~n468 & ~n1035;
  assign n1037 = n91 & n228;
  assign n1038 = n51 & ~n1037;
  assign n1039 = ~n244 & ~n1038;
  assign n1040 = n1036 & n1039;
  assign n1041 = n1034 & n1040;
  assign n1042 = n1031 & n1041;
  assign n1043 = n1009 & n1042;
  assign n1424 = ~n575 & n1043;
  assign n1425 = ~n956 & n1424;
  assign n1426 = n575 & n956;
  assign n1427 = ~n1425 & ~n1426;
  assign n1044 = ~n956 & ~n1043;
  assign n1045 = n575 & n1044;
  assign n1046 = n956 & n1043;
  assign n1433 = ~n1045 & ~n1046;
  assign n1491 = ~n1079 & ~n1433;
  assign n1492 = n1427 & ~n1491;
  assign n1649 = n956 & ~n1492;
  assign n968 = ~x22 & ~n28;
  assign n969 = n968 ^ x5;
  assign n1490 = ~n786 & n969;
  assign n1650 = ~n1490 & ~n1491;
  assign n1651 = ~n1649 & ~n1650;
  assign n1652 = ~n1425 & n1651;
  assign n1825 = ~n1647 & n1652;
  assign n747 = ~n699 & n746;
  assign n748 = ~n745 & ~n747;
  assign n1503 = n699 ^ n308;
  assign n1643 = ~n748 & ~n1503;
  assign n753 = n743 ^ n518;
  assign n1644 = n864 ^ n699;
  assign n1645 = n753 & ~n1644;
  assign n1646 = ~n1643 & ~n1645;
  assign n1826 = n1647 ^ n1426;
  assign n1827 = ~n1651 & n1826;
  assign n1828 = ~n1646 & ~n1827;
  assign n1829 = ~n1825 & ~n1828;
  assign n1830 = n1646 & ~n1647;
  assign n1831 = n1425 & ~n1830;
  assign n1832 = n1829 & ~n1831;
  assign n1675 = n812 ^ n315;
  assign n1818 = ~n967 & ~n1675;
  assign n1819 = n812 ^ n308;
  assign n1820 = n858 & ~n1819;
  assign n1821 = ~n1818 & ~n1820;
  assign n309 = ~x22 & ~n31;
  assign n310 = n309 ^ x8;
  assign n1811 = ~n310 & ~n786;
  assign n1812 = n1068 & ~n1811;
  assign n1813 = ~n312 & n1070;
  assign n1814 = ~n310 & ~n800;
  assign n1815 = ~n1813 & ~n1814;
  assign n1816 = ~n1812 & n1815;
  assign n1809 = n1427 & ~n1647;
  assign n1810 = n1809 ^ n1425;
  assign n1817 = n1816 ^ n1810;
  assign n1822 = n1821 ^ n1817;
  assign n1804 = ~n748 & ~n1644;
  assign n1805 = n989 ^ n699;
  assign n1806 = n753 & n1805;
  assign n1807 = ~n1804 & ~n1806;
  assign n754 = x6 & ~x22;
  assign n755 = ~n749 & ~n754;
  assign n756 = n755 ^ x7;
  assign n1802 = ~n756 & ~n786;
  assign n576 = ~n188 & ~n366;
  assign n578 = ~n463 & ~n577;
  assign n579 = n576 & n578;
  assign n580 = ~n195 & ~n220;
  assign n581 = n557 & n580;
  assign n582 = n579 & n581;
  assign n583 = n347 & n582;
  assign n585 = n165 & ~n584;
  assign n586 = ~n353 & ~n585;
  assign n587 = ~n398 & n586;
  assign n588 = ~n394 & n587;
  assign n590 = ~n496 & ~n589;
  assign n591 = n427 & n590;
  assign n592 = n588 & n591;
  assign n593 = n583 & n592;
  assign n594 = ~n244 & ~n264;
  assign n596 = ~n280 & ~n322;
  assign n597 = ~n595 & n596;
  assign n598 = n594 & n597;
  assign n599 = n179 & n598;
  assign n601 = ~n40 & ~n164;
  assign n602 = ~n170 & n601;
  assign n603 = ~n485 & ~n602;
  assign n604 = ~n600 & n603;
  assign n605 = n599 & n604;
  assign n405 = n101 & ~n404;
  assign n606 = ~n289 & ~n405;
  assign n607 = ~n334 & ~n382;
  assign n608 = n606 & n607;
  assign n611 = n609 & n610;
  assign n612 = n608 & n611;
  assign n614 = n116 & n512;
  assign n615 = n130 & ~n614;
  assign n616 = ~n613 & ~n615;
  assign n618 = n51 & ~n617;
  assign n619 = n85 & ~n123;
  assign n620 = ~n618 & ~n619;
  assign n621 = n616 & n620;
  assign n622 = n458 & n621;
  assign n623 = n612 & n622;
  assign n624 = n605 & n623;
  assign n625 = n593 & n624;
  assign n626 = ~n575 & ~n625;
  assign n1212 = ~n518 & ~n626;
  assign n628 = n575 & n625;
  assign n1798 = n628 & ~n1079;
  assign n1799 = n1212 & ~n1798;
  assign n627 = n518 & n626;
  assign n1800 = n627 & ~n1079;
  assign n1801 = ~n1799 & ~n1800;
  assign n1803 = n1802 ^ n1801;
  assign n1808 = n1807 ^ n1803;
  assign n1823 = n1822 ^ n1808;
  assign n629 = ~n518 & n628;
  assign n630 = ~n627 & ~n629;
  assign n1499 = n989 ^ n518;
  assign n1683 = ~n630 & n1499;
  assign n633 = n625 ^ n575;
  assign n1684 = n1079 ^ n518;
  assign n1685 = n633 & n1684;
  assign n1686 = ~n1683 & ~n1685;
  assign n1069 = n786 & n1068;
  assign n1678 = ~n310 & n1070;
  assign n1679 = n756 & n1072;
  assign n1680 = n1679 ^ n786;
  assign n1681 = ~n1678 & n1680;
  assign n1682 = ~n1069 & n1681;
  assign n1687 = n1686 ^ n1682;
  assign n1495 = n812 ^ n312;
  assign n1674 = ~n967 & ~n1495;
  assign n1676 = n858 & ~n1675;
  assign n1677 = ~n1674 & ~n1676;
  assign n1795 = n1686 ^ n1677;
  assign n1796 = n1687 & n1795;
  assign n1797 = n1796 ^ n1677;
  assign n1824 = n1823 ^ n1797;
  assign n1833 = n1832 ^ n1824;
  assign n1688 = n1687 ^ n1677;
  assign n1418 = n699 ^ n315;
  assign n1502 = ~n748 & ~n1418;
  assign n1504 = n753 & ~n1503;
  assign n1505 = ~n1502 & ~n1504;
  assign n1414 = n864 ^ n518;
  assign n1498 = ~n630 & ~n1414;
  assign n1500 = n633 & n1499;
  assign n1501 = ~n1498 & ~n1500;
  assign n1506 = n1505 ^ n1501;
  assign n1410 = n812 ^ n310;
  assign n1494 = ~n967 & ~n1410;
  assign n1496 = n858 & ~n1495;
  assign n1497 = ~n1494 & ~n1496;
  assign n1671 = n1505 ^ n1497;
  assign n1672 = ~n1506 & n1671;
  assign n1673 = n1672 ^ n1497;
  assign n1689 = n1688 ^ n1673;
  assign n1481 = ~n756 & n1134;
  assign n1482 = n750 & n1072;
  assign n1483 = n1482 ^ n786;
  assign n1484 = ~n1481 & n1483;
  assign n1112 = n699 ^ n312;
  assign n1417 = ~n748 & ~n1112;
  assign n1419 = n753 & ~n1418;
  assign n1420 = ~n1417 & ~n1419;
  assign n1108 = n518 ^ n308;
  assign n1413 = ~n630 & ~n1108;
  assign n1415 = n633 & ~n1414;
  assign n1416 = ~n1413 & ~n1415;
  assign n1421 = n1420 ^ n1416;
  assign n1104 = n812 ^ n756;
  assign n1409 = ~n967 & n1104;
  assign n1411 = n858 & ~n1410;
  assign n1412 = ~n1409 & ~n1411;
  assign n1478 = n1420 ^ n1412;
  assign n1479 = ~n1421 & n1478;
  assign n1480 = n1479 ^ n1412;
  assign n1485 = n1484 ^ n1480;
  assign n1428 = n1079 & ~n1427;
  assign n1247 = ~n575 & ~n1044;
  assign n1429 = ~n1043 & ~n1247;
  assign n1430 = ~n1079 & ~n1424;
  assign n1431 = ~n1429 & n1430;
  assign n1432 = ~n1428 & ~n1431;
  assign n1434 = ~n989 & ~n1433;
  assign n1435 = n1432 & ~n1434;
  assign n1056 = ~x22 & ~n27;
  assign n1057 = n1056 ^ x4;
  assign n1423 = ~n786 & n1057;
  assign n1436 = n1435 ^ n1423;
  assign n1468 = n1423 ^ n956;
  assign n1469 = ~n1043 & ~n1468;
  assign n1470 = n1469 ^ n956;
  assign n1471 = ~n1436 & ~n1470;
  assign n1472 = ~n989 & n1045;
  assign n1473 = ~n1423 & ~n1472;
  assign n1474 = n989 & n1424;
  assign n1475 = n956 & ~n1474;
  assign n1476 = ~n1473 & ~n1475;
  assign n1477 = ~n1471 & ~n1476;
  assign n1668 = n1484 ^ n1477;
  assign n1669 = n1485 & ~n1668;
  assign n1670 = n1669 ^ n1480;
  assign n1792 = n1673 ^ n1670;
  assign n1793 = n1689 & n1792;
  assign n1794 = n1793 ^ n1670;
  assign n1834 = n1833 ^ n1794;
  assign n1653 = ~n1426 & ~n1652;
  assign n1648 = n1647 ^ n1646;
  assign n1654 = n1653 ^ n1648;
  assign n1507 = n1506 ^ n1497;
  assign n1493 = n1492 ^ n1490;
  assign n1508 = n1507 ^ n1493;
  assign n1446 = n750 & n1134;
  assign n1447 = n969 & n1072;
  assign n1448 = n1447 ^ n786;
  assign n1449 = ~n1446 & n1448;
  assign n1047 = ~n575 & n1046;
  assign n1048 = ~n1045 & ~n1047;
  assign n1087 = n864 ^ n575;
  assign n1097 = ~n1048 & ~n1087;
  assign n1051 = n1043 ^ n956;
  assign n1098 = n989 ^ n575;
  assign n1099 = n1051 & n1098;
  assign n1100 = ~n1097 & ~n1099;
  assign n859 = ~x22 & ~n26;
  assign n860 = n859 ^ x3;
  assign n1095 = ~n786 & n860;
  assign n1442 = n1100 ^ n1095;
  assign n876 = ~n567 & n875;
  assign n878 = ~n359 & n877;
  assign n880 = ~n216 & ~n272;
  assign n881 = n879 & n880;
  assign n882 = n878 & n881;
  assign n883 = n662 & n882;
  assign n884 = n101 & ~n506;
  assign n885 = ~n264 & ~n884;
  assign n886 = ~n274 & n885;
  assign n887 = ~n299 & ~n613;
  assign n889 = ~n137 & ~n888;
  assign n890 = n887 & ~n889;
  assign n891 = n886 & n890;
  assign n892 = n883 & n891;
  assign n893 = n78 & ~n111;
  assign n894 = ~n40 & ~n893;
  assign n895 = ~n100 & ~n894;
  assign n896 = ~n601 & ~n893;
  assign n897 = n146 & ~n896;
  assign n898 = ~n895 & ~n897;
  assign n899 = n130 & ~n317;
  assign n900 = ~n418 & ~n899;
  assign n901 = ~n898 & n900;
  assign n902 = n765 & n901;
  assign n903 = n892 & n902;
  assign n904 = n876 & n903;
  assign n1093 = n904 & ~n1079;
  assign n1094 = ~n956 & ~n1093;
  assign n1443 = n1100 ^ n1094;
  assign n1444 = ~n1442 & n1443;
  assign n1445 = n1444 ^ n1095;
  assign n1450 = n1449 ^ n1445;
  assign n980 = n699 ^ n310;
  assign n1111 = ~n748 & ~n980;
  assign n1113 = n753 & ~n1112;
  assign n1114 = ~n1111 & ~n1113;
  assign n976 = n518 ^ n315;
  assign n1107 = ~n630 & ~n976;
  assign n1109 = n633 & ~n1108;
  assign n1110 = ~n1107 & ~n1109;
  assign n1115 = n1114 ^ n1110;
  assign n972 = n812 ^ n750;
  assign n1103 = ~n967 & ~n972;
  assign n1105 = n858 & n1104;
  assign n1106 = ~n1103 & ~n1105;
  assign n1439 = n1114 ^ n1106;
  assign n1440 = ~n1115 & n1439;
  assign n1441 = n1440 ^ n1106;
  assign n1487 = n1449 ^ n1441;
  assign n1488 = ~n1450 & ~n1487;
  assign n1489 = n1488 ^ n1445;
  assign n1640 = n1507 ^ n1489;
  assign n1641 = n1508 & ~n1640;
  assign n1642 = n1641 ^ n1489;
  assign n1655 = n1654 ^ n1642;
  assign n1509 = n1508 ^ n1489;
  assign n1486 = n1485 ^ n1477;
  assign n1510 = n1509 ^ n1486;
  assign n1422 = n1421 ^ n1412;
  assign n1437 = n1436 ^ n1422;
  assign n1080 = ~n904 & ~n1079;
  assign n1081 = n1080 ^ n956;
  assign n1082 = n904 & ~n989;
  assign n1083 = ~n1081 & ~n1082;
  assign n1128 = ~n786 & n1083;
  assign n1121 = ~n786 & ~n1057;
  assign n1122 = n1068 & ~n1121;
  assign n1123 = n786 & ~n969;
  assign n1124 = n1123 ^ n1057;
  assign n1125 = n800 & ~n1124;
  assign n1126 = n1125 ^ n1057;
  assign n1127 = ~n1122 & n1126;
  assign n1129 = n1128 ^ n1127;
  assign n757 = n756 ^ n699;
  assign n979 = ~n748 & n757;
  assign n981 = n753 & ~n980;
  assign n982 = ~n979 & ~n981;
  assign n634 = n518 ^ n312;
  assign n975 = ~n630 & ~n634;
  assign n977 = n633 & ~n976;
  assign n978 = ~n975 & ~n977;
  assign n983 = n982 ^ n978;
  assign n970 = n969 ^ n812;
  assign n971 = ~n967 & ~n970;
  assign n973 = n858 & ~n972;
  assign n974 = ~n971 & ~n973;
  assign n1118 = n982 ^ n974;
  assign n1119 = ~n983 & n1118;
  assign n1120 = n1119 ^ n974;
  assign n1406 = n1128 ^ n1120;
  assign n1407 = ~n1129 & ~n1406;
  assign n1408 = n1407 ^ n1120;
  assign n1465 = n1422 ^ n1408;
  assign n1466 = n1437 & n1465;
  assign n1467 = n1466 ^ n1408;
  assign n1637 = n1509 ^ n1467;
  assign n1638 = ~n1510 & n1637;
  assign n1639 = n1638 ^ n1467;
  assign n1784 = n1642 ^ n1639;
  assign n1785 = n1655 & ~n1784;
  assign n1786 = n1785 ^ n1639;
  assign n1511 = n1510 ^ n1467;
  assign n1451 = n1450 ^ n1441;
  assign n1438 = n1437 ^ n1408;
  assign n1452 = n1451 ^ n1438;
  assign n1130 = n1129 ^ n1120;
  assign n1116 = n1115 ^ n1106;
  assign n1096 = n1095 ^ n1094;
  assign n1101 = n1100 ^ n1096;
  assign n1084 = n1083 ^ n786;
  assign n1071 = ~n1057 & n1070;
  assign n1073 = ~n860 & n1072;
  assign n1074 = n1073 ^ n786;
  assign n1075 = ~n1071 & n1074;
  assign n1076 = ~n1069 & n1075;
  assign n1085 = n1084 ^ n1076;
  assign n1052 = n575 ^ n308;
  assign n1086 = ~n1048 & ~n1052;
  assign n1088 = n1051 & ~n1087;
  assign n1089 = ~n1086 & ~n1088;
  assign n1090 = n1089 ^ n1084;
  assign n1091 = n1085 & n1090;
  assign n1092 = n1091 ^ n1089;
  assign n1102 = n1101 ^ n1092;
  assign n1117 = n1116 ^ n1102;
  assign n1131 = n1130 ^ n1117;
  assign n984 = n983 ^ n974;
  assign n751 = n750 ^ n699;
  assign n752 = ~n748 & ~n751;
  assign n758 = n753 & n757;
  assign n759 = ~n752 & ~n758;
  assign n631 = n518 ^ n310;
  assign n632 = ~n630 & ~n631;
  assign n635 = n633 & ~n634;
  assign n636 = ~n632 & ~n635;
  assign n760 = n759 ^ n636;
  assign n861 = n858 & n860;
  assign n862 = n857 & ~n861;
  assign n905 = n864 & ~n904;
  assign n957 = n956 ^ n905;
  assign n958 = n308 & n904;
  assign n959 = ~n957 & ~n958;
  assign n960 = n862 & n959;
  assign n961 = n960 ^ n636;
  assign n962 = n760 & n961;
  assign n963 = n962 ^ n759;
  assign n985 = n984 ^ n963;
  assign n1049 = n575 ^ n315;
  assign n1050 = ~n1048 & ~n1049;
  assign n1053 = n1051 & ~n1052;
  assign n1054 = ~n1050 & ~n1053;
  assign n986 = n864 & n904;
  assign n990 = ~n904 & ~n989;
  assign n991 = n990 ^ n956;
  assign n992 = ~n986 & ~n991;
  assign n1055 = n1054 ^ n992;
  assign n1058 = n1057 ^ n812;
  assign n1059 = ~n967 & ~n1058;
  assign n1060 = n858 & ~n970;
  assign n1061 = ~n1059 & ~n1060;
  assign n1062 = n1061 ^ n1054;
  assign n1063 = n1055 & n1062;
  assign n1064 = n1063 ^ n1061;
  assign n1065 = n1064 ^ n984;
  assign n1066 = n985 & ~n1065;
  assign n1067 = n1066 ^ n963;
  assign n1453 = n1130 ^ n1067;
  assign n1454 = ~n1131 & n1453;
  assign n1455 = n1454 ^ n1067;
  assign n1456 = n1455 ^ n1451;
  assign n1457 = ~n1452 & ~n1456;
  assign n1458 = n1457 ^ n1455;
  assign n1132 = n1131 ^ n1067;
  assign n1133 = n1064 ^ n985;
  assign n1136 = n960 ^ n760;
  assign n1135 = n860 & n1134;
  assign n1137 = n1136 ^ n1135;
  assign n1142 = n756 ^ n518;
  assign n1143 = ~n630 & n1142;
  assign n1144 = ~n631 & n633;
  assign n1145 = ~n1143 & ~n1144;
  assign n1138 = n575 ^ n312;
  assign n1139 = ~n1048 & ~n1138;
  assign n1140 = ~n1049 & n1051;
  assign n1141 = ~n1139 & ~n1140;
  assign n1146 = n1145 ^ n1141;
  assign n1147 = n969 ^ n699;
  assign n1148 = ~n748 & ~n1147;
  assign n1149 = ~n751 & n753;
  assign n1150 = ~n1148 & ~n1149;
  assign n1151 = n1150 ^ n1145;
  assign n1152 = ~n1146 & n1151;
  assign n1153 = n1152 ^ n1150;
  assign n1154 = n1153 ^ n1135;
  assign n1155 = n1137 & n1154;
  assign n1156 = n1155 ^ n1136;
  assign n1157 = ~n1133 & n1156;
  assign n1158 = n1132 & ~n1157;
  assign n1200 = n750 ^ n575;
  assign n1201 = ~n1048 & ~n1200;
  assign n1202 = n756 ^ n575;
  assign n1203 = n1051 & n1202;
  assign n1204 = ~n1201 & ~n1203;
  assign n1195 = n1057 ^ n518;
  assign n1196 = ~n630 & ~n1195;
  assign n1197 = n969 ^ n518;
  assign n1198 = n633 & ~n1197;
  assign n1199 = ~n1196 & ~n1198;
  assign n1205 = n1204 ^ n1199;
  assign n1191 = n312 & ~n904;
  assign n1192 = n1191 ^ n956;
  assign n1193 = n310 & n904;
  assign n1194 = ~n1192 & ~n1193;
  assign n1206 = n1205 ^ n1194;
  assign n1207 = n627 & n860;
  assign n1208 = n633 & ~n1195;
  assign n1209 = ~n1207 & ~n1208;
  assign n1210 = n629 & ~n860;
  assign n1211 = n1209 & ~n1210;
  assign n1213 = n633 & n860;
  assign n1214 = n1212 & ~n1213;
  assign n1215 = ~n1211 & n1214;
  assign n1216 = n969 ^ n575;
  assign n1217 = ~n1048 & ~n1216;
  assign n1218 = n1051 & ~n1200;
  assign n1219 = ~n1217 & ~n1218;
  assign n1220 = ~n756 & n904;
  assign n1221 = n956 ^ n310;
  assign n1222 = n1221 ^ n1193;
  assign n1223 = ~n1220 & ~n1222;
  assign n1231 = ~n1219 & n1223;
  assign n1229 = n753 & n860;
  assign n1224 = n1223 ^ n1219;
  assign n1225 = n1211 & ~n1214;
  assign n1226 = n1225 ^ n1223;
  assign n1227 = ~n1224 & n1226;
  assign n1228 = n1227 ^ n1219;
  assign n1230 = n1229 ^ n1228;
  assign n1232 = n1231 ^ n1230;
  assign n1233 = ~n1215 & n1232;
  assign n1234 = n1233 ^ n1231;
  assign n1235 = n1206 & ~n1234;
  assign n1236 = n1214 ^ n1211;
  assign n1237 = n1236 ^ n1224;
  assign n1242 = n1057 ^ n575;
  assign n1243 = ~n1048 & ~n1242;
  assign n1244 = n1051 & ~n1216;
  assign n1245 = ~n1243 & ~n1244;
  assign n1238 = n750 & n904;
  assign n1239 = n956 ^ n756;
  assign n1240 = n1239 ^ n1220;
  assign n1241 = ~n1238 & n1240;
  assign n1246 = n1245 ^ n1241;
  assign n1248 = n860 & ~n1046;
  assign n1249 = n1247 & ~n1248;
  assign n1250 = n904 & n969;
  assign n1251 = n956 ^ n750;
  assign n1252 = n1251 ^ n1238;
  assign n1253 = ~n1250 & ~n1252;
  assign n1254 = n1249 & n1253;
  assign n1255 = n1254 ^ n1241;
  assign n1256 = ~n1246 & ~n1255;
  assign n1257 = n1256 ^ n1245;
  assign n1258 = n1237 & ~n1257;
  assign n1259 = ~n1235 & ~n1258;
  assign n1260 = ~n1213 & ~n1249;
  assign n1261 = ~n1246 & ~n1260;
  assign n1262 = ~n1253 & ~n1261;
  assign n1263 = ~n860 & n1047;
  assign n1264 = n1051 & ~n1242;
  assign n1265 = ~n1263 & ~n1264;
  assign n1266 = n860 & n1045;
  assign n1267 = n1265 & ~n1266;
  assign n1268 = n1246 & n1267;
  assign n1269 = ~n1249 & n1268;
  assign n1270 = ~n1262 & ~n1269;
  assign n1271 = ~n1246 & ~n1267;
  assign n1272 = ~n1213 & ~n1271;
  assign n1273 = n1270 & ~n1272;
  assign n1274 = ~n860 & n1057;
  assign n1275 = ~n956 & ~n1274;
  assign n1276 = n904 & n1057;
  assign n1277 = n1275 & ~n1276;
  assign n1278 = n860 & ~n1043;
  assign n1279 = ~n904 & n969;
  assign n1280 = ~n1278 & ~n1279;
  assign n1281 = n1277 & n1280;
  assign n1282 = n956 & n1279;
  assign n1283 = n1278 & n1282;
  assign n1284 = ~n1281 & ~n1283;
  assign n1285 = ~n1273 & n1284;
  assign n1286 = ~n1268 & ~n1272;
  assign n1287 = ~n1253 & ~n1286;
  assign n1288 = n1241 & ~n1245;
  assign n1289 = ~n1237 & ~n1288;
  assign n1290 = n1246 & n1260;
  assign n1291 = ~n1289 & ~n1290;
  assign n1292 = ~n1287 & n1291;
  assign n1293 = ~n1285 & n1292;
  assign n1294 = n1259 & ~n1293;
  assign n1295 = ~n1206 & n1234;
  assign n1296 = ~n1294 & ~n1295;
  assign n1297 = n1215 & n1231;
  assign n1298 = ~n1228 & n1229;
  assign n1299 = ~n1297 & ~n1298;
  assign n1300 = n1199 ^ n1194;
  assign n1301 = n1205 & n1300;
  assign n1302 = n1301 ^ n1204;
  assign n1303 = ~n1299 & ~n1302;
  assign n1304 = ~n1296 & ~n1303;
  assign n1305 = n1299 & n1302;
  assign n1175 = n750 ^ n518;
  assign n1176 = ~n630 & ~n1175;
  assign n1177 = n633 & n1142;
  assign n1178 = ~n1176 & ~n1177;
  assign n1170 = n575 ^ n310;
  assign n1171 = ~n1048 & ~n1170;
  assign n1172 = n1051 & ~n1138;
  assign n1173 = ~n1171 & ~n1172;
  assign n1166 = n308 & ~n904;
  assign n1167 = n1166 ^ n956;
  assign n1168 = n315 & n904;
  assign n1169 = ~n1167 & ~n1168;
  assign n1174 = n1173 ^ n1169;
  assign n1334 = n1178 ^ n1174;
  assign n1327 = ~n860 & n1326;
  assign n1328 = ~n747 & ~n1327;
  assign n1329 = n315 & ~n904;
  assign n1330 = n1329 ^ n956;
  assign n1331 = n312 & n904;
  assign n1332 = ~n1330 & ~n1331;
  assign n1333 = ~n1328 & n1332;
  assign n1335 = n1334 ^ n1333;
  assign n1314 = n1057 ^ n699;
  assign n1322 = ~n748 & ~n1314;
  assign n1323 = n753 & ~n1147;
  assign n1324 = ~n1322 & ~n1323;
  assign n1325 = n1324 ^ n861;
  assign n1336 = n1335 ^ n1325;
  assign n1309 = ~n630 & ~n1197;
  assign n1310 = n633 & ~n1175;
  assign n1311 = ~n1309 & ~n1310;
  assign n1306 = ~n1048 & n1202;
  assign n1307 = n1051 & ~n1170;
  assign n1308 = ~n1306 & ~n1307;
  assign n1312 = n1311 ^ n1308;
  assign n1313 = n745 & n860;
  assign n1315 = n753 & ~n1314;
  assign n1316 = ~n1313 & ~n1315;
  assign n1317 = n747 & ~n860;
  assign n1318 = n1316 & ~n1317;
  assign n1319 = n1318 ^ n1308;
  assign n1320 = n1312 & ~n1319;
  assign n1321 = n1320 ^ n1311;
  assign n1337 = n1336 ^ n1321;
  assign n1338 = n1318 ^ n1312;
  assign n1339 = n1332 ^ n1328;
  assign n1340 = ~n1338 & ~n1339;
  assign n1341 = ~n1337 & ~n1340;
  assign n1342 = ~n1305 & ~n1341;
  assign n1343 = ~n1304 & n1342;
  assign n1344 = n1337 & n1340;
  assign n1345 = ~n1343 & ~n1344;
  assign n1346 = ~n1305 & n1337;
  assign n1347 = ~n1296 & ~n1346;
  assign n1348 = ~n1303 & ~n1337;
  assign n1349 = n1338 & n1339;
  assign n1350 = ~n1348 & ~n1349;
  assign n1351 = ~n1347 & n1350;
  assign n1352 = n1345 & ~n1351;
  assign n1353 = n1150 ^ n1146;
  assign n1354 = n1352 & n1353;
  assign n1355 = n1321 & ~n1334;
  assign n1356 = n1333 ^ n1324;
  assign n1357 = n1325 & ~n1356;
  assign n1358 = n1357 ^ n1333;
  assign n1359 = n1355 & ~n1358;
  assign n1360 = ~n1321 & n1334;
  assign n1361 = ~n861 & n1324;
  assign n1362 = ~n1333 & n1361;
  assign n1363 = ~n1360 & n1362;
  assign n1364 = ~n1359 & ~n1363;
  assign n1179 = n1178 ^ n1169;
  assign n1180 = ~n1174 & n1179;
  assign n1181 = n1180 ^ n1173;
  assign n1160 = n860 & n964;
  assign n1161 = n858 & ~n1058;
  assign n1162 = ~n1160 & ~n1161;
  assign n1163 = ~n860 & n966;
  assign n1164 = n1162 & ~n1163;
  assign n1159 = n959 ^ n862;
  assign n1165 = n1164 ^ n1159;
  assign n1365 = n1181 ^ n1165;
  assign n1366 = ~n1364 & ~n1365;
  assign n1187 = n1153 ^ n1137;
  assign n1185 = n1061 ^ n1055;
  assign n1182 = n1181 ^ n1164;
  assign n1183 = n1165 & n1182;
  assign n1184 = n1183 ^ n1181;
  assign n1186 = n1185 ^ n1184;
  assign n1367 = n1187 ^ n1186;
  assign n1368 = ~n1366 & n1367;
  assign n1369 = n1358 & n1360;
  assign n1370 = n861 & ~n1324;
  assign n1371 = n1333 & n1370;
  assign n1372 = ~n1355 & n1371;
  assign n1373 = ~n1369 & ~n1372;
  assign n1374 = n1365 & ~n1373;
  assign n1375 = ~n1368 & ~n1374;
  assign n1376 = ~n1354 & ~n1375;
  assign n1377 = n1364 & n1365;
  assign n1378 = n1373 & ~n1377;
  assign n1379 = ~n1367 & n1378;
  assign n1380 = ~n1353 & ~n1379;
  assign n1381 = ~n1352 & n1380;
  assign n1382 = n1367 & ~n1378;
  assign n1383 = ~n1381 & ~n1382;
  assign n1384 = ~n1376 & n1383;
  assign n1188 = n1187 ^ n1185;
  assign n1189 = ~n1186 & n1188;
  assign n1190 = n1189 ^ n1184;
  assign n1385 = n1384 ^ n1190;
  assign n1386 = n1089 ^ n1085;
  assign n1387 = n1386 ^ n1190;
  assign n1388 = n1385 & n1387;
  assign n1389 = n1388 ^ n1384;
  assign n1390 = ~n1158 & ~n1389;
  assign n1391 = n1190 & ~n1386;
  assign n1392 = ~n1132 & ~n1391;
  assign n1393 = n1384 & ~n1392;
  assign n1394 = ~n1190 & n1386;
  assign n1395 = n1132 & ~n1394;
  assign n1396 = n1133 & ~n1156;
  assign n1397 = ~n1395 & ~n1396;
  assign n1398 = ~n1393 & n1397;
  assign n1399 = ~n1132 & n1157;
  assign n1400 = ~n1398 & ~n1399;
  assign n1401 = ~n1390 & n1400;
  assign n1402 = n1116 ^ n1101;
  assign n1403 = n1102 & ~n1402;
  assign n1404 = n1403 ^ n1092;
  assign n1657 = n1401 & n1404;
  assign n1658 = ~n1458 & ~n1657;
  assign n1659 = n1511 & ~n1658;
  assign n1660 = ~n1401 & ~n1404;
  assign n1460 = n1455 ^ n1438;
  assign n1461 = ~n1452 & n1460;
  assign n1661 = n1511 ^ n1451;
  assign n1662 = n1461 & ~n1661;
  assign n1663 = n1662 ^ n1511;
  assign n1664 = ~n1660 & n1663;
  assign n1665 = n1458 & n1657;
  assign n1666 = ~n1664 & ~n1665;
  assign n1667 = ~n1659 & n1666;
  assign n1690 = n1689 ^ n1670;
  assign n1880 = ~n1667 & ~n1690;
  assign n1881 = ~n1786 & ~n1880;
  assign n1882 = ~n1834 & ~n1881;
  assign n1883 = n1667 & n1690;
  assign n1788 = n1655 & n1784;
  assign n1884 = n1834 ^ n1654;
  assign n1885 = n1788 & ~n1884;
  assign n1886 = n1885 ^ n1834;
  assign n1887 = ~n1883 & ~n1886;
  assign n1888 = n1786 & n1880;
  assign n1889 = ~n1887 & ~n1888;
  assign n1890 = ~n1882 & n1889;
  assign n1891 = n1832 ^ n1794;
  assign n1892 = n1833 & n1891;
  assign n1893 = n1892 ^ n1794;
  assign n1902 = n1821 ^ n1810;
  assign n1903 = n1817 & n1902;
  assign n1904 = n1903 ^ n1821;
  assign n1898 = n756 ^ n310;
  assign n1899 = ~n786 & ~n1898;
  assign n1900 = n1899 ^ n1212;
  assign n1894 = n1807 ^ n1802;
  assign n1895 = n1807 ^ n1801;
  assign n1896 = n1894 & ~n1895;
  assign n1897 = n1896 ^ n1802;
  assign n1901 = n1900 ^ n1897;
  assign n1905 = n1904 ^ n1901;
  assign n2069 = n1893 & n1905;
  assign n2070 = n1890 & ~n2069;
  assign n2071 = ~n1893 & ~n1905;
  assign n1915 = ~n748 & n1805;
  assign n1916 = n1079 ^ n699;
  assign n1917 = n753 & n1916;
  assign n1918 = ~n1915 & ~n1917;
  assign n1910 = n800 & n1697;
  assign n1911 = n1910 ^ n312;
  assign n1912 = ~n1068 & n1911;
  assign n1913 = ~n312 & ~n786;
  assign n1914 = ~n1912 & ~n1913;
  assign n1919 = n1918 ^ n1914;
  assign n1906 = ~n967 & ~n1819;
  assign n1908 = n858 & ~n1907;
  assign n1909 = ~n1906 & ~n1908;
  assign n1920 = n1919 ^ n1909;
  assign n1921 = n1808 ^ n1797;
  assign n1922 = ~n1823 & ~n1921;
  assign n1923 = n1922 ^ n1822;
  assign n1924 = n1920 & ~n1923;
  assign n1966 = n310 & ~n756;
  assign n1967 = n1212 & ~n1966;
  assign n1968 = ~n310 & n756;
  assign n1969 = ~n786 & ~n1968;
  assign n1970 = ~n1967 & n1969;
  assign n1960 = ~n308 & n1070;
  assign n1961 = ~n1069 & ~n1960;
  assign n1962 = n1068 ^ n800;
  assign n1963 = n315 & ~n1962;
  assign n1964 = n1963 ^ n800;
  assign n1965 = n1961 & n1964;
  assign n1971 = n1970 ^ n1965;
  assign n1957 = n1918 ^ n1909;
  assign n1958 = ~n1919 & n1957;
  assign n1959 = n1958 ^ n1909;
  assign n1972 = n1971 ^ n1959;
  assign n1956 = n1955 ^ n1949;
  assign n1973 = n1972 ^ n1956;
  assign n1943 = n1904 ^ n1897;
  assign n1944 = ~n1901 & n1943;
  assign n1945 = n1944 ^ n1904;
  assign n1974 = n1973 ^ n1945;
  assign n2072 = ~n1924 & ~n1974;
  assign n2073 = ~n2071 & ~n2072;
  assign n2074 = ~n2070 & n2073;
  assign n2075 = n1924 & n1974;
  assign n2076 = ~n2074 & ~n2075;
  assign n2077 = n1974 & ~n2071;
  assign n2078 = n1890 & ~n2077;
  assign n1934 = ~n1920 & n1923;
  assign n2079 = ~n1974 & ~n2069;
  assign n2080 = ~n1934 & ~n2079;
  assign n2081 = ~n2078 & n2080;
  assign n2082 = n2076 & ~n2081;
  assign n2060 = n1970 ^ n1959;
  assign n2061 = ~n1971 & ~n2060;
  assign n2062 = n2061 ^ n1959;
  assign n2059 = n2058 ^ n2049;
  assign n2063 = n2062 ^ n2059;
  assign n2045 = ~n786 & n1697;
  assign n2046 = n2045 ^ n1326;
  assign n2306 = n2062 ^ n2046;
  assign n2307 = n2063 & ~n2306;
  assign n2308 = n2307 ^ n2059;
  assign n2065 = n1972 ^ n1945;
  assign n2066 = ~n1973 & n2065;
  assign n2067 = n2066 ^ n1945;
  assign n2302 = n2059 & n2062;
  assign n2303 = n2046 & n2302;
  assign n2311 = ~n2067 & ~n2303;
  assign n2312 = n2308 & ~n2311;
  assign n2299 = ~n2059 & ~n2062;
  assign n2300 = ~n2046 & n2299;
  assign n2301 = ~n2067 & n2300;
  assign n2381 = ~n2301 & n2337;
  assign n2382 = ~n2312 & ~n2381;
  assign n2383 = ~n2082 & ~n2382;
  assign n2309 = n2067 & ~n2300;
  assign n2310 = ~n2308 & ~n2309;
  assign n2304 = n2067 & n2303;
  assign n2384 = ~n2304 & ~n2337;
  assign n2385 = ~n2310 & ~n2384;
  assign n2386 = ~n2383 & ~n2385;
  assign n2461 = n2424 ^ n2386;
  assign n2462 = ~n2425 & ~n2461;
  assign n2463 = n2462 ^ n2386;
  assign n2471 = n2470 ^ n2463;
  assign n1570 = ~n164 & ~n813;
  assign n1571 = ~n137 & ~n1570;
  assign n1572 = n111 & n130;
  assign n1573 = ~n1571 & ~n1572;
  assign n1574 = ~n1542 & n1573;
  assign n1575 = n504 & n1574;
  assign n1576 = n586 & n928;
  assign n1577 = ~n253 & ~n447;
  assign n1578 = n1576 & n1577;
  assign n1579 = n1575 & n1578;
  assign n1580 = ~n374 & ~n428;
  assign n1581 = n439 & n1580;
  assign n1582 = ~n399 & ~n672;
  assign n1583 = n1581 & n1582;
  assign n1584 = n1579 & n1583;
  assign n2448 = ~n343 & ~n366;
  assign n2449 = ~n273 & n2448;
  assign n2450 = ~n322 & ~n523;
  assign n2451 = ~n212 & n2450;
  assign n2452 = n2449 & n2451;
  assign n2453 = n209 & n2452;
  assign n2454 = n1584 & n2453;
  assign n1523 = ~n245 & ~n919;
  assign n2024 = n78 & n140;
  assign n2025 = n51 & ~n2024;
  assign n2026 = n1591 & ~n2025;
  assign n2027 = n1523 & n2026;
  assign n2028 = ~n539 & ~n688;
  assign n2029 = n880 & n2028;
  assign n2030 = n2027 & n2029;
  assign n2455 = n182 & ~n293;
  assign n2001 = n85 & ~n706;
  assign n2002 = ~n423 & ~n2001;
  assign n2456 = n729 & n2002;
  assign n2457 = n2455 & n2456;
  assign n2458 = n479 & n2457;
  assign n2459 = n2030 & n2458;
  assign n2460 = n2454 & n2459;
  assign n2472 = n2471 ^ n2460;
  assign n2426 = n2425 ^ n2386;
  assign n2305 = ~n2301 & ~n2304;
  assign n2313 = n2312 ^ n2310;
  assign n2314 = ~n2082 & n2313;
  assign n2315 = n2314 ^ n2310;
  assign n2316 = n2305 & ~n2315;
  assign n2338 = n2337 ^ n2316;
  assign n1998 = ~n85 & n211;
  assign n1999 = ~n78 & ~n1998;
  assign n2000 = n1581 & ~n1999;
  assign n2003 = n57 & ~n159;
  assign n2004 = n2002 & ~n2003;
  assign n2005 = n130 & ~n149;
  assign n2006 = n2004 & ~n2005;
  assign n2007 = n638 & n2006;
  assign n2008 = n2000 & n2007;
  assign n2009 = ~n262 & ~n366;
  assign n2010 = n260 & n2009;
  assign n2011 = n570 & n2010;
  assign n2012 = n2008 & n2011;
  assign n1589 = ~n424 & ~n485;
  assign n1590 = ~n358 & n1589;
  assign n1524 = ~n672 & ~n728;
  assign n2277 = n50 & n680;
  assign n2278 = n1524 & ~n2277;
  assign n2279 = ~n355 & ~n380;
  assign n2280 = n2278 & n2279;
  assign n2281 = n1590 & n2280;
  assign n2282 = n101 & ~n801;
  assign n2283 = n840 & ~n2282;
  assign n2284 = n2281 & n2283;
  assign n2285 = n658 & n2284;
  assign n2286 = ~n367 & n650;
  assign n2287 = ~n200 & ~n769;
  assign n2288 = n2286 & n2287;
  assign n2289 = n648 & n2288;
  assign n2290 = ~n188 & ~n410;
  assign n2291 = ~n242 & ~n341;
  assign n2292 = n2290 & n2291;
  assign n279 = ~n129 & ~n278;
  assign n2293 = n279 & n551;
  assign n2294 = n2292 & n2293;
  assign n2295 = ~n825 & n2294;
  assign n2296 = n2289 & n2295;
  assign n2297 = n2285 & n2296;
  assign n2298 = n2012 & n2297;
  assign n2339 = n2338 ^ n2298;
  assign n2064 = n2063 ^ n2046;
  assign n2068 = n2067 ^ n2064;
  assign n2083 = n2082 ^ n2068;
  assign n2013 = n101 & ~n171;
  assign n2014 = ~n181 & ~n2013;
  assign n2015 = n2012 & n2014;
  assign n292 = ~n286 & n291;
  assign n2016 = n56 & ~n116;
  assign n2017 = ~n687 & ~n2016;
  assign n2018 = n369 & n2017;
  assign n2019 = n292 & n2018;
  assign n395 = ~n242 & ~n394;
  assign n2020 = ~n57 & n395;
  assign n2021 = ~n779 & ~n2020;
  assign n2022 = ~n345 & ~n2021;
  assign n2023 = n2019 & n2022;
  assign n2031 = ~n40 & ~n344;
  assign n2032 = n681 & ~n2031;
  assign n2033 = ~n50 & ~n221;
  assign n2034 = ~n2032 & ~n2033;
  assign n2035 = ~n330 & ~n2034;
  assign n2036 = n165 & ~n949;
  assign n2037 = ~n689 & ~n2036;
  assign n2038 = ~n1572 & n2037;
  assign n2039 = n100 & ~n155;
  assign n2040 = n2038 & ~n2039;
  assign n2041 = n2035 & n2040;
  assign n2042 = n2030 & n2041;
  assign n2043 = n2023 & n2042;
  assign n2044 = n2015 & n2043;
  assign n2084 = n2083 ^ n2044;
  assign n1925 = n1905 & n1924;
  assign n1926 = ~n1893 & ~n1925;
  assign n1927 = n1923 ^ n1920;
  assign n1928 = n1923 ^ n1905;
  assign n1929 = n1927 & ~n1928;
  assign n1930 = n1929 ^ n1905;
  assign n1931 = ~n1926 & n1930;
  assign n1932 = ~n1890 & n1931;
  assign n1933 = n1905 ^ n1893;
  assign n1935 = ~n1905 & n1934;
  assign n1936 = ~n1925 & ~n1935;
  assign n1937 = ~n1933 & ~n1936;
  assign n1938 = ~n1932 & ~n1937;
  assign n1939 = ~n1893 & ~n1930;
  assign n1940 = ~n1935 & ~n1939;
  assign n1941 = n1890 & ~n1940;
  assign n1942 = n1938 & ~n1941;
  assign n1975 = n1974 ^ n1942;
  assign n231 = n226 & ~n230;
  assign n232 = n223 & n231;
  assign n246 = ~n244 & ~n245;
  assign n247 = ~n242 & n246;
  assign n248 = n241 & n247;
  assign n249 = n232 & n248;
  assign n250 = ~n215 & n249;
  assign n1625 = ~n152 & ~n397;
  assign n1856 = ~n170 & ~n1625;
  assign n1857 = ~n140 & n813;
  assign n1858 = ~n1856 & ~n1857;
  assign n1859 = ~n367 & n1858;
  assign n1860 = ~n274 & ~n519;
  assign n1861 = ~n577 & n1860;
  assign n1862 = n1859 & n1861;
  assign n1863 = ~n92 & ~n366;
  assign n1864 = ~n468 & n1863;
  assign n1865 = ~n111 & n236;
  assign n1866 = ~n165 & n1865;
  assign n1867 = ~n826 & ~n1866;
  assign n1868 = ~n418 & ~n998;
  assign n1869 = ~n424 & n1868;
  assign n1870 = ~n399 & n1869;
  assign n1871 = ~n1867 & n1870;
  assign n1872 = n1864 & n1871;
  assign n1873 = n1862 & n1872;
  assign n1874 = ~n79 & n1017;
  assign n1875 = ~n343 & ~n1874;
  assign n1876 = ~n372 & n1875;
  assign n1877 = n1873 & n1876;
  assign n1878 = n556 & n1877;
  assign n1879 = n250 & n1878;
  assign n1976 = n1975 ^ n1879;
  assign n1986 = n1933 ^ n1927;
  assign n1987 = n1986 ^ n1890;
  assign n429 = n51 & ~n255;
  assign n430 = ~n428 & ~n429;
  assign n431 = ~n91 & n100;
  assign n432 = n137 & ~n431;
  assign n433 = ~n211 & ~n432;
  assign n434 = n430 & ~n433;
  assign n435 = n427 & n434;
  assign n1977 = n435 & n1522;
  assign n1978 = n165 & ~n779;
  assign n1979 = ~n563 & ~n1978;
  assign n1980 = n360 & n1979;
  assign n1981 = n534 & n1980;
  assign n1982 = n587 & n1981;
  assign n1983 = n1977 & n1982;
  assign n1984 = n134 & n583;
  assign n1985 = n1983 & n1984;
  assign n1988 = n1987 ^ n1985;
  assign n1691 = n1690 ^ n1667;
  assign n1787 = n1786 ^ n1690;
  assign n1789 = n1788 ^ n1787;
  assign n1790 = ~n1691 & n1789;
  assign n1791 = n1790 ^ n1788;
  assign n1835 = n1834 ^ n1791;
  assign n400 = ~n396 & ~n399;
  assign n1623 = n400 & ~n672;
  assign n1762 = ~n183 & ~n264;
  assign n1763 = ~n92 & ~n286;
  assign n1764 = n1762 & n1763;
  assign n1768 = ~n600 & n1767;
  assign n1769 = n1764 & n1768;
  assign n1770 = n1623 & n1769;
  assign n1771 = n554 & n1770;
  assign n1772 = ~n272 & ~n497;
  assign n1773 = ~n258 & n1772;
  assign n1774 = ~n341 & ~n358;
  assign n1775 = n1773 & n1774;
  assign n1550 = ~n69 & n130;
  assign n1776 = ~n244 & ~n1550;
  assign n1777 = n1775 & n1776;
  assign n1778 = ~n359 & ~n645;
  assign n1779 = ~n197 & n1778;
  assign n1780 = n448 & n1779;
  assign n1781 = n1777 & n1780;
  assign n1782 = n1771 & n1781;
  assign n1783 = n1761 & n1782;
  assign n1836 = n1835 ^ n1783;
  assign n1656 = n1655 ^ n1639;
  assign n1692 = n1691 ^ n1656;
  assign n1585 = n165 & ~n617;
  assign n1586 = ~n288 & ~n1585;
  assign n1587 = ~n679 & n1586;
  assign n1588 = n1514 & n1587;
  assign n1592 = n551 & n1591;
  assign n1593 = n1590 & n1592;
  assign n1594 = n1588 & n1593;
  assign n1624 = n719 & n1623;
  assign n1626 = ~n361 & ~n1625;
  assign n1627 = ~n728 & ~n1626;
  assign n1628 = n1624 & n1627;
  assign n318 = ~n165 & n317;
  assign n319 = ~n83 & n137;
  assign n320 = ~n318 & ~n319;
  assign n321 = ~n316 & ~n320;
  assign n324 = n130 & ~n323;
  assign n326 = n57 & ~n325;
  assign n327 = ~n324 & ~n326;
  assign n328 = ~n322 & n327;
  assign n329 = n321 & n328;
  assign n1629 = n111 & n1017;
  assign n1630 = ~n418 & ~n1629;
  assign n1631 = ~n195 & n1630;
  assign n1632 = n586 & n1631;
  assign n1633 = n329 & n1632;
  assign n1634 = n1628 & n1633;
  assign n1635 = n1594 & n1634;
  assign n1636 = n517 & n1635;
  assign n1693 = n1692 ^ n1636;
  assign n1558 = n1455 ^ n1452;
  assign n1405 = n1404 ^ n1401;
  assign n1559 = n1558 ^ n1405;
  assign n1525 = n164 & ~n170;
  assign n1526 = n1524 & ~n1525;
  assign n1527 = n1523 & n1526;
  assign n1528 = ~n428 & ~n687;
  assign n1529 = n83 & ~n204;
  assign n1530 = ~n844 & ~n1529;
  assign n1531 = n1528 & n1530;
  assign n1532 = ~n56 & n146;
  assign n1533 = ~n40 & n116;
  assign n1534 = ~n50 & n1533;
  assign n1535 = ~n1532 & ~n1534;
  assign n1536 = n40 & n91;
  assign n1537 = n1535 & ~n1536;
  assign n1538 = n100 & ~n140;
  assign n1539 = ~n1537 & ~n1538;
  assign n1540 = n1531 & n1539;
  assign n1541 = n1527 & n1540;
  assign n1544 = ~n424 & ~n497;
  assign n1545 = ~n1032 & n1544;
  assign n1546 = n1543 & n1545;
  assign n1547 = ~n188 & ~n237;
  assign n1548 = n400 & n1547;
  assign n1549 = n1546 & n1548;
  assign n1551 = ~n367 & ~n1550;
  assign n1552 = n57 & ~n404;
  assign n1553 = n1551 & ~n1552;
  assign n1554 = n736 & n1553;
  assign n1555 = n1549 & n1554;
  assign n1556 = n1541 & n1555;
  assign n1557 = n1522 & n1556;
  assign n1560 = n1559 ^ n1557;
  assign n1561 = n1156 ^ n1133;
  assign n1563 = n1386 ^ n1384;
  assign n1564 = n1387 & n1563;
  assign n1562 = n1389 ^ n1133;
  assign n1565 = n1564 ^ n1562;
  assign n1566 = n1561 & ~n1565;
  assign n1567 = n1566 ^ n1564;
  assign n1568 = n1567 ^ n1132;
  assign n1569 = ~n58 & ~n926;
  assign n1595 = n100 & ~n146;
  assign n1596 = n56 & ~n201;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = ~n330 & n1597;
  assign n1599 = n481 & n1598;
  assign n1600 = n265 & n936;
  assign n1601 = n1599 & n1600;
  assign n1602 = n516 & n548;
  assign n1603 = n1601 & n1602;
  assign n1604 = n1594 & n1603;
  assign n1605 = n1584 & n1604;
  assign n1606 = ~n1569 & n1605;
  assign n1607 = n1568 & n1606;
  assign n1608 = n1607 ^ n1557;
  assign n1609 = ~n1560 & ~n1608;
  assign n1610 = n1609 ^ n1559;
  assign n1459 = n1458 ^ n1404;
  assign n1462 = n1461 ^ n1459;
  assign n1463 = ~n1405 & ~n1462;
  assign n1464 = n1463 ^ n1461;
  assign n1512 = n1511 ^ n1464;
  assign n1619 = n1610 ^ n1512;
  assign n333 = ~n330 & n332;
  assign n335 = ~n129 & ~n334;
  assign n337 = ~n237 & ~n336;
  assign n338 = n335 & n337;
  assign n339 = n333 & n338;
  assign n282 = ~n280 & ~n281;
  assign n348 = n282 & n347;
  assign n349 = n339 & n348;
  assign n350 = n329 & n349;
  assign n392 = n371 & n391;
  assign n393 = n350 & n392;
  assign n401 = n395 & n400;
  assign n406 = ~n238 & ~n286;
  assign n407 = ~n405 & n406;
  assign n408 = n403 & n407;
  assign n409 = n401 & n408;
  assign n412 = ~n410 & ~n411;
  assign n414 = ~n221 & ~n272;
  assign n415 = ~n413 & n414;
  assign n416 = n412 & n415;
  assign n417 = n409 & n416;
  assign n436 = n421 & n435;
  assign n437 = n417 & n436;
  assign n438 = n393 & n437;
  assign n1620 = n1610 ^ n438;
  assign n1621 = ~n1619 & n1620;
  assign n1622 = n1621 ^ n1512;
  assign n1749 = n1692 ^ n1622;
  assign n1750 = ~n1693 & n1749;
  assign n1751 = n1750 ^ n1622;
  assign n1989 = n1783 ^ n1751;
  assign n1990 = ~n1836 & ~n1989;
  assign n1991 = n1990 ^ n1835;
  assign n1992 = n1991 ^ n1987;
  assign n1993 = n1988 & n1992;
  assign n1994 = n1993 ^ n1991;
  assign n1995 = n1994 ^ n1975;
  assign n1996 = n1976 & n1995;
  assign n1997 = n1996 ^ n1994;
  assign n2274 = n2083 ^ n1997;
  assign n2275 = ~n2084 & ~n2274;
  assign n2276 = n2275 ^ n1997;
  assign n2378 = n2338 ^ n2276;
  assign n2379 = n2339 & n2378;
  assign n2380 = n2379 ^ n2276;
  assign n2427 = n2426 ^ n2380;
  assign n2362 = ~n286 & ~n293;
  assign n2363 = ~n595 & n2362;
  assign n2364 = ~n216 & n356;
  assign n2365 = n2363 & n2364;
  assign n2366 = n111 & ~n888;
  assign n2367 = ~n497 & ~n693;
  assign n2368 = ~n2366 & n2367;
  assign n2369 = n260 & n2368;
  assign n2370 = n2365 & n2369;
  assign n2371 = n383 & n726;
  assign n2372 = n514 & n2371;
  assign n2373 = n832 & n2372;
  assign n2374 = n2370 & n2373;
  assign n2375 = n939 & n2374;
  assign n2376 = n622 & ~n687;
  assign n2377 = n2375 & n2376;
  assign n2445 = n2426 ^ n2377;
  assign n2446 = ~n2427 & ~n2445;
  assign n2447 = n2446 ^ n2380;
  assign n2499 = n2471 ^ n2447;
  assign n2500 = ~n2472 & ~n2499;
  assign n2501 = n2500 ^ n2447;
  assign n2518 = n2517 ^ n2501;
  assign n2519 = n989 & n2230;
  assign n2520 = ~n1079 & ~n2519;
  assign n2521 = ~n786 & n2520;
  assign n2522 = ~n2464 & ~n2521;
  assign n2528 = n2469 & ~n2522;
  assign n2523 = ~n989 & ~n2230;
  assign n2524 = ~n786 & n2523;
  assign n2529 = n800 & ~n1079;
  assign n2530 = n2524 & n2529;
  assign n2531 = ~n2528 & ~n2530;
  assign n2532 = n2463 & ~n2531;
  assign n2824 = n2532 ^ n2517;
  assign n2825 = ~n2518 & ~n2824;
  assign n2826 = n2825 ^ n2501;
  assign n2928 = n2823 & ~n2826;
  assign n294 = n128 & ~n165;
  assign n295 = n78 & ~n130;
  assign n296 = ~n294 & ~n295;
  assign n297 = ~n293 & ~n296;
  assign n300 = ~n298 & ~n299;
  assign n301 = n297 & n300;
  assign n2903 = ~n380 & n1582;
  assign n2904 = n994 & n1528;
  assign n2905 = n2903 & n2904;
  assign n2906 = ~n288 & ~n539;
  assign n2907 = ~n769 & n2906;
  assign n2908 = n2905 & n2907;
  assign n2909 = n301 & n2908;
  assign n2910 = n460 & n2909;
  assign n2911 = ~n112 & ~n413;
  assign n2912 = ~n259 & n2911;
  assign n2913 = ~n195 & ~n239;
  assign n2914 = ~n242 & n1868;
  assign n2915 = n2913 & n2914;
  assign n2916 = n2912 & n2915;
  assign n2917 = n128 & n236;
  assign n2918 = ~n912 & ~n2917;
  assign n2919 = n2916 & ~n2918;
  assign n2920 = ~n569 & ~n646;
  assign n2921 = n57 & ~n323;
  assign n2922 = ~n92 & ~n2921;
  assign n2923 = n2920 & n2922;
  assign n2924 = n2456 & n2923;
  assign n2925 = n2919 & n2924;
  assign n2926 = n501 & n2925;
  assign n2927 = n2910 & n2926;
  assign n2929 = n2928 ^ n2927;
  assign n3051 = x1 & ~n2929;
  assign n2430 = ~x1 & x2;
  assign n2827 = n2826 ^ n2823;
  assign n3052 = n2430 & n2827;
  assign n3053 = ~x0 & ~n3052;
  assign n3054 = ~n3051 & n3053;
  assign n3028 = x2 ^ x1;
  assign n2473 = n2472 ^ n2447;
  assign n2486 = n2377 & n2427;
  assign n2487 = n2380 & ~n2426;
  assign n2488 = ~n2472 & ~n2487;
  assign n2489 = ~n2486 & ~n2488;
  assign n2340 = n2339 ^ n2276;
  assign n2085 = n2084 ^ n1997;
  assign n2086 = n1994 ^ n1976;
  assign n2087 = n1991 ^ n1988;
  assign n1513 = n1512 ^ n438;
  assign n1611 = n1610 ^ n1513;
  assign n1612 = n1607 ^ n1560;
  assign n1613 = n1611 & n1612;
  assign n1694 = n1693 ^ n1622;
  assign n1746 = ~n1613 & n1694;
  assign n1837 = n1836 ^ n1751;
  assign n2088 = ~n1746 & n1837;
  assign n2089 = n2087 & ~n2088;
  assign n2090 = ~n2086 & ~n2089;
  assign n2341 = ~n2085 & ~n2090;
  assign n2490 = ~n2340 & ~n2341;
  assign n2491 = ~n2489 & ~n2490;
  assign n2492 = n2473 & ~n2491;
  assign n2525 = n2522 & ~n2524;
  assign n2526 = n2525 ^ n2463;
  assign n2527 = n2470 & n2526;
  assign n2533 = n2532 ^ n2527;
  assign n2534 = n2518 & ~n2533;
  assign n2535 = n2534 ^ n2532;
  assign n3001 = ~n2492 & ~n2535;
  assign n3002 = ~n2823 & n2826;
  assign n3003 = ~n3001 & n3002;
  assign n3004 = n2927 & ~n3003;
  assign n2896 = ~n2501 & n2517;
  assign n2897 = n2527 & n2896;
  assign n2428 = n2427 ^ n2377;
  assign n1614 = n1606 ^ n1568;
  assign n1615 = n1612 & ~n1614;
  assign n1616 = ~n1611 & ~n1615;
  assign n1747 = ~n1616 & ~n1694;
  assign n2091 = ~n1747 & ~n1837;
  assign n2092 = ~n2087 & ~n2091;
  assign n2093 = n2086 & ~n2092;
  assign n2342 = n2085 & ~n2093;
  assign n2493 = n2340 & ~n2342;
  assign n2494 = n2428 & ~n2493;
  assign n2495 = ~n2473 & ~n2494;
  assign n3010 = n2495 & ~n2826;
  assign n3011 = ~n2897 & ~n3010;
  assign n3012 = ~n2823 & ~n3011;
  assign n3013 = n2823 & n2826;
  assign n2898 = n2501 & ~n2517;
  assign n2899 = ~n2527 & n2898;
  assign n3014 = ~n2495 & n2899;
  assign n3015 = n3013 & ~n3014;
  assign n3016 = ~n3012 & ~n3015;
  assign n3017 = ~n2927 & ~n2928;
  assign n3055 = ~n3001 & ~n3017;
  assign n3056 = n3016 & ~n3055;
  assign n3057 = ~n3004 & ~n3056;
  assign n3058 = n3028 & n3057;
  assign n2985 = n2927 & n2928;
  assign n2967 = ~n158 & n164;
  assign n2968 = ~n569 & ~n2967;
  assign n2969 = n432 & n2968;
  assign n2970 = ~n778 & n2969;
  assign n2971 = n486 & n557;
  assign n2972 = n2970 & n2971;
  assign n2973 = ~n353 & n720;
  assign n2974 = ~n385 & ~n1572;
  assign n2975 = n414 & n2974;
  assign n2976 = n2973 & n2975;
  assign n2977 = n2972 & n2976;
  assign n2978 = n2294 & n2977;
  assign n2979 = n430 & n1028;
  assign n2980 = ~n199 & ~n545;
  assign n2981 = n2979 & n2980;
  assign n2982 = n765 & n2981;
  assign n2983 = n806 & n2982;
  assign n2984 = n2978 & n2983;
  assign n3034 = n2985 ^ n2984;
  assign n3059 = n3058 ^ n3034;
  assign n3060 = x0 & n3059;
  assign n3061 = ~n3054 & ~n3060;
  assign n2431 = x22 ^ x2;
  assign n2432 = ~n2430 & n2431;
  assign n2433 = ~n26 & ~n2432;
  assign n2434 = x0 & ~x22;
  assign n2435 = x2 & n2434;
  assign n2436 = n2433 & ~n2435;
  assign n3062 = n3061 ^ n2436;
  assign n2484 = n2436 ^ n860;
  assign n2541 = n2493 ^ n2490;
  assign n2542 = ~n2428 & n2541;
  assign n2543 = n2542 ^ n2493;
  assign n2544 = ~n2473 & ~n2543;
  assign n2545 = n2484 & ~n2544;
  assign n2546 = n969 & ~n2545;
  assign n2437 = ~n860 & ~n2436;
  assign n2547 = n1057 & n2428;
  assign n2548 = n969 & ~n1057;
  assign n2549 = ~n2340 & n2548;
  assign n2550 = ~n2547 & ~n2549;
  assign n2551 = n2437 & ~n2550;
  assign n2440 = n860 & n2436;
  assign n2474 = ~n1057 & n2440;
  assign n2552 = n2428 & n2474;
  assign n2441 = ~n969 & n1057;
  assign n2442 = n2440 & n2441;
  assign n2553 = ~n2340 & n2442;
  assign n2554 = ~n2552 & ~n2553;
  assign n2555 = ~n2551 & n2554;
  assign n2556 = n2546 & n2555;
  assign n2557 = ~n969 & ~n2555;
  assign n2558 = ~n969 & n2484;
  assign n2559 = n2473 & ~n2543;
  assign n2560 = n2558 & n2559;
  assign n2561 = n2473 ^ n1057;
  assign n2562 = n2484 & n2543;
  assign n2563 = n2561 & n2562;
  assign n2564 = ~n2560 & ~n2563;
  assign n2565 = ~n2557 & n2564;
  assign n2566 = ~n2556 & n2565;
  assign n1855 = n969 ^ n750;
  assign n2124 = ~n2089 & ~n2092;
  assign n2125 = ~n2086 & ~n2124;
  assign n2126 = n1855 & n2125;
  assign n2098 = n750 & n969;
  assign n2097 = ~n750 & ~n969;
  assign n2099 = n2098 ^ n2097;
  assign n2100 = n756 & n2099;
  assign n2101 = n2100 ^ n2097;
  assign n2127 = ~n2087 & n2101;
  assign n2103 = n2100 ^ n2098;
  assign n2104 = ~n1898 & n2103;
  assign n2128 = n1837 & n2104;
  assign n2129 = ~n2127 & ~n2128;
  assign n2130 = ~n2126 & n2129;
  assign n2131 = ~n310 & ~n2130;
  assign n2132 = n2086 & ~n2124;
  assign n2133 = n1855 & ~n2132;
  assign n2134 = n310 & n2129;
  assign n2135 = ~n2133 & n2134;
  assign n2136 = n1855 & n2124;
  assign n2137 = n2086 ^ n756;
  assign n2138 = n2136 & n2137;
  assign n2139 = ~n2135 & ~n2138;
  assign n2140 = ~n2131 & n2139;
  assign n313 = n312 ^ n310;
  assign n1700 = n315 ^ n308;
  assign n1714 = n1560 & n1614;
  assign n1715 = n1700 & n1714;
  assign n1716 = n1715 ^ n1611;
  assign n1717 = n313 & n1716;
  assign n1698 = ~n313 & n1697;
  assign n1718 = n1612 & n1698;
  assign n1701 = n312 ^ n308;
  assign n1702 = n1700 & n1701;
  assign n1703 = ~n313 & n1702;
  assign n1719 = ~n1614 & n1703;
  assign n1720 = ~n1718 & ~n1719;
  assign n1721 = ~n1717 & n1720;
  assign n1722 = ~n1560 & n1614;
  assign n1723 = n310 & n312;
  assign n1724 = ~n1614 & n1723;
  assign n1725 = ~n315 & n1724;
  assign n1726 = n1725 ^ n1723;
  assign n1727 = ~n1722 & ~n1726;
  assign n1728 = ~n310 & ~n312;
  assign n1729 = n315 & ~n1614;
  assign n1730 = n1728 & ~n1729;
  assign n1731 = n1727 & ~n1730;
  assign n1732 = n308 & ~n1731;
  assign n1733 = n1721 & n1732;
  assign n1735 = ~n1614 & n1734;
  assign n1617 = ~n1613 & ~n1616;
  assign n1618 = n315 & n1617;
  assign n1695 = n1694 ^ n1618;
  assign n1696 = n313 & ~n1695;
  assign n1699 = n1611 & n1698;
  assign n1704 = n1612 & n1703;
  assign n1705 = ~n1699 & ~n1704;
  assign n1706 = ~n1696 & n1705;
  assign n1707 = ~n308 & ~n1706;
  assign n1708 = ~n315 & n1617;
  assign n1709 = n1708 ^ n1694;
  assign n1710 = n313 & ~n1709;
  assign n1711 = n308 & n1705;
  assign n1712 = ~n1710 & n1711;
  assign n1713 = ~n1707 & ~n1712;
  assign n2120 = n1735 ^ n1713;
  assign n2119 = n1712 & ~n1735;
  assign n2121 = n2120 ^ n2119;
  assign n2122 = n1733 & n2121;
  assign n2123 = n2122 ^ n2120;
  assign n2141 = n2140 ^ n2123;
  assign n2198 = n308 & n1731;
  assign n2199 = n2198 ^ n1721;
  assign n2145 = ~n310 & ~n1617;
  assign n2146 = n1855 & ~n2145;
  assign n2147 = n756 & n1617;
  assign n2148 = n2147 ^ n1694;
  assign n2149 = n2146 & ~n2148;
  assign n2150 = ~n1617 & n1694;
  assign n2151 = n1855 & ~n2150;
  assign n2152 = n1611 & n2101;
  assign n2153 = n1612 & n2104;
  assign n2154 = ~n2152 & ~n2153;
  assign n2155 = ~n310 & n2154;
  assign n2156 = ~n2151 & n2155;
  assign n2157 = ~n2149 & ~n2156;
  assign n2158 = n310 & ~n2154;
  assign n2159 = n2157 & ~n2158;
  assign n2160 = n1714 & ~n1898;
  assign n2161 = n2160 ^ n1611;
  assign n2162 = n1855 & n2161;
  assign n2163 = n1612 & n2101;
  assign n2164 = ~n1614 & n2104;
  assign n2165 = ~n2163 & ~n2164;
  assign n2166 = ~n2162 & n2165;
  assign n2167 = n1612 & n1855;
  assign n2168 = n1614 & ~n2167;
  assign n2169 = ~n2103 & ~n2168;
  assign n2170 = n310 & ~n2169;
  assign n2171 = n2166 & n2170;
  assign n2172 = n313 & ~n1614;
  assign n2173 = ~n2171 & ~n2172;
  assign n2174 = n2159 & ~n2173;
  assign n2142 = n313 & n1612;
  assign n2143 = ~n1724 & ~n2142;
  assign n2144 = n2143 ^ n1729;
  assign n2175 = n2174 ^ n2144;
  assign n1748 = ~n1746 & ~n1747;
  assign n2176 = n1837 ^ n1748;
  assign n2177 = ~n756 & n1855;
  assign n2178 = n2176 & n2177;
  assign n2179 = ~n1694 & n2101;
  assign n2180 = n1611 & n2104;
  assign n2181 = ~n2179 & ~n2180;
  assign n2182 = ~n1966 & n2181;
  assign n2183 = n756 & n1855;
  assign n2184 = n1837 & n2183;
  assign n2185 = n2182 & ~n2184;
  assign n2186 = ~n2178 & n2185;
  assign n2187 = ~n1837 & n2181;
  assign n2188 = n310 & ~n2187;
  assign n2189 = ~n2186 & ~n2188;
  assign n2190 = n1855 & n2176;
  assign n2191 = n310 & ~n2177;
  assign n2192 = n2181 & n2191;
  assign n2193 = ~n2190 & n2192;
  assign n2194 = ~n2189 & ~n2193;
  assign n2195 = n2194 ^ n2144;
  assign n2196 = ~n2175 & ~n2195;
  assign n2197 = n2196 ^ n2174;
  assign n2200 = n2199 ^ n2197;
  assign n2201 = ~n2088 & ~n2091;
  assign n2202 = ~n2087 & ~n2201;
  assign n2203 = n1855 & n2202;
  assign n2204 = n1837 & n2101;
  assign n2205 = ~n1694 & n2104;
  assign n2206 = ~n2204 & ~n2205;
  assign n2207 = ~n2203 & n2206;
  assign n2208 = n310 & ~n2207;
  assign n2209 = n2087 & ~n2201;
  assign n2210 = n1855 & ~n2209;
  assign n2211 = ~n310 & n2206;
  assign n2212 = ~n2210 & n2211;
  assign n2213 = n1855 & n2201;
  assign n2214 = n2087 ^ n756;
  assign n2215 = n2213 & ~n2214;
  assign n2216 = ~n2212 & ~n2215;
  assign n2217 = ~n2208 & n2216;
  assign n2218 = n2217 ^ n2199;
  assign n2219 = n2200 & ~n2218;
  assign n2220 = n2219 ^ n2217;
  assign n2221 = n2220 ^ n2140;
  assign n2222 = ~n2141 & ~n2221;
  assign n2223 = n2222 ^ n2220;
  assign n2094 = ~n2090 & ~n2093;
  assign n2095 = n2085 & ~n2094;
  assign n2096 = n1855 & n2095;
  assign n2102 = ~n2086 & n2101;
  assign n2105 = ~n2087 & n2104;
  assign n2106 = ~n2102 & ~n2105;
  assign n2107 = ~n2096 & n2106;
  assign n2108 = ~n310 & ~n2107;
  assign n2109 = ~n2085 & ~n2094;
  assign n2110 = n1855 & ~n2109;
  assign n2111 = n310 & n2106;
  assign n2112 = ~n2110 & n2111;
  assign n2113 = n1855 & n2094;
  assign n2114 = n2085 ^ n756;
  assign n2115 = n2113 & ~n2114;
  assign n2116 = ~n2112 & ~n2115;
  assign n2117 = ~n2108 & n2116;
  assign n1838 = n313 & n1837;
  assign n1839 = ~n1748 & n1838;
  assign n1840 = ~n1694 & n1698;
  assign n1841 = n1611 & n1703;
  assign n1842 = ~n1840 & ~n1841;
  assign n1843 = ~n1839 & n1842;
  assign n1844 = ~n308 & ~n1843;
  assign n1845 = n313 & n1748;
  assign n1846 = n308 & n1842;
  assign n1847 = ~n1845 & n1846;
  assign n1848 = ~n1838 & n1847;
  assign n1849 = n1837 ^ n315;
  assign n1850 = n1845 & n1849;
  assign n1851 = ~n1848 & ~n1850;
  assign n1852 = ~n1844 & n1851;
  assign n1738 = n1612 & n1734;
  assign n1742 = ~n989 & ~n1614;
  assign n1739 = n308 & n864;
  assign n1740 = n1739 ^ n989;
  assign n1741 = ~n1614 & ~n1740;
  assign n1743 = n1742 ^ n1741;
  assign n1744 = ~n1738 & ~n1743;
  assign n1745 = n1744 ^ n1742;
  assign n1853 = n1852 ^ n1745;
  assign n1736 = ~n1733 & ~n1735;
  assign n1737 = ~n1713 & ~n1736;
  assign n1854 = n1853 ^ n1737;
  assign n2118 = n2117 ^ n1854;
  assign n2540 = n2223 ^ n2118;
  assign n2567 = n2566 ^ n2540;
  assign n2569 = ~n2490 & ~n2493;
  assign n2570 = n2428 & ~n2569;
  assign n2571 = n969 & n2484;
  assign n2572 = n2570 & n2571;
  assign n2475 = n1057 & n2437;
  assign n2476 = ~n2474 & ~n2475;
  assign n2573 = ~n2340 & ~n2476;
  assign n2485 = n1057 ^ n969;
  assign n2574 = n1057 & ~n2440;
  assign n2575 = ~n1057 & ~n2437;
  assign n2576 = ~n2574 & ~n2575;
  assign n2577 = n2485 & n2576;
  assign n2578 = n2085 & n2577;
  assign n2579 = ~n2573 & ~n2578;
  assign n2580 = n969 & ~n2579;
  assign n2581 = ~n2572 & ~n2580;
  assign n2582 = n2428 ^ n1057;
  assign n2583 = n2484 & n2569;
  assign n2584 = ~n2582 & n2583;
  assign n2585 = n2581 & ~n2584;
  assign n2586 = ~n2428 & ~n2569;
  assign n2587 = n2484 & ~n2586;
  assign n2588 = ~n969 & n2579;
  assign n2589 = ~n2587 & n2588;
  assign n2590 = n2585 & ~n2589;
  assign n2568 = n2220 ^ n2141;
  assign n2591 = n2590 ^ n2568;
  assign n2343 = ~n2341 & ~n2342;
  assign n2351 = n2340 & ~n2343;
  assign n2593 = ~n2351 & n2484;
  assign n2594 = n2085 & ~n2476;
  assign n2595 = ~n2086 & n2577;
  assign n2596 = ~n2594 & ~n2595;
  assign n2597 = n969 & n2596;
  assign n2598 = ~n2593 & n2597;
  assign n2599 = n2343 & n2484;
  assign n2600 = n2340 ^ n1057;
  assign n2601 = n2599 & ~n2600;
  assign n2602 = ~n2598 & ~n2601;
  assign n2344 = ~n2340 & ~n2343;
  assign n2603 = n2344 & n2558;
  assign n2604 = ~n969 & ~n2596;
  assign n2605 = ~n2603 & ~n2604;
  assign n2606 = n2602 & n2605;
  assign n2592 = n2217 ^ n2200;
  assign n2607 = n2606 ^ n2592;
  assign n2609 = n2095 & n2571;
  assign n2610 = ~n2086 & ~n2476;
  assign n2611 = ~n2087 & n2577;
  assign n2612 = ~n2610 & ~n2611;
  assign n2613 = n969 & ~n2612;
  assign n2614 = ~n2609 & ~n2613;
  assign n2615 = ~n2109 & n2484;
  assign n2616 = ~n969 & n2612;
  assign n2617 = ~n2615 & n2616;
  assign n2618 = n2614 & ~n2617;
  assign n2619 = n2094 & n2484;
  assign n2620 = n2085 ^ n1057;
  assign n2621 = n2619 & ~n2620;
  assign n2622 = n2618 & ~n2621;
  assign n2608 = n2194 ^ n2175;
  assign n2623 = n2622 ^ n2608;
  assign n2627 = ~n2087 & ~n2476;
  assign n2628 = n1837 & n2577;
  assign n2629 = ~n2627 & ~n2628;
  assign n2630 = n969 & n2629;
  assign n2631 = n2124 & n2630;
  assign n2632 = ~n2558 & ~n2631;
  assign n2633 = n1057 & n2124;
  assign n2634 = ~n2086 & ~n2633;
  assign n2635 = ~n2632 & n2634;
  assign n2636 = ~n2132 & n2484;
  assign n2637 = n2630 & ~n2636;
  assign n2638 = n2086 & n2124;
  assign n2639 = n1057 & n2484;
  assign n2640 = n2638 & n2639;
  assign n2641 = ~n969 & ~n2629;
  assign n2642 = ~n2640 & ~n2641;
  assign n2643 = ~n2637 & n2642;
  assign n2644 = ~n2635 & n2643;
  assign n2624 = n2173 ^ n2159;
  assign n2625 = n2171 & n2172;
  assign n2626 = n2624 & ~n2625;
  assign n2645 = n2644 ^ n2626;
  assign n2648 = n2202 & n2558;
  assign n2649 = n1837 & ~n2476;
  assign n2650 = ~n1694 & n2577;
  assign n2651 = ~n2649 & ~n2650;
  assign n2652 = ~n969 & ~n2651;
  assign n2653 = ~n2648 & ~n2652;
  assign n2654 = n2087 ^ n1057;
  assign n2655 = n2201 & n2484;
  assign n2656 = ~n2654 & n2655;
  assign n2657 = n2653 & ~n2656;
  assign n2658 = ~n2209 & n2484;
  assign n2659 = n969 & n2651;
  assign n2660 = ~n2658 & n2659;
  assign n2661 = n2657 & ~n2660;
  assign n2646 = n310 & n2169;
  assign n2647 = n2646 ^ n2166;
  assign n2662 = n2661 ^ n2647;
  assign n2667 = n1617 & n2485;
  assign n2668 = n2667 ^ n1694;
  assign n2669 = n2484 & ~n2668;
  assign n2670 = n1611 & ~n2476;
  assign n2671 = n1612 & n2577;
  assign n2672 = ~n2670 & ~n2671;
  assign n2673 = ~n2669 & n2672;
  assign n2674 = n1714 & n2485;
  assign n2675 = n2674 ^ n1611;
  assign n2676 = n2484 & ~n2675;
  assign n2677 = n1057 ^ n860;
  assign n2678 = n1612 & n2677;
  assign n2679 = n969 ^ n860;
  assign n2680 = ~n2677 & n2679;
  assign n2681 = ~n1614 & n2680;
  assign n2682 = ~n2484 & ~n2681;
  assign n2683 = ~n2678 & n2682;
  assign n2684 = ~n2676 & ~n2683;
  assign n2685 = ~n1722 & ~n2576;
  assign n2686 = n969 & ~n2685;
  assign n2687 = ~n2684 & n2686;
  assign n2688 = n2673 & ~n2687;
  assign n2689 = ~n750 & n969;
  assign n2690 = ~n1614 & n2689;
  assign n2691 = n2688 & ~n2690;
  assign n2692 = n750 & ~n969;
  assign n2693 = ~n1614 & n2692;
  assign n2694 = ~n2673 & ~n2693;
  assign n2695 = ~n2691 & ~n2694;
  assign n2664 = ~n1614 & n2098;
  assign n2665 = ~n2167 & ~n2664;
  assign n2663 = ~n756 & ~n1614;
  assign n2666 = n2665 ^ n2663;
  assign n2696 = n2695 ^ n2666;
  assign n2701 = n1748 & n2485;
  assign n2702 = n2701 ^ n969;
  assign n2703 = n2702 ^ n1837;
  assign n2697 = ~n1694 & n2677;
  assign n2698 = n1611 & n2680;
  assign n2699 = ~n2697 & ~n2698;
  assign n2700 = n2699 ^ n969;
  assign n2704 = n2703 ^ n2700;
  assign n2705 = ~n2484 & ~n2704;
  assign n2706 = n2705 ^ n2703;
  assign n2707 = n2706 ^ n2666;
  assign n2708 = ~n2696 & n2707;
  assign n2709 = n2708 ^ n2695;
  assign n2710 = n2709 ^ n2647;
  assign n2711 = n2662 & n2710;
  assign n2712 = n2711 ^ n2661;
  assign n2713 = n2712 ^ n2626;
  assign n2714 = n2645 & ~n2713;
  assign n2715 = n2714 ^ n2644;
  assign n2716 = n2715 ^ n2608;
  assign n2717 = n2623 & n2716;
  assign n2718 = n2717 ^ n2622;
  assign n2719 = n2718 ^ n2592;
  assign n2720 = n2607 & n2719;
  assign n2721 = n2720 ^ n2606;
  assign n2722 = n2721 ^ n2568;
  assign n2723 = n2591 & n2722;
  assign n2724 = n2723 ^ n2590;
  assign n2725 = n2724 ^ n2566;
  assign n2726 = ~n2567 & ~n2725;
  assign n2727 = n2726 ^ n2724;
  assign n2429 = n969 & ~n2428;
  assign n2438 = ~n1057 & n2437;
  assign n2439 = ~n2429 & n2438;
  assign n2443 = ~n2428 & n2442;
  assign n2444 = ~n2439 & ~n2443;
  assign n2478 = ~n2437 & ~n2474;
  assign n2479 = ~n969 & ~n2478;
  assign n2477 = n969 & ~n2476;
  assign n2480 = n2479 ^ n2477;
  assign n2481 = n2473 & n2480;
  assign n2482 = n2481 ^ n2479;
  assign n2483 = n2444 & ~n2482;
  assign n2496 = ~n2492 & ~n2495;
  assign n2497 = n2485 & n2496;
  assign n2498 = n2497 ^ n969;
  assign n2536 = n2535 ^ n2498;
  assign n2537 = n2484 & ~n2536;
  assign n2538 = n2483 & ~n2537;
  assign n2345 = n1855 & n2344;
  assign n2346 = n2085 & n2101;
  assign n2347 = ~n2086 & n2104;
  assign n2348 = ~n2346 & ~n2347;
  assign n2349 = ~n2345 & n2348;
  assign n2350 = n310 & ~n2349;
  assign n2352 = n1855 & ~n2351;
  assign n2353 = ~n310 & n2348;
  assign n2354 = ~n2352 & n2353;
  assign n2355 = n1855 & n2343;
  assign n2356 = n2340 ^ n756;
  assign n2357 = n2355 & ~n2356;
  assign n2358 = ~n2354 & ~n2357;
  assign n2359 = ~n2350 & n2358;
  assign n2253 = n1698 & n1837;
  assign n2254 = ~n1694 & n1703;
  assign n2255 = ~n2253 & ~n2254;
  assign n2256 = ~n308 & n2255;
  assign n2257 = n2201 & n2256;
  assign n2258 = n308 & n313;
  assign n2259 = ~n2257 & ~n2258;
  assign n2260 = ~n315 & n2201;
  assign n2261 = ~n2087 & ~n2260;
  assign n2262 = ~n2259 & n2261;
  assign n2263 = n313 & ~n2209;
  assign n2264 = n2256 & ~n2263;
  assign n2265 = n313 & ~n315;
  assign n2266 = n2087 & n2265;
  assign n2267 = n2201 & n2266;
  assign n2268 = n308 & ~n2255;
  assign n2269 = ~n2267 & ~n2268;
  assign n2270 = ~n2264 & n2269;
  assign n2271 = ~n2262 & n2270;
  assign n2240 = n1714 & n2239;
  assign n2241 = n2240 ^ n1611;
  assign n2242 = n1734 & n2241;
  assign n2234 = n989 & n1739;
  assign n2243 = ~n989 & n2230;
  assign n2244 = ~n2234 & ~n2243;
  assign n2245 = n1612 & ~n2244;
  assign n2231 = ~n1079 & n2230;
  assign n2246 = n1079 & n1739;
  assign n2247 = ~n2231 & ~n2246;
  assign n2248 = n2239 & ~n2247;
  assign n2249 = ~n1614 & n2248;
  assign n2250 = ~n2245 & ~n2249;
  assign n2251 = ~n2242 & n2250;
  assign n2232 = ~n1742 & n2231;
  assign n2233 = ~n1722 & ~n2232;
  assign n2235 = ~n1614 & n2234;
  assign n2236 = n2235 ^ n1739;
  assign n2237 = n2233 & ~n2236;
  assign n2238 = ~n1079 & n2237;
  assign n2252 = n2251 ^ n2238;
  assign n2272 = n2271 ^ n2252;
  assign n2227 = n1745 ^ n1737;
  assign n2228 = n1853 & n2227;
  assign n2229 = n2228 ^ n1852;
  assign n2273 = n2272 ^ n2229;
  assign n2360 = n2359 ^ n2273;
  assign n2224 = n2223 ^ n2117;
  assign n2225 = n2118 & ~n2224;
  assign n2226 = n2225 ^ n2223;
  assign n2361 = n2360 ^ n2226;
  assign n2539 = n2538 ^ n2361;
  assign n3063 = n2727 ^ n2539;
  assign n3064 = n3062 & n3063;
  assign n2804 = n2535 ^ n2473;
  assign n2805 = ~n2496 & n2804;
  assign n2900 = ~n2897 & ~n2899;
  assign n2901 = n2900 ^ n2823;
  assign n2902 = ~n2805 & n2901;
  assign n2930 = n2929 ^ n2902;
  assign n3039 = x22 ^ x1;
  assign n3040 = x0 & n3039;
  assign n3242 = ~n2930 & n3040;
  assign n3025 = x1 & ~x2;
  assign n3031 = ~x0 & x1;
  assign n3243 = ~n3025 & ~n3031;
  assign n3244 = ~n2827 & ~n3243;
  assign n3245 = n2430 & ~n2535;
  assign n3246 = ~x0 & ~n3245;
  assign n3247 = ~n3244 & n3246;
  assign n3248 = ~n3028 & ~n3031;
  assign n3249 = ~n2929 & n3248;
  assign n3250 = ~n3247 & ~n3249;
  assign n3251 = n2433 & n3250;
  assign n3252 = ~n3242 & n3251;
  assign n3253 = n2435 & n2930;
  assign n3254 = n3252 & ~n3253;
  assign n3026 = x0 & x22;
  assign n3027 = n3025 & n3026;
  assign n3255 = ~n2930 & n3027;
  assign n3168 = ~n25 & n2432;
  assign n3256 = n3168 & ~n3250;
  assign n3257 = ~n3255 & ~n3256;
  assign n3258 = ~n3254 & n3257;
  assign n3066 = n2535 ^ n2431;
  assign n3067 = x1 & ~n3066;
  assign n3068 = n2430 & ~n2473;
  assign n3069 = ~x0 & ~n3068;
  assign n3070 = ~n3067 & n3069;
  assign n3072 = n2805 & n3028;
  assign n3071 = n2827 ^ n2436;
  assign n3073 = n3072 ^ n3071;
  assign n3074 = x0 & ~n3073;
  assign n3075 = ~n3070 & ~n3074;
  assign n3065 = n2721 ^ n2591;
  assign n3076 = n3075 ^ n3065;
  assign n3078 = x1 & n2473;
  assign n3079 = n2428 & n2430;
  assign n3080 = ~x0 & ~n3079;
  assign n3081 = ~n3078 & n3080;
  assign n3082 = n2496 & n3028;
  assign n3083 = n3082 ^ n2535;
  assign n3084 = x0 & ~n3083;
  assign n3085 = ~n3081 & ~n3084;
  assign n3086 = n3085 ^ n2436;
  assign n3077 = n2718 ^ n2607;
  assign n3087 = n3086 ^ n3077;
  assign n3089 = n2543 & n3028;
  assign n3090 = n3089 ^ n2473;
  assign n3091 = x0 & n3090;
  assign n3092 = n2428 & n3031;
  assign n3035 = ~x0 & n2430;
  assign n3093 = ~n2340 & n3035;
  assign n3094 = ~n3092 & ~n3093;
  assign n3095 = ~n3091 & n3094;
  assign n3096 = n3095 ^ n2436;
  assign n3088 = n2715 ^ n2623;
  assign n3097 = n3096 ^ n3088;
  assign n3098 = n2709 ^ n2662;
  assign n3100 = n2094 & n3028;
  assign n3101 = n3100 ^ n2085;
  assign n3102 = x0 & n3101;
  assign n3103 = ~n2086 & n3031;
  assign n3104 = ~n2087 & n3035;
  assign n3105 = ~n3103 & ~n3104;
  assign n3106 = ~n3102 & n3105;
  assign n3107 = n3106 ^ n2436;
  assign n3099 = n2706 ^ n2696;
  assign n3108 = n3107 ^ n3099;
  assign n3029 = x0 & ~n3028;
  assign n3115 = ~n2086 & n3029;
  assign n3116 = ~n2087 & n3031;
  assign n3117 = n1837 & n3035;
  assign n3118 = ~n3116 & ~n3117;
  assign n3119 = ~n3115 & n3118;
  assign n3120 = n2436 & n3119;
  assign n3121 = n2124 ^ n2086;
  assign n3122 = n3040 & ~n3121;
  assign n3123 = n3120 & ~n3122;
  assign n3124 = n2432 & ~n3119;
  assign n3125 = n2430 & n2434;
  assign n3126 = ~n3027 & ~n3125;
  assign n3127 = ~n3121 & ~n3126;
  assign n3128 = ~n3124 & ~n3127;
  assign n3129 = ~n3123 & n3128;
  assign n3111 = n2688 ^ n750;
  assign n3109 = n969 & ~n2687;
  assign n3110 = n3109 ^ n2673;
  assign n3112 = n3111 ^ n3110;
  assign n3113 = n1614 & n3112;
  assign n3114 = n3113 ^ n3111;
  assign n3130 = n3129 ^ n3114;
  assign n3151 = n1612 & n2484;
  assign n3176 = n1614 & ~n3151;
  assign n3177 = n969 & ~n2576;
  assign n3178 = ~n3176 & n3177;
  assign n3179 = n3178 ^ n2684;
  assign n3147 = n1612 & ~n2437;
  assign n3148 = n2574 & ~n3147;
  assign n3149 = ~n2474 & ~n3148;
  assign n3150 = ~n1614 & ~n3149;
  assign n3152 = n1057 & ~n1614;
  assign n3153 = n3151 & ~n3152;
  assign n3154 = ~n3150 & ~n3153;
  assign n3131 = n1617 & n3028;
  assign n3132 = n3131 ^ n1694;
  assign n3133 = x0 & ~n3132;
  assign n3134 = n1611 & n3031;
  assign n3135 = n1612 & n3035;
  assign n3136 = ~n3134 & ~n3135;
  assign n3137 = ~n3133 & n3136;
  assign n3140 = ~n1611 & n1722;
  assign n3141 = ~n860 & ~n1614;
  assign n3142 = ~n3140 & ~n3141;
  assign n3143 = n2436 & ~n3142;
  assign n3138 = n860 & ~n2436;
  assign n3139 = ~n1614 & n3138;
  assign n3144 = n3143 ^ n3139;
  assign n3145 = ~n3137 & n3144;
  assign n3146 = n3145 ^ n3143;
  assign n3155 = n3154 ^ n3146;
  assign n3156 = x0 & ~n1837;
  assign n3157 = n1694 & n3031;
  assign n3158 = ~n1611 & n2430;
  assign n3159 = x0 & n3028;
  assign n3160 = ~n3158 & ~n3159;
  assign n3161 = ~n3157 & n3160;
  assign n3162 = ~n3156 & n3161;
  assign n3163 = n2433 & ~n3162;
  assign n3164 = n3040 ^ n2435;
  assign n3165 = n2176 & n3164;
  assign n3166 = n3165 ^ n2435;
  assign n3167 = n3163 & ~n3166;
  assign n3169 = n3162 & n3168;
  assign n3170 = n2176 & n3027;
  assign n3171 = ~n3169 & ~n3170;
  assign n3172 = ~n3167 & n3171;
  assign n3173 = n3172 ^ n3154;
  assign n3174 = ~n3155 & ~n3173;
  assign n3175 = n3174 ^ n3146;
  assign n3180 = n3179 ^ n3175;
  assign n3181 = ~n2087 & n3029;
  assign n3182 = n1837 & n3031;
  assign n3183 = ~n1694 & n3035;
  assign n3184 = ~n3182 & ~n3183;
  assign n3185 = ~n3181 & n3184;
  assign n3186 = n2436 & n3185;
  assign n3187 = n2201 ^ n2087;
  assign n3188 = n3159 & ~n3187;
  assign n3189 = n3186 & ~n3188;
  assign n3190 = n2432 & ~n3185;
  assign n3191 = ~n3126 & ~n3187;
  assign n3192 = ~n3190 & ~n3191;
  assign n3193 = ~n3189 & n3192;
  assign n3194 = n3193 ^ n3179;
  assign n3195 = n3180 & n3194;
  assign n3196 = n3195 ^ n3175;
  assign n3197 = n3196 ^ n3114;
  assign n3198 = n3130 & n3197;
  assign n3199 = n3198 ^ n3129;
  assign n3200 = n3199 ^ n3099;
  assign n3201 = n3108 & ~n3200;
  assign n3202 = n3201 ^ n3107;
  assign n3203 = n3098 & ~n3202;
  assign n3204 = n2343 & n3028;
  assign n3205 = n3204 ^ n2340;
  assign n3206 = x0 & n3205;
  assign n3207 = x1 & n2085;
  assign n3208 = ~n2086 & n2430;
  assign n3209 = ~x0 & ~n3208;
  assign n3210 = ~n3207 & n3209;
  assign n3211 = ~n3206 & ~n3210;
  assign n3212 = n3211 ^ n2436;
  assign n3213 = n2712 ^ n2645;
  assign n3214 = n2569 & n3028;
  assign n3215 = n3214 ^ n2428;
  assign n3216 = x0 & n3215;
  assign n3217 = ~n2340 & n3031;
  assign n3218 = n2085 & n3035;
  assign n3219 = ~n3217 & ~n3218;
  assign n3220 = ~n3216 & n3219;
  assign n3221 = n3220 ^ n3211;
  assign n3222 = ~n3213 & ~n3221;
  assign n3223 = ~n3212 & n3222;
  assign n3224 = n3223 ^ n3212;
  assign n3225 = ~n3203 & ~n3224;
  assign n3226 = n3220 ^ n2436;
  assign n3227 = n3226 ^ n3213;
  assign n3228 = ~n3098 & n3202;
  assign n3229 = n3228 ^ n3226;
  assign n3230 = n3227 & ~n3229;
  assign n3231 = n3230 ^ n3213;
  assign n3232 = ~n3225 & ~n3231;
  assign n3233 = n3232 ^ n3088;
  assign n3234 = n3097 & n3233;
  assign n3235 = n3234 ^ n3096;
  assign n3236 = n3235 ^ n3077;
  assign n3237 = n3087 & n3236;
  assign n3238 = n3237 ^ n3086;
  assign n3239 = n3238 ^ n3065;
  assign n3240 = ~n3076 & n3239;
  assign n3241 = n3240 ^ n3075;
  assign n3259 = n3258 ^ n3241;
  assign n3260 = n2724 ^ n2567;
  assign n3261 = n3260 ^ n3258;
  assign n3262 = ~n3259 & n3261;
  assign n3263 = n3262 ^ n3241;
  assign n3264 = ~n3064 & ~n3263;
  assign n3387 = ~n382 & ~n523;
  assign n3388 = ~n394 & n3387;
  assign n3389 = n2363 & n3388;
  assign n3390 = n1862 & n3389;
  assign n3391 = ~n264 & ~n411;
  assign n3392 = n3390 & n3391;
  assign n3393 = ~n259 & n3392;
  assign n3394 = ~n422 & ~n485;
  assign n3395 = ~n180 & n3394;
  assign n3396 = n84 & ~n149;
  assign n3397 = n400 & ~n3396;
  assign n3398 = n3395 & n3397;
  assign n3399 = n1777 & n3398;
  assign n3400 = n118 & ~n199;
  assign n3401 = n333 & n3400;
  assign n3402 = n3399 & n3401;
  assign n3403 = n85 & ~n174;
  assign n3404 = n2510 & ~n3403;
  assign n3405 = n724 & n3404;
  assign n3406 = n3402 & n3405;
  assign n3407 = n3393 & n3406;
  assign n3408 = n3263 & ~n3407;
  assign n3409 = ~n57 & ~n471;
  assign n3410 = ~n419 & n3409;
  assign n3411 = n155 & n176;
  assign n3412 = ~n3410 & ~n3411;
  assign n3413 = n1007 & ~n3412;
  assign n275 = ~n273 & ~n274;
  assign n276 = ~n272 & n275;
  assign n3414 = ~n131 & ~n424;
  assign n3415 = n276 & n3414;
  assign n3416 = n1754 & n3415;
  assign n3417 = n3413 & n3416;
  assign n3418 = ~n316 & ~n341;
  assign n3419 = n736 & n3418;
  assign n3420 = n3417 & n3419;
  assign n3421 = ~n188 & ~n372;
  assign n3422 = n2911 & n3421;
  assign n3423 = n609 & n3422;
  assign n3424 = n140 & ~n152;
  assign n3425 = ~n130 & n3424;
  assign n3426 = ~n708 & ~n3425;
  assign n3427 = ~n345 & ~n3426;
  assign n3428 = n3423 & n3427;
  assign n3429 = n1527 & n3428;
  assign n3430 = ~n180 & ~n418;
  assign n3431 = n57 & ~n174;
  assign n3432 = ~n505 & ~n3431;
  assign n3433 = n3430 & n3432;
  assign n3434 = n282 & n664;
  assign n3435 = n3433 & n3434;
  assign n3436 = ~n200 & ~n649;
  assign n3437 = n101 & ~n779;
  assign n3438 = ~n2277 & ~n3437;
  assign n3439 = n3436 & n3438;
  assign n3440 = n3435 & n3439;
  assign n3441 = n3429 & n3440;
  assign n3442 = n3420 & n3441;
  assign n3443 = n3408 & ~n3442;
  assign n3444 = n3064 & ~n3443;
  assign n3445 = n3063 ^ n3062;
  assign n3446 = ~n3444 & ~n3445;
  assign n3447 = ~n3264 & ~n3446;
  assign n3267 = n3034 ^ n2431;
  assign n3268 = x1 & n3267;
  assign n3269 = n2430 & n2929;
  assign n3270 = ~x0 & ~n3269;
  assign n3271 = ~n3268 & n3270;
  assign n2986 = n2984 & n2985;
  assign n2952 = n91 & n2809;
  assign n2953 = n50 & ~n2952;
  assign n2954 = n806 & ~n2953;
  assign n2955 = n97 & n317;
  assign n2956 = ~n56 & ~n165;
  assign n2957 = ~n2955 & ~n2956;
  assign n2958 = ~n385 & ~n488;
  assign n2959 = ~n2957 & n2958;
  assign n2960 = n51 & ~n793;
  assign n2961 = ~n523 & ~n2960;
  assign n2962 = n360 & n2961;
  assign n2963 = n2959 & n2962;
  assign n2964 = n798 & n2963;
  assign n2965 = n774 & n2964;
  assign n2966 = n2954 & n2965;
  assign n3032 = n2986 ^ n2966;
  assign n3275 = n3032 ^ x22;
  assign n3005 = n2928 & n3001;
  assign n3006 = ~n2984 & ~n3005;
  assign n3007 = ~n3004 & n3006;
  assign n3018 = n3016 & n3017;
  assign n3019 = n2984 & ~n3018;
  assign n3272 = ~n3007 & ~n3019;
  assign n3273 = n3028 & ~n3272;
  assign n3274 = n3273 ^ x1;
  assign n3276 = n3275 ^ n3274;
  assign n3277 = x0 & ~n3276;
  assign n3278 = ~n3271 & ~n3277;
  assign n2794 = n1057 & n2535;
  assign n2795 = ~n2548 & ~n2794;
  assign n2796 = n2438 & ~n2473;
  assign n2797 = n2796 ^ n2437;
  assign n2798 = ~n2795 & n2797;
  assign n2799 = n2474 & n2535;
  assign n2800 = n2442 & n2473;
  assign n2801 = ~n2799 & ~n2800;
  assign n2802 = ~n2798 & n2801;
  assign n2803 = n969 & ~n2802;
  assign n2828 = n2827 ^ n1057;
  assign n2829 = n2484 & ~n2828;
  assign n2830 = n2805 & n2829;
  assign n2831 = ~n2803 & ~n2830;
  assign n2832 = ~n2805 & n2827;
  assign n2833 = n2571 & n2832;
  assign n2834 = n2831 & ~n2833;
  assign n2835 = ~n969 & n2802;
  assign n2836 = ~n2805 & ~n2827;
  assign n2837 = n2484 & ~n2836;
  assign n2838 = n2835 & ~n2837;
  assign n2839 = n2834 & ~n2838;
  assign n2777 = n1855 & n2570;
  assign n2778 = n2101 & ~n2340;
  assign n2779 = n2085 & n2104;
  assign n2780 = ~n2778 & ~n2779;
  assign n2781 = ~n2777 & n2780;
  assign n2782 = n310 & ~n2781;
  assign n2783 = n1855 & ~n2586;
  assign n2784 = ~n310 & n2780;
  assign n2785 = ~n2783 & n2784;
  assign n2786 = n2428 ^ n756;
  assign n2787 = n1855 & n2569;
  assign n2788 = n2786 & n2787;
  assign n2789 = ~n2785 & ~n2788;
  assign n2790 = ~n2782 & n2789;
  assign n2761 = n313 & ~n2132;
  assign n2762 = n1698 & ~n2087;
  assign n2763 = n1703 & n1837;
  assign n2764 = ~n2762 & ~n2763;
  assign n2765 = ~n308 & n2764;
  assign n2766 = ~n2761 & n2765;
  assign n2767 = n2125 & n2258;
  assign n2768 = n308 & ~n2764;
  assign n2769 = ~n2767 & ~n2768;
  assign n2770 = ~n2766 & n2769;
  assign n2771 = n313 & n2124;
  assign n2772 = n2086 ^ n315;
  assign n2773 = n2771 & n2772;
  assign n2774 = n2770 & ~n2773;
  assign n2737 = n1617 & n2239;
  assign n2738 = n2737 ^ n1694;
  assign n2739 = n1734 & n2738;
  assign n2740 = ~n989 & n1611;
  assign n2741 = n989 & ~n1079;
  assign n2742 = n1612 & n2741;
  assign n2743 = n2230 & ~n2742;
  assign n2744 = ~n2740 & n2743;
  assign n2745 = n989 & n1611;
  assign n2746 = ~n989 & n1079;
  assign n2747 = n1612 & n2746;
  assign n2748 = n1739 & ~n2747;
  assign n2749 = ~n2745 & n2748;
  assign n2750 = ~n2744 & ~n2749;
  assign n2751 = ~n2739 & n2750;
  assign n2752 = ~n2237 & n2251;
  assign n2753 = ~n1079 & n1614;
  assign n2757 = ~n2752 & n2753;
  assign n2754 = n2753 ^ n1614;
  assign n2755 = ~n2752 & ~n2754;
  assign n2756 = n2755 ^ n1614;
  assign n2758 = n2757 ^ n2756;
  assign n2759 = ~n2751 & n2758;
  assign n2760 = n2759 ^ n2757;
  assign n2775 = n2774 ^ n2760;
  assign n2734 = n2252 ^ n2229;
  assign n2735 = ~n2272 & ~n2734;
  assign n2736 = n2735 ^ n2271;
  assign n2776 = n2775 ^ n2736;
  assign n2791 = n2790 ^ n2776;
  assign n2731 = n2273 ^ n2226;
  assign n2732 = n2360 & ~n2731;
  assign n2733 = n2732 ^ n2359;
  assign n2792 = n2791 ^ n2733;
  assign n2728 = n2727 ^ n2361;
  assign n2729 = n2539 & ~n2728;
  assign n2730 = n2729 ^ n2538;
  assign n2793 = n2792 ^ n2730;
  assign n3266 = n2839 ^ n2793;
  assign n3448 = n3278 ^ n3266;
  assign n3449 = ~n3447 & ~n3448;
  assign n3450 = ~n3064 & n3442;
  assign n3451 = n3448 & ~n3450;
  assign n3265 = ~n3062 & ~n3063;
  assign n3452 = n3265 & ~n3408;
  assign n3453 = n3451 & ~n3452;
  assign n3454 = n3264 & n3407;
  assign n3455 = n3453 & ~n3454;
  assign n3456 = ~n3449 & ~n3455;
  assign n3457 = ~n3407 & n3445;
  assign n3458 = ~n3408 & n3442;
  assign n3459 = ~n3457 & n3458;
  assign n3460 = ~n3456 & ~n3459;
  assign n3461 = ~n137 & ~n250;
  assign n3462 = ~n281 & ~n1550;
  assign n3463 = ~n343 & ~n769;
  assign n3464 = n3462 & n3463;
  assign n3465 = n580 & n3464;
  assign n3466 = n1860 & n2980;
  assign n3467 = n101 & ~n2809;
  assign n3468 = ~n468 & ~n3467;
  assign n3469 = ~n78 & n84;
  assign n3470 = ~n497 & ~n3469;
  assign n3471 = ~n288 & n3470;
  assign n3472 = n3468 & n3471;
  assign n3473 = n3466 & n3472;
  assign n3474 = n3465 & n3473;
  assign n3475 = n443 & n3474;
  assign n3476 = ~n3461 & n3475;
  assign n3477 = n391 & ~n410;
  assign n3478 = ~n183 & ~n539;
  assign n3479 = n57 & ~n170;
  assign n3480 = ~n463 & ~n3479;
  assign n3481 = n3478 & n3480;
  assign n3482 = n2923 & n3481;
  assign n3483 = n697 & n3482;
  assign n3484 = n297 & n2511;
  assign n3485 = ~n353 & n715;
  assign n3486 = n846 & n3485;
  assign n3487 = n2286 & n3486;
  assign n3488 = n3484 & n3487;
  assign n3489 = n3483 & n3488;
  assign n3490 = n3477 & n3489;
  assign n3491 = n3476 & n3490;
  assign n3492 = n3460 & ~n3491;
  assign n3279 = n3266 & ~n3278;
  assign n3280 = ~n3265 & ~n3279;
  assign n3281 = ~n3264 & n3280;
  assign n3282 = ~n3266 & n3278;
  assign n3283 = ~n3281 & ~n3282;
  assign n3008 = n2966 & ~n2986;
  assign n3009 = ~n3007 & n3008;
  assign n3020 = n3019 ^ n2986;
  assign n3021 = n2966 & ~n3020;
  assign n3022 = n3021 ^ n3019;
  assign n3023 = ~n3009 & n3022;
  assign n2987 = n2966 & n2986;
  assign n2988 = ~n278 & n2954;
  assign n2989 = n78 & n361;
  assign n2990 = n164 & ~n2989;
  assign n2991 = ~n288 & ~n2990;
  assign n2992 = ~n456 & n2991;
  assign n2993 = n255 & n776;
  assign n2994 = ~n81 & n2993;
  assign n2995 = n50 & ~n2994;
  assign n2996 = n1776 & ~n2995;
  assign n2997 = n2992 & n2996;
  assign n2998 = n783 & n2997;
  assign n2999 = n2988 & n2998;
  assign n3000 = ~n2987 & ~n2999;
  assign n3024 = n3023 ^ n3000;
  assign n3030 = n3000 & n3029;
  assign n3033 = n3031 & ~n3032;
  assign n3036 = ~n3034 & n3035;
  assign n3037 = ~n3033 & ~n3036;
  assign n3038 = ~n3030 & n3037;
  assign n3041 = n2433 & ~n3040;
  assign n3042 = n3038 & n3041;
  assign n3043 = ~n3027 & ~n3042;
  assign n3044 = n3024 & ~n3043;
  assign n3045 = n2432 & ~n3038;
  assign n3046 = ~n3044 & ~n3045;
  assign n3047 = n2436 & n3038;
  assign n3048 = ~n3024 & n3047;
  assign n3049 = n3046 & ~n3048;
  assign n2931 = ~n2485 & n2929;
  assign n2932 = n2931 ^ n969;
  assign n2933 = n2484 & n2932;
  assign n2934 = ~n2930 & n2933;
  assign n2935 = n2902 & ~n2929;
  assign n2936 = n2639 & n2935;
  assign n2937 = ~n2934 & ~n2936;
  assign n2938 = ~n2902 & n2929;
  assign n2939 = n2558 & ~n2938;
  assign n2940 = n2440 & n2794;
  assign n2941 = ~n2476 & n2827;
  assign n2942 = ~n2940 & ~n2941;
  assign n2943 = ~n969 & ~n2942;
  assign n2944 = n2438 & n2535;
  assign n2945 = n969 & ~n2944;
  assign n2946 = ~n2941 & n2945;
  assign n2947 = ~n2943 & ~n2946;
  assign n2948 = ~n2939 & n2947;
  assign n2949 = n2937 & ~n2948;
  assign n2880 = n1855 & n2559;
  assign n2881 = n2101 & n2428;
  assign n2882 = n2104 & ~n2340;
  assign n2883 = ~n2881 & ~n2882;
  assign n2884 = ~n2880 & n2883;
  assign n2885 = n310 & ~n2884;
  assign n2886 = n1855 & ~n2544;
  assign n2887 = ~n310 & n2883;
  assign n2888 = ~n2886 & n2887;
  assign n2889 = n1855 & n2543;
  assign n2890 = n2473 ^ n756;
  assign n2891 = n2889 & n2890;
  assign n2892 = ~n2888 & ~n2891;
  assign n2893 = ~n2885 & n2892;
  assign n2864 = n313 & n2095;
  assign n2865 = n1698 & ~n2086;
  assign n2866 = n1703 & ~n2087;
  assign n2867 = ~n2865 & ~n2866;
  assign n2868 = ~n2864 & n2867;
  assign n2869 = ~n308 & ~n2868;
  assign n2870 = n313 & ~n2109;
  assign n2871 = n308 & n2867;
  assign n2872 = ~n2870 & n2871;
  assign n2873 = n313 & n2094;
  assign n2874 = n2085 ^ n315;
  assign n2875 = n2873 & n2874;
  assign n2876 = ~n2872 & ~n2875;
  assign n2877 = ~n2869 & n2876;
  assign n2856 = n1748 & n2239;
  assign n2857 = n2856 ^ n1837;
  assign n2858 = n1734 & n2857;
  assign n2859 = ~n1694 & ~n2244;
  assign n2860 = n1611 & n2248;
  assign n2861 = ~n2859 & ~n2860;
  assign n2862 = ~n2858 & n2861;
  assign n2849 = ~n1079 & ~n1614;
  assign n2850 = ~n2752 & ~n2849;
  assign n2851 = ~n2751 & ~n2850;
  assign n2852 = n2851 ^ n1612;
  assign n2853 = ~n2851 & ~n2852;
  assign n2854 = n1079 & n2853;
  assign n2855 = n2854 ^ n2852;
  assign n2863 = n2862 ^ n2855;
  assign n2878 = n2877 ^ n2863;
  assign n2846 = n2760 ^ n2736;
  assign n2847 = ~n2775 & n2846;
  assign n2848 = n2847 ^ n2774;
  assign n2879 = n2878 ^ n2848;
  assign n2894 = n2893 ^ n2879;
  assign n2843 = n2776 ^ n2733;
  assign n2844 = ~n2791 & n2843;
  assign n2845 = n2844 ^ n2790;
  assign n2895 = n2894 ^ n2845;
  assign n2950 = n2949 ^ n2895;
  assign n2840 = n2839 ^ n2730;
  assign n2841 = n2793 & n2840;
  assign n2842 = n2841 ^ n2839;
  assign n2951 = n2950 ^ n2842;
  assign n3050 = n3049 ^ n2951;
  assign n3493 = n3283 ^ n3050;
  assign n3494 = n3492 & ~n3493;
  assign n3495 = ~n3460 & n3491;
  assign n3496 = n3493 & n3495;
  assign n3497 = ~n3494 & ~n3496;
  assign n3358 = x1 & n3000;
  assign n3359 = n2430 & ~n3032;
  assign n3360 = ~x0 & ~n3359;
  assign n3361 = ~n3358 & n3360;
  assign n3376 = n2999 & n3022;
  assign n3377 = n3000 & ~n3009;
  assign n3378 = ~n3376 & ~n3377;
  assign n3379 = n3028 & n3378;
  assign n3362 = n243 & n506;
  assign n3363 = n57 & ~n3362;
  assign n3364 = ~n129 & ~n644;
  assign n3365 = n100 & ~n116;
  assign n3366 = n3364 & ~n3365;
  assign n3367 = ~n3363 & n3366;
  assign n3368 = ~n287 & ~n424;
  assign n3369 = n3367 & n3368;
  assign n3370 = ~n354 & ~n545;
  assign n3371 = n162 & n3370;
  assign n3372 = n100 & ~n2994;
  assign n3373 = n3371 & ~n3372;
  assign n3374 = n3369 & n3373;
  assign n3375 = n1027 & n3374;
  assign n3380 = n3379 ^ n3375;
  assign n3381 = x0 & n3380;
  assign n3382 = ~n3361 & ~n3381;
  assign n3383 = n3382 ^ n2436;
  assign n3339 = ~n2496 & n2535;
  assign n3340 = n1855 & n3339;
  assign n3341 = n2101 & n2473;
  assign n3342 = n2104 & n2428;
  assign n3343 = ~n3341 & ~n3342;
  assign n3344 = ~n3340 & n3343;
  assign n3345 = n310 & ~n3344;
  assign n3346 = ~n2496 & ~n2535;
  assign n3347 = n1855 & ~n3346;
  assign n3348 = ~n310 & n3343;
  assign n3349 = ~n3347 & n3348;
  assign n3350 = n1855 & n2496;
  assign n3351 = n2535 ^ n756;
  assign n3352 = n3350 & n3351;
  assign n3353 = ~n3349 & ~n3352;
  assign n3354 = ~n3345 & n3353;
  assign n3322 = n313 & n2344;
  assign n3323 = n1698 & n2085;
  assign n3324 = n1703 & ~n2086;
  assign n3325 = ~n3323 & ~n3324;
  assign n3326 = ~n3322 & n3325;
  assign n3327 = ~n308 & ~n3326;
  assign n3328 = n313 & ~n2351;
  assign n3329 = n308 & n3325;
  assign n3330 = ~n3328 & n3329;
  assign n3331 = n313 & n2343;
  assign n3332 = n2340 ^ n315;
  assign n3333 = n3331 & ~n3332;
  assign n3334 = ~n3330 & ~n3333;
  assign n3335 = ~n3327 & n3334;
  assign n3316 = n2862 ^ n2851;
  assign n3317 = n2852 & ~n3316;
  assign n3318 = n3317 ^ n1612;
  assign n3319 = n3318 ^ n1611;
  assign n3320 = ~n1079 & ~n3319;
  assign n3309 = n2201 & n2239;
  assign n3310 = n3309 ^ n2087;
  assign n3311 = n1734 & ~n3310;
  assign n3312 = n1837 & ~n2244;
  assign n3313 = ~n1694 & n2248;
  assign n3314 = ~n3312 & ~n3313;
  assign n3315 = ~n3311 & n3314;
  assign n3321 = n3320 ^ n3315;
  assign n3336 = n3335 ^ n3321;
  assign n3306 = n2863 ^ n2848;
  assign n3307 = ~n2878 & ~n3306;
  assign n3308 = n3307 ^ n2877;
  assign n3337 = n3336 ^ n3308;
  assign n3303 = n2893 ^ n2845;
  assign n3304 = n2894 & n3303;
  assign n3305 = n3304 ^ n2845;
  assign n3338 = n3337 ^ n3305;
  assign n3355 = n3354 ^ n3338;
  assign n3300 = n2949 ^ n2842;
  assign n3301 = n2950 & n3300;
  assign n3302 = n3301 ^ n2842;
  assign n3356 = n3355 ^ n3302;
  assign n3287 = n2485 & n3057;
  assign n3288 = n3287 ^ n969;
  assign n3289 = n3288 ^ n3034;
  assign n3290 = n2484 & n3289;
  assign n3291 = n969 & ~n2827;
  assign n3292 = n2438 & ~n3291;
  assign n3293 = n2442 & ~n2827;
  assign n3294 = ~n3292 & ~n3293;
  assign n3295 = n2479 & n2929;
  assign n3296 = n3294 & ~n3295;
  assign n3297 = n2477 & ~n2929;
  assign n3298 = n3296 & ~n3297;
  assign n3299 = ~n3290 & n3298;
  assign n3357 = n3356 ^ n3299;
  assign n3384 = n3383 ^ n3357;
  assign n3284 = n3283 ^ n3049;
  assign n3285 = ~n3050 & n3284;
  assign n3286 = n3285 ^ n3283;
  assign n3385 = n3384 ^ n3286;
  assign n277 = ~n271 & n276;
  assign n283 = ~n195 & n282;
  assign n284 = n279 & n283;
  assign n285 = n277 & n284;
  assign n302 = n292 & n301;
  assign n303 = n285 & n302;
  assign n304 = n270 & n303;
  assign n305 = n250 & n304;
  assign n306 = n187 & n305;
  assign n3386 = n3385 ^ n306;
  assign n3498 = n3497 ^ n3386;
  assign n3637 = x23 ^ x22;
  assign n3638 = n3637 ^ n306;
  assign n3639 = ~n3386 & n3638;
  assign n3640 = n3639 ^ n3385;
  assign n3641 = n3496 & ~n3640;
  assign n3642 = n306 & ~n3385;
  assign n3643 = ~n3637 & n3642;
  assign n3644 = n3643 ^ n3640;
  assign n3645 = ~n3494 & n3644;
  assign n3646 = n3645 ^ n3640;
  assign n3647 = ~n3641 & ~n3646;
  assign n3648 = ~n306 & n3385;
  assign n3649 = ~n3496 & n3648;
  assign n3650 = n3637 & n3649;
  assign n3651 = n3647 & ~n3650;
  assign n3607 = n2430 & n3000;
  assign n3608 = x1 & ~n3375;
  assign n3609 = ~x0 & ~n3608;
  assign n3610 = ~n3607 & n3609;
  assign n3626 = ~n3375 & ~n3376;
  assign n3627 = n3375 & ~n3377;
  assign n3628 = ~n3626 & ~n3627;
  assign n3629 = n3028 & n3628;
  assign n3514 = ~n289 & ~n569;
  assign n3515 = ~n485 & n3514;
  assign n3611 = n152 & ~n1004;
  assign n3612 = n3515 & ~n3611;
  assign n3613 = n891 & n3612;
  assign n3614 = n132 & n1514;
  assign n3615 = n3613 & n3614;
  assign n3616 = n617 & n706;
  assign n3617 = n130 & ~n3616;
  assign n3618 = n791 & ~n3617;
  assign n3619 = ~n331 & n2367;
  assign n3620 = ~n463 & n3619;
  assign n3621 = ~n447 & n3620;
  assign n3622 = n3618 & n3621;
  assign n3623 = n725 & n3622;
  assign n3624 = n3615 & n3623;
  assign n3625 = n437 & n3624;
  assign n3630 = n3629 ^ n3625;
  assign n3631 = x0 & n3630;
  assign n3632 = ~n3610 & ~n3631;
  assign n3633 = n3632 ^ n2436;
  assign n3589 = ~n3032 & ~n3272;
  assign n3590 = n2571 & n3589;
  assign n3591 = ~n2476 & ~n3034;
  assign n3592 = n2577 & ~n2929;
  assign n3593 = ~n3591 & ~n3592;
  assign n3594 = n969 & ~n3593;
  assign n3595 = ~n3590 & ~n3594;
  assign n3596 = n2484 & n3272;
  assign n3597 = n3032 ^ n1057;
  assign n3598 = n3596 & n3597;
  assign n3599 = n3595 & ~n3598;
  assign n3600 = n3032 & ~n3272;
  assign n3601 = n2484 & ~n3600;
  assign n3602 = ~n969 & n3593;
  assign n3603 = ~n3601 & n3602;
  assign n3604 = n3599 & ~n3603;
  assign n3573 = n1855 & n2832;
  assign n3574 = n2101 & n2535;
  assign n3575 = n2104 & n2473;
  assign n3576 = ~n3574 & ~n3575;
  assign n3577 = ~n3573 & n3576;
  assign n3578 = ~n310 & ~n3577;
  assign n3579 = n1855 & ~n2836;
  assign n3580 = n310 & n3576;
  assign n3581 = ~n3579 & n3580;
  assign n3582 = n2827 ^ n756;
  assign n3583 = n1855 & ~n3582;
  assign n3584 = n2805 & n3583;
  assign n3585 = ~n3581 & ~n3584;
  assign n3586 = ~n3578 & n3585;
  assign n3557 = n2258 & n2570;
  assign n3558 = n1698 & ~n2340;
  assign n3559 = n1703 & n2085;
  assign n3560 = ~n3558 & ~n3559;
  assign n3561 = n308 & ~n3560;
  assign n3562 = ~n3557 & ~n3561;
  assign n3563 = n313 & ~n2586;
  assign n3564 = ~n308 & n3560;
  assign n3565 = ~n3563 & n3564;
  assign n3566 = n3562 & ~n3565;
  assign n3567 = n2428 ^ n315;
  assign n3568 = n313 & n2569;
  assign n3569 = ~n3567 & n3568;
  assign n3570 = n3566 & ~n3569;
  assign n3549 = n1611 & n3318;
  assign n3550 = ~n3315 & ~n3549;
  assign n3551 = ~n1611 & ~n3318;
  assign n3552 = ~n1079 & ~n3551;
  assign n3553 = ~n3550 & n3552;
  assign n3554 = n3553 ^ n1694;
  assign n3555 = ~n1079 & n3554;
  assign n3534 = n2124 & n2239;
  assign n3535 = n3534 ^ n2086;
  assign n3536 = n1734 & n3535;
  assign n3537 = n1837 & n2741;
  assign n3538 = n2230 & ~n3537;
  assign n3539 = ~n2087 & n2234;
  assign n3540 = n3539 ^ n1739;
  assign n3541 = ~n3538 & ~n3540;
  assign n3542 = ~n308 & ~n2087;
  assign n3543 = n308 & n1079;
  assign n3544 = n1837 & n3543;
  assign n3545 = ~n3542 & ~n3544;
  assign n3546 = ~n989 & ~n3545;
  assign n3547 = ~n3541 & ~n3546;
  assign n3548 = ~n3536 & ~n3547;
  assign n3556 = n3555 ^ n3548;
  assign n3571 = n3570 ^ n3556;
  assign n3531 = n3321 ^ n3308;
  assign n3532 = n3336 & ~n3531;
  assign n3533 = n3532 ^ n3335;
  assign n3572 = n3571 ^ n3533;
  assign n3587 = n3586 ^ n3572;
  assign n3528 = n3354 ^ n3305;
  assign n3529 = n3338 & n3528;
  assign n3530 = n3529 ^ n3354;
  assign n3588 = n3587 ^ n3530;
  assign n3605 = n3604 ^ n3588;
  assign n3525 = n3355 ^ n3299;
  assign n3526 = ~n3356 & n3525;
  assign n3527 = n3526 ^ n3302;
  assign n3606 = n3605 ^ n3527;
  assign n3634 = n3633 ^ n3606;
  assign n3522 = n3383 ^ n3286;
  assign n3523 = n3384 & ~n3522;
  assign n3524 = n3523 ^ n3286;
  assign n3635 = n3634 ^ n3524;
  assign n3499 = ~n424 & ~n563;
  assign n3500 = n85 & ~n793;
  assign n3501 = ~n600 & ~n3500;
  assign n3502 = n3499 & n3501;
  assign n3503 = n297 & n3502;
  assign n3504 = n57 & ~n2917;
  assign n3505 = ~n998 & ~n3504;
  assign n3506 = n3387 & n3505;
  assign n3507 = n3503 & n3506;
  assign n3508 = n2041 & n3507;
  assign n3509 = n260 & ~n447;
  assign n3510 = ~n372 & ~n453;
  assign n3511 = n3509 & n3510;
  assign n3512 = n3508 & n3511;
  assign n3513 = n3474 & n3512;
  assign n3516 = n2958 & n3515;
  assign n3517 = n3484 & n3516;
  assign n3518 = ~n344 & ~n3517;
  assign n3519 = ~n428 & ~n919;
  assign n3520 = ~n3518 & n3519;
  assign n3521 = n3513 & n3520;
  assign n3636 = n3635 ^ n3521;
  assign n3652 = n3651 ^ n3636;
  assign n3655 = n3491 ^ n3460;
  assign n3656 = n3493 ^ n3491;
  assign n3657 = ~n3655 & ~n3656;
  assign n3658 = n3657 ^ n3460;
  assign n3665 = ~n3642 & n3658;
  assign n3666 = ~n3494 & n3665;
  assign n3667 = n3636 & ~n3648;
  assign n3668 = ~n3666 & n3667;
  assign n3669 = n3496 ^ n3385;
  assign n3670 = n3636 ^ n306;
  assign n3671 = n3386 & n3670;
  assign n3672 = n3669 & n3671;
  assign n3673 = n3672 ^ n3636;
  assign n3674 = ~n3668 & n3673;
  assign n3653 = n3636 & ~n3642;
  assign n3654 = n3494 & ~n3653;
  assign n3659 = ~n3386 & ~n3496;
  assign n3660 = ~n3658 & n3659;
  assign n3661 = ~n3654 & ~n3660;
  assign n3662 = n3494 & n3648;
  assign n3663 = ~n3636 & ~n3662;
  assign n3664 = ~n3661 & ~n3663;
  assign n3677 = ~n3637 & ~n3664;
  assign n3678 = ~n3674 & ~n3677;
  assign n3675 = n3637 & ~n3674;
  assign n3676 = ~n3664 & ~n3675;
  assign n3679 = n3678 ^ n3676;
  assign n3803 = ~n3521 & ~n3635;
  assign n3804 = ~n3648 & ~n3803;
  assign n3805 = ~n3665 & n3804;
  assign n3806 = n3521 & n3635;
  assign n3807 = ~n3805 & ~n3806;
  assign n3786 = n3625 ^ n2431;
  assign n3787 = x1 & n3786;
  assign n3788 = n2430 & n3375;
  assign n3789 = ~x0 & ~n3788;
  assign n3790 = ~n3787 & n3789;
  assign n3791 = n3627 ^ n3626;
  assign n3792 = ~n3625 & n3791;
  assign n3793 = n3792 ^ n3626;
  assign n3794 = n3028 & ~n3793;
  assign n3795 = n3794 ^ x1;
  assign n3796 = n3795 ^ x22;
  assign n3797 = x0 & n3796;
  assign n3798 = ~n3790 & ~n3797;
  assign n3763 = ~n3000 & ~n3023;
  assign n3764 = n2484 & ~n3763;
  assign n3765 = n1057 & ~n3032;
  assign n3766 = n2548 & ~n3034;
  assign n3767 = ~n3765 & ~n3766;
  assign n3768 = n2437 & ~n3767;
  assign n3769 = n2474 & ~n3032;
  assign n3770 = n2442 & ~n3034;
  assign n3771 = ~n3769 & ~n3770;
  assign n3772 = ~n3768 & n3771;
  assign n3773 = n969 & n3772;
  assign n3774 = ~n3764 & n3773;
  assign n3775 = ~n3000 & n3023;
  assign n3776 = n2639 & n3775;
  assign n3777 = ~n969 & ~n3772;
  assign n3778 = ~n3776 & ~n3777;
  assign n3779 = ~n3774 & n3778;
  assign n3780 = n3023 & n3773;
  assign n3781 = ~n2558 & ~n3780;
  assign n3782 = n1057 & n3023;
  assign n3783 = n3000 & ~n3782;
  assign n3784 = ~n3781 & n3783;
  assign n3785 = n3779 & ~n3784;
  assign n3799 = n3798 ^ n3785;
  assign n3738 = n2827 ^ n310;
  assign n3739 = n2097 & n3738;
  assign n3740 = ~n756 & ~n2098;
  assign n3741 = ~n756 & ~n2535;
  assign n3742 = ~n310 & n3741;
  assign n3743 = ~n3740 & ~n3742;
  assign n3744 = ~n3739 & ~n3743;
  assign n3745 = ~n310 & n2098;
  assign n3746 = n2827 & n3745;
  assign n3747 = n310 & n2097;
  assign n3748 = ~n2535 & n3747;
  assign n3749 = n756 & ~n3748;
  assign n3750 = ~n3746 & n3749;
  assign n3751 = ~n3744 & ~n3750;
  assign n3752 = n310 & ~n2827;
  assign n3753 = n2098 & n3752;
  assign n3754 = ~n3751 & ~n3753;
  assign n3755 = ~n1898 & n2902;
  assign n3756 = n3755 ^ n310;
  assign n3757 = n3756 ^ n2929;
  assign n3758 = n1855 & ~n3757;
  assign n3759 = n3754 & ~n3758;
  assign n3722 = n313 & ~n2544;
  assign n3723 = n1698 & n2428;
  assign n3724 = n1703 & ~n2340;
  assign n3725 = ~n3723 & ~n3724;
  assign n3726 = ~n308 & n3725;
  assign n3727 = ~n3722 & n3726;
  assign n3728 = n2258 & n2559;
  assign n3729 = n308 & ~n3725;
  assign n3730 = ~n3728 & ~n3729;
  assign n3731 = ~n3727 & n3730;
  assign n3732 = n2473 ^ n315;
  assign n3733 = n313 & n2543;
  assign n3734 = ~n3732 & n3733;
  assign n3735 = n3731 & ~n3734;
  assign n3716 = n3553 ^ n3548;
  assign n3717 = ~n3554 & n3716;
  assign n3718 = n3717 ^ n1694;
  assign n3719 = n3718 ^ n1837;
  assign n3720 = ~n1079 & n3719;
  assign n3709 = n2094 & n2239;
  assign n3710 = n3709 ^ n2085;
  assign n3711 = n1734 & n3710;
  assign n3712 = ~n2086 & ~n2244;
  assign n3713 = ~n2087 & n2248;
  assign n3714 = ~n3712 & ~n3713;
  assign n3715 = ~n3711 & n3714;
  assign n3721 = n3720 ^ n3715;
  assign n3736 = n3735 ^ n3721;
  assign n3706 = n3556 ^ n3533;
  assign n3707 = n3571 & n3706;
  assign n3708 = n3707 ^ n3570;
  assign n3737 = n3736 ^ n3708;
  assign n3760 = n3759 ^ n3737;
  assign n3703 = n3572 ^ n3530;
  assign n3704 = n3587 & n3703;
  assign n3705 = n3704 ^ n3586;
  assign n3761 = n3760 ^ n3705;
  assign n3700 = n3604 ^ n3527;
  assign n3701 = ~n3605 & n3700;
  assign n3702 = n3701 ^ n3527;
  assign n3762 = n3761 ^ n3702;
  assign n3800 = n3799 ^ n3762;
  assign n3697 = n3633 ^ n3524;
  assign n3698 = ~n3634 & ~n3697;
  assign n3699 = n3698 ^ n3524;
  assign n3801 = n3800 ^ n3699;
  assign n3680 = n174 & n236;
  assign n3681 = n130 & ~n3680;
  assign n3682 = ~n2277 & ~n3681;
  assign n3683 = ~n216 & ~n358;
  assign n3684 = n3682 & n3683;
  assign n3685 = ~n298 & ~n998;
  assign n3686 = n815 & n3685;
  assign n3687 = n3684 & n3686;
  assign n3688 = ~n381 & ~n844;
  assign n3689 = n146 & n228;
  assign n3690 = n165 & ~n3689;
  assign n3691 = ~n271 & ~n343;
  assign n3692 = ~n3690 & n3691;
  assign n3693 = n3688 & n3692;
  assign n3694 = n3687 & n3693;
  assign n3695 = n718 & n3694;
  assign n3696 = n3393 & n3695;
  assign n3802 = n3801 ^ n3696;
  assign n3808 = n3807 ^ n3802;
  assign n3809 = n3679 & ~n3808;
  assign n3810 = n3809 ^ n3678;
  assign n3945 = n3807 ^ n3801;
  assign n3946 = ~n3802 & ~n3945;
  assign n3947 = n3946 ^ n3807;
  assign n3948 = n3675 & n3947;
  assign n3949 = n3696 & n3801;
  assign n3950 = ~n3807 & n3949;
  assign n3951 = n3674 & n3950;
  assign n3952 = ~n3948 & ~n3951;
  assign n3953 = ~n3696 & ~n3801;
  assign n3954 = n3807 & n3953;
  assign n3955 = ~n3677 & n3954;
  assign n3956 = n3952 & ~n3955;
  assign n3957 = ~n3637 & ~n3947;
  assign n3958 = n3664 & ~n3950;
  assign n3959 = n3957 & ~n3958;
  assign n3960 = n3956 & ~n3959;
  assign n3926 = ~n3702 & n3761;
  assign n3927 = ~n3785 & n3798;
  assign n3928 = ~n3699 & n3927;
  assign n3929 = ~n3926 & n3928;
  assign n3930 = n3785 & ~n3798;
  assign n3931 = n3702 & ~n3761;
  assign n3932 = n3930 & ~n3931;
  assign n3933 = n3699 & n3932;
  assign n3934 = ~n3929 & ~n3933;
  assign n3935 = n3798 ^ n3699;
  assign n3936 = n3799 & ~n3935;
  assign n3937 = n3936 ^ n3699;
  assign n3938 = n3937 ^ n3761;
  assign n3939 = n3937 ^ n3702;
  assign n3940 = ~n3938 & n3939;
  assign n3941 = n3934 & n3940;
  assign n3942 = n3941 ^ n3934;
  assign n3907 = ~n3625 & ~n3627;
  assign n3908 = x1 & n3907;
  assign n3909 = x2 & n3627;
  assign n3910 = ~n3908 & ~n3909;
  assign n3911 = n3026 & ~n3910;
  assign n3912 = x2 & x22;
  assign n3913 = x1 & n3912;
  assign n3914 = ~n3625 & ~n3913;
  assign n3915 = ~n3035 & ~n3912;
  assign n3916 = ~n3914 & ~n3915;
  assign n3917 = ~x2 & ~x22;
  assign n3918 = n3031 & n3917;
  assign n3919 = ~n3916 & ~n3918;
  assign n3920 = ~n3911 & n3919;
  assign n3921 = n2434 & ~n3908;
  assign n3922 = x2 & ~n3907;
  assign n3923 = n3921 & ~n3922;
  assign n3924 = n3920 & ~n3923;
  assign n3880 = ~n3375 & ~n3378;
  assign n3881 = n2484 & n3880;
  assign n3882 = n1057 & ~n3000;
  assign n3883 = ~n1057 & n3032;
  assign n3884 = ~n969 & n2438;
  assign n3885 = n3884 ^ n2437;
  assign n3886 = ~n3883 & n3885;
  assign n3887 = ~n3882 & n3886;
  assign n3888 = n2474 & n3000;
  assign n3889 = n2442 & ~n3032;
  assign n3890 = ~n3888 & ~n3889;
  assign n3891 = ~n3887 & n3890;
  assign n3892 = ~n969 & n3891;
  assign n3893 = ~n3881 & ~n3892;
  assign n3894 = ~n2558 & ~n3893;
  assign n3895 = n2571 & n3378;
  assign n3896 = ~n3892 & ~n3895;
  assign n3897 = n1057 & n3378;
  assign n3898 = n3375 & ~n3897;
  assign n3899 = ~n3896 & n3898;
  assign n3900 = n2639 & ~n3375;
  assign n3901 = n3378 & n3900;
  assign n3902 = n969 & ~n3891;
  assign n3903 = ~n3901 & ~n3902;
  assign n3904 = ~n3899 & n3903;
  assign n3905 = ~n3894 & n3904;
  assign n3860 = n2929 ^ n310;
  assign n3861 = n2098 & n3860;
  assign n3862 = n2097 & ~n3752;
  assign n3863 = ~n3861 & ~n3862;
  assign n3864 = n756 & ~n3863;
  assign n3865 = ~n2929 & n3747;
  assign n3866 = ~n2827 & n3745;
  assign n3867 = ~n3865 & ~n3866;
  assign n3868 = ~n756 & ~n3867;
  assign n3869 = ~n310 & n2097;
  assign n3870 = n2929 & n3869;
  assign n3871 = ~n3868 & ~n3870;
  assign n3872 = ~n3864 & n3871;
  assign n3873 = ~n1898 & n3057;
  assign n3874 = n3873 ^ n310;
  assign n3875 = n3874 ^ n3034;
  assign n3876 = n1855 & n3875;
  assign n3877 = n3872 & ~n3876;
  assign n3845 = n313 & n3339;
  assign n3846 = n1698 & n2473;
  assign n3847 = n1703 & n2428;
  assign n3848 = ~n3846 & ~n3847;
  assign n3849 = ~n3845 & n3848;
  assign n3850 = ~n308 & ~n3849;
  assign n3851 = n313 & ~n3346;
  assign n3852 = n308 & n3848;
  assign n3853 = ~n3851 & n3852;
  assign n3854 = n2535 ^ n315;
  assign n3855 = n2496 & n3854;
  assign n3856 = n313 & n3855;
  assign n3857 = ~n3853 & ~n3856;
  assign n3858 = ~n3850 & n3857;
  assign n3841 = ~n1079 & n2087;
  assign n3836 = n1837 & n3715;
  assign n3837 = n3718 & ~n3836;
  assign n3838 = ~n1837 & ~n3715;
  assign n3839 = ~n1079 & ~n3838;
  assign n3840 = ~n3837 & n3839;
  assign n3842 = n3841 ^ n3840;
  assign n3829 = n2239 & n2343;
  assign n3830 = n3829 ^ n2340;
  assign n3831 = n1734 & ~n3830;
  assign n3832 = n2085 & ~n2244;
  assign n3833 = ~n2086 & n2248;
  assign n3834 = ~n3832 & ~n3833;
  assign n3835 = ~n3831 & n3834;
  assign n3843 = n3842 ^ n3835;
  assign n3826 = n3721 ^ n3708;
  assign n3827 = ~n3736 & n3826;
  assign n3828 = n3827 ^ n3735;
  assign n3844 = n3843 ^ n3828;
  assign n3859 = n3858 ^ n3844;
  assign n3878 = n3877 ^ n3859;
  assign n3823 = n3759 ^ n3705;
  assign n3824 = ~n3760 & n3823;
  assign n3825 = n3824 ^ n3705;
  assign n3879 = n3878 ^ n3825;
  assign n3906 = n3905 ^ n3879;
  assign n3925 = n3924 ^ n3906;
  assign n3943 = n3942 ^ n3925;
  assign n3811 = n1517 & n3510;
  assign n3812 = ~n129 & ~n293;
  assign n3813 = n3811 & n3812;
  assign n3814 = ~n422 & ~n589;
  assign n3815 = ~n355 & n3814;
  assign n3816 = n571 & n3815;
  assign n3817 = n3813 & n3816;
  assign n3818 = n2030 & n3817;
  assign n3819 = n638 & n3439;
  assign n3820 = n470 & n3819;
  assign n3821 = n3818 & n3820;
  assign n3822 = n876 & n3821;
  assign n3944 = n3943 ^ n3822;
  assign n3961 = n3960 ^ n3944;
  assign n3967 = n3822 & ~n3943;
  assign n3968 = n3947 & ~n3967;
  assign n3969 = ~n3822 & n3943;
  assign n3970 = n3674 & ~n3954;
  assign n3971 = ~n3969 & n3970;
  assign n3972 = n3968 & n3971;
  assign n3973 = n3944 & n3951;
  assign n3974 = ~n3972 & ~n3973;
  assign n3962 = ~n3947 & ~n3950;
  assign n3963 = ~n3944 & ~n3962;
  assign n3964 = n3664 & ~n3963;
  assign n3965 = n3944 & ~n3954;
  assign n3966 = n3964 & ~n3965;
  assign n3977 = ~n3637 & ~n3966;
  assign n3978 = n3974 & ~n3977;
  assign n3975 = n3637 & n3974;
  assign n3976 = ~n3966 & ~n3975;
  assign n3979 = n3978 ^ n3976;
  assign n4082 = ~n3968 & ~n3969;
  assign n4074 = ~n3925 & ~n3928;
  assign n4075 = ~n3926 & ~n3933;
  assign n4076 = ~n4074 & n4075;
  assign n4077 = ~n3925 & ~n3931;
  assign n4078 = ~n3937 & ~n4077;
  assign n4079 = ~n4076 & ~n4078;
  assign n4052 = n3625 & ~n3628;
  assign n4053 = n2484 & ~n4052;
  assign n4054 = n2474 & ~n3375;
  assign n4055 = ~n2442 & ~n4054;
  assign n4056 = ~n3882 & ~n4055;
  assign n4057 = n2475 & ~n3375;
  assign n4058 = ~n4056 & ~n4057;
  assign n4059 = n2438 & n3000;
  assign n4060 = n969 & ~n4059;
  assign n4061 = n4058 & n4060;
  assign n4062 = ~n4053 & n4061;
  assign n4063 = ~n3625 & ~n3628;
  assign n4064 = n2558 & n4063;
  assign n4065 = n3625 ^ n1057;
  assign n4066 = n2484 & ~n4065;
  assign n4067 = n3628 & n4066;
  assign n4068 = ~n969 & ~n4058;
  assign n4069 = ~n4067 & ~n4068;
  assign n4070 = ~n4064 & n4069;
  assign n4071 = ~n4062 & n4070;
  assign n4036 = n1855 & n3589;
  assign n4037 = n2101 & ~n3034;
  assign n4038 = n2104 & ~n2929;
  assign n4039 = ~n4037 & ~n4038;
  assign n4040 = ~n4036 & n4039;
  assign n4041 = n310 & ~n4040;
  assign n4042 = n1855 & ~n3600;
  assign n4043 = ~n310 & n4039;
  assign n4044 = ~n4042 & n4043;
  assign n4045 = n1855 & n3272;
  assign n4046 = n3032 ^ n756;
  assign n4047 = n4045 & ~n4046;
  assign n4048 = ~n4044 & ~n4047;
  assign n4049 = ~n4041 & n4048;
  assign n4019 = n2827 ^ n315;
  assign n4020 = n313 & ~n4019;
  assign n4021 = n2805 & n4020;
  assign n4022 = n1698 & n2535;
  assign n4023 = n1703 & n2473;
  assign n4024 = ~n4022 & ~n4023;
  assign n4025 = n308 & ~n4024;
  assign n4026 = ~n4021 & ~n4025;
  assign n4027 = n2258 & n2832;
  assign n4028 = n4026 & ~n4027;
  assign n4029 = n313 & ~n2836;
  assign n4030 = ~n308 & n4024;
  assign n4031 = ~n4029 & n4030;
  assign n4032 = n4028 & ~n4031;
  assign n4004 = n1734 & n2570;
  assign n4005 = ~n2244 & ~n2340;
  assign n4006 = n2085 & n2248;
  assign n4007 = ~n4005 & ~n4006;
  assign n4008 = ~n4004 & n4007;
  assign n4009 = ~n1079 & ~n4008;
  assign n4010 = n1734 & ~n2586;
  assign n4011 = n1079 & n4007;
  assign n4012 = ~n4010 & n4011;
  assign n4013 = n2428 ^ n989;
  assign n4014 = n1734 & n2569;
  assign n4015 = n4013 & n4014;
  assign n4016 = ~n4012 & ~n4015;
  assign n4017 = ~n4009 & n4016;
  assign n4018 = n4017 ^ n2436;
  assign n4033 = n4032 ^ n4018;
  assign n3998 = n3840 ^ n2087;
  assign n3999 = n3840 ^ n3835;
  assign n4000 = ~n3998 & ~n3999;
  assign n4001 = n4000 ^ n2087;
  assign n4002 = n4001 ^ n2086;
  assign n4003 = ~n1079 & n4002;
  assign n4034 = n4033 ^ n4003;
  assign n3995 = n3858 ^ n3828;
  assign n3996 = n3844 & ~n3995;
  assign n3997 = n3996 ^ n3858;
  assign n4035 = n4034 ^ n3997;
  assign n4050 = n4049 ^ n4035;
  assign n3992 = n3859 ^ n3825;
  assign n3993 = n3878 & n3992;
  assign n3994 = n3993 ^ n3877;
  assign n4051 = n4050 ^ n3994;
  assign n4072 = n4071 ^ n4051;
  assign n3989 = n3924 ^ n3905;
  assign n3990 = n3906 & ~n3989;
  assign n3991 = n3990 ^ n3924;
  assign n4073 = n4072 ^ n3991;
  assign n4080 = n4079 ^ n4073;
  assign n3980 = n564 & n721;
  assign n3981 = ~n92 & n2504;
  assign n3982 = n3980 & n3981;
  assign n3983 = n152 & ~n2809;
  assign n3984 = n840 & ~n3983;
  assign n3985 = n3982 & n3984;
  assign n3986 = n612 & n3985;
  assign n3987 = n1541 & n3986;
  assign n3988 = n517 & n3987;
  assign n4081 = n4080 ^ n3988;
  assign n4083 = n4082 ^ n4081;
  assign n4084 = n3979 & ~n4083;
  assign n4085 = n4084 ^ n3978;
  assign n4233 = n3988 & ~n4080;
  assign n4234 = n4082 & n4233;
  assign n4235 = ~n3977 & ~n4234;
  assign n4236 = ~n4082 & ~n4233;
  assign n4237 = ~n3988 & n4080;
  assign n4238 = ~n4236 & ~n4237;
  assign n4239 = ~n3975 & n4238;
  assign n4240 = ~n4235 & n4239;
  assign n4241 = ~n4082 & n4237;
  assign n4242 = ~n3977 & n4241;
  assign n4243 = n3975 & ~n4238;
  assign n4244 = ~n4242 & ~n4243;
  assign n4245 = ~n4240 & n4244;
  assign n4209 = ~n3991 & ~n4071;
  assign n4210 = n4079 & ~n4209;
  assign n4211 = ~n3994 & n4050;
  assign n4212 = n3994 & ~n4050;
  assign n4213 = n4071 & ~n4212;
  assign n4214 = n3991 & n4213;
  assign n4215 = ~n4211 & ~n4214;
  assign n4216 = n4210 & ~n4215;
  assign n4222 = ~n4071 & n4212;
  assign n4217 = n4071 ^ n4050;
  assign n4218 = n4217 ^ n3994;
  assign n4219 = n4211 & ~n4218;
  assign n4220 = n4219 ^ n4218;
  assign n4221 = ~n3991 & ~n4220;
  assign n4223 = n4222 ^ n4221;
  assign n4224 = ~n4079 & n4223;
  assign n4225 = n4071 & n4211;
  assign n4226 = n4225 ^ n4222;
  assign n4227 = n3991 & n4226;
  assign n4228 = n4227 ^ n4222;
  assign n4229 = ~n4224 & ~n4228;
  assign n4230 = ~n4216 & n4229;
  assign n4193 = ~n2440 & n2575;
  assign n4194 = n3793 & n4193;
  assign n4195 = ~n2476 & ~n3625;
  assign n4196 = n969 & ~n4195;
  assign n4197 = ~n1057 & ~n2436;
  assign n4198 = ~n3375 & n4197;
  assign n4199 = n4196 & ~n4198;
  assign n4200 = ~n2484 & ~n4199;
  assign n4201 = ~n4194 & ~n4200;
  assign n4202 = ~n3793 & ~n4196;
  assign n4203 = n4201 & ~n4202;
  assign n4204 = n2442 & ~n3375;
  assign n4205 = ~n4195 & ~n4204;
  assign n4206 = ~n969 & ~n4205;
  assign n4207 = ~n4203 & ~n4206;
  assign n4176 = n3000 & ~n3023;
  assign n4177 = n1855 & n4176;
  assign n4178 = n2101 & ~n3032;
  assign n4179 = n2104 & ~n3034;
  assign n4180 = ~n4178 & ~n4179;
  assign n4181 = ~n4177 & n4180;
  assign n4182 = ~n310 & ~n4181;
  assign n4183 = n1855 & ~n3763;
  assign n4184 = n310 & n4180;
  assign n4185 = ~n4183 & n4184;
  assign n4186 = n3000 ^ n756;
  assign n4187 = n1855 & ~n4186;
  assign n4188 = n3023 & n4187;
  assign n4189 = ~n4185 & ~n4188;
  assign n4190 = ~n4182 & n4189;
  assign n4136 = ~n1079 & ~n2086;
  assign n4165 = n4018 & n4032;
  assign n4166 = ~n4136 & n4165;
  assign n4167 = n4018 ^ n2086;
  assign n4168 = ~n4001 & ~n4167;
  assign n4169 = ~n4032 & ~n4168;
  assign n4170 = ~n2086 & ~n4018;
  assign n4171 = n4001 & ~n4170;
  assign n4172 = ~n1079 & ~n4171;
  assign n4173 = ~n4169 & n4172;
  assign n4174 = ~n4166 & ~n4173;
  assign n4142 = ~n315 & n2935;
  assign n4143 = n313 & n315;
  assign n4144 = n2929 & n4143;
  assign n4145 = n4144 ^ n313;
  assign n4146 = ~n2938 & n4145;
  assign n4147 = ~n4142 & n4146;
  assign n4148 = n1698 & n2827;
  assign n4149 = n1703 & n2535;
  assign n4150 = ~n4148 & ~n4149;
  assign n4151 = n308 & n4150;
  assign n4152 = ~n4147 & n4151;
  assign n4153 = n315 & n2902;
  assign n4154 = ~n308 & ~n2929;
  assign n4155 = n313 & n4154;
  assign n4156 = ~n4153 & n4155;
  assign n4157 = ~n308 & ~n4150;
  assign n4158 = ~n308 & n4143;
  assign n4159 = n2929 & n4158;
  assign n4160 = n2902 & n4159;
  assign n4161 = ~n4157 & ~n4160;
  assign n4162 = ~n4156 & n4161;
  assign n4163 = ~n4152 & n4162;
  assign n4126 = ~n2436 & n4017;
  assign n4127 = ~n2086 & n4126;
  assign n4128 = ~n1079 & n2085;
  assign n4129 = ~n4127 & n4128;
  assign n4130 = n2436 & ~n4017;
  assign n4131 = n2086 & n4130;
  assign n4132 = n4129 & ~n4131;
  assign n4133 = n1079 & n4130;
  assign n4134 = ~n4132 & ~n4133;
  assign n4135 = ~n2085 & n4131;
  assign n4137 = ~n2085 & n4136;
  assign n4138 = n4126 & n4137;
  assign n4139 = ~n4135 & ~n4138;
  assign n4140 = n4134 & n4139;
  assign n4105 = n1734 & ~n2544;
  assign n4106 = ~n1079 & ~n4105;
  assign n4107 = n989 & n2428;
  assign n4108 = ~n2340 & n2746;
  assign n4109 = ~n4107 & ~n4108;
  assign n4110 = n1739 & ~n4109;
  assign n4111 = ~n989 & ~n2428;
  assign n4112 = n2231 & ~n2340;
  assign n4113 = ~n2243 & ~n4112;
  assign n4114 = ~n4111 & ~n4113;
  assign n4115 = ~n4110 & ~n4114;
  assign n4116 = n4106 & n4115;
  assign n4117 = n1079 & ~n4115;
  assign n4118 = n1079 & n1734;
  assign n4119 = n2559 & n4118;
  assign n4120 = n2473 ^ n989;
  assign n4121 = n1734 & n2543;
  assign n4122 = ~n4120 & n4121;
  assign n4123 = ~n4119 & ~n4122;
  assign n4124 = ~n4117 & n4123;
  assign n4125 = ~n4116 & n4124;
  assign n4141 = n4140 ^ n4125;
  assign n4164 = n4163 ^ n4141;
  assign n4175 = n4174 ^ n4164;
  assign n4191 = n4190 ^ n4175;
  assign n4102 = n4049 ^ n4034;
  assign n4103 = n4035 & n4102;
  assign n4104 = n4103 ^ n4049;
  assign n4192 = n4191 ^ n4104;
  assign n4208 = n4207 ^ n4192;
  assign n4231 = n4230 ^ n4208;
  assign n4086 = ~n51 & n128;
  assign n4087 = ~n85 & n146;
  assign n4088 = ~n4086 & ~n4087;
  assign n4089 = ~n238 & ~n4088;
  assign n4090 = ~n164 & n219;
  assign n4091 = ~n341 & n4090;
  assign n4092 = ~n768 & ~n4091;
  assign n4093 = n4089 & ~n4092;
  assign n4094 = n1876 & n4093;
  assign n4095 = ~n286 & n360;
  assign n4096 = n226 & n3478;
  assign n4097 = n4095 & n4096;
  assign n4098 = n4094 & n4097;
  assign n4099 = n3622 & n4098;
  assign n4100 = n3520 & n4099;
  assign n4101 = n2925 & n4100;
  assign n4232 = n4231 ^ n4101;
  assign n4246 = n4245 ^ n4232;
  assign n4368 = ~n4238 & ~n4241;
  assign n4369 = n4368 ^ n4234;
  assign n4370 = n4232 & n4369;
  assign n4371 = n4370 ^ n4368;
  assign n4372 = ~n3974 & n4371;
  assign n4373 = n3637 & ~n4372;
  assign n4374 = ~n4232 & n4236;
  assign n4375 = n3966 & ~n4234;
  assign n4376 = ~n4374 & n4375;
  assign n4377 = n4232 ^ n4082;
  assign n4378 = ~n4237 & n4377;
  assign n4379 = n4378 ^ n4082;
  assign n4380 = n4376 & ~n4379;
  assign n4381 = ~n4373 & ~n4380;
  assign n4355 = n3991 & n4071;
  assign n4356 = ~n4208 & ~n4212;
  assign n4357 = ~n4355 & ~n4356;
  assign n4358 = ~n4210 & n4357;
  assign n4359 = n4208 & ~n4214;
  assign n4360 = n4079 & ~n4359;
  assign n4361 = ~n4208 & ~n4209;
  assign n4362 = ~n4211 & ~n4361;
  assign n4363 = ~n4360 & n4362;
  assign n4364 = ~n4358 & ~n4363;
  assign n4342 = ~n1057 & n3907;
  assign n4343 = n4342 ^ n3627;
  assign n4344 = ~n2440 & n4343;
  assign n4345 = n969 & n3627;
  assign n4346 = n4344 & ~n4345;
  assign n4347 = n2437 ^ n969;
  assign n4348 = n2437 ^ n1057;
  assign n4349 = ~n4347 & n4348;
  assign n4350 = ~n3625 & n4349;
  assign n4351 = n4350 ^ n969;
  assign n4352 = ~n4346 & n4351;
  assign n4339 = n4207 ^ n4191;
  assign n4340 = n4192 & n4339;
  assign n4341 = n4340 ^ n4207;
  assign n4353 = n4352 ^ n4341;
  assign n4322 = n1855 & n3880;
  assign n4323 = n2101 & n3000;
  assign n4324 = n2104 & ~n3032;
  assign n4325 = ~n4323 & ~n4324;
  assign n4326 = ~n4322 & n4325;
  assign n4327 = ~n310 & ~n4326;
  assign n4328 = n3375 & ~n3378;
  assign n4329 = n1855 & ~n4328;
  assign n4330 = n310 & n4325;
  assign n4331 = ~n4329 & n4330;
  assign n4332 = n3375 ^ n756;
  assign n4333 = n1855 & n4332;
  assign n4334 = n3378 & n4333;
  assign n4335 = ~n4331 & ~n4334;
  assign n4336 = ~n4327 & n4335;
  assign n4305 = n313 & ~n3034;
  assign n4306 = ~n3057 & n4305;
  assign n4307 = n1698 & ~n2929;
  assign n4308 = n1703 & n2827;
  assign n4309 = ~n4307 & ~n4308;
  assign n4310 = ~n4306 & n4309;
  assign n4311 = ~n308 & ~n4310;
  assign n4312 = n313 & n3057;
  assign n4314 = n308 & n4309;
  assign n4315 = ~n4305 & n4314;
  assign n4313 = n3034 ^ n315;
  assign n4316 = n4315 ^ n4313;
  assign n4317 = n4312 & ~n4316;
  assign n4318 = n4317 ^ n4315;
  assign n4319 = ~n4311 & ~n4318;
  assign n4291 = n4127 & n4128;
  assign n4292 = ~n4135 & ~n4291;
  assign n4293 = n2340 & ~n4292;
  assign n4294 = n2085 & ~n2086;
  assign n4295 = n4017 & n4294;
  assign n4296 = ~n1079 & ~n2340;
  assign n4297 = ~n4295 & n4296;
  assign n4298 = ~n4135 & n4297;
  assign n4299 = n2436 & n4128;
  assign n4300 = ~n2340 & n4299;
  assign n4301 = ~n4133 & ~n4300;
  assign n4302 = ~n4298 & n4301;
  assign n4303 = ~n4293 & n4302;
  assign n4274 = ~n1079 & n2473;
  assign n4275 = n2243 & n4274;
  assign n4276 = n2246 & n4111;
  assign n4277 = ~n1079 & ~n2428;
  assign n4278 = n2519 & ~n4277;
  assign n4279 = ~n4276 & ~n4278;
  assign n4280 = ~n4275 & n4279;
  assign n4281 = n2473 ^ n1079;
  assign n4282 = n1079 & n2230;
  assign n4283 = ~n2234 & ~n4282;
  assign n4284 = n4281 & ~n4283;
  assign n4285 = n4280 & ~n4284;
  assign n4286 = n2239 & ~n2496;
  assign n4287 = n4286 ^ n989;
  assign n4288 = n4287 ^ n2535;
  assign n4289 = n1734 & n4288;
  assign n4290 = n4285 & ~n4289;
  assign n4304 = n4303 ^ n4290;
  assign n4320 = n4319 ^ n4304;
  assign n4271 = n4163 ^ n4140;
  assign n4272 = ~n4141 & n4271;
  assign n4273 = n4272 ^ n4163;
  assign n4321 = n4320 ^ n4273;
  assign n4337 = n4336 ^ n4321;
  assign n4268 = n4190 ^ n4174;
  assign n4269 = ~n4175 & n4268;
  assign n4270 = n4269 ^ n4190;
  assign n4338 = n4337 ^ n4270;
  assign n4354 = n4353 ^ n4338;
  assign n4365 = n4364 ^ n4354;
  assign n4250 = ~n40 & ~n141;
  assign n4251 = n236 & ~n4250;
  assign n4252 = ~n196 & ~n4251;
  assign n4253 = n3510 & ~n4252;
  assign n4254 = n3515 & n4253;
  assign n4255 = n226 & ~n380;
  assign n4256 = n1523 & n4255;
  assign n4257 = n416 & n4256;
  assign n4258 = n4254 & n4257;
  assign n4259 = ~n180 & ~n577;
  assign n4260 = n1515 & n4259;
  assign n4261 = n472 & n4260;
  assign n4262 = ~n237 & ~n278;
  assign n4263 = n2958 & n4262;
  assign n4264 = n4261 & n4263;
  assign n4265 = n4258 & n4264;
  assign n4266 = n1531 & n4265;
  assign n4267 = n3476 & n4266;
  assign n4366 = n4365 ^ n4267;
  assign n4247 = n4238 ^ n4231;
  assign n4248 = n4232 & ~n4247;
  assign n4249 = n4248 ^ n4238;
  assign n4367 = n4366 ^ n4249;
  assign n4382 = n4381 ^ n4367;
  assign n4481 = n4372 & ~n4380;
  assign n4482 = n4367 & n4481;
  assign n4483 = ~n4367 & n4380;
  assign n4484 = ~n3637 & ~n4483;
  assign n4485 = ~n4482 & ~n4484;
  assign n4462 = ~n4270 & n4337;
  assign n4463 = ~n4352 & ~n4462;
  assign n4464 = n4270 & ~n4337;
  assign n4465 = ~n4463 & ~n4464;
  assign n4466 = ~n4352 & n4464;
  assign n4467 = ~n4341 & ~n4466;
  assign n4468 = ~n4465 & ~n4467;
  assign n4469 = n4364 & n4468;
  assign n4470 = n4352 & n4462;
  assign n4471 = ~n4466 & ~n4470;
  assign n4472 = n4353 & ~n4471;
  assign n4473 = ~n4469 & ~n4472;
  assign n4474 = ~n4341 & n4465;
  assign n4475 = ~n4470 & ~n4474;
  assign n4476 = ~n4364 & ~n4475;
  assign n4477 = n4473 & ~n4476;
  assign n4433 = ~n2244 & n2535;
  assign n4434 = n2248 & n2473;
  assign n4435 = ~n4433 & ~n4434;
  assign n4436 = n2239 & n2805;
  assign n4437 = n4436 ^ n2827;
  assign n4438 = n1734 & n4437;
  assign n4439 = n4435 & ~n4438;
  assign n4440 = ~n4128 & ~n4136;
  assign n4441 = ~n4296 & n4440;
  assign n4442 = ~n4017 & n4441;
  assign n4443 = n2436 & n4442;
  assign n4444 = n2428 & ~n4443;
  assign n4445 = n4439 & ~n4444;
  assign n4446 = ~n2340 & ~n2436;
  assign n4447 = n4295 & n4446;
  assign n4448 = ~n4445 & ~n4447;
  assign n4449 = ~n4277 & ~n4443;
  assign n4450 = ~n4439 & n4449;
  assign n4451 = n4448 & ~n4450;
  assign n4452 = ~n2428 & n4447;
  assign n4453 = n1079 & ~n4130;
  assign n4454 = ~n4452 & ~n4453;
  assign n4455 = n4439 & ~n4454;
  assign n4456 = ~n4451 & ~n4455;
  assign n4457 = n4456 ^ n969;
  assign n4430 = n4319 ^ n4303;
  assign n4431 = n4304 & n4430;
  assign n4432 = n4431 ^ n4319;
  assign n4458 = n4457 ^ n4432;
  assign n4413 = n313 & ~n3600;
  assign n4414 = n1698 & ~n3034;
  assign n4415 = n1703 & ~n2929;
  assign n4416 = ~n4414 & ~n4415;
  assign n4417 = ~n308 & n4416;
  assign n4418 = ~n4413 & n4417;
  assign n4419 = n308 & ~n4416;
  assign n4420 = n3032 & n3272;
  assign n4421 = n2265 & n4420;
  assign n4422 = ~n4419 & ~n4421;
  assign n4423 = ~n4418 & n4422;
  assign n4424 = n3272 & n4417;
  assign n4425 = ~n2258 & ~n4424;
  assign n4426 = ~n315 & n3272;
  assign n4427 = ~n3032 & ~n4426;
  assign n4428 = ~n4425 & n4427;
  assign n4429 = n4423 & ~n4428;
  assign n4459 = n4458 ^ n4429;
  assign n4410 = n4336 ^ n4320;
  assign n4411 = n4321 & ~n4410;
  assign n4412 = n4411 ^ n4336;
  assign n4460 = n4459 ^ n4412;
  assign n4396 = n1855 & n4063;
  assign n4397 = n2104 & n3000;
  assign n4398 = n2101 & ~n3375;
  assign n4399 = ~n4397 & ~n4398;
  assign n4400 = ~n4396 & n4399;
  assign n4401 = n310 & ~n4400;
  assign n4402 = n1855 & ~n4052;
  assign n4403 = ~n310 & n4399;
  assign n4404 = ~n4402 & n4403;
  assign n4405 = n3625 ^ n756;
  assign n4406 = n1855 & ~n4405;
  assign n4407 = n3628 & n4406;
  assign n4408 = ~n4404 & ~n4407;
  assign n4409 = ~n4401 & n4408;
  assign n4461 = n4460 ^ n4409;
  assign n4478 = n4477 ^ n4461;
  assign n4386 = ~n140 & ~n3428;
  assign n4387 = ~n91 & n397;
  assign n4388 = n457 & ~n4387;
  assign n4389 = ~n495 & ~n512;
  assign n4390 = n4388 & ~n4389;
  assign n4391 = n2973 & n4089;
  assign n4392 = n4390 & n4391;
  assign n4393 = n4258 & n4392;
  assign n4394 = ~n4386 & n4393;
  assign n4395 = n2015 & n4394;
  assign n4479 = n4478 ^ n4395;
  assign n4383 = n4365 ^ n4249;
  assign n4384 = ~n4366 & n4383;
  assign n4385 = n4384 ^ n4249;
  assign n4480 = n4479 ^ n4385;
  assign n4486 = n4485 ^ n4480;
  assign n4609 = ~n4480 & n4482;
  assign n4610 = n3637 & ~n4609;
  assign n4611 = n4480 & n4483;
  assign n4612 = ~n4610 & ~n4611;
  assign n4590 = n57 & ~n795;
  assign n4591 = n816 & ~n4590;
  assign n4592 = n78 & n2809;
  assign n4593 = n85 & ~n4592;
  assign n4594 = n4591 & ~n4593;
  assign n4595 = n1574 & n4594;
  assign n4596 = n3477 & n4595;
  assign n4597 = n836 & n1515;
  assign n4598 = n335 & n2914;
  assign n4599 = n4597 & n4598;
  assign n4600 = ~n146 & n165;
  assign n4601 = n56 & ~n97;
  assign n4602 = ~n4600 & ~n4601;
  assign n4603 = ~n1550 & n4602;
  assign n4604 = n604 & n4603;
  assign n4605 = n4599 & n4604;
  assign n4606 = n4596 & n4605;
  assign n4607 = n3420 & n4606;
  assign n4575 = ~n4461 & ~n4462;
  assign n4576 = n4364 ^ n4341;
  assign n4577 = n4353 & n4576;
  assign n4578 = n4577 ^ n4364;
  assign n4579 = ~n4575 & ~n4578;
  assign n4580 = n4341 & n4463;
  assign n4581 = n4461 & ~n4580;
  assign n4582 = n4364 & ~n4581;
  assign n4583 = ~n4341 & n4352;
  assign n4584 = ~n4461 & ~n4583;
  assign n4585 = ~n4464 & ~n4584;
  assign n4586 = ~n4582 & n4585;
  assign n4587 = ~n4579 & ~n4586;
  assign n4554 = ~n315 & n3000;
  assign n4555 = ~n4176 & ~n4554;
  assign n4556 = n313 & ~n4555;
  assign n4557 = n1698 & ~n3032;
  assign n4558 = n1703 & ~n3034;
  assign n4559 = ~n4557 & ~n4558;
  assign n4560 = ~n4556 & n4559;
  assign n4561 = ~n308 & ~n4560;
  assign n4562 = n3023 & n4554;
  assign n4563 = n313 & ~n4562;
  assign n4564 = ~n315 & n3775;
  assign n4565 = n4564 ^ n3000;
  assign n4566 = n4563 & n4565;
  assign n4567 = n308 & n4559;
  assign n4568 = ~n4566 & n4567;
  assign n4569 = n3775 & n4158;
  assign n4570 = ~n4568 & ~n4569;
  assign n4571 = ~n4561 & n4570;
  assign n4529 = n2428 & ~n2436;
  assign n4530 = n4439 & ~n4529;
  assign n4531 = n4295 & n4296;
  assign n4532 = n2436 & ~n4442;
  assign n4533 = ~n4531 & ~n4532;
  assign n4534 = n2428 & ~n4533;
  assign n4535 = ~n4530 & ~n4534;
  assign n4536 = ~n1079 & ~n4535;
  assign n4537 = n1079 & ~n4439;
  assign n4538 = ~n4531 & ~n4537;
  assign n4539 = ~n2436 & ~n4538;
  assign n4540 = ~n4536 & ~n4539;
  assign n4541 = n969 & ~n4540;
  assign n4542 = ~n4533 & n4537;
  assign n4543 = ~n4541 & ~n4542;
  assign n4544 = ~n2428 & ~n4533;
  assign n4545 = ~n4537 & ~n4544;
  assign n4546 = n2436 & ~n4545;
  assign n4547 = ~n1079 & n4529;
  assign n4548 = n4533 & ~n4547;
  assign n4549 = n4439 & ~n4548;
  assign n4550 = ~n4546 & ~n4549;
  assign n4551 = ~n969 & ~n4550;
  assign n4552 = n4543 & ~n4551;
  assign n4513 = n1734 & ~n2929;
  assign n4514 = ~n2902 & n4513;
  assign n4515 = ~n2244 & n2827;
  assign n4516 = n2248 & n2535;
  assign n4517 = ~n4515 & ~n4516;
  assign n4518 = ~n4514 & n4517;
  assign n4519 = ~n1079 & ~n4518;
  assign n4520 = n2929 ^ n989;
  assign n4521 = n1734 & ~n4520;
  assign n4522 = n2902 & n4521;
  assign n4523 = ~n4519 & ~n4522;
  assign n4524 = n1734 & ~n2938;
  assign n4525 = n1079 & n4517;
  assign n4526 = ~n4524 & n4525;
  assign n4527 = n4523 & ~n4526;
  assign n4507 = n969 & n2436;
  assign n4508 = n2428 & ~n4507;
  assign n4509 = ~n1079 & n4508;
  assign n4510 = ~n969 & ~n2436;
  assign n4511 = ~n4509 & ~n4510;
  assign n4512 = n4511 ^ n4274;
  assign n4528 = n4527 ^ n4512;
  assign n4553 = n4552 ^ n4528;
  assign n4572 = n4571 ^ n4553;
  assign n4504 = n4459 ^ n4409;
  assign n4505 = n4460 & n4504;
  assign n4506 = n4505 ^ n4412;
  assign n4573 = n4572 ^ n4506;
  assign n4493 = n1855 & n3793;
  assign n4494 = n756 & n4493;
  assign n4495 = n2101 & ~n3625;
  assign n4496 = n2104 & ~n3375;
  assign n4497 = ~n4495 & ~n4496;
  assign n4498 = n310 & ~n4497;
  assign n4499 = ~n4494 & ~n4498;
  assign n4500 = ~n310 & n4497;
  assign n4501 = ~n4493 & n4500;
  assign n4502 = n4499 & ~n4501;
  assign n4490 = n4457 ^ n4429;
  assign n4491 = ~n4458 & ~n4490;
  assign n4492 = n4491 ^ n4432;
  assign n4503 = n4502 ^ n4492;
  assign n4574 = n4573 ^ n4503;
  assign n4588 = n4587 ^ n4574;
  assign n4487 = n4478 ^ n4385;
  assign n4488 = n4479 & ~n4487;
  assign n4489 = n4488 ^ n4385;
  assign n4589 = n4588 ^ n4489;
  assign n4608 = n4607 ^ n4589;
  assign n4613 = n4612 ^ n4608;
  assign n4693 = ~n4607 & n4610;
  assign n4694 = ~n3637 & ~n4611;
  assign n4695 = ~n4588 & ~n4694;
  assign n4696 = ~n4693 & ~n4695;
  assign n4697 = n4607 & ~n4610;
  assign n4698 = ~n4489 & ~n4697;
  assign n4699 = ~n4696 & n4698;
  assign n4700 = ~n4588 & ~n4607;
  assign n4701 = n4610 & n4700;
  assign n4702 = n4588 & n4607;
  assign n4703 = n4694 & n4702;
  assign n4704 = ~n4701 & ~n4703;
  assign n4705 = ~n4699 & n4704;
  assign n4706 = ~n4610 & n4702;
  assign n4707 = n4694 & ~n4700;
  assign n4708 = ~n4706 & ~n4707;
  assign n4709 = n4489 & ~n4708;
  assign n4710 = n4705 & ~n4709;
  assign n4674 = n4506 & ~n4572;
  assign n4675 = ~n4492 & n4502;
  assign n4681 = n4674 & ~n4675;
  assign n4677 = ~n4506 & n4572;
  assign n4678 = n4492 & ~n4502;
  assign n4682 = ~n4677 & n4678;
  assign n4683 = ~n4681 & ~n4682;
  assign n4676 = ~n4674 & n4675;
  assign n4679 = n4677 & ~n4678;
  assign n4680 = ~n4676 & ~n4679;
  assign n4684 = n4683 ^ n4680;
  assign n4685 = ~n4587 & n4684;
  assign n4686 = n4685 ^ n4683;
  assign n4687 = n4572 ^ n4502;
  assign n4688 = n4503 & ~n4687;
  assign n4689 = n4573 & n4688;
  assign n4690 = n4686 & ~n4689;
  assign n4657 = n313 & n3880;
  assign n4658 = n1698 & n3000;
  assign n4659 = n1703 & ~n3032;
  assign n4660 = ~n4658 & ~n4659;
  assign n4661 = ~n4657 & n4660;
  assign n4662 = ~n308 & ~n4661;
  assign n4663 = n313 & ~n4328;
  assign n4664 = n308 & n4660;
  assign n4665 = ~n4663 & n4664;
  assign n4666 = n3375 ^ n315;
  assign n4667 = n313 & ~n4666;
  assign n4668 = n3378 & n4667;
  assign n4669 = ~n4665 & ~n4668;
  assign n4670 = ~n4662 & n4669;
  assign n4653 = n4527 ^ n4274;
  assign n4654 = n4527 ^ n4511;
  assign n4655 = ~n4653 & n4654;
  assign n4656 = n4655 ^ n4274;
  assign n4671 = n4670 ^ n4656;
  assign n4639 = n2741 & n2827;
  assign n4640 = n2230 & ~n4639;
  assign n4641 = n2234 & ~n2929;
  assign n4642 = n4641 ^ n1739;
  assign n4643 = ~n4640 & ~n4642;
  assign n4644 = n2827 & n3543;
  assign n4645 = ~n4154 & ~n4644;
  assign n4646 = ~n989 & ~n4645;
  assign n4647 = ~n4643 & ~n4646;
  assign n4648 = n2239 & n3057;
  assign n4649 = n4648 ^ n3034;
  assign n4650 = n1734 & n4649;
  assign n4651 = ~n4647 & ~n4650;
  assign n4638 = ~n1079 & ~n2804;
  assign n4652 = n4651 ^ n4638;
  assign n4672 = n4671 ^ n4652;
  assign n4626 = n756 & n3907;
  assign n4627 = n4626 ^ n3627;
  assign n4628 = ~n2098 & n4627;
  assign n4629 = n310 & n3627;
  assign n4630 = n4628 & ~n4629;
  assign n4631 = n2097 ^ n310;
  assign n4632 = n2097 ^ n756;
  assign n4633 = ~n4631 & ~n4632;
  assign n4634 = ~n3625 & n4633;
  assign n4635 = n4634 ^ n310;
  assign n4636 = ~n4630 & n4635;
  assign n4623 = n4571 ^ n4552;
  assign n4624 = n4553 & n4623;
  assign n4625 = n4624 ^ n4571;
  assign n4637 = n4636 ^ n4625;
  assign n4673 = n4672 ^ n4637;
  assign n4691 = n4690 ^ n4673;
  assign n4614 = ~n595 & n1860;
  assign n4615 = ~n281 & ~n374;
  assign n4616 = n720 & n4615;
  assign n4617 = n4614 & n4616;
  assign n4618 = n3506 & n4617;
  assign n4619 = n459 & n4263;
  assign n4620 = n4618 & n4619;
  assign n4621 = n3483 & n4620;
  assign n4622 = n437 & n4621;
  assign n4692 = n4691 ^ n4622;
  assign n4711 = n4710 ^ n4692;
  assign n4793 = n4607 ^ n4588;
  assign n4794 = n4489 & ~n4793;
  assign n4795 = n4611 & ~n4794;
  assign n4796 = n4692 & ~n4700;
  assign n4797 = n4795 & ~n4796;
  assign n4786 = ~n4489 & ~n4702;
  assign n4798 = ~n4692 & n4786;
  assign n4799 = n4797 & ~n4798;
  assign n4800 = ~n3637 & ~n4799;
  assign n4801 = n4692 & ~n4702;
  assign n4802 = n4609 & ~n4801;
  assign n4803 = ~n4692 & ~n4700;
  assign n4804 = n4803 ^ n4793;
  assign n4805 = ~n4489 & ~n4804;
  assign n4806 = n4805 ^ n4803;
  assign n4807 = n4802 & ~n4806;
  assign n4808 = ~n4800 & ~n4807;
  assign n4787 = ~n4622 & n4691;
  assign n4788 = ~n4700 & ~n4787;
  assign n4789 = ~n4786 & n4788;
  assign n4790 = n4622 & ~n4691;
  assign n4791 = ~n4789 & ~n4790;
  assign n4774 = ~n4673 & ~n4675;
  assign n4775 = ~n4681 & ~n4774;
  assign n4776 = ~n4673 & ~n4677;
  assign n4777 = ~n4682 & ~n4776;
  assign n4778 = n4775 & n4777;
  assign n4779 = n4587 & ~n4778;
  assign n4780 = n4678 & ~n4775;
  assign n4781 = ~n4676 & n4776;
  assign n4782 = ~n4780 & ~n4781;
  assign n4783 = ~n4779 & n4782;
  assign n4758 = n313 & ~n4052;
  assign n4759 = n1703 & n3000;
  assign n4760 = n1698 & ~n3375;
  assign n4761 = ~n4759 & ~n4760;
  assign n4762 = ~n308 & n4761;
  assign n4763 = ~n4758 & n4762;
  assign n4764 = n2258 & n4063;
  assign n4765 = n3625 ^ n315;
  assign n4766 = n313 & n4765;
  assign n4767 = n3628 & n4766;
  assign n4768 = n308 & ~n4761;
  assign n4769 = ~n4767 & ~n4768;
  assign n4770 = ~n4764 & n4769;
  assign n4771 = ~n4763 & n4770;
  assign n4755 = n4672 ^ n4636;
  assign n4756 = n4637 & ~n4755;
  assign n4757 = n4756 ^ n4672;
  assign n4772 = n4771 ^ n4757;
  assign n4749 = n2827 ^ n2473;
  assign n4750 = ~n1079 & n4749;
  assign n4751 = n4750 ^ n310;
  assign n4743 = n4651 ^ n1079;
  assign n4744 = n4743 ^ n2535;
  assign n4745 = n4651 ^ n2473;
  assign n4746 = n2804 & n4745;
  assign n4747 = ~n4744 & n4746;
  assign n4748 = n4747 ^ n4743;
  assign n4752 = n4751 ^ n4748;
  assign n4723 = n3034 ^ n1079;
  assign n4724 = n2230 & n4723;
  assign n4725 = n2246 & n2929;
  assign n4726 = n4725 ^ n1739;
  assign n4727 = ~n4724 & ~n4726;
  assign n4728 = ~n989 & ~n4727;
  assign n4729 = n2246 & ~n3034;
  assign n4730 = ~n1079 & n2929;
  assign n4731 = n2230 & n4730;
  assign n4732 = ~n4729 & ~n4731;
  assign n4733 = n989 & ~n4732;
  assign n4734 = ~n1079 & n1739;
  assign n4735 = n3034 & n4734;
  assign n4736 = ~n4733 & ~n4735;
  assign n4737 = ~n4728 & n4736;
  assign n4738 = n2239 & ~n3272;
  assign n4739 = n4738 ^ n989;
  assign n4740 = n4739 ^ n3032;
  assign n4741 = n1734 & n4740;
  assign n4742 = n4737 & ~n4741;
  assign n4753 = n4752 ^ n4742;
  assign n4720 = n4656 ^ n4652;
  assign n4721 = n4671 & ~n4720;
  assign n4722 = n4721 ^ n4670;
  assign n4754 = n4753 ^ n4722;
  assign n4773 = n4772 ^ n4754;
  assign n4784 = n4783 ^ n4773;
  assign n4712 = n83 & ~n251;
  assign n4713 = n275 & ~n4712;
  assign n4714 = ~n503 & ~n1552;
  assign n4715 = n4713 & n4714;
  assign n4716 = n3517 & n4715;
  assign n4717 = n853 & n4716;
  assign n4718 = n939 & n3440;
  assign n4719 = n4717 & n4718;
  assign n4785 = n4784 ^ n4719;
  assign n4792 = n4791 ^ n4785;
  assign n4809 = n4808 ^ n4792;
  assign n4879 = n4792 & n4799;
  assign n4880 = ~n3637 & ~n4879;
  assign n4881 = ~n4792 & n4807;
  assign n4882 = ~n4880 & ~n4881;
  assign n4859 = n4771 ^ n4722;
  assign n4860 = ~n4754 & ~n4859;
  assign n4861 = n4860 ^ n4771;
  assign n4862 = ~n4757 & n4861;
  assign n4863 = ~n4722 & ~n4753;
  assign n4864 = n4771 & n4863;
  assign n4865 = ~n4862 & ~n4864;
  assign n4866 = n4783 & ~n4865;
  assign n4867 = n4722 & n4753;
  assign n4868 = ~n4771 & n4867;
  assign n4869 = ~n4864 & ~n4868;
  assign n4870 = n4772 & ~n4869;
  assign n4871 = ~n4866 & ~n4870;
  assign n4872 = ~n4757 & ~n4868;
  assign n4873 = ~n4861 & ~n4872;
  assign n4874 = ~n4783 & n4873;
  assign n4875 = n4871 & ~n4874;
  assign n4842 = n1734 & ~n3763;
  assign n4843 = ~n2244 & ~n3032;
  assign n4844 = n2248 & ~n3034;
  assign n4845 = ~n4843 & ~n4844;
  assign n4846 = ~n1079 & n4845;
  assign n4847 = ~n4842 & n4846;
  assign n4848 = n4118 & n4176;
  assign n4849 = n3000 ^ n989;
  assign n4850 = n1734 & ~n4849;
  assign n4851 = n3023 & n4850;
  assign n4852 = n1079 & ~n4845;
  assign n4853 = ~n4851 & ~n4852;
  assign n4854 = ~n4848 & n4853;
  assign n4855 = ~n4847 & n4854;
  assign n4835 = n2473 ^ n310;
  assign n4836 = ~n4749 & ~n4835;
  assign n4837 = n4836 ^ n310;
  assign n4838 = n2929 & n4837;
  assign n4839 = ~n1079 & ~n4838;
  assign n4840 = ~n2929 & ~n4837;
  assign n4841 = n4839 & ~n4840;
  assign n4856 = n4855 ^ n4841;
  assign n4832 = n4751 ^ n4742;
  assign n4833 = n4752 & ~n4832;
  assign n4834 = n4833 ^ n4748;
  assign n4857 = n4856 ^ n4834;
  assign n4822 = n313 & n3793;
  assign n4823 = n1698 & ~n3625;
  assign n4824 = n1703 & ~n3375;
  assign n4825 = ~n4823 & ~n4824;
  assign n4826 = n308 & n4825;
  assign n4827 = ~n4822 & n4826;
  assign n4828 = n3793 & n4143;
  assign n4829 = ~n308 & ~n4825;
  assign n4830 = ~n4828 & ~n4829;
  assign n4831 = ~n4827 & n4830;
  assign n4858 = n4857 ^ n4831;
  assign n4876 = n4875 ^ n4858;
  assign n4813 = n544 & n3369;
  assign n4814 = n51 & ~n149;
  assign n4815 = n56 & ~n236;
  assign n4816 = ~n4814 & ~n4815;
  assign n4817 = ~n797 & n4816;
  assign n4818 = n564 & n610;
  assign n4819 = n4817 & n4818;
  assign n4820 = n4813 & n4819;
  assign n4821 = n835 & n4820;
  assign n4877 = n4876 ^ n4821;
  assign n4810 = n4791 ^ n4784;
  assign n4811 = ~n4785 & ~n4810;
  assign n4812 = n4811 ^ n4791;
  assign n4878 = n4877 ^ n4812;
  assign n4883 = n4882 ^ n4878;
  assign n4970 = ~n4878 & n4879;
  assign n4971 = ~n3637 & ~n4970;
  assign n4972 = n4878 & n4881;
  assign n4973 = ~n4971 & ~n4972;
  assign n4956 = ~n538 & ~n826;
  assign n4957 = ~n293 & ~n413;
  assign n4958 = ~n539 & n4957;
  assign n4959 = ~n4956 & n4958;
  assign n4960 = n164 & ~n219;
  assign n4961 = ~n441 & ~n4960;
  assign n4962 = n1763 & n4961;
  assign n4963 = n571 & n4962;
  assign n4964 = n3693 & n4963;
  assign n4965 = n2296 & n4964;
  assign n4966 = n1759 & n4965;
  assign n4967 = n4959 & n4966;
  assign n4927 = n4840 & ~n4855;
  assign n4928 = ~n3034 & ~n4927;
  assign n4929 = n4837 & n4855;
  assign n4930 = n4730 & n4929;
  assign n4931 = n4928 & ~n4930;
  assign n4932 = n4839 & ~n4927;
  assign n4933 = n2929 & ~n4855;
  assign n4934 = n3034 & ~n4933;
  assign n4935 = ~n4932 & n4934;
  assign n4936 = ~n4931 & ~n4935;
  assign n4937 = n1079 & ~n4855;
  assign n4938 = ~n4936 & ~n4937;
  assign n4939 = n4856 ^ n4831;
  assign n4940 = ~n4857 & n4939;
  assign n4941 = n4940 ^ n4834;
  assign n4942 = ~n4938 & n4941;
  assign n4943 = ~n1079 & ~n4840;
  assign n4944 = ~n4929 & n4943;
  assign n4945 = ~n4730 & n4855;
  assign n4946 = ~n3034 & ~n4945;
  assign n4947 = ~n4944 & n4946;
  assign n4948 = ~n1079 & n4927;
  assign n4949 = ~n4839 & n4855;
  assign n4950 = n3034 & ~n4949;
  assign n4951 = ~n4948 & n4950;
  assign n4952 = ~n4947 & ~n4951;
  assign n4953 = ~n4941 & n4952;
  assign n4954 = ~n4942 & ~n4953;
  assign n4913 = ~n4757 & n4771;
  assign n4914 = ~n4783 & ~n4913;
  assign n4915 = n4757 & ~n4771;
  assign n4916 = ~n4858 & ~n4863;
  assign n4917 = ~n4915 & ~n4916;
  assign n4918 = ~n4914 & n4917;
  assign n4919 = ~n4863 & n4915;
  assign n4920 = n4858 & ~n4919;
  assign n4921 = ~n4783 & ~n4920;
  assign n4922 = ~n4858 & ~n4913;
  assign n4923 = ~n4867 & ~n4922;
  assign n4924 = ~n4921 & n4923;
  assign n4925 = ~n4918 & ~n4924;
  assign n4898 = n1734 & ~n4328;
  assign n4899 = ~n2244 & n3000;
  assign n4900 = n2248 & ~n3032;
  assign n4901 = ~n4899 & ~n4900;
  assign n4902 = ~n1079 & n4901;
  assign n4903 = ~n4898 & n4902;
  assign n4904 = n3880 & n4118;
  assign n4905 = n3375 ^ n989;
  assign n4906 = n1734 & n4905;
  assign n4907 = n3378 & n4906;
  assign n4908 = n1079 & ~n4901;
  assign n4909 = ~n4907 & ~n4908;
  assign n4910 = ~n4904 & n4909;
  assign n4911 = ~n4903 & n4910;
  assign n4887 = ~n315 & n3907;
  assign n4888 = n4887 ^ n3627;
  assign n4889 = ~n1723 & n4888;
  assign n4890 = n308 & n3627;
  assign n4891 = n4889 & ~n4890;
  assign n4892 = n1728 ^ n315;
  assign n4893 = n1728 ^ n308;
  assign n4894 = n4892 & ~n4893;
  assign n4895 = ~n3625 & n4894;
  assign n4896 = n4895 ^ n308;
  assign n4897 = ~n4891 & n4896;
  assign n4912 = n4911 ^ n4897;
  assign n4926 = n4925 ^ n4912;
  assign n4955 = n4954 ^ n4926;
  assign n4968 = n4967 ^ n4955;
  assign n4884 = n4876 ^ n4812;
  assign n4885 = n4877 & n4884;
  assign n4886 = n4885 ^ n4812;
  assign n4969 = n4968 ^ n4886;
  assign n4974 = n4973 ^ n4969;
  assign n5062 = ~n4969 & n4970;
  assign n5063 = ~n3637 & ~n5062;
  assign n5064 = n4969 & n4972;
  assign n5065 = ~n5063 & ~n5064;
  assign n4994 = ~n4925 & ~n4942;
  assign n4995 = ~n4953 & n4994;
  assign n5028 = ~n1079 & n4928;
  assign n5029 = ~n4949 & ~n5028;
  assign n5001 = n3625 ^ n989;
  assign n5002 = n3628 & n5001;
  assign n5003 = ~n4052 & ~n5002;
  assign n5004 = n2519 & n3000;
  assign n5005 = ~n2244 & ~n3375;
  assign n5006 = ~n1079 & ~n5005;
  assign n5007 = ~n5004 & n5006;
  assign n5008 = ~n5003 & n5007;
  assign n5009 = n1079 & ~n3000;
  assign n5010 = n1739 & ~n5009;
  assign n5011 = n3375 ^ n1079;
  assign n5012 = n2230 & n5011;
  assign n5013 = ~n989 & ~n5012;
  assign n5014 = ~n5010 & n5013;
  assign n5015 = n2231 & ~n3000;
  assign n5016 = n2246 & ~n3375;
  assign n5017 = n989 & ~n5016;
  assign n5018 = ~n5015 & n5017;
  assign n5019 = ~n5014 & ~n5018;
  assign n5020 = ~n1079 & n3375;
  assign n5021 = n1739 & n5020;
  assign n5022 = ~n5019 & ~n5021;
  assign n5023 = ~n5008 & n5022;
  assign n5024 = ~n4063 & ~n5002;
  assign n5025 = n4118 & ~n5024;
  assign n5026 = n5023 & ~n5025;
  assign n4996 = ~n3032 & ~n3034;
  assign n4997 = n2966 & n3034;
  assign n4998 = ~n1079 & ~n4997;
  assign n4999 = ~n4996 & n4998;
  assign n5000 = n4999 ^ n308;
  assign n5027 = n5026 ^ n5000;
  assign n5030 = n5029 ^ n5027;
  assign n5031 = ~n4953 & ~n5030;
  assign n5032 = n4925 & ~n5031;
  assign n5033 = ~n4995 & ~n5032;
  assign n5034 = ~n4942 & n5030;
  assign n5035 = n4897 & ~n4911;
  assign n5036 = ~n5034 & ~n5035;
  assign n5037 = ~n5033 & n5036;
  assign n5038 = ~n4925 & ~n5030;
  assign n5039 = ~n4953 & n5030;
  assign n5040 = ~n4897 & n4911;
  assign n5041 = n5039 & ~n5040;
  assign n5042 = n5030 ^ n4953;
  assign n5043 = n5035 ^ n5030;
  assign n5044 = ~n5042 & ~n5043;
  assign n5045 = n5044 ^ n4953;
  assign n5046 = ~n5041 & ~n5045;
  assign n5047 = ~n5038 & n5046;
  assign n5048 = ~n4995 & n5047;
  assign n5049 = n4994 & ~n5030;
  assign n5050 = n5040 & n5049;
  assign n5051 = ~n5048 & ~n5050;
  assign n5052 = ~n5037 & n5051;
  assign n5053 = n4994 & n5035;
  assign n5054 = n4925 & ~n4954;
  assign n5055 = ~n5039 & ~n5040;
  assign n5056 = ~n5054 & n5055;
  assign n5057 = ~n5053 & ~n5056;
  assign n5058 = ~n5049 & ~n5057;
  assign n5059 = n5052 & ~n5058;
  assign n4978 = n942 & n3427;
  assign n4979 = ~n340 & ~n563;
  assign n4980 = ~n92 & ~n326;
  assign n4981 = n4979 & n4980;
  assign n4982 = n4978 & n4981;
  assign n4983 = ~n190 & ~n361;
  assign n4984 = n130 & ~n776;
  assign n4985 = ~n585 & ~n4984;
  assign n4986 = ~n4983 & n4985;
  assign n4987 = ~n380 & ~n485;
  assign n4988 = ~n2960 & n4987;
  assign n4989 = n4986 & n4988;
  assign n4990 = n4982 & n4989;
  assign n4991 = n209 & n4990;
  assign n4992 = n3392 & n4991;
  assign n4993 = n3520 & n4992;
  assign n5060 = n5059 ^ n4993;
  assign n4975 = n4955 ^ n4886;
  assign n4976 = n4968 & n4975;
  assign n4977 = n4976 ^ n4886;
  assign n5061 = n5060 ^ n4977;
  assign n5066 = n5065 ^ n5061;
  assign n5115 = n5061 & n5062;
  assign n5116 = ~n3637 & ~n5115;
  assign n5117 = ~n5061 & n5064;
  assign n5118 = ~n5116 & ~n5117;
  assign n5103 = ~n5034 & n5040;
  assign n5104 = ~n5031 & ~n5103;
  assign n5105 = ~n4925 & n5104;
  assign n5106 = n5034 & ~n5040;
  assign n5107 = n5042 & ~n5043;
  assign n5108 = n5107 ^ n4953;
  assign n5109 = ~n5106 & ~n5108;
  assign n5110 = ~n5105 & n5109;
  assign n5111 = ~n5053 & n5110;
  assign n5089 = n2239 & n3793;
  assign n5090 = n1734 & ~n5089;
  assign n5091 = n989 & ~n3625;
  assign n5092 = n2746 & ~n3375;
  assign n5093 = n1739 & ~n5092;
  assign n5094 = ~n5091 & n5093;
  assign n5095 = n2243 & n3625;
  assign n5096 = ~n1079 & ~n3375;
  assign n5097 = n2519 & ~n5096;
  assign n5098 = ~n5095 & ~n5097;
  assign n5099 = ~n5094 & n5098;
  assign n5100 = ~n5090 & n5099;
  assign n5085 = ~n308 & ~n4997;
  assign n5086 = ~n4996 & ~n5085;
  assign n5087 = n5086 ^ n3000;
  assign n5088 = ~n1079 & n5087;
  assign n5101 = n5100 ^ n5088;
  assign n5082 = n5029 ^ n5026;
  assign n5083 = ~n5027 & ~n5082;
  assign n5084 = n5083 ^ n5029;
  assign n5102 = n5101 ^ n5084;
  assign n5112 = n5111 ^ n5102;
  assign n5070 = ~n453 & ~n728;
  assign n5071 = n1763 & n5070;
  assign n5072 = n83 & ~n4592;
  assign n5073 = n5071 & ~n5072;
  assign n5074 = ~n225 & ~n2277;
  assign n5075 = n332 & n5074;
  assign n5076 = n2958 & n5075;
  assign n5077 = n5073 & n5076;
  assign n5078 = n347 & n5077;
  assign n5079 = n883 & n5078;
  assign n5080 = n1584 & n2376;
  assign n5081 = n5079 & n5080;
  assign n5113 = n5112 ^ n5081;
  assign n5067 = n5059 ^ n4977;
  assign n5068 = ~n5060 & ~n5067;
  assign n5069 = n5068 ^ n4977;
  assign n5114 = n5113 ^ n5069;
  assign n5119 = n5118 ^ n5114;
  assign n5186 = n5114 & n5117;
  assign n5187 = n3637 & ~n5186;
  assign n5188 = ~n5114 & n5115;
  assign n5189 = ~n5187 & ~n5188;
  assign n5171 = ~n237 & n576;
  assign n5172 = n1009 & n5171;
  assign n5173 = ~n195 & ~n200;
  assign n5174 = n5074 & n5173;
  assign n5175 = n57 & ~n639;
  assign n5176 = ~n595 & ~n5175;
  assign n5177 = ~n405 & n5176;
  assign n5178 = n5174 & n5177;
  assign n5179 = n3400 & n5178;
  assign n5180 = n918 & n5179;
  assign n5181 = n1771 & n5180;
  assign n5182 = n5172 & n5181;
  assign n5183 = n4959 & n5182;
  assign n5123 = n5111 ^ n5084;
  assign n5124 = n5102 & ~n5123;
  assign n5125 = n5124 ^ n5111;
  assign n5132 = n1734 & n3627;
  assign n5133 = n2239 & n2244;
  assign n5134 = ~n3625 & n5133;
  assign n5135 = ~n5132 & n5134;
  assign n5126 = n1079 & n5100;
  assign n5128 = n3000 & n5086;
  assign n5129 = ~n1079 & ~n5128;
  assign n5127 = n5088 & n5100;
  assign n5130 = n5129 ^ n5127;
  assign n5131 = ~n5126 & ~n5130;
  assign n5152 = ~n1079 & ~n3000;
  assign n5153 = ~n5096 & ~n5152;
  assign n5154 = ~n5131 & n5153;
  assign n5139 = n3000 & n5096;
  assign n5155 = ~n5130 & n5139;
  assign n5156 = ~n5154 & ~n5155;
  assign n5157 = ~n5135 & ~n5156;
  assign n5140 = n5130 & n5139;
  assign n5136 = ~n3000 & n3375;
  assign n5158 = n1079 & ~n5100;
  assign n5159 = ~n5136 & ~n5158;
  assign n5160 = ~n5140 & n5159;
  assign n5161 = n5135 & ~n5160;
  assign n5141 = n5086 & n5100;
  assign n5162 = ~n1079 & n5141;
  assign n5142 = ~n3000 & ~n5135;
  assign n5163 = ~n3375 & n5142;
  assign n5164 = ~n5158 & n5163;
  assign n5165 = ~n5162 & n5164;
  assign n5166 = ~n5161 & ~n5165;
  assign n5167 = ~n5157 & n5166;
  assign n5137 = n5135 & ~n5136;
  assign n5138 = ~n5131 & n5137;
  assign n5143 = n5020 & n5142;
  assign n5144 = ~n5141 & n5143;
  assign n5145 = ~n5140 & ~n5144;
  assign n5146 = ~n5138 & n5145;
  assign n5147 = n3375 ^ n3000;
  assign n5148 = ~n1079 & n5147;
  assign n5149 = ~n5135 & ~n5148;
  assign n5150 = n5131 & n5149;
  assign n5151 = n5146 & ~n5150;
  assign n5168 = n5167 ^ n5151;
  assign n5169 = ~n5125 & n5168;
  assign n5170 = n5169 ^ n5167;
  assign n5184 = n5183 ^ n5170;
  assign n5120 = n5112 ^ n5069;
  assign n5121 = n5113 & n5120;
  assign n5122 = n5121 ^ n5069;
  assign n5185 = n5184 ^ n5122;
  assign n5190 = n5189 ^ n5185;
  assign n5223 = ~n5185 & n5188;
  assign n5224 = ~n3637 & ~n5223;
  assign n5225 = n5185 & n5186;
  assign n5226 = ~n5224 & ~n5225;
  assign n5212 = n3375 & n5135;
  assign n5213 = ~n5131 & n5212;
  assign n5214 = n5148 & ~n5213;
  assign n5215 = ~n5131 & ~n5137;
  assign n5216 = ~n5214 & n5215;
  assign n5217 = n5125 & ~n5216;
  assign n5218 = n5131 & ~n5149;
  assign n5219 = ~n5217 & ~n5218;
  assign n5205 = n1079 & ~n5135;
  assign n5206 = n989 & n3375;
  assign n5207 = n5015 & n5206;
  assign n5208 = n3000 & ~n5020;
  assign n5209 = n3625 & ~n5208;
  assign n5210 = ~n5207 & ~n5209;
  assign n5211 = ~n5205 & n5210;
  assign n5220 = n5219 ^ n5211;
  assign n5194 = ~n57 & n2297;
  assign n5195 = ~n318 & ~n5194;
  assign n5196 = ~n471 & ~n2277;
  assign n5197 = ~n687 & n5196;
  assign n5198 = n3391 & n5197;
  assign n5199 = n2914 & n5198;
  assign n5200 = n3465 & n5199;
  assign n5201 = n4981 & n5200;
  assign n5202 = n3405 & n5201;
  assign n5203 = n556 & n5202;
  assign n5204 = ~n5195 & n5203;
  assign n5221 = n5220 ^ n5204;
  assign n5191 = n5170 ^ n5122;
  assign n5192 = n5184 & n5191;
  assign n5193 = n5192 ^ n5122;
  assign n5222 = n5221 ^ n5193;
  assign n5227 = n5226 ^ n5222;
  assign n5243 = ~n5222 & n5225;
  assign n5244 = n3637 & ~n5243;
  assign n5245 = n5222 & n5223;
  assign n5246 = ~n5244 & ~n5245;
  assign n5231 = n490 & n2455;
  assign n5232 = n4987 & n5231;
  assign n5233 = ~n224 & ~n505;
  assign n5234 = n2511 & n5233;
  assign n5235 = ~n111 & n379;
  assign n5236 = ~n826 & ~n5235;
  assign n5237 = n551 & ~n5236;
  assign n5238 = n5234 & n5237;
  assign n5239 = n5232 & n5238;
  assign n5240 = n698 & n5239;
  assign n5241 = n2925 & n5240;
  assign n5228 = n5220 ^ n5193;
  assign n5229 = ~n5221 & ~n5228;
  assign n5230 = n5229 ^ n5193;
  assign n5242 = n5241 ^ n5230;
  assign n5247 = n5246 ^ n5242;
  assign n5257 = n5245 ^ n5230;
  assign n5258 = n5242 & n5257;
  assign n5259 = n5258 ^ n5245;
  assign n5260 = ~n3637 & ~n5259;
  assign n5261 = ~n5230 & n5241;
  assign n5262 = n5243 & n5261;
  assign n5263 = n5230 & ~n5241;
  assign n5264 = n5244 & n5263;
  assign n5265 = ~n5262 & ~n5264;
  assign n5266 = ~n5260 & n5265;
  assign n5248 = n194 & n588;
  assign n5249 = ~n618 & n815;
  assign n5250 = n3463 & n3812;
  assign n5251 = n5249 & n5250;
  assign n5252 = n1013 & n5251;
  assign n5253 = n5248 & n5252;
  assign n5254 = n391 & n5253;
  assign n5255 = n910 & n5254;
  assign n5256 = n3417 & n5255;
  assign n5267 = n5266 ^ n5256;
  assign n5279 = ~n5256 & ~n5263;
  assign n5280 = n5243 & ~n5279;
  assign n5281 = ~n5242 & n5245;
  assign n5282 = ~n5280 & ~n5281;
  assign n5283 = n5256 & ~n5262;
  assign n5284 = ~n5282 & ~n5283;
  assign n5285 = n3637 & ~n5284;
  assign n5277 = ~n5256 & n5259;
  assign n5268 = n130 & ~n2917;
  assign n5269 = n420 & ~n5268;
  assign n5270 = n148 & n165;
  assign n5271 = ~n299 & ~n5270;
  assign n5272 = n5269 & n5271;
  assign n5273 = n4089 & n5272;
  assign n5274 = n2812 & n5273;
  assign n5275 = n536 & n5274;
  assign n5276 = n5172 & n5275;
  assign n5278 = n5277 ^ n5276;
  assign n5286 = n5285 ^ n5278;
  assign n5297 = ~n5276 & n5277;
  assign n5298 = n5285 & n5297;
  assign n5299 = n5276 & ~n5277;
  assign n5300 = n5284 & n5299;
  assign n5301 = ~n3637 & ~n5297;
  assign n5302 = ~n5300 & ~n5301;
  assign n5303 = ~n5298 & n5302;
  assign n5287 = ~n85 & ~n672;
  assign n5288 = ~n262 & n5287;
  assign n5289 = ~n216 & n5288;
  assign n5290 = n137 & n584;
  assign n5291 = ~n351 & ~n5290;
  assign n5292 = n5289 & ~n5291;
  assign n5293 = n4096 & n5292;
  assign n5294 = ~n2953 & n5293;
  assign n5295 = n593 & n5294;
  assign n5296 = n4596 & n5295;
  assign n5304 = n5303 ^ n5296;
  assign n5311 = ~n5296 & n5298;
  assign n5312 = n5277 ^ n3637;
  assign n5313 = n5296 ^ n5276;
  assign n5314 = n5278 & ~n5313;
  assign n5315 = n5312 & n5314;
  assign n5316 = n5315 ^ n3637;
  assign n5317 = ~n5285 & ~n5316;
  assign n5318 = ~n5311 & ~n5317;
  assign n5305 = ~n56 & n170;
  assign n5306 = ~n699 & ~n5305;
  assign n5307 = ~n464 & ~n644;
  assign n5308 = n786 & n5307;
  assign n5309 = n2988 & n5308;
  assign n5310 = ~n5306 & n5309;
  assign n5319 = n5318 ^ n5310;
  assign n5323 = ~n5276 & ~n5296;
  assign n5324 = ~n5310 & n5323;
  assign n5320 = n5310 ^ n5296;
  assign n5321 = ~n5313 & ~n5320;
  assign n5322 = ~n5277 & n5321;
  assign n5325 = n5324 ^ n5322;
  assign n5326 = n5284 & n5325;
  assign n5327 = n1070 & ~n2995;
  assign n5328 = n5277 & n5324;
  assign n5329 = n5328 ^ n5277;
  assign n5330 = ~n5327 & ~n5329;
  assign n5331 = n5330 ^ n5277;
  assign n5332 = n5326 & n5331;
  assign n5333 = n5328 ^ n5327;
  assign n5334 = ~n3637 & ~n5333;
  assign n5335 = ~n5332 & ~n5334;
  assign n5336 = n3637 & n5333;
  assign n5337 = ~n5326 & n5336;
  assign n5338 = n5335 & ~n5337;
  assign n5339 = ~x21 & ~x22;
  assign n5340 = n1070 & n5339;
  assign n5341 = ~n5327 & n5328;
  assign n5342 = n5285 ^ n3637;
  assign n5343 = n5341 & ~n5342;
  assign n5344 = n5343 ^ n3637;
  assign n5345 = ~n5340 & ~n5344;
  assign n5346 = n5327 & ~n5328;
  assign n5347 = ~n5339 & n5346;
  assign n5348 = n5326 & n5347;
  assign n5349 = ~n5345 & ~n5348;
  assign n5350 = n3637 & ~n5348;
  assign y0 = ~n3498;
  assign y1 = n3652;
  assign y2 = ~n3810;
  assign y3 = ~n3961;
  assign y4 = ~n4085;
  assign y5 = ~n4246;
  assign y6 = n4382;
  assign y7 = n4486;
  assign y8 = n4613;
  assign y9 = ~n4711;
  assign y10 = n4809;
  assign y11 = ~n4883;
  assign y12 = ~n4974;
  assign y13 = n5066;
  assign y14 = ~n5119;
  assign y15 = n5190;
  assign y16 = n5227;
  assign y17 = n5247;
  assign y18 = ~n5267;
  assign y19 = ~n5286;
  assign y20 = ~n5304;
  assign y21 = ~n5319;
  assign y22 = ~n5338;
  assign y23 = n5349;
  assign y24 = n5350;
endmodule
