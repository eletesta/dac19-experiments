module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63;
  wire n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356;
  assign n833 = x70 ^ x32;
  assign n834 = x75 ^ x58;
  assign n835 = n833 & n834;
  assign n836 = x74 ^ x0;
  assign n837 = x72 ^ x16;
  assign n838 = n836 & n837;
  assign n839 = x71 ^ x24;
  assign n840 = x73 ^ x8;
  assign n841 = ~n839 & n840;
  assign n842 = n838 & n841;
  assign n843 = n835 & n842;
  assign n844 = ~n833 & n834;
  assign n845 = n836 & ~n837;
  assign n846 = n839 & ~n840;
  assign n847 = n845 & n846;
  assign n848 = n839 & n840;
  assign n849 = ~n836 & ~n837;
  assign n850 = n848 & n849;
  assign n851 = ~n847 & ~n850;
  assign n852 = n844 & ~n851;
  assign n853 = ~n839 & ~n840;
  assign n854 = n838 & n853;
  assign n855 = n841 & n849;
  assign n856 = ~n854 & ~n855;
  assign n857 = n844 & ~n856;
  assign n858 = ~n833 & ~n834;
  assign n859 = n842 & n858;
  assign n860 = n833 & ~n834;
  assign n861 = n845 & n848;
  assign n862 = ~n836 & n837;
  assign n863 = n848 & n862;
  assign n864 = ~n861 & ~n863;
  assign n865 = n860 & ~n864;
  assign n866 = ~n859 & ~n865;
  assign n867 = ~n857 & n866;
  assign n868 = n841 & n862;
  assign n869 = n858 & n868;
  assign n870 = n849 & n853;
  assign n871 = ~n842 & ~n870;
  assign n872 = n860 & ~n871;
  assign n873 = ~n869 & ~n872;
  assign n874 = n845 & n853;
  assign n875 = n858 & n874;
  assign n876 = n853 & n862;
  assign n877 = n841 & n845;
  assign n878 = ~n876 & ~n877;
  assign n879 = n835 & ~n878;
  assign n880 = ~n875 & ~n879;
  assign n881 = n846 & n862;
  assign n882 = n838 & n846;
  assign n883 = ~n881 & ~n882;
  assign n884 = n851 & ~n868;
  assign n885 = n883 & n884;
  assign n886 = n835 & ~n885;
  assign n887 = n840 ^ n836;
  assign n888 = n839 ^ n837;
  assign n889 = ~n887 & ~n888;
  assign n890 = n844 & n889;
  assign n891 = ~n886 & ~n890;
  assign n892 = n858 & n876;
  assign n893 = n846 & n849;
  assign n894 = n856 & ~n893;
  assign n895 = ~n882 & n894;
  assign n896 = n860 & ~n895;
  assign n897 = n839 & n887;
  assign n898 = n858 & n897;
  assign n899 = ~n896 & ~n898;
  assign n900 = ~n892 & n899;
  assign n901 = n891 & n900;
  assign n902 = n880 & n901;
  assign n903 = n873 & n902;
  assign n904 = n867 & n903;
  assign n905 = ~n852 & n904;
  assign n906 = ~n843 & n905;
  assign n907 = n906 ^ x27;
  assign n908 = n907 ^ x129;
  assign n909 = x93 ^ x28;
  assign n910 = x88 ^ x2;
  assign n911 = n909 & ~n910;
  assign n912 = x90 ^ x52;
  assign n913 = x91 ^ x44;
  assign n914 = ~n912 & ~n913;
  assign n915 = x89 ^ x60;
  assign n916 = x92 ^ x36;
  assign n917 = ~n915 & ~n916;
  assign n918 = n914 & n917;
  assign n919 = n911 & n918;
  assign n920 = ~n909 & ~n910;
  assign n921 = n912 & n913;
  assign n922 = n915 & ~n916;
  assign n923 = n921 & n922;
  assign n924 = ~n912 & n913;
  assign n925 = n915 & n916;
  assign n926 = n924 & n925;
  assign n927 = ~n923 & ~n926;
  assign n928 = n920 & ~n927;
  assign n929 = ~n919 & ~n928;
  assign n930 = n909 & n910;
  assign n931 = ~n915 & n916;
  assign n932 = n921 & n931;
  assign n933 = n930 & n932;
  assign n934 = n912 & ~n913;
  assign n935 = n925 & n934;
  assign n936 = ~n923 & ~n935;
  assign n937 = n911 & ~n936;
  assign n938 = ~n933 & ~n937;
  assign n939 = n918 & n930;
  assign n940 = n917 & n921;
  assign n941 = n914 & n931;
  assign n942 = ~n940 & ~n941;
  assign n943 = n911 & ~n942;
  assign n944 = ~n939 & ~n943;
  assign n945 = n917 & n924;
  assign n946 = n930 & n945;
  assign n947 = ~n920 & ~n930;
  assign n948 = n931 & n934;
  assign n949 = ~n941 & ~n948;
  assign n950 = ~n947 & ~n949;
  assign n951 = ~n946 & ~n950;
  assign n952 = n924 & n931;
  assign n953 = n922 & n924;
  assign n954 = ~n926 & ~n953;
  assign n955 = ~n952 & n954;
  assign n956 = n911 & ~n955;
  assign n957 = n914 & n922;
  assign n958 = ~n940 & ~n957;
  assign n959 = n922 & n934;
  assign n960 = n921 & n925;
  assign n961 = ~n959 & ~n960;
  assign n962 = n958 & n961;
  assign n963 = n920 & ~n962;
  assign n964 = ~n956 & ~n963;
  assign n965 = n914 & n925;
  assign n966 = ~n909 & n910;
  assign n967 = ~n926 & ~n959;
  assign n968 = ~n966 & n967;
  assign n969 = ~n965 & n968;
  assign n970 = ~n932 & ~n965;
  assign n971 = n917 & n934;
  assign n972 = ~n952 & ~n971;
  assign n973 = ~n948 & ~n953;
  assign n974 = ~n960 & n973;
  assign n975 = n972 & n974;
  assign n976 = n930 & ~n967;
  assign n977 = n975 & ~n976;
  assign n978 = n970 & n977;
  assign n979 = ~n957 & n978;
  assign n980 = ~n969 & ~n979;
  assign n981 = n910 & n980;
  assign n982 = n964 & ~n981;
  assign n983 = n951 & n982;
  assign n984 = n944 & n983;
  assign n985 = n938 & n984;
  assign n986 = n929 & n985;
  assign n987 = n986 ^ x1;
  assign n988 = n987 ^ x124;
  assign n989 = ~n908 & n988;
  assign n990 = x82 ^ x34;
  assign n991 = x87 ^ x60;
  assign n992 = ~n990 & ~n991;
  assign n993 = x86 ^ x2;
  assign n994 = x83 ^ x26;
  assign n995 = x84 ^ x18;
  assign n996 = x85 ^ x10;
  assign n997 = n995 & n996;
  assign n998 = n994 & n997;
  assign n999 = ~n993 & n998;
  assign n1000 = n995 & ~n996;
  assign n1001 = ~n993 & ~n994;
  assign n1002 = n1000 & n1001;
  assign n1003 = ~n999 & ~n1002;
  assign n1004 = n993 & n994;
  assign n1005 = n1000 & n1004;
  assign n1006 = ~n995 & n996;
  assign n1007 = n994 & n1006;
  assign n1008 = ~n1005 & ~n1007;
  assign n1009 = ~n993 & n997;
  assign n1010 = ~n995 & ~n996;
  assign n1011 = ~n1001 & ~n1004;
  assign n1012 = n1010 & n1011;
  assign n1013 = ~n1009 & ~n1012;
  assign n1014 = n1008 & n1013;
  assign n1015 = n1003 & n1014;
  assign n1016 = n992 & n1015;
  assign n1017 = n991 & ~n1003;
  assign n1018 = n990 & n991;
  assign n1019 = ~n994 & n1010;
  assign n1020 = n995 & n1004;
  assign n1021 = n993 & n1006;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = ~n1019 & n1022;
  assign n1024 = n1018 & ~n1023;
  assign n1025 = ~n1017 & ~n1024;
  assign n1026 = ~n1016 & n1025;
  assign n1027 = ~n990 & n991;
  assign n1028 = n993 & n1000;
  assign n1029 = n996 ^ n994;
  assign n1030 = n996 ^ n995;
  assign n1031 = n1029 & ~n1030;
  assign n1032 = n1031 ^ n1006;
  assign n1033 = n993 & n1032;
  assign n1034 = n1033 ^ n1006;
  assign n1035 = ~n1028 & ~n1034;
  assign n1036 = n1027 & ~n1035;
  assign n1037 = n990 & ~n991;
  assign n1038 = n993 & n997;
  assign n1039 = ~n994 & n1006;
  assign n1040 = ~n993 & n1000;
  assign n1041 = n993 & n1010;
  assign n1042 = ~n997 & ~n1041;
  assign n1043 = n994 & ~n1042;
  assign n1044 = ~n1040 & ~n1043;
  assign n1045 = ~n1039 & n1044;
  assign n1046 = ~n1038 & n1045;
  assign n1047 = n1037 & n1046;
  assign n1048 = ~n1036 & ~n1047;
  assign n1049 = n1026 & n1048;
  assign n1050 = n1049 ^ x51;
  assign n1051 = n1050 ^ x126;
  assign n1052 = x67 ^ x40;
  assign n1053 = x66 ^ x48;
  assign n1054 = n1052 & n1053;
  assign n1055 = x65 ^ x56;
  assign n1056 = x68 ^ x32;
  assign n1057 = n1055 & ~n1056;
  assign n1058 = n1054 & n1057;
  assign n1059 = x69 ^ x24;
  assign n1060 = x64 ^ x6;
  assign n1061 = n1059 & n1060;
  assign n1062 = n1052 & ~n1053;
  assign n1063 = n1057 & n1062;
  assign n1064 = n1061 & n1063;
  assign n1065 = n1059 & ~n1060;
  assign n1066 = ~n1055 & n1056;
  assign n1067 = n1054 & n1066;
  assign n1068 = n1065 & n1067;
  assign n1069 = ~n1064 & ~n1068;
  assign n1070 = n1055 & n1056;
  assign n1071 = ~n1052 & n1053;
  assign n1072 = n1070 & n1071;
  assign n1073 = n1061 & n1072;
  assign n1074 = ~n1052 & ~n1053;
  assign n1075 = n1057 & n1074;
  assign n1076 = n1061 & n1075;
  assign n1078 = ~n1053 & ~n1055;
  assign n1077 = ~n1052 & n1056;
  assign n1079 = n1078 ^ n1077;
  assign n1080 = n1065 & n1079;
  assign n1081 = ~n1059 & ~n1060;
  assign n1082 = n1057 & n1071;
  assign n1083 = n1054 & n1070;
  assign n1084 = ~n1063 & ~n1083;
  assign n1085 = ~n1082 & n1084;
  assign n1086 = n1081 & ~n1085;
  assign n1087 = n1075 & n1081;
  assign n1088 = n1062 & n1066;
  assign n1089 = n1081 & n1088;
  assign n1090 = ~n1055 & ~n1056;
  assign n1091 = n1071 & n1090;
  assign n1092 = n1054 & n1090;
  assign n1093 = ~n1067 & ~n1088;
  assign n1094 = ~n1092 & n1093;
  assign n1095 = ~n1091 & n1094;
  assign n1096 = n1061 & ~n1095;
  assign n1097 = n1066 & n1074;
  assign n1098 = ~n1091 & ~n1097;
  assign n1099 = n1081 & ~n1098;
  assign n1100 = ~n1059 & n1060;
  assign n1101 = n1066 & n1071;
  assign n1102 = n1074 & n1090;
  assign n1103 = ~n1101 & ~n1102;
  assign n1104 = n1062 & n1070;
  assign n1105 = ~n1083 & ~n1092;
  assign n1106 = ~n1104 & n1105;
  assign n1107 = n1103 & n1106;
  assign n1108 = ~n1097 & n1107;
  assign n1109 = ~n1082 & n1108;
  assign n1110 = n1100 & ~n1109;
  assign n1111 = ~n1099 & ~n1110;
  assign n1112 = ~n1096 & n1111;
  assign n1113 = ~n1089 & n1112;
  assign n1114 = ~n1087 & n1113;
  assign n1115 = ~n1086 & n1114;
  assign n1116 = ~n1080 & n1115;
  assign n1117 = ~n1076 & n1116;
  assign n1118 = ~n1073 & n1117;
  assign n1119 = n1069 & n1118;
  assign n1120 = ~n1058 & n1119;
  assign n1121 = n1120 ^ x59;
  assign n1122 = n1121 ^ x125;
  assign n1123 = n1051 & n1122;
  assign n1124 = x100 ^ x4;
  assign n1125 = x105 ^ x30;
  assign n1126 = n1124 & n1125;
  assign n1127 = x101 ^ x62;
  assign n1128 = x103 ^ x46;
  assign n1129 = ~n1127 & ~n1128;
  assign n1130 = x102 ^ x54;
  assign n1131 = x104 ^ x38;
  assign n1132 = ~n1130 & n1131;
  assign n1133 = n1129 & n1132;
  assign n1134 = n1126 & n1133;
  assign n1135 = ~n1124 & n1125;
  assign n1136 = ~n1127 & n1128;
  assign n1137 = ~n1130 & ~n1131;
  assign n1138 = n1136 & n1137;
  assign n1139 = n1135 & n1138;
  assign n1140 = ~n1134 & ~n1139;
  assign n1141 = n1127 & ~n1128;
  assign n1142 = n1132 & n1141;
  assign n1143 = n1130 & ~n1131;
  assign n1144 = n1141 & n1143;
  assign n1145 = ~n1142 & ~n1144;
  assign n1146 = n1135 & ~n1145;
  assign n1147 = n1127 & n1128;
  assign n1148 = ~n1131 & n1147;
  assign n1149 = n1126 & n1148;
  assign n1150 = n1136 & n1143;
  assign n1151 = ~n1133 & ~n1150;
  assign n1152 = n1135 & ~n1151;
  assign n1153 = ~n1149 & ~n1152;
  assign n1154 = ~n1146 & n1153;
  assign n1155 = n1130 & n1131;
  assign n1156 = n1129 & n1155;
  assign n1157 = n1135 & n1156;
  assign n1158 = n1137 & n1141;
  assign n1159 = ~n1124 & ~n1125;
  assign n1160 = ~n1126 & ~n1159;
  assign n1161 = n1158 & ~n1160;
  assign n1162 = ~n1157 & ~n1161;
  assign n1163 = n1141 & n1155;
  assign n1164 = n1126 & n1163;
  assign n1165 = n1135 & n1147;
  assign n1166 = n1143 & n1165;
  assign n1167 = n1136 & n1155;
  assign n1168 = n1135 & n1167;
  assign n1169 = ~n1166 & ~n1168;
  assign n1170 = n1124 & ~n1125;
  assign n1171 = n1137 & n1147;
  assign n1172 = n1132 & n1136;
  assign n1173 = n1129 & n1143;
  assign n1174 = ~n1172 & ~n1173;
  assign n1175 = ~n1171 & n1174;
  assign n1176 = ~n1142 & ~n1150;
  assign n1177 = ~n1163 & n1176;
  assign n1178 = n1175 & n1177;
  assign n1179 = ~n1133 & n1178;
  assign n1180 = ~n1167 & n1179;
  assign n1181 = n1170 & n1180;
  assign n1182 = ~n1150 & n1174;
  assign n1183 = n1126 & ~n1182;
  assign n1184 = ~n1138 & ~n1156;
  assign n1185 = ~n1132 & ~n1143;
  assign n1186 = n1147 & n1185;
  assign n1187 = n1151 & ~n1186;
  assign n1188 = ~n1163 & n1187;
  assign n1189 = n1184 & n1188;
  assign n1190 = n1159 & ~n1189;
  assign n1191 = ~n1183 & ~n1190;
  assign n1192 = ~n1181 & n1191;
  assign n1193 = n1169 & n1192;
  assign n1194 = ~n1164 & n1193;
  assign n1195 = n1162 & n1194;
  assign n1196 = n1154 & n1195;
  assign n1197 = n1140 & n1196;
  assign n1198 = n1197 ^ x35;
  assign n1199 = n1198 ^ x128;
  assign n1200 = x99 ^ x62;
  assign n1201 = x94 ^ x36;
  assign n1202 = n1200 & ~n1201;
  assign n1203 = x96 ^ x20;
  assign n1204 = x95 ^ x28;
  assign n1205 = ~n1203 & ~n1204;
  assign n1206 = x98 ^ x4;
  assign n1207 = x97 ^ x12;
  assign n1208 = n1206 & ~n1207;
  assign n1209 = n1205 & n1208;
  assign n1210 = ~n1206 & ~n1207;
  assign n1211 = n1203 & ~n1204;
  assign n1212 = n1210 & n1211;
  assign n1213 = ~n1209 & ~n1212;
  assign n1214 = n1203 & n1204;
  assign n1215 = ~n1206 & n1207;
  assign n1216 = n1214 & n1215;
  assign n1217 = n1204 & n1208;
  assign n1218 = n1203 & n1217;
  assign n1219 = ~n1216 & ~n1218;
  assign n1220 = n1213 & n1219;
  assign n1221 = n1202 & ~n1220;
  assign n1222 = ~n1200 & ~n1201;
  assign n1223 = n1208 & n1211;
  assign n1224 = n1222 & n1223;
  assign n1225 = n1205 & n1210;
  assign n1226 = n1202 & n1225;
  assign n1227 = ~n1224 & ~n1226;
  assign n1228 = n1205 & n1215;
  assign n1229 = n1222 & n1228;
  assign n1230 = n1200 & n1201;
  assign n1231 = n1206 & n1207;
  assign n1232 = n1211 & n1231;
  assign n1233 = ~n1228 & ~n1232;
  assign n1234 = n1230 & ~n1233;
  assign n1235 = ~n1229 & ~n1234;
  assign n1236 = n1205 & n1231;
  assign n1237 = ~n1201 & n1236;
  assign n1238 = n1211 & n1215;
  assign n1239 = ~n1222 & ~n1230;
  assign n1240 = n1238 & ~n1239;
  assign n1241 = ~n1237 & ~n1240;
  assign n1242 = n1209 & n1230;
  assign n1243 = ~n1203 & n1204;
  assign n1244 = n1210 & n1243;
  assign n1245 = n1231 & n1243;
  assign n1246 = ~n1244 & ~n1245;
  assign n1247 = n1202 & ~n1246;
  assign n1248 = n1210 & n1214;
  assign n1249 = ~n1203 & n1217;
  assign n1250 = ~n1248 & ~n1249;
  assign n1251 = n1246 & n1250;
  assign n1252 = n1230 & ~n1251;
  assign n1253 = n1214 & n1231;
  assign n1254 = ~n1200 & n1201;
  assign n1255 = ~n1253 & ~n1254;
  assign n1256 = n1215 & n1243;
  assign n1257 = ~n1218 & ~n1248;
  assign n1258 = ~n1256 & n1257;
  assign n1259 = n1255 & n1258;
  assign n1260 = ~n1200 & ~n1259;
  assign n1261 = ~n1252 & ~n1260;
  assign n1262 = ~n1222 & n1246;
  assign n1263 = n1230 & ~n1250;
  assign n1264 = n1262 & ~n1263;
  assign n1265 = n1213 & n1264;
  assign n1266 = n1233 & n1265;
  assign n1267 = ~n1253 & n1266;
  assign n1268 = ~n1216 & n1267;
  assign n1269 = ~n1261 & ~n1268;
  assign n1270 = ~n1247 & ~n1269;
  assign n1271 = ~n1242 & n1270;
  assign n1272 = n1241 & n1271;
  assign n1273 = n1235 & n1272;
  assign n1274 = n1227 & n1273;
  assign n1275 = ~n1221 & n1274;
  assign n1276 = n1275 ^ x43;
  assign n1277 = n1276 ^ x127;
  assign n1278 = n1199 & n1277;
  assign n1279 = n1123 & n1278;
  assign n1280 = n989 & n1279;
  assign n1281 = n1051 & ~n1122;
  assign n1282 = ~n1199 & n1277;
  assign n1283 = n1281 & n1282;
  assign n1284 = n908 & n988;
  assign n1285 = ~n908 & ~n988;
  assign n1286 = ~n1284 & ~n1285;
  assign n1287 = n1283 & ~n1286;
  assign n1288 = n908 & ~n988;
  assign n1289 = ~n1051 & n1122;
  assign n1290 = n1278 & n1289;
  assign n1291 = n1288 & n1290;
  assign n1292 = n1278 & n1281;
  assign n1293 = n1284 & n1292;
  assign n1294 = n1199 & ~n1277;
  assign n1295 = n1289 & n1294;
  assign n1296 = n1285 & n1295;
  assign n1297 = ~n1293 & ~n1296;
  assign n1298 = ~n1291 & n1297;
  assign n1299 = ~n1287 & n1298;
  assign n1300 = n1285 & n1292;
  assign n1301 = n1123 & n1294;
  assign n1302 = ~n1290 & ~n1301;
  assign n1303 = n989 & ~n1302;
  assign n1304 = ~n1300 & ~n1303;
  assign n1305 = ~n1199 & ~n1277;
  assign n1306 = n1123 & n1305;
  assign n1307 = ~n1285 & n1306;
  assign n1308 = ~n1051 & ~n1122;
  assign n1309 = n1278 & n1308;
  assign n1310 = n1289 & n1305;
  assign n1311 = ~n1051 & n1282;
  assign n1312 = n1122 & n1311;
  assign n1313 = ~n1301 & ~n1312;
  assign n1314 = ~n1310 & n1313;
  assign n1315 = ~n1309 & n1314;
  assign n1316 = ~n1286 & ~n1315;
  assign n1317 = ~n1307 & ~n1316;
  assign n1318 = n1305 & n1308;
  assign n1319 = n1284 & n1318;
  assign n1320 = ~n1279 & ~n1295;
  assign n1321 = n1288 & ~n1320;
  assign n1322 = ~n1319 & ~n1321;
  assign n1323 = n1281 & n1305;
  assign n1324 = n1285 & n1323;
  assign n1325 = n1294 & n1308;
  assign n1326 = ~n1122 & n1311;
  assign n1327 = n1281 & n1294;
  assign n1328 = ~n1326 & ~n1327;
  assign n1329 = ~n1325 & n1328;
  assign n1330 = ~n1318 & n1329;
  assign n1331 = ~n1288 & n1330;
  assign n1332 = n1123 & n1282;
  assign n1333 = ~n1323 & ~n1325;
  assign n1334 = ~n989 & n1333;
  assign n1335 = ~n1326 & n1334;
  assign n1336 = ~n1332 & n1335;
  assign n1337 = ~n1331 & ~n1336;
  assign n1338 = n1286 & n1337;
  assign n1339 = ~n1324 & ~n1338;
  assign n1340 = n1322 & n1339;
  assign n1341 = n1317 & n1340;
  assign n1342 = n1304 & n1341;
  assign n1343 = n1299 & n1342;
  assign n1344 = ~n1280 & n1343;
  assign n1345 = n1344 ^ x2;
  assign n1346 = n1345 ^ x184;
  assign n1347 = ~n1023 & n1037;
  assign n1348 = ~n1015 & n1027;
  assign n1349 = ~n1347 & ~n1348;
  assign n1350 = n992 & ~n1035;
  assign n1351 = n1018 & ~n1046;
  assign n1352 = ~n1350 & ~n1351;
  assign n1353 = n1349 & n1352;
  assign n1354 = n1003 & n1353;
  assign n1355 = n1354 ^ x57;
  assign n1356 = n1355 ^ x159;
  assign n1357 = n850 & n858;
  assign n1358 = n835 & n881;
  assign n1359 = n844 & n868;
  assign n1360 = ~n1358 & ~n1359;
  assign n1361 = ~n1357 & n1360;
  assign n1362 = n838 & n848;
  assign n1363 = n834 ^ n833;
  assign n1364 = n1362 & ~n1363;
  assign n1365 = ~n855 & ~n893;
  assign n1366 = ~n874 & n1365;
  assign n1367 = n835 & ~n1366;
  assign n1368 = ~n1364 & ~n1367;
  assign n1369 = n858 & ~n895;
  assign n1370 = ~n854 & ~n870;
  assign n1371 = n864 & n1370;
  assign n1372 = ~n882 & n1371;
  assign n1373 = n844 & ~n1372;
  assign n1374 = ~n847 & n883;
  assign n1375 = ~n863 & n1374;
  assign n1376 = n878 & n1375;
  assign n1377 = n860 & ~n1376;
  assign n1378 = ~n1373 & ~n1377;
  assign n1379 = ~n1369 & n1378;
  assign n1380 = n1368 & n1379;
  assign n1381 = n880 & n1380;
  assign n1382 = n873 & n1381;
  assign n1383 = n1361 & n1382;
  assign n1384 = ~n852 & n1383;
  assign n1385 = ~n843 & n1384;
  assign n1386 = n1385 ^ x39;
  assign n1387 = n1386 ^ x154;
  assign n1388 = ~n1356 & n1387;
  assign n1389 = x78 ^ x50;
  assign n1390 = x80 ^ x34;
  assign n1391 = ~n1389 & ~n1390;
  assign n1392 = x79 ^ x42;
  assign n1393 = x77 ^ x58;
  assign n1394 = n1392 & ~n1393;
  assign n1395 = n1391 & n1394;
  assign n1396 = ~n1392 & n1393;
  assign n1397 = n1391 & n1396;
  assign n1398 = x81 ^ x26;
  assign n1399 = x76 ^ x0;
  assign n1400 = n1398 & ~n1399;
  assign n1401 = ~n1398 & n1399;
  assign n1402 = ~n1400 & ~n1401;
  assign n1403 = n1397 & n1402;
  assign n1404 = n1389 & n1390;
  assign n1405 = ~n1392 & ~n1393;
  assign n1406 = n1404 & n1405;
  assign n1407 = n1400 & n1406;
  assign n1408 = n1396 & n1404;
  assign n1409 = n1402 & n1408;
  assign n1410 = ~n1407 & ~n1409;
  assign n1411 = ~n1403 & n1410;
  assign n1412 = n1398 & n1399;
  assign n1413 = ~n1389 & n1390;
  assign n1414 = n1394 & n1413;
  assign n1415 = n1391 & n1405;
  assign n1416 = ~n1414 & ~n1415;
  assign n1417 = n1412 & ~n1416;
  assign n1418 = n1392 & n1393;
  assign n1419 = n1404 & n1418;
  assign n1420 = n1391 & n1418;
  assign n1421 = ~n1419 & ~n1420;
  assign n1422 = n1400 & ~n1421;
  assign n1423 = ~n1417 & ~n1422;
  assign n1424 = ~n1402 & ~n1416;
  assign n1425 = n1389 & ~n1390;
  assign n1426 = n1405 & n1425;
  assign n1427 = n1401 & n1426;
  assign n1428 = n1396 & n1413;
  assign n1429 = n1396 & n1425;
  assign n1430 = ~n1428 & ~n1429;
  assign n1431 = n1400 & ~n1430;
  assign n1432 = ~n1427 & ~n1431;
  assign n1433 = ~n1398 & ~n1399;
  assign n1434 = n1405 & n1413;
  assign n1435 = n1394 & n1404;
  assign n1436 = ~n1428 & ~n1435;
  assign n1437 = ~n1434 & n1436;
  assign n1438 = n1421 & n1437;
  assign n1439 = n1433 & ~n1438;
  assign n1440 = n1394 & n1425;
  assign n1441 = ~n1406 & ~n1440;
  assign n1442 = ~n1395 & n1441;
  assign n1443 = ~n1419 & n1442;
  assign n1444 = n1412 & ~n1443;
  assign n1445 = n1413 & n1418;
  assign n1446 = n1430 & ~n1445;
  assign n1447 = ~n1435 & n1446;
  assign n1448 = n1401 & ~n1447;
  assign n1449 = ~n1444 & ~n1448;
  assign n1450 = ~n1439 & n1449;
  assign n1451 = n1432 & n1450;
  assign n1452 = ~n1424 & n1451;
  assign n1453 = n1423 & n1452;
  assign n1454 = n1411 & n1453;
  assign n1455 = ~n1395 & n1454;
  assign n1456 = n1455 ^ x23;
  assign n1457 = n1456 ^ x156;
  assign n1458 = n1061 & ~n1103;
  assign n1459 = n1062 & n1090;
  assign n1460 = ~n1101 & ~n1459;
  assign n1461 = n1081 & ~n1460;
  assign n1462 = ~n1458 & ~n1461;
  assign n1463 = n1060 & n1067;
  assign n1464 = ~n1058 & ~n1104;
  assign n1465 = ~n1072 & ~n1082;
  assign n1466 = n1464 & n1465;
  assign n1467 = n1065 & ~n1466;
  assign n1468 = ~n1463 & ~n1467;
  assign n1469 = n1462 & n1468;
  assign n1470 = ~n1061 & ~n1081;
  assign n1471 = n1092 & ~n1470;
  assign n1472 = ~n1075 & n1098;
  assign n1473 = n1100 & ~n1472;
  assign n1474 = n1081 & ~n1465;
  assign n1475 = ~n1076 & ~n1474;
  assign n1476 = n1070 & n1074;
  assign n1477 = n1061 & n1476;
  assign n1478 = n1083 & ~n1470;
  assign n1479 = ~n1477 & ~n1478;
  assign n1480 = ~n1097 & ~n1459;
  assign n1481 = ~n1092 & n1480;
  assign n1482 = n1065 & ~n1481;
  assign n1483 = ~n1082 & n1464;
  assign n1484 = ~n1063 & n1483;
  assign n1485 = n1100 & ~n1484;
  assign n1486 = ~n1482 & ~n1485;
  assign n1487 = n1479 & n1486;
  assign n1488 = n1475 & n1487;
  assign n1489 = ~n1087 & n1488;
  assign n1490 = n1069 & n1489;
  assign n1491 = ~n1473 & n1490;
  assign n1492 = ~n1471 & n1491;
  assign n1493 = n1469 & n1492;
  assign n1494 = ~n1089 & n1493;
  assign n1495 = n1494 ^ x15;
  assign n1496 = n1495 ^ x157;
  assign n1497 = ~n1457 & n1496;
  assign n1498 = n1135 & n1172;
  assign n1499 = n1155 & n1165;
  assign n1500 = ~n1164 & ~n1499;
  assign n1501 = ~n1142 & ~n1167;
  assign n1502 = n1126 & ~n1501;
  assign n1503 = n1126 & n1173;
  assign n1504 = n1137 & n1165;
  assign n1505 = ~n1503 & ~n1504;
  assign n1506 = n1135 & n1173;
  assign n1507 = n1159 & n1180;
  assign n1508 = ~n1506 & ~n1507;
  assign n1509 = n1129 & n1137;
  assign n1510 = ~n1156 & ~n1509;
  assign n1511 = n1124 & ~n1510;
  assign n1512 = ~n1144 & n1188;
  assign n1513 = n1170 & ~n1512;
  assign n1514 = ~n1511 & ~n1513;
  assign n1515 = n1508 & n1514;
  assign n1516 = n1505 & n1515;
  assign n1517 = ~n1502 & n1516;
  assign n1518 = n1500 & n1517;
  assign n1519 = n1154 & n1518;
  assign n1520 = ~n1498 & n1519;
  assign n1521 = n1520 ^ x7;
  assign n1522 = n1521 ^ x158;
  assign n1523 = n1202 & n1238;
  assign n1524 = ~n1213 & ~n1239;
  assign n1525 = ~n1523 & ~n1524;
  assign n1526 = ~n1236 & ~n1253;
  assign n1527 = n1250 & n1526;
  assign n1528 = n1219 & n1527;
  assign n1529 = n1202 & ~n1528;
  assign n1530 = ~n1232 & ~n1256;
  assign n1531 = ~n1244 & n1530;
  assign n1532 = n1255 & n1531;
  assign n1533 = ~n1230 & n1532;
  assign n1534 = n1219 & ~n1256;
  assign n1535 = ~n1244 & n1534;
  assign n1536 = n1230 & ~n1535;
  assign n1537 = n1206 ^ n1203;
  assign n1538 = n1537 ^ n1204;
  assign n1539 = n1538 ^ n1207;
  assign n1540 = ~n1204 & n1539;
  assign n1541 = ~n1206 & n1540;
  assign n1542 = n1541 ^ n1538;
  assign n1543 = n1254 & ~n1542;
  assign n1544 = ~n1536 & ~n1543;
  assign n1545 = ~n1222 & n1544;
  assign n1546 = ~n1533 & ~n1545;
  assign n1547 = ~n1529 & ~n1546;
  assign n1548 = n1525 & n1547;
  assign n1549 = n1235 & n1548;
  assign n1550 = n1227 & n1549;
  assign n1551 = n1550 ^ x31;
  assign n1552 = n1551 ^ x155;
  assign n1553 = n1522 & n1552;
  assign n1554 = n1497 & n1553;
  assign n1555 = n1388 & n1554;
  assign n1556 = n1356 & ~n1387;
  assign n1557 = n1457 & n1496;
  assign n1558 = n1553 & n1557;
  assign n1559 = ~n1457 & ~n1496;
  assign n1560 = ~n1522 & n1552;
  assign n1561 = n1559 & n1560;
  assign n1562 = ~n1558 & ~n1561;
  assign n1563 = n1556 & ~n1562;
  assign n1564 = n1356 & n1387;
  assign n1565 = n1522 & ~n1552;
  assign n1566 = n1557 & n1565;
  assign n1567 = ~n1522 & ~n1552;
  assign n1568 = n1497 & n1567;
  assign n1569 = ~n1566 & ~n1568;
  assign n1570 = n1564 & ~n1569;
  assign n1571 = ~n1563 & ~n1570;
  assign n1572 = ~n1552 & n1559;
  assign n1573 = ~n1522 & n1572;
  assign n1574 = n1388 & n1573;
  assign n1575 = n1553 & n1559;
  assign n1576 = n1564 & n1575;
  assign n1577 = n1497 & n1560;
  assign n1578 = n1388 & n1577;
  assign n1579 = ~n1576 & ~n1578;
  assign n1580 = ~n1574 & n1579;
  assign n1581 = ~n1356 & ~n1387;
  assign n1582 = n1577 & n1581;
  assign n1583 = n1557 & n1567;
  assign n1584 = n1556 & n1583;
  assign n1585 = ~n1582 & ~n1584;
  assign n1586 = n1457 & ~n1496;
  assign n1587 = n1553 & n1586;
  assign n1588 = ~n1561 & ~n1587;
  assign n1589 = n1388 & ~n1588;
  assign n1590 = n1557 & n1560;
  assign n1591 = ~n1587 & ~n1590;
  assign n1592 = n1556 & ~n1591;
  assign n1593 = ~n1589 & ~n1592;
  assign n1594 = ~n1558 & ~n1575;
  assign n1595 = n1581 & ~n1594;
  assign n1596 = n1567 & n1586;
  assign n1597 = n1565 & n1586;
  assign n1598 = ~n1566 & ~n1597;
  assign n1599 = ~n1596 & n1598;
  assign n1600 = n1388 & ~n1599;
  assign n1601 = ~n1595 & ~n1600;
  assign n1602 = n1387 ^ n1356;
  assign n1603 = n1560 & n1586;
  assign n1604 = ~n1602 & n1603;
  assign n1605 = ~n1554 & ~n1596;
  assign n1606 = n1564 & ~n1605;
  assign n1607 = n1522 & n1572;
  assign n1608 = ~n1597 & ~n1607;
  assign n1609 = ~n1577 & n1608;
  assign n1610 = n1556 & ~n1609;
  assign n1611 = ~n1567 & ~n1581;
  assign n1612 = n1497 & n1565;
  assign n1613 = ~n1583 & ~n1612;
  assign n1614 = ~n1572 & n1613;
  assign n1615 = ~n1611 & ~n1614;
  assign n1616 = ~n1602 & n1615;
  assign n1617 = ~n1610 & ~n1616;
  assign n1618 = ~n1606 & n1617;
  assign n1619 = ~n1604 & n1618;
  assign n1620 = n1601 & n1619;
  assign n1621 = n1593 & n1620;
  assign n1622 = n1585 & n1621;
  assign n1623 = n1580 & n1622;
  assign n1624 = n1571 & n1623;
  assign n1625 = ~n1555 & n1624;
  assign n1626 = n1625 ^ x28;
  assign n1627 = n1626 ^ x189;
  assign n1628 = ~n1346 & n1627;
  assign n1629 = n1400 & n1426;
  assign n1630 = n1402 & n1445;
  assign n1631 = ~n1629 & ~n1630;
  assign n1632 = n1401 & n1419;
  assign n1633 = n1400 & n1434;
  assign n1634 = ~n1632 & ~n1633;
  assign n1635 = n1397 & ~n1398;
  assign n1636 = n1408 & n1412;
  assign n1637 = ~n1635 & ~n1636;
  assign n1638 = n1401 & ~n1441;
  assign n1639 = ~n1424 & ~n1638;
  assign n1640 = n1637 & n1639;
  assign n1641 = ~n1400 & ~n1430;
  assign n1642 = n1418 & n1425;
  assign n1643 = ~n1408 & ~n1642;
  assign n1644 = n1421 & n1643;
  assign n1645 = n1400 & ~n1644;
  assign n1646 = n1433 & ~n1442;
  assign n1647 = ~n1406 & ~n1415;
  assign n1648 = ~n1395 & n1647;
  assign n1649 = n1412 & ~n1648;
  assign n1650 = n1399 ^ n1398;
  assign n1651 = n1435 & ~n1650;
  assign n1652 = ~n1649 & ~n1651;
  assign n1653 = ~n1646 & n1652;
  assign n1654 = ~n1645 & n1653;
  assign n1655 = ~n1641 & n1654;
  assign n1656 = n1640 & n1655;
  assign n1657 = n1634 & n1656;
  assign n1658 = n1631 & n1657;
  assign n1659 = n1658 ^ x17;
  assign n1660 = n1659 ^ x120;
  assign n1661 = x111 ^ x56;
  assign n1662 = x106 ^ x38;
  assign n1663 = n1661 & n1662;
  assign n1664 = x109 ^ x14;
  assign n1665 = x108 ^ x22;
  assign n1666 = ~n1664 & n1665;
  assign n1667 = x110 ^ x6;
  assign n1668 = x107 ^ x30;
  assign n1669 = ~n1667 & n1668;
  assign n1670 = n1666 & n1669;
  assign n1671 = n1663 & n1670;
  assign n1672 = n1667 & n1668;
  assign n1673 = n1666 & n1672;
  assign n1674 = ~n1661 & ~n1662;
  assign n1675 = ~n1663 & ~n1674;
  assign n1676 = n1673 & ~n1675;
  assign n1677 = n1664 & ~n1665;
  assign n1678 = n1672 & n1677;
  assign n1679 = n1664 & n1665;
  assign n1680 = n1669 & n1679;
  assign n1681 = ~n1678 & ~n1680;
  assign n1682 = n1663 & ~n1681;
  assign n1683 = ~n1676 & ~n1682;
  assign n1684 = ~n1661 & n1662;
  assign n1685 = ~n1664 & ~n1665;
  assign n1686 = n1669 & n1685;
  assign n1687 = ~n1673 & ~n1686;
  assign n1688 = n1684 & ~n1687;
  assign n1689 = n1672 & n1679;
  assign n1690 = n1669 & n1677;
  assign n1691 = ~n1689 & ~n1690;
  assign n1692 = ~n1670 & n1691;
  assign n1693 = n1674 & ~n1692;
  assign n1694 = ~n1688 & ~n1693;
  assign n1695 = n1661 & ~n1662;
  assign n1696 = n1667 & ~n1668;
  assign n1697 = n1679 & n1696;
  assign n1698 = ~n1667 & ~n1668;
  assign n1699 = n1685 & n1698;
  assign n1700 = ~n1697 & ~n1699;
  assign n1701 = n1666 & n1696;
  assign n1702 = n1679 & n1698;
  assign n1703 = ~n1701 & ~n1702;
  assign n1704 = n1700 & n1703;
  assign n1705 = n1695 & ~n1704;
  assign n1706 = n1677 & n1696;
  assign n1707 = n1663 & n1706;
  assign n1708 = ~n1691 & n1695;
  assign n1709 = ~n1707 & ~n1708;
  assign n1710 = ~n1674 & ~n1684;
  assign n1711 = ~n1697 & ~n1706;
  assign n1712 = ~n1710 & ~n1711;
  assign n1713 = n1672 & n1685;
  assign n1714 = ~n1670 & ~n1713;
  assign n1715 = n1695 & ~n1714;
  assign n1716 = ~n1712 & ~n1715;
  assign n1717 = n1685 & n1696;
  assign n1718 = n1666 & n1698;
  assign n1719 = ~n1717 & ~n1718;
  assign n1720 = ~n1675 & ~n1719;
  assign n1721 = n1663 & n1699;
  assign n1722 = n1677 & n1698;
  assign n1723 = ~n1680 & ~n1722;
  assign n1724 = ~n1713 & n1723;
  assign n1725 = ~n1699 & n1724;
  assign n1726 = n1684 & ~n1725;
  assign n1727 = ~n1721 & ~n1726;
  assign n1728 = ~n1720 & n1727;
  assign n1729 = n1716 & n1728;
  assign n1730 = n1709 & n1729;
  assign n1731 = ~n1705 & n1730;
  assign n1732 = n1694 & n1731;
  assign n1733 = n1683 & n1732;
  assign n1734 = ~n1671 & n1733;
  assign n1735 = n1734 ^ x25;
  assign n1736 = n1735 ^ x119;
  assign n1737 = ~n1660 & n1736;
  assign n1738 = n987 ^ x122;
  assign n1739 = ~n1133 & ~n1173;
  assign n1740 = n1159 & ~n1739;
  assign n1741 = n1170 & ~n1184;
  assign n1742 = ~n1740 & ~n1741;
  assign n1743 = n1160 & n1509;
  assign n1744 = n1170 & n1172;
  assign n1745 = n1125 ^ n1124;
  assign n1746 = ~n1177 & n1745;
  assign n1747 = n1147 & ~n1185;
  assign n1748 = ~n1138 & ~n1747;
  assign n1749 = n1126 & ~n1748;
  assign n1750 = ~n1746 & ~n1749;
  assign n1751 = n1143 & n1147;
  assign n1752 = n1170 & n1751;
  assign n1753 = n1130 & n1148;
  assign n1754 = n1753 ^ n1147;
  assign n1755 = ~n1144 & ~n1754;
  assign n1756 = ~n1167 & n1755;
  assign n1757 = n1159 & ~n1756;
  assign n1758 = ~n1752 & ~n1757;
  assign n1759 = n1750 & n1758;
  assign n1760 = ~n1744 & n1759;
  assign n1761 = ~n1743 & n1760;
  assign n1762 = n1742 & n1761;
  assign n1763 = n1162 & n1762;
  assign n1764 = ~n1502 & n1763;
  assign n1765 = n1505 & n1764;
  assign n1766 = n1140 & n1765;
  assign n1767 = ~n1498 & n1766;
  assign n1768 = n1767 ^ x9;
  assign n1769 = n1768 ^ x121;
  assign n1770 = n1738 & n1769;
  assign n1771 = n1737 & n1770;
  assign n1772 = n1222 & n1238;
  assign n1773 = ~n1201 & n1244;
  assign n1774 = ~n1772 & ~n1773;
  assign n1775 = ~n1209 & ~n1223;
  assign n1776 = ~n1239 & ~n1775;
  assign n1777 = n1233 & ~n1236;
  assign n1778 = ~n1212 & ~n1216;
  assign n1779 = n1250 & n1778;
  assign n1780 = n1777 & n1779;
  assign n1781 = n1202 & ~n1780;
  assign n1782 = ~n1776 & ~n1781;
  assign n1783 = ~n1225 & ~n1228;
  assign n1784 = n1230 & ~n1783;
  assign n1785 = ~n1245 & n1258;
  assign n1786 = n1200 & n1785;
  assign n1787 = ~n1230 & n1534;
  assign n1788 = ~n1245 & n1787;
  assign n1789 = ~n1239 & ~n1788;
  assign n1790 = n1527 & n1531;
  assign n1791 = ~n1212 & n1790;
  assign n1792 = n1254 & ~n1791;
  assign n1793 = ~n1789 & ~n1792;
  assign n1794 = ~n1786 & ~n1793;
  assign n1795 = ~n1784 & ~n1794;
  assign n1796 = n1782 & n1795;
  assign n1797 = n1774 & n1796;
  assign n1798 = n1797 ^ x33;
  assign n1799 = n1798 ^ x118;
  assign n1800 = n1121 ^ x123;
  assign n1801 = ~n1799 & ~n1800;
  assign n1802 = n1771 & n1801;
  assign n1803 = n1799 & ~n1800;
  assign n1804 = n1660 & n1736;
  assign n1805 = n1738 & ~n1769;
  assign n1806 = n1804 & n1805;
  assign n1807 = n1803 & n1806;
  assign n1808 = ~n1802 & ~n1807;
  assign n1809 = ~n1799 & n1800;
  assign n1810 = ~n1738 & ~n1769;
  assign n1811 = n1804 & n1810;
  assign n1812 = n1809 & n1811;
  assign n1813 = n1660 & ~n1736;
  assign n1814 = n1805 & n1813;
  assign n1815 = n1799 & n1800;
  assign n1816 = ~n1801 & ~n1815;
  assign n1817 = n1814 & ~n1816;
  assign n1818 = ~n1812 & ~n1817;
  assign n1819 = ~n1738 & n1769;
  assign n1820 = n1737 & n1819;
  assign n1821 = ~n1806 & ~n1820;
  assign n1822 = n1801 & ~n1821;
  assign n1823 = n1771 & n1815;
  assign n1824 = n1737 & n1805;
  assign n1825 = ~n1811 & ~n1824;
  assign n1826 = n1803 & ~n1825;
  assign n1827 = ~n1823 & ~n1826;
  assign n1828 = ~n1822 & n1827;
  assign n1829 = n1813 & n1819;
  assign n1830 = n1815 & n1829;
  assign n1831 = ~n1660 & ~n1736;
  assign n1832 = n1810 & n1831;
  assign n1833 = n1815 & n1832;
  assign n1834 = n1804 & n1819;
  assign n1835 = n1809 & n1834;
  assign n1836 = n1805 & n1831;
  assign n1837 = n1815 & n1836;
  assign n1838 = ~n1835 & ~n1837;
  assign n1839 = n1815 & ~n1825;
  assign n1840 = n1799 & n1834;
  assign n1841 = n1770 & n1804;
  assign n1842 = n1819 & n1831;
  assign n1843 = ~n1736 & n1805;
  assign n1844 = ~n1842 & ~n1843;
  assign n1845 = ~n1832 & n1844;
  assign n1846 = ~n1841 & n1845;
  assign n1847 = ~n1771 & n1846;
  assign n1848 = n1809 & ~n1847;
  assign n1849 = n1737 & n1810;
  assign n1850 = n1770 & n1831;
  assign n1851 = n1810 & n1813;
  assign n1852 = ~n1850 & ~n1851;
  assign n1853 = ~n1832 & n1852;
  assign n1854 = ~n1849 & n1853;
  assign n1855 = n1801 & ~n1854;
  assign n1856 = n1769 & n1803;
  assign n1857 = ~n1736 & n1856;
  assign n1858 = ~n1855 & ~n1857;
  assign n1859 = ~n1848 & n1858;
  assign n1860 = ~n1840 & n1859;
  assign n1861 = ~n1839 & n1860;
  assign n1862 = n1838 & n1861;
  assign n1863 = ~n1833 & n1862;
  assign n1864 = ~n1830 & n1863;
  assign n1865 = n1828 & n1864;
  assign n1866 = n1818 & n1865;
  assign n1867 = n1808 & n1866;
  assign n1868 = n1867 ^ x52;
  assign n1869 = n1868 ^ x186;
  assign n1870 = ~n1470 & n1476;
  assign n1871 = n1084 & n1465;
  assign n1872 = n1100 & ~n1871;
  assign n1873 = ~n1870 & ~n1872;
  assign n1874 = n1061 & n1082;
  assign n1875 = ~n1058 & ~n1072;
  assign n1876 = n1081 & ~n1875;
  assign n1877 = ~n1874 & ~n1876;
  assign n1878 = ~n1075 & n1103;
  assign n1879 = n1065 & ~n1878;
  assign n1880 = ~n1083 & n1483;
  assign n1881 = n1065 & ~n1880;
  assign n1882 = n1094 & ~n1097;
  assign n1883 = n1100 & ~n1882;
  assign n1884 = ~n1881 & ~n1883;
  assign n1885 = n1061 & ~n1460;
  assign n1886 = ~n1088 & n1460;
  assign n1887 = ~n1092 & n1886;
  assign n1888 = ~n1081 & n1887;
  assign n1889 = ~n1095 & ~n1888;
  assign n1890 = ~n1885 & ~n1889;
  assign n1891 = ~n1470 & ~n1890;
  assign n1892 = n1884 & ~n1891;
  assign n1893 = ~n1879 & n1892;
  assign n1894 = n1877 & n1893;
  assign n1895 = n1873 & n1894;
  assign n1896 = ~n1073 & n1895;
  assign n1897 = ~n1087 & n1896;
  assign n1898 = n1069 & n1897;
  assign n1899 = n1898 ^ x61;
  assign n1900 = n1899 ^ x135;
  assign n1968 = n930 & ~n936;
  assign n1969 = ~n918 & ~n948;
  assign n1970 = n966 & ~n1969;
  assign n1971 = ~n1968 & ~n1970;
  assign n1972 = ~n945 & ~n952;
  assign n1973 = ~n948 & n1972;
  assign n1974 = n930 & ~n1973;
  assign n1975 = ~n940 & n961;
  assign n1976 = n954 & n1975;
  assign n1977 = n966 & ~n1976;
  assign n1978 = ~n1974 & ~n1977;
  assign n1979 = n910 & n957;
  assign n1980 = ~n947 & n965;
  assign n1981 = ~n1979 & ~n1980;
  assign n1982 = ~n932 & ~n959;
  assign n1983 = ~n941 & ~n971;
  assign n1984 = ~n945 & n1983;
  assign n1985 = n1982 & n1984;
  assign n1986 = n920 & ~n1985;
  assign n1987 = n958 & n975;
  assign n1988 = n911 & ~n1987;
  assign n1989 = ~n1986 & ~n1988;
  assign n1990 = n1981 & n1989;
  assign n1991 = n1978 & n1990;
  assign n1992 = n1971 & n1991;
  assign n1993 = n929 & n1992;
  assign n1994 = ~n933 & n1993;
  assign n1995 = n1994 ^ x19;
  assign n1996 = n1995 ^ x132;
  assign n1901 = n1420 & n1433;
  assign n1902 = n1402 & n1428;
  assign n1903 = ~n1901 & ~n1902;
  assign n1904 = n1412 & ~n1421;
  assign n1905 = ~n1398 & n1445;
  assign n1906 = ~n1429 & ~n1642;
  assign n1907 = ~n1402 & ~n1906;
  assign n1908 = ~n1415 & ~n1420;
  assign n1909 = ~n1445 & n1908;
  assign n1910 = ~n1440 & n1909;
  assign n1911 = n1400 & ~n1910;
  assign n1912 = ~n1907 & ~n1911;
  assign n1913 = ~n1434 & n1648;
  assign n1914 = n1401 & ~n1913;
  assign n1915 = ~n1395 & ~n1397;
  assign n1916 = ~n1433 & n1915;
  assign n1917 = ~n1414 & ~n1440;
  assign n1918 = ~n1412 & n1917;
  assign n1919 = ~n1916 & ~n1918;
  assign n1920 = ~n1426 & ~n1919;
  assign n1921 = ~n1435 & n1920;
  assign n1922 = n1402 & ~n1921;
  assign n1923 = ~n1914 & ~n1922;
  assign n1924 = n1912 & n1923;
  assign n1925 = ~n1905 & n1924;
  assign n1926 = ~n1904 & n1925;
  assign n1927 = n1903 & n1926;
  assign n1928 = n1410 & n1927;
  assign n1929 = n1634 & n1928;
  assign n1930 = n1929 ^ x3;
  assign n1931 = n1930 ^ x134;
  assign n1933 = ~n1699 & ~n1701;
  assign n1934 = n1663 & ~n1933;
  assign n1935 = n1663 & n1722;
  assign n1936 = ~n1673 & ~n1678;
  assign n1937 = n1695 & ~n1936;
  assign n1938 = ~n1935 & ~n1937;
  assign n1939 = n1703 & n1719;
  assign n1940 = n1674 & ~n1939;
  assign n1941 = ~n1702 & ~n1717;
  assign n1942 = n1700 & n1941;
  assign n1943 = n1684 & ~n1942;
  assign n1944 = n1695 & ~n1939;
  assign n1945 = n1674 & n1678;
  assign n1946 = ~n1680 & ~n1686;
  assign n1947 = n1663 & ~n1946;
  assign n1948 = ~n1945 & ~n1947;
  assign n1949 = ~n1689 & n1948;
  assign n1950 = ~n1675 & ~n1949;
  assign n1951 = ~n1684 & ~n1686;
  assign n1952 = n1674 & n1686;
  assign n1953 = n1714 & ~n1952;
  assign n1954 = ~n1673 & n1953;
  assign n1955 = ~n1951 & ~n1954;
  assign n1956 = ~n1690 & ~n1955;
  assign n1957 = ~n1710 & ~n1956;
  assign n1958 = ~n1950 & ~n1957;
  assign n1959 = ~n1944 & n1958;
  assign n1960 = ~n1671 & n1959;
  assign n1961 = ~n1943 & n1960;
  assign n1962 = ~n1940 & n1961;
  assign n1963 = n1938 & n1962;
  assign n1964 = n1709 & n1963;
  assign n1965 = ~n1934 & n1964;
  assign n1966 = n1965 ^ x11;
  assign n1967 = n1966 ^ x133;
  assign n2007 = ~n1931 & n1967;
  assign n1932 = n1198 ^ x130;
  assign n1997 = n907 ^ x131;
  assign n2032 = n1932 & ~n1997;
  assign n2033 = ~n2007 & n2032;
  assign n2034 = ~n1996 & n2033;
  assign n2010 = n1967 ^ n1931;
  assign n2011 = n1997 & ~n2010;
  assign n2006 = n1996 & ~n1997;
  assign n2035 = n2006 & n2007;
  assign n2036 = ~n2011 & ~n2035;
  assign n2037 = n1932 & ~n2036;
  assign n1998 = n1996 & n1997;
  assign n2038 = n1998 & n2010;
  assign n2008 = ~n1932 & n2007;
  assign n2039 = n1931 & n2006;
  assign n2040 = ~n1967 & n1997;
  assign n2041 = ~n2039 & ~n2040;
  assign n2042 = ~n1932 & ~n2041;
  assign n2043 = ~n2008 & ~n2042;
  assign n2044 = ~n2038 & ~n2043;
  assign n2045 = ~n2037 & ~n2044;
  assign n2046 = ~n2034 & n2045;
  assign n2000 = ~n1996 & n1997;
  assign n2001 = n1967 & n2000;
  assign n1999 = ~n1967 & n1998;
  assign n2002 = n2001 ^ n1999;
  assign n2003 = n1932 & n2002;
  assign n2004 = n2003 ^ n2001;
  assign n2005 = ~n1931 & n2004;
  assign n2009 = n2006 & n2008;
  assign n2012 = ~n1996 & n2011;
  assign n2013 = ~n2000 & ~n2006;
  assign n2014 = n1931 & ~n1967;
  assign n2015 = n2013 & n2014;
  assign n2016 = ~n2012 & ~n2015;
  assign n2017 = n1996 ^ n1931;
  assign n2018 = ~n1967 & ~n2017;
  assign n2019 = n2016 & ~n2018;
  assign n2020 = ~n1932 & ~n2019;
  assign n2021 = ~n2009 & ~n2020;
  assign n2022 = n2000 & n2014;
  assign n2023 = n1931 & n1967;
  assign n2024 = n1996 & n2023;
  assign n2025 = n2014 ^ n1996;
  assign n2026 = ~n1997 & ~n2025;
  assign n2027 = ~n2024 & ~n2026;
  assign n2028 = ~n2022 & n2027;
  assign n2029 = n1932 & ~n2028;
  assign n2030 = n2021 & ~n2029;
  assign n2031 = ~n2005 & n2030;
  assign n2047 = n2046 ^ n2031;
  assign n2048 = n1900 & ~n2047;
  assign n2049 = n2048 ^ n2046;
  assign n2050 = n2049 ^ x36;
  assign n2051 = n2050 ^ x188;
  assign n2052 = n1735 ^ x117;
  assign n2053 = n1521 ^ x112;
  assign n2054 = n2052 & n2053;
  assign n2055 = n1355 ^ x113;
  assign n2056 = n1798 ^ x116;
  assign n2057 = n2055 & n2056;
  assign n2058 = n835 & n868;
  assign n2059 = n858 & ~n883;
  assign n2060 = ~n2058 & ~n2059;
  assign n2061 = n858 & ~n864;
  assign n2062 = ~n882 & ~n1362;
  assign n2063 = n834 & ~n2062;
  assign n2064 = n844 & ~n1366;
  assign n2065 = ~n842 & n1366;
  assign n2066 = n858 & ~n2065;
  assign n2067 = ~n2064 & ~n2066;
  assign n2068 = ~n870 & ~n877;
  assign n2069 = ~n874 & n2068;
  assign n2070 = ~n861 & n2069;
  assign n2071 = n835 & ~n2070;
  assign n2072 = ~n881 & ~n893;
  assign n2073 = ~n842 & n2072;
  assign n2074 = n884 & n1370;
  assign n2075 = n2073 & n2074;
  assign n2076 = n860 & ~n2075;
  assign n2077 = ~n2071 & ~n2076;
  assign n2078 = n2067 & n2077;
  assign n2079 = ~n852 & n2078;
  assign n2080 = ~n2063 & n2079;
  assign n2081 = ~n2061 & n2080;
  assign n2082 = n1360 & n2081;
  assign n2083 = n2060 & n2082;
  assign n2084 = n2083 ^ x49;
  assign n2085 = n2084 ^ x114;
  assign n2086 = ~n947 & ~n972;
  assign n2087 = n920 & ~n1976;
  assign n2088 = ~n2086 & ~n2087;
  assign n2089 = ~n911 & n965;
  assign n2090 = n973 & n1982;
  assign n2091 = ~n935 & n2090;
  assign n2092 = ~n957 & n2091;
  assign n2093 = n911 & ~n2092;
  assign n2094 = n927 & ~n960;
  assign n2095 = ~n966 & n2094;
  assign n2096 = ~n935 & n1973;
  assign n2097 = ~n926 & n2096;
  assign n2098 = n958 & n2097;
  assign n2099 = ~n930 & n2098;
  assign n2100 = ~n2095 & ~n2099;
  assign n2101 = n910 & n2100;
  assign n2102 = ~n2093 & ~n2101;
  assign n2103 = ~n2089 & n2102;
  assign n2104 = n2088 & n2103;
  assign n2105 = n944 & n2104;
  assign n2106 = ~n933 & n2105;
  assign n2107 = n2106 ^ x41;
  assign n2108 = n2107 ^ x115;
  assign n2109 = n2085 & n2108;
  assign n2110 = n2057 & n2109;
  assign n2111 = n2054 & n2110;
  assign n2112 = n2052 & ~n2053;
  assign n2113 = ~n2085 & n2108;
  assign n2114 = ~n2055 & ~n2056;
  assign n2115 = n2113 & n2114;
  assign n2116 = n2112 & n2115;
  assign n2117 = ~n2111 & ~n2116;
  assign n2118 = n2055 & ~n2056;
  assign n2119 = ~n2085 & ~n2108;
  assign n2120 = n2118 & n2119;
  assign n2121 = n2054 & n2120;
  assign n2122 = n2109 & n2118;
  assign n2123 = n2085 & ~n2108;
  assign n2124 = n2118 & n2123;
  assign n2125 = n2057 & n2119;
  assign n2126 = ~n2124 & ~n2125;
  assign n2127 = ~n2122 & n2126;
  assign n2128 = n2112 & ~n2127;
  assign n2129 = ~n2121 & ~n2128;
  assign n2130 = n2114 & n2123;
  assign n2131 = n2054 & n2130;
  assign n2132 = ~n2052 & n2053;
  assign n2133 = ~n2055 & n2056;
  assign n2134 = n2119 & n2133;
  assign n2135 = n2132 & n2134;
  assign n2136 = ~n2131 & ~n2135;
  assign n2137 = n2113 & n2133;
  assign n2138 = n2132 & n2137;
  assign n2139 = n2054 & n2134;
  assign n2140 = ~n2138 & ~n2139;
  assign n2141 = ~n2052 & ~n2053;
  assign n2142 = n2134 & n2141;
  assign n2143 = n2123 & n2133;
  assign n2144 = n2112 & n2143;
  assign n2145 = ~n2142 & ~n2144;
  assign n2146 = n2109 & n2114;
  assign n2147 = n2141 & n2146;
  assign n2148 = n2057 & n2113;
  assign n2149 = n2109 & n2133;
  assign n2150 = n2114 & n2119;
  assign n2151 = ~n2149 & ~n2150;
  assign n2152 = ~n2148 & n2151;
  assign n2153 = ~n2122 & n2152;
  assign n2154 = n2054 & ~n2153;
  assign n2155 = ~n2147 & ~n2154;
  assign n2156 = ~n2130 & ~n2143;
  assign n2157 = ~n2052 & ~n2156;
  assign n2158 = n2113 & n2118;
  assign n2159 = n2057 & n2123;
  assign n2160 = ~n2149 & ~n2159;
  assign n2161 = ~n2158 & n2160;
  assign n2162 = n2112 & ~n2161;
  assign n2163 = n2141 & n2158;
  assign n2164 = ~n2124 & ~n2148;
  assign n2165 = ~n2110 & n2164;
  assign n2166 = n2141 & ~n2165;
  assign n2167 = ~n2120 & ~n2159;
  assign n2168 = ~n2122 & n2167;
  assign n2169 = ~n2110 & n2168;
  assign n2170 = n2132 & ~n2169;
  assign n2171 = ~n2166 & ~n2170;
  assign n2172 = ~n2163 & n2171;
  assign n2173 = ~n2162 & n2172;
  assign n2174 = ~n2157 & n2173;
  assign n2175 = n2155 & n2174;
  assign n2176 = n2145 & n2175;
  assign n2177 = n2140 & n2176;
  assign n2178 = n2136 & n2177;
  assign n2179 = n2129 & n2178;
  assign n2180 = n2117 & n2179;
  assign n2181 = n2180 ^ x60;
  assign n2182 = n2181 ^ x185;
  assign n2183 = n2051 & ~n2182;
  assign n2184 = ~n1869 & n2183;
  assign n2185 = n1628 & n2184;
  assign n2186 = n1346 & ~n1627;
  assign n2187 = ~n993 & n1006;
  assign n2188 = n994 & n1000;
  assign n2189 = ~n2187 & ~n2188;
  assign n2190 = ~n994 & ~n1042;
  assign n2191 = n2189 & ~n2190;
  assign n2192 = ~n1038 & n2191;
  assign n2193 = n1027 & ~n2192;
  assign n2194 = ~n1004 & n1006;
  assign n2195 = n1010 & ~n1011;
  assign n2196 = ~n2194 & ~n2195;
  assign n2197 = ~n999 & n2196;
  assign n2198 = ~n1028 & n2197;
  assign n2199 = n1037 & ~n2198;
  assign n2200 = ~n2193 & ~n2199;
  assign n2201 = n1006 & ~n1011;
  assign n2202 = ~n1019 & ~n2201;
  assign n2203 = ~n998 & n2202;
  assign n2204 = ~n1028 & n2203;
  assign n2205 = n992 & n2204;
  assign n2206 = ~n994 & n995;
  assign n2207 = n993 & n2206;
  assign n2208 = ~n993 & n1010;
  assign n2209 = ~n2201 & ~n2208;
  assign n2210 = ~n2207 & n2209;
  assign n2211 = n1003 & n2210;
  assign n2212 = n1018 & ~n2211;
  assign n2213 = ~n2205 & ~n2212;
  assign n2214 = n2200 & n2213;
  assign n2215 = n2214 ^ x37;
  assign n2216 = n2215 ^ x142;
  assign n2217 = n910 & ~n954;
  assign n2218 = ~n935 & n961;
  assign n2219 = ~n965 & n2218;
  assign n2220 = n920 & ~n2219;
  assign n2221 = n970 & n972;
  assign n2222 = n958 & n2221;
  assign n2223 = n911 & ~n2222;
  assign n2224 = ~n923 & n970;
  assign n2225 = ~n945 & n2224;
  assign n2226 = n966 & ~n2225;
  assign n2227 = ~n2223 & ~n2226;
  assign n2228 = n920 & n941;
  assign n2229 = ~n920 & n1984;
  assign n2230 = ~n957 & n1972;
  assign n2231 = ~n930 & n2230;
  assign n2232 = ~n2229 & ~n2231;
  assign n2233 = ~n947 & n2232;
  assign n2234 = ~n2228 & ~n2233;
  assign n2235 = n2227 & n2234;
  assign n2236 = n938 & n2235;
  assign n2237 = ~n2220 & n2236;
  assign n2238 = ~n2217 & n2237;
  assign n2239 = n1971 & n2238;
  assign n2240 = n2239 ^ x63;
  assign n2241 = n2240 ^ x147;
  assign n2242 = ~n2216 & n2241;
  assign n2243 = ~n1670 & ~n1718;
  assign n2244 = n1695 & ~n2243;
  assign n2245 = n1662 & n1713;
  assign n2246 = ~n1675 & ~n1681;
  assign n2247 = ~n2245 & ~n2246;
  assign n2248 = n1663 & n1702;
  assign n2249 = ~n1697 & ~n1722;
  assign n2250 = n1703 & n2249;
  assign n2251 = n1691 & n2250;
  assign n2252 = ~n1686 & n2251;
  assign n2253 = n1684 & ~n2252;
  assign n2254 = ~n2248 & ~n2253;
  assign n2255 = n2247 & n2254;
  assign n2256 = n1695 & ~n1711;
  assign n2257 = ~n1675 & n1722;
  assign n2258 = n1663 & n1718;
  assign n2259 = ~n1706 & n1719;
  assign n2260 = n1674 & ~n2259;
  assign n2261 = ~n2258 & ~n2260;
  assign n2262 = ~n2257 & n2261;
  assign n2263 = ~n1934 & n2262;
  assign n2264 = ~n1662 & ~n1687;
  assign n2265 = n2263 & ~n2264;
  assign n2266 = ~n2256 & n2265;
  assign n2267 = n2255 & n2266;
  assign n2268 = ~n1708 & n2267;
  assign n2269 = ~n2244 & n2268;
  assign n2270 = n2269 ^ x29;
  assign n2271 = n2270 ^ x143;
  assign n2272 = n1060 & ~n1098;
  assign n2273 = ~n1088 & ~n1102;
  assign n2274 = n1100 & ~n2273;
  assign n2275 = n1061 & ~n1105;
  assign n2276 = n1464 & n1480;
  assign n2277 = ~n1067 & n2276;
  assign n2278 = n1081 & ~n2277;
  assign n2279 = ~n2275 & ~n2278;
  assign n2280 = ~n1058 & n1084;
  assign n2281 = ~n1476 & n2280;
  assign n2282 = n1100 & ~n2281;
  assign n2283 = n1094 & n1871;
  assign n2284 = ~n1102 & n2283;
  assign n2285 = n1065 & ~n2284;
  assign n2286 = ~n2282 & ~n2285;
  assign n2287 = n2279 & n2286;
  assign n2288 = ~n2274 & n2287;
  assign n2289 = ~n2272 & n2288;
  assign n2290 = ~n1885 & n2289;
  assign n2291 = n1475 & n2290;
  assign n2292 = ~n1073 & n2291;
  assign n2293 = ~n1089 & n2292;
  assign n2294 = n2293 ^ x13;
  assign n2295 = n2294 ^ x145;
  assign n2296 = n2271 & ~n2295;
  assign n2297 = n1395 & n1401;
  assign n2298 = n1406 & n1433;
  assign n2299 = ~n2297 & ~n2298;
  assign n2300 = ~n1398 & n1434;
  assign n2301 = n1402 & n1426;
  assign n2302 = ~n2300 & ~n2301;
  assign n2303 = n2299 & n2302;
  assign n2304 = ~n1400 & n1435;
  assign n2305 = n1397 & n1400;
  assign n2306 = ~n1402 & n1440;
  assign n2307 = ~n1395 & ~n1434;
  assign n2308 = n1400 & ~n2307;
  assign n2309 = ~n2306 & ~n2308;
  assign n2310 = n1402 & n1642;
  assign n2311 = n1421 & n1430;
  assign n2312 = n1401 & ~n2311;
  assign n2313 = ~n2310 & ~n2312;
  assign n2314 = n2309 & n2313;
  assign n2315 = n1631 & n2314;
  assign n2316 = n1411 & n2315;
  assign n2317 = ~n2305 & n2316;
  assign n2318 = ~n2304 & n2317;
  assign n2319 = n2303 & n2318;
  assign n2320 = n1423 & n2319;
  assign n2321 = n2320 ^ x5;
  assign n2322 = n2321 ^ x146;
  assign n2323 = n1124 & n1150;
  assign n2324 = n1135 & n1163;
  assign n2325 = ~n2323 & ~n2324;
  assign n2326 = ~n1158 & ~n1167;
  assign n2327 = n1160 & ~n2326;
  assign n2328 = ~n1138 & ~n1172;
  assign n2329 = n1159 & ~n2328;
  assign n2330 = ~n2327 & ~n2329;
  assign n2331 = ~n1167 & ~n1509;
  assign n2332 = n1126 & ~n2331;
  assign n2333 = ~n1142 & ~n1186;
  assign n2334 = n1170 & ~n2333;
  assign n2335 = ~n1144 & ~n1159;
  assign n2336 = ~n1158 & ~n1163;
  assign n2337 = ~n1126 & n2336;
  assign n2338 = ~n2335 & ~n2337;
  assign n2339 = ~n1747 & ~n2338;
  assign n2340 = ~n1160 & ~n2339;
  assign n2341 = ~n2334 & ~n2340;
  assign n2342 = ~n2332 & n2341;
  assign n2343 = n2330 & n2342;
  assign n2344 = n2325 & n2343;
  assign n2345 = ~n1146 & n2344;
  assign n2346 = n1500 & n2345;
  assign n2347 = n1742 & n2346;
  assign n2348 = ~n1498 & n2347;
  assign n2349 = n1140 & n2348;
  assign n2350 = n2349 ^ x21;
  assign n2351 = n2350 ^ x144;
  assign n2352 = n2322 & ~n2351;
  assign n2353 = n2296 & n2352;
  assign n2354 = n2271 & n2295;
  assign n2355 = ~n2322 & ~n2351;
  assign n2356 = n2354 & n2355;
  assign n2357 = ~n2353 & ~n2356;
  assign n2358 = n2242 & ~n2357;
  assign n2359 = ~n2271 & n2295;
  assign n2360 = n2355 & n2359;
  assign n2361 = n2242 & n2360;
  assign n2362 = n2216 & ~n2241;
  assign n2363 = ~n2271 & ~n2295;
  assign n2364 = ~n2322 & n2351;
  assign n2365 = n2363 & n2364;
  assign n2366 = n2362 & n2365;
  assign n2367 = n2216 & n2241;
  assign n2368 = ~n2216 & ~n2241;
  assign n2369 = ~n2367 & ~n2368;
  assign n2370 = n2355 & n2363;
  assign n2371 = ~n2369 & n2370;
  assign n2372 = ~n2366 & ~n2371;
  assign n2373 = ~n2361 & n2372;
  assign n2374 = n2354 & n2364;
  assign n2375 = n2367 & n2374;
  assign n2376 = n2322 & n2351;
  assign n2377 = n2363 & n2376;
  assign n2378 = ~n2369 & n2377;
  assign n2379 = ~n2375 & ~n2378;
  assign n2380 = ~n2353 & ~n2374;
  assign n2381 = n2368 & ~n2380;
  assign n2382 = n2296 & n2376;
  assign n2383 = n2242 & n2382;
  assign n2384 = n2368 & n2382;
  assign n2385 = n2352 & n2359;
  assign n2386 = ~n2370 & ~n2385;
  assign n2387 = ~n2377 & n2386;
  assign n2388 = ~n2374 & n2387;
  assign n2389 = n2242 & ~n2388;
  assign n2390 = ~n2384 & ~n2389;
  assign n2391 = n2359 & n2376;
  assign n2392 = ~n2241 & n2391;
  assign n2393 = n2359 & n2364;
  assign n2394 = ~n2385 & ~n2393;
  assign n2395 = n2296 & n2364;
  assign n2396 = n2296 & n2355;
  assign n2397 = ~n2395 & ~n2396;
  assign n2398 = n2357 & n2397;
  assign n2399 = n2394 & n2398;
  assign n2400 = n2362 & ~n2399;
  assign n2401 = n2352 & n2363;
  assign n2402 = ~n2360 & ~n2401;
  assign n2403 = ~n2395 & n2402;
  assign n2404 = n2367 & ~n2403;
  assign n2405 = n2352 & n2354;
  assign n2406 = n2354 & n2376;
  assign n2407 = n2367 & n2406;
  assign n2408 = n2356 & n2368;
  assign n2409 = ~n2407 & ~n2408;
  assign n2410 = ~n2405 & n2409;
  assign n2411 = ~n2369 & ~n2410;
  assign n2412 = ~n2404 & ~n2411;
  assign n2413 = ~n2400 & n2412;
  assign n2414 = ~n2392 & n2413;
  assign n2415 = n2390 & n2414;
  assign n2416 = ~n2383 & n2415;
  assign n2417 = ~n2381 & n2416;
  assign n2418 = n2379 & n2417;
  assign n2419 = n2373 & n2418;
  assign n2420 = ~n2358 & n2419;
  assign n2421 = n2420 ^ x44;
  assign n2422 = n2421 ^ x187;
  assign n2423 = ~n1869 & n2182;
  assign n2424 = n2051 & n2423;
  assign n2425 = n2422 & n2424;
  assign n2426 = ~n2182 & n2422;
  assign n2427 = ~n2051 & n2426;
  assign n2428 = n1869 & n2427;
  assign n2429 = n1869 & n2051;
  assign n2430 = ~n2182 & n2429;
  assign n2431 = ~n2422 & n2430;
  assign n2432 = ~n2428 & ~n2431;
  assign n2433 = ~n2425 & n2432;
  assign n2434 = n2186 & ~n2433;
  assign n2435 = ~n2185 & ~n2434;
  assign n2436 = ~n1869 & n2427;
  assign n2437 = ~n1628 & ~n2186;
  assign n2438 = n2436 & ~n2437;
  assign n2439 = n1346 & n1627;
  assign n2440 = ~n2422 & n2424;
  assign n2441 = ~n2051 & ~n2422;
  assign n2442 = n2423 & n2441;
  assign n2443 = ~n2051 & n2182;
  assign n2444 = n1869 & n2443;
  assign n2445 = n2422 & n2444;
  assign n2446 = n2182 & n2429;
  assign n2447 = ~n2422 & n2446;
  assign n2448 = ~n2445 & ~n2447;
  assign n2449 = ~n2442 & n2448;
  assign n2450 = ~n2440 & n2449;
  assign n2451 = n2439 & ~n2450;
  assign n2452 = ~n2438 & ~n2451;
  assign n2453 = n2435 & n2452;
  assign n2454 = ~n1346 & n2428;
  assign n2455 = ~n1346 & ~n1627;
  assign n2456 = ~n2182 & n2441;
  assign n2457 = n1869 & n2456;
  assign n2458 = n2426 & n2429;
  assign n2459 = ~n1869 & n2456;
  assign n2460 = ~n2458 & ~n2459;
  assign n2461 = ~n2457 & n2460;
  assign n2462 = n2455 & ~n2461;
  assign n2463 = n1628 & n2457;
  assign n2464 = ~n2439 & ~n2463;
  assign n2465 = n2051 & n2426;
  assign n2466 = ~n1869 & n2465;
  assign n2467 = ~n2436 & ~n2459;
  assign n2468 = ~n2463 & n2467;
  assign n2469 = ~n2466 & n2468;
  assign n2470 = ~n2431 & n2469;
  assign n2471 = ~n2464 & ~n2470;
  assign n2472 = ~n2051 & n2423;
  assign n2473 = n2422 & n2472;
  assign n2474 = n2422 & n2446;
  assign n2475 = ~n2442 & ~n2474;
  assign n2476 = ~n2473 & n2475;
  assign n2477 = n1628 & ~n2476;
  assign n2478 = ~n2186 & ~n2455;
  assign n2479 = n2182 & n2441;
  assign n2480 = n1869 & n2479;
  assign n2481 = n2475 & ~n2480;
  assign n2482 = ~n2447 & n2481;
  assign n2483 = ~n2455 & n2482;
  assign n2484 = ~n2440 & ~n2480;
  assign n2485 = ~n2425 & n2484;
  assign n2486 = ~n2473 & n2485;
  assign n2487 = ~n2186 & n2486;
  assign n2488 = ~n2483 & ~n2487;
  assign n2489 = ~n2478 & n2488;
  assign n2490 = ~n2477 & ~n2489;
  assign n2491 = ~n2471 & n2490;
  assign n2492 = ~n2462 & n2491;
  assign n2493 = ~n2454 & n2492;
  assign n2494 = n2453 & n2493;
  assign n2495 = n2494 ^ n987;
  assign n2496 = n2495 ^ x220;
  assign n2497 = n2110 & n2112;
  assign n2498 = n2122 & n2132;
  assign n2499 = n2054 & ~n2156;
  assign n2500 = ~n2498 & ~n2499;
  assign n2501 = ~n2497 & n2500;
  assign n2502 = n2122 & n2141;
  assign n2503 = n2125 & n2132;
  assign n2504 = ~n2502 & ~n2503;
  assign n2505 = n2115 & n2132;
  assign n2506 = n2054 & n2158;
  assign n2507 = n2145 & ~n2506;
  assign n2508 = ~n2505 & n2507;
  assign n2509 = n2054 & n2146;
  assign n2510 = ~n2137 & ~n2146;
  assign n2511 = n2167 & n2510;
  assign n2512 = n2141 & ~n2511;
  assign n2513 = ~n2509 & ~n2512;
  assign n2514 = ~n2130 & n2160;
  assign n2515 = n2132 & ~n2514;
  assign n2516 = ~n2134 & n2152;
  assign n2517 = n2112 & ~n2516;
  assign n2518 = ~n2515 & ~n2517;
  assign n2519 = n2513 & n2518;
  assign n2520 = ~n2121 & n2519;
  assign n2521 = n2140 & n2520;
  assign n2522 = n2508 & n2521;
  assign n2523 = n2504 & n2522;
  assign n2524 = n2501 & n2523;
  assign n2525 = ~n2163 & n2524;
  assign n2526 = n2117 & n2525;
  assign n2527 = ~n2124 & n2526;
  assign n2528 = n2527 ^ x58;
  assign n2529 = n2528 ^ x171;
  assign n2530 = n2242 & n2370;
  assign n2531 = ~n2381 & ~n2530;
  assign n2532 = n2362 & n2405;
  assign n2533 = n2353 & n2367;
  assign n2534 = ~n2532 & ~n2533;
  assign n2535 = ~n2374 & ~n2396;
  assign n2536 = n2216 & ~n2535;
  assign n2537 = ~n2356 & n2397;
  assign n2538 = ~n2362 & n2537;
  assign n2539 = ~n2242 & ~n2362;
  assign n2540 = ~n2391 & ~n2395;
  assign n2541 = ~n2242 & n2540;
  assign n2542 = ~n2539 & ~n2541;
  assign n2543 = n2362 & ~n2386;
  assign n2544 = ~n2542 & ~n2543;
  assign n2545 = ~n2538 & ~n2544;
  assign n2546 = ~n2536 & ~n2545;
  assign n2547 = ~n2391 & n2394;
  assign n2548 = n2242 & ~n2547;
  assign n2549 = n2351 ^ n2322;
  assign n2550 = n2363 & n2549;
  assign n2551 = ~n2393 & ~n2550;
  assign n2552 = ~n2368 & n2551;
  assign n2553 = ~n2367 & n2403;
  assign n2554 = ~n2552 & ~n2553;
  assign n2555 = ~n2377 & ~n2554;
  assign n2556 = ~n2406 & n2555;
  assign n2557 = ~n2369 & ~n2556;
  assign n2558 = ~n2548 & ~n2557;
  assign n2559 = n2546 & n2558;
  assign n2560 = n2534 & n2559;
  assign n2561 = ~n2408 & n2560;
  assign n2562 = n2531 & n2561;
  assign n2563 = n2241 ^ n2216;
  assign n2564 = n2382 & n2563;
  assign n2565 = n2562 & ~n2564;
  assign n2566 = n2565 ^ x32;
  assign n2567 = n2566 ^ x166;
  assign n2568 = n2529 & ~n2567;
  assign n2569 = n2270 ^ x141;
  assign n2570 = n1930 ^ x136;
  assign n2571 = ~n2569 & ~n2570;
  assign n2572 = n2215 ^ x140;
  assign n2573 = n855 & ~n1363;
  assign n2574 = n834 & n847;
  assign n2575 = ~n2573 & ~n2574;
  assign n2576 = n864 & ~n874;
  assign n2577 = n835 & ~n2576;
  assign n2578 = n878 & ~n1362;
  assign n2579 = n858 & ~n2578;
  assign n2580 = ~n2577 & ~n2579;
  assign n2581 = n851 & ~n853;
  assign n2582 = n860 & ~n2581;
  assign n2583 = ~n861 & n2073;
  assign n2584 = n844 & ~n2583;
  assign n2585 = ~n2582 & ~n2584;
  assign n2586 = n2580 & n2585;
  assign n2587 = n2575 & n2586;
  assign n2588 = n2060 & n2587;
  assign n2589 = n1361 & n2588;
  assign n2590 = n867 & n2589;
  assign n2591 = ~n843 & n2590;
  assign n2592 = n2591 ^ x53;
  assign n2593 = n2592 ^ x138;
  assign n2594 = n2572 & n2593;
  assign n2595 = ~n1201 & n1217;
  assign n2596 = n1202 & ~n1530;
  assign n2597 = ~n2595 & ~n2596;
  assign n2598 = n1222 & n1236;
  assign n2599 = ~n1223 & ~n1238;
  assign n2600 = n1230 & ~n2599;
  assign n2601 = ~n1248 & n1777;
  assign n2602 = ~n1225 & n2601;
  assign n2603 = n1219 & n2602;
  assign n2604 = n1239 & n2603;
  assign n2605 = ~n1244 & n2604;
  assign n2606 = ~n1256 & n1262;
  assign n2607 = ~n1787 & ~n2606;
  assign n2608 = n1255 & ~n2607;
  assign n2609 = ~n2605 & ~n2608;
  assign n2610 = ~n2600 & ~n2609;
  assign n2611 = ~n2598 & n2610;
  assign n2612 = n2597 & n2611;
  assign n2613 = ~n1221 & n2612;
  assign n2614 = n1525 & n2613;
  assign n2615 = n2614 ^ x45;
  assign n2616 = n2615 ^ x139;
  assign n2617 = n1899 ^ x137;
  assign n2618 = ~n2616 & n2617;
  assign n2619 = n2594 & n2618;
  assign n2620 = ~n2572 & ~n2593;
  assign n2621 = n2618 & n2620;
  assign n2622 = ~n2619 & ~n2621;
  assign n2623 = n2571 & ~n2622;
  assign n2624 = ~n2569 & n2570;
  assign n2625 = ~n2572 & n2593;
  assign n2626 = n2618 & n2625;
  assign n2627 = n2572 & ~n2593;
  assign n2628 = n2618 & n2627;
  assign n2629 = ~n2626 & ~n2628;
  assign n2630 = n2624 & ~n2629;
  assign n2631 = ~n2623 & ~n2630;
  assign n2632 = n2569 & ~n2570;
  assign n2633 = ~n2616 & ~n2617;
  assign n2634 = n2620 & n2633;
  assign n2635 = n2616 & ~n2617;
  assign n2636 = n2627 & n2635;
  assign n2637 = ~n2634 & ~n2636;
  assign n2638 = n2632 & ~n2637;
  assign n2639 = n2569 & n2570;
  assign n2640 = n2625 & n2633;
  assign n2641 = n2639 & n2640;
  assign n2642 = n2616 & n2617;
  assign n2643 = n2627 & n2642;
  assign n2644 = n2571 & n2643;
  assign n2645 = n2625 & n2642;
  assign n2646 = ~n2619 & ~n2645;
  assign n2647 = n2624 & ~n2646;
  assign n2648 = ~n2644 & ~n2647;
  assign n2649 = ~n2641 & n2648;
  assign n2650 = ~n2638 & n2649;
  assign n2651 = n2594 & n2633;
  assign n2652 = n2632 & n2651;
  assign n2653 = n2594 & n2635;
  assign n2654 = ~n2651 & ~n2653;
  assign n2655 = n2571 & ~n2654;
  assign n2656 = ~n2652 & ~n2655;
  assign n2657 = n2632 & n2643;
  assign n2658 = n2636 & n2639;
  assign n2659 = ~n2657 & ~n2658;
  assign n2660 = n2625 & n2635;
  assign n2661 = n2627 & n2633;
  assign n2662 = ~n2660 & ~n2661;
  assign n2663 = n2571 & ~n2662;
  assign n2664 = n2620 & n2635;
  assign n2665 = ~n2653 & ~n2664;
  assign n2666 = ~n2628 & n2665;
  assign n2667 = ~n2645 & n2666;
  assign n2668 = n2632 & ~n2667;
  assign n2669 = ~n2663 & ~n2668;
  assign n2670 = n2620 & n2642;
  assign n2671 = ~n2569 & n2670;
  assign n2672 = ~n2640 & ~n2653;
  assign n2673 = ~n2636 & n2672;
  assign n2674 = n2624 & ~n2673;
  assign n2675 = n2594 & n2642;
  assign n2676 = n2629 & ~n2675;
  assign n2677 = ~n2621 & n2676;
  assign n2678 = ~n2664 & n2677;
  assign n2679 = ~n2661 & n2678;
  assign n2680 = n2639 & ~n2679;
  assign n2681 = ~n2674 & ~n2680;
  assign n2682 = ~n2671 & n2681;
  assign n2683 = n2669 & n2682;
  assign n2684 = n2659 & n2683;
  assign n2685 = n2656 & n2684;
  assign n2686 = n2650 & n2685;
  assign n2687 = n2631 & n2686;
  assign n2688 = n2687 ^ x0;
  assign n2689 = n2688 ^ x170;
  assign n2690 = n1561 & n1581;
  assign n2691 = ~n1356 & n1558;
  assign n2692 = n1556 & n1568;
  assign n2693 = ~n2691 & ~n2692;
  assign n2694 = ~n2690 & n2693;
  assign n2695 = ~n1590 & ~n1603;
  assign n2696 = n1564 & ~n2695;
  assign n2697 = n1388 & n1568;
  assign n2698 = n1581 & ~n1613;
  assign n2699 = ~n2697 & ~n2698;
  assign n2700 = n1388 & n1603;
  assign n2701 = ~n1387 & ~n1591;
  assign n2702 = ~n2700 & ~n2701;
  assign n2703 = ~n1356 & ~n1608;
  assign n2704 = ~n1568 & ~n1607;
  assign n2705 = ~n1558 & n2704;
  assign n2706 = n1613 & n2705;
  assign n2707 = n1564 & ~n2706;
  assign n2708 = ~n1554 & n1599;
  assign n2709 = ~n1561 & n2708;
  assign n2710 = n1556 & ~n2709;
  assign n2711 = ~n2707 & ~n2710;
  assign n2712 = ~n2703 & n2711;
  assign n2713 = n2702 & n2712;
  assign n2714 = n2699 & n2713;
  assign n2715 = ~n2696 & n2714;
  assign n2716 = n1580 & n2715;
  assign n2717 = n2694 & n2716;
  assign n2718 = ~n1555 & n2717;
  assign n2719 = n2718 ^ x24;
  assign n2720 = n2719 ^ x167;
  assign n2721 = ~n2689 & n2720;
  assign n2722 = n1037 & ~n2211;
  assign n2723 = n992 & ~n2192;
  assign n2724 = ~n2722 & ~n2723;
  assign n2725 = n1018 & n2198;
  assign n2726 = n1027 & ~n2204;
  assign n2727 = ~n2725 & ~n2726;
  assign n2728 = n2724 & n2727;
  assign n2729 = n2728 ^ x55;
  assign n2730 = n2729 ^ x150;
  assign n2731 = n1386 ^ x152;
  assign n2732 = n2730 & ~n2731;
  assign n2733 = n2240 ^ x149;
  assign n2734 = n1674 & ~n2249;
  assign n2735 = n1665 ^ n1664;
  assign n2736 = n1696 & n2735;
  assign n2737 = n1681 & ~n2736;
  assign n2738 = ~n1689 & n2737;
  assign n2739 = ~n1699 & n2738;
  assign n2740 = n1695 & ~n2739;
  assign n2741 = ~n2734 & ~n2740;
  assign n2742 = ~n1675 & ~n1941;
  assign n2743 = n1711 & n1719;
  assign n2744 = n1684 & ~n2743;
  assign n2745 = n1687 & ~n1690;
  assign n2746 = ~n1713 & n2745;
  assign n2747 = n1674 & ~n2746;
  assign n2748 = n1663 & n1678;
  assign n2749 = ~n1688 & ~n2748;
  assign n2750 = n1691 & n2749;
  assign n2751 = n1662 & ~n2750;
  assign n2752 = ~n2747 & ~n2751;
  assign n2753 = ~n2744 & n2752;
  assign n2754 = ~n2742 & n2753;
  assign n2755 = n2741 & n2754;
  assign n2756 = ~n2244 & n2755;
  assign n2757 = ~n1671 & n2756;
  assign n2758 = ~n1934 & n2757;
  assign n2759 = n2758 ^ x47;
  assign n2760 = n2759 ^ x151;
  assign n2761 = n2733 & ~n2760;
  assign n2762 = n2732 & n2761;
  assign n2763 = n2321 ^ x148;
  assign n2764 = n1551 ^ x153;
  assign n2765 = n2763 & n2764;
  assign n2766 = n2762 & n2765;
  assign n2767 = ~n2733 & n2760;
  assign n2768 = ~n2730 & ~n2731;
  assign n2769 = n2767 & n2768;
  assign n2770 = ~n2763 & n2764;
  assign n2771 = n2769 & n2770;
  assign n2772 = ~n2766 & ~n2771;
  assign n2773 = ~n2730 & n2731;
  assign n2774 = n2761 & n2773;
  assign n2775 = n2733 & n2760;
  assign n2776 = n2732 & n2775;
  assign n2777 = ~n2774 & ~n2776;
  assign n2778 = n2770 & ~n2777;
  assign n2779 = n2768 & n2775;
  assign n2780 = ~n2774 & ~n2779;
  assign n2781 = ~n2769 & n2780;
  assign n2782 = n2763 & ~n2764;
  assign n2783 = ~n2781 & n2782;
  assign n2784 = ~n2778 & ~n2783;
  assign n2785 = n2730 & n2731;
  assign n2786 = n2761 & n2785;
  assign n2787 = ~n2763 & ~n2764;
  assign n2788 = n2786 & ~n2787;
  assign n2789 = ~n2733 & ~n2760;
  assign n2790 = n2785 & n2789;
  assign n2791 = n2767 & n2773;
  assign n2792 = n2768 & n2789;
  assign n2793 = ~n2791 & ~n2792;
  assign n2794 = ~n2790 & n2793;
  assign n2795 = ~n2762 & n2794;
  assign n2796 = n2787 & ~n2795;
  assign n2797 = n2773 & n2789;
  assign n2798 = n2767 & n2785;
  assign n2799 = n2732 & n2767;
  assign n2800 = n2732 & n2789;
  assign n2801 = ~n2799 & ~n2800;
  assign n2802 = ~n2798 & n2801;
  assign n2803 = ~n2797 & n2802;
  assign n2804 = ~n2770 & ~n2782;
  assign n2805 = ~n2803 & ~n2804;
  assign n2806 = n2775 & n2785;
  assign n2807 = n2761 & n2768;
  assign n2808 = ~n2806 & ~n2807;
  assign n2809 = n2773 & n2775;
  assign n2810 = ~n2776 & ~n2809;
  assign n2811 = n2808 & n2810;
  assign n2812 = n2787 & ~n2811;
  assign n2813 = n2733 ^ n2730;
  assign n2814 = n2813 ^ n2731;
  assign n2815 = n2814 ^ n2760;
  assign n2816 = n2761 & ~n2815;
  assign n2817 = n2816 ^ n2815;
  assign n2818 = n2765 & ~n2817;
  assign n2819 = ~n2812 & ~n2818;
  assign n2820 = ~n2805 & n2819;
  assign n2821 = ~n2796 & n2820;
  assign n2822 = ~n2788 & n2821;
  assign n2823 = n2784 & n2822;
  assign n2824 = n2772 & n2823;
  assign n2825 = n2824 ^ x8;
  assign n2826 = n2825 ^ x169;
  assign n2827 = n989 & n1332;
  assign n2828 = n1283 & n1288;
  assign n2829 = n989 & n1325;
  assign n2830 = ~n1295 & ~n1306;
  assign n2831 = n1284 & ~n2830;
  assign n2832 = ~n2829 & ~n2831;
  assign n2833 = ~n2828 & n2832;
  assign n2834 = ~n2827 & n2833;
  assign n2835 = n1288 & n1301;
  assign n2836 = ~n1279 & ~n1312;
  assign n2837 = n1285 & ~n2836;
  assign n2838 = ~n2835 & ~n2837;
  assign n2839 = n989 & ~n1313;
  assign n2840 = ~n1310 & n1328;
  assign n2841 = ~n1290 & n2840;
  assign n2842 = n1284 & ~n2841;
  assign n2843 = n1288 & ~n2836;
  assign n2844 = ~n1318 & ~n1332;
  assign n2845 = ~n1309 & ~n1327;
  assign n2846 = n2844 & n2845;
  assign n2847 = n1285 & ~n2846;
  assign n2848 = ~n1318 & ~n1323;
  assign n2849 = ~n1288 & n2848;
  assign n2850 = ~n1334 & ~n2849;
  assign n2851 = ~n1309 & ~n2850;
  assign n2852 = n1286 & ~n2851;
  assign n2853 = ~n2847 & ~n2852;
  assign n2854 = ~n2843 & n2853;
  assign n2855 = ~n2842 & n2854;
  assign n2856 = ~n2839 & n2855;
  assign n2857 = n2838 & n2856;
  assign n2858 = n1299 & n2857;
  assign n2859 = n2834 & n2858;
  assign n2860 = ~n1280 & n2859;
  assign n2861 = n2860 ^ x16;
  assign n2862 = n2861 ^ x168;
  assign n2863 = n2826 & n2862;
  assign n2864 = n2721 & n2863;
  assign n2865 = n2568 & n2864;
  assign n2866 = ~n2529 & ~n2567;
  assign n2867 = ~n2689 & ~n2720;
  assign n2868 = n2863 & n2867;
  assign n2869 = n2866 & n2868;
  assign n2870 = n2529 & n2567;
  assign n2871 = ~n2826 & ~n2862;
  assign n2872 = n2867 & n2871;
  assign n2873 = n2870 & n2872;
  assign n2874 = ~n2869 & ~n2873;
  assign n2875 = ~n2865 & n2874;
  assign n2876 = ~n2826 & n2862;
  assign n2877 = n2867 & n2876;
  assign n2878 = n2870 & n2877;
  assign n2879 = n2721 & n2871;
  assign n2880 = n2568 & n2879;
  assign n2881 = ~n2878 & ~n2880;
  assign n2882 = n2689 & n2720;
  assign n2883 = n2826 & ~n2862;
  assign n2884 = n2882 & n2883;
  assign n2885 = n2568 & n2884;
  assign n2886 = ~n2529 & n2567;
  assign n2887 = n2689 & ~n2720;
  assign n2888 = n2863 & n2887;
  assign n2889 = n2867 & n2883;
  assign n2890 = ~n2888 & ~n2889;
  assign n2891 = n2886 & ~n2890;
  assign n2892 = ~n2885 & ~n2891;
  assign n2893 = n2720 & n2876;
  assign n2894 = n2689 & n2893;
  assign n2895 = n2568 & n2894;
  assign n2896 = n2866 & n2872;
  assign n2897 = ~n2895 & ~n2896;
  assign n2898 = n2876 & n2887;
  assign n2899 = ~n2872 & ~n2898;
  assign n2900 = n2886 & ~n2899;
  assign n2901 = n2871 & n2882;
  assign n2902 = n2886 & n2901;
  assign n2903 = n2866 & n2901;
  assign n2904 = n2870 & n2884;
  assign n2905 = ~n2903 & ~n2904;
  assign n2906 = ~n2866 & ~n2870;
  assign n2907 = n2883 & n2887;
  assign n2908 = n2871 & n2887;
  assign n2909 = n2721 & n2883;
  assign n2910 = ~n2894 & ~n2909;
  assign n2911 = ~n2908 & n2910;
  assign n2912 = ~n2907 & n2911;
  assign n2913 = ~n2864 & n2912;
  assign n2914 = ~n2906 & ~n2913;
  assign n2915 = n2863 & n2882;
  assign n2916 = n2886 & n2915;
  assign n2917 = n2568 & n2898;
  assign n2918 = ~n2916 & ~n2917;
  assign n2919 = ~n2689 & n2893;
  assign n2920 = ~n2909 & ~n2919;
  assign n2921 = n2886 & ~n2920;
  assign n2922 = ~n2877 & n2890;
  assign n2923 = n2568 & ~n2922;
  assign n2924 = ~n2921 & ~n2923;
  assign n2925 = n2918 & n2924;
  assign n2926 = ~n2914 & n2925;
  assign n2927 = n2905 & n2926;
  assign n2928 = ~n2902 & n2927;
  assign n2929 = ~n2900 & n2928;
  assign n2930 = n2897 & n2929;
  assign n2931 = n2892 & n2930;
  assign n2932 = n2881 & n2931;
  assign n2933 = n2875 & n2932;
  assign n2934 = n2933 ^ n907;
  assign n2935 = n2934 ^ x225;
  assign n2936 = n2496 & n2935;
  assign n2937 = n2356 & n2362;
  assign n2938 = ~n2543 & ~n2937;
  assign n2939 = n2367 & n2395;
  assign n2940 = ~n2365 & ~n2391;
  assign n2941 = n2242 & ~n2940;
  assign n2942 = ~n2939 & ~n2941;
  assign n2943 = n2242 & n2405;
  assign n2944 = n2396 & ~n2539;
  assign n2945 = ~n2943 & ~n2944;
  assign n2946 = ~n2241 & n2401;
  assign n2947 = ~n2369 & ~n2394;
  assign n2948 = ~n2357 & n2367;
  assign n2949 = ~n2947 & ~n2948;
  assign n2950 = ~n2946 & n2949;
  assign n2951 = n2362 & n2406;
  assign n2952 = ~n2374 & ~n2405;
  assign n2953 = ~n2395 & n2952;
  assign n2954 = n2368 & ~n2953;
  assign n2955 = ~n2951 & ~n2954;
  assign n2956 = n2950 & n2955;
  assign n2957 = n2945 & n2956;
  assign n2958 = n2379 & n2957;
  assign n2959 = n2942 & n2958;
  assign n2960 = ~n2564 & n2959;
  assign n2961 = n2938 & n2960;
  assign n2962 = n2373 & n2961;
  assign n2963 = ~n2358 & n2962;
  assign n2964 = n2963 ^ x30;
  assign n2965 = n2964 ^ x201;
  assign n2966 = ~n1285 & n1332;
  assign n2967 = ~n1286 & ~n2848;
  assign n2968 = ~n2966 & ~n2967;
  assign n2969 = n1286 & n1310;
  assign n2970 = ~n1306 & ~n1325;
  assign n2971 = n1285 & ~n2970;
  assign n2972 = ~n2969 & ~n2971;
  assign n2973 = ~n1309 & ~n1326;
  assign n2974 = n1284 & ~n2973;
  assign n2975 = ~n1278 & ~n1311;
  assign n2976 = ~n1288 & n2975;
  assign n2977 = ~n1292 & ~n1309;
  assign n2978 = n989 & ~n2977;
  assign n2979 = n1329 & ~n2978;
  assign n2980 = ~n2976 & ~n2979;
  assign n2981 = n1286 & n2980;
  assign n2982 = ~n2974 & ~n2981;
  assign n2983 = n2972 & n2982;
  assign n2984 = n2968 & n2983;
  assign n2985 = n1304 & n2984;
  assign n2986 = n2838 & n2985;
  assign n2987 = n1298 & n2986;
  assign n2988 = n2833 & n2987;
  assign n2989 = n2988 ^ x4;
  assign n2990 = n2989 ^ x196;
  assign n2991 = n2965 & n2990;
  assign n2992 = n2624 & n2643;
  assign n2993 = n2639 & ~n2662;
  assign n2994 = ~n2992 & ~n2993;
  assign n2995 = ~n2660 & n2677;
  assign n2996 = n2632 & ~n2995;
  assign n2997 = ~n2670 & ~n2675;
  assign n2998 = ~n2626 & n2997;
  assign n2999 = ~n2643 & n2998;
  assign n3000 = ~n2651 & n2999;
  assign n3001 = n2639 & ~n3000;
  assign n3002 = ~n2996 & ~n3001;
  assign n3003 = n2629 & ~n2664;
  assign n3004 = ~n2634 & n3003;
  assign n3005 = ~n2621 & n3004;
  assign n3006 = n2571 & ~n3005;
  assign n3007 = n2637 & n2997;
  assign n3008 = ~n2661 & n3007;
  assign n3009 = n2624 & ~n3008;
  assign n3010 = ~n3006 & ~n3009;
  assign n3011 = n3002 & n3010;
  assign n3012 = n2994 & n3011;
  assign n3013 = n2656 & n3012;
  assign n3014 = n2650 & n3013;
  assign n3015 = n3014 ^ x62;
  assign n3016 = n3015 ^ x197;
  assign n3017 = n1522 & n1559;
  assign n3018 = ~n1566 & ~n3017;
  assign n3019 = ~n1603 & n3018;
  assign n3020 = n1556 & ~n3019;
  assign n3021 = ~n1554 & ~n1573;
  assign n3022 = ~n1597 & n3021;
  assign n3023 = n1581 & ~n3022;
  assign n3024 = ~n3020 & ~n3023;
  assign n3025 = n1588 & ~n1590;
  assign n3026 = n1564 & ~n3025;
  assign n3027 = ~n1596 & ~n1612;
  assign n3028 = ~n1602 & ~n3027;
  assign n3029 = n1608 & n1613;
  assign n3030 = n1388 & ~n3029;
  assign n3031 = ~n3028 & ~n3030;
  assign n3032 = ~n3026 & n3031;
  assign n3033 = n3024 & n3032;
  assign n3034 = n1579 & n3033;
  assign n3035 = n1593 & n3034;
  assign n3036 = ~n1570 & n3035;
  assign n3037 = n1585 & n3036;
  assign n3038 = n2694 & n3037;
  assign n3039 = n3038 ^ x46;
  assign n3040 = n3039 ^ x199;
  assign n3041 = n3016 & n3040;
  assign n3042 = ~n1900 & n2047;
  assign n3043 = n3042 ^ n2046;
  assign n3044 = n3043 ^ x54;
  assign n3045 = n3044 ^ x198;
  assign n3046 = n1809 & ~n1821;
  assign n3047 = ~n1830 & ~n3046;
  assign n3048 = ~n1829 & ~n1836;
  assign n3049 = n1801 & ~n3048;
  assign n3050 = ~n1833 & ~n3049;
  assign n3051 = n1771 & n1799;
  assign n3052 = n1803 & n1834;
  assign n3053 = ~n3051 & ~n3052;
  assign n3054 = n1815 & ~n1852;
  assign n3055 = n1821 & ~n1842;
  assign n3056 = n1801 & ~n3055;
  assign n3057 = ~n1841 & ~n1849;
  assign n3058 = ~n1816 & ~n3057;
  assign n3059 = n1770 & n1813;
  assign n3060 = ~n1842 & ~n3059;
  assign n3061 = ~n1836 & n3060;
  assign n3062 = ~n1834 & n3061;
  assign n3063 = n1809 & ~n3062;
  assign n3064 = ~n3058 & ~n3063;
  assign n3065 = ~n3056 & n3064;
  assign n3066 = n1816 & n1824;
  assign n3067 = n1853 & ~n3059;
  assign n3068 = ~n1820 & n3067;
  assign n3069 = n1803 & ~n3068;
  assign n3070 = ~n3066 & ~n3069;
  assign n3071 = n3065 & n3070;
  assign n3072 = n1818 & n3071;
  assign n3073 = ~n3054 & n3072;
  assign n3074 = n3053 & n3073;
  assign n3075 = n3050 & n3074;
  assign n3076 = n3047 & n3075;
  assign n3077 = n3076 ^ x38;
  assign n3078 = n3077 ^ x200;
  assign n3079 = ~n3045 & ~n3078;
  assign n3080 = n3041 & n3079;
  assign n3081 = ~n3045 & n3078;
  assign n3082 = n3016 & ~n3040;
  assign n3083 = n3081 & n3082;
  assign n3084 = ~n3080 & ~n3083;
  assign n3085 = n2991 & ~n3084;
  assign n3086 = n2965 & ~n2990;
  assign n3087 = n3079 & n3082;
  assign n3088 = n3045 & n3078;
  assign n3089 = n3082 & n3088;
  assign n3090 = ~n3087 & ~n3089;
  assign n3091 = n3086 & ~n3090;
  assign n3092 = ~n3085 & ~n3091;
  assign n3093 = n3045 & ~n3078;
  assign n3094 = n3082 & n3093;
  assign n3095 = ~n2965 & ~n2990;
  assign n3096 = n3094 & n3095;
  assign n3097 = ~n3016 & ~n3040;
  assign n3098 = n3079 & n3097;
  assign n3099 = n2991 & n3098;
  assign n3100 = n3078 ^ n3045;
  assign n3101 = n3041 & n3100;
  assign n3102 = n3095 & n3101;
  assign n3103 = ~n3099 & ~n3102;
  assign n3104 = ~n3016 & n3040;
  assign n3105 = n3081 & n3104;
  assign n3106 = n3086 & n3105;
  assign n3107 = n3083 & n3095;
  assign n3108 = ~n3106 & ~n3107;
  assign n3109 = n3079 & n3104;
  assign n3110 = n3088 & n3097;
  assign n3111 = ~n3109 & ~n3110;
  assign n3112 = n3093 & n3104;
  assign n3113 = n3081 & n3097;
  assign n3114 = ~n3112 & ~n3113;
  assign n3115 = n3111 & n3114;
  assign n3116 = ~n2990 & ~n3115;
  assign n3117 = n3041 & n3093;
  assign n3118 = n3088 & n3104;
  assign n3119 = ~n3094 & ~n3118;
  assign n3120 = n3111 & n3119;
  assign n3121 = ~n3117 & n3120;
  assign n3122 = n2991 & ~n3121;
  assign n3123 = ~n3116 & ~n3122;
  assign n3124 = n3080 & n3086;
  assign n3125 = ~n2965 & n2990;
  assign n3126 = ~n3098 & ~n3118;
  assign n3127 = ~n3110 & n3126;
  assign n3128 = ~n3089 & ~n3117;
  assign n3129 = ~n3105 & n3128;
  assign n3130 = n3127 & n3129;
  assign n3131 = ~n3083 & n3130;
  assign n3132 = ~n3109 & n3131;
  assign n3133 = n3125 & n3132;
  assign n3134 = ~n3124 & ~n3133;
  assign n3135 = n3123 & n3134;
  assign n3136 = n3108 & n3135;
  assign n3137 = n3103 & n3136;
  assign n3138 = ~n3096 & n3137;
  assign n3139 = n3092 & n3138;
  assign n3140 = n3139 ^ n1198;
  assign n3141 = n3140 ^ x224;
  assign n3142 = n2765 & n2776;
  assign n3143 = ~n2786 & ~n2807;
  assign n3144 = n2770 & ~n3143;
  assign n3145 = n2765 & ~n2780;
  assign n3146 = ~n3144 & ~n3145;
  assign n3147 = ~n3142 & n3146;
  assign n3148 = ~n2769 & ~n2790;
  assign n3149 = n2765 & ~n3148;
  assign n3150 = ~n2790 & ~n2799;
  assign n3151 = ~n2762 & n3150;
  assign n3152 = n2787 & ~n3151;
  assign n3153 = ~n3149 & ~n3152;
  assign n3154 = ~n2792 & ~n2798;
  assign n3155 = n2765 & ~n3154;
  assign n3156 = ~n2786 & n2793;
  assign n3157 = n3148 & n3156;
  assign n3158 = n2777 & n3157;
  assign n3159 = ~n2798 & n3158;
  assign n3160 = n2782 & n3159;
  assign n3161 = ~n3155 & ~n3160;
  assign n3162 = ~n2779 & n3150;
  assign n3163 = ~n2791 & n3162;
  assign n3164 = ~n2797 & n3163;
  assign n3165 = n2770 & ~n3164;
  assign n3166 = n2777 & ~n2809;
  assign n3167 = ~n2797 & n3166;
  assign n3168 = ~n2769 & n3167;
  assign n3169 = n2787 & ~n3168;
  assign n3170 = ~n3165 & ~n3169;
  assign n3171 = n3161 & n3170;
  assign n3172 = n2772 & n3171;
  assign n3173 = n3153 & n3172;
  assign n3174 = n3147 & n3173;
  assign n3175 = n3174 ^ x34;
  assign n3176 = n3175 ^ x178;
  assign n3177 = n2181 ^ x183;
  assign n3178 = ~n3176 & n3177;
  assign n3179 = n1345 ^ x182;
  assign n3180 = ~n2622 & n2639;
  assign n3181 = n2632 & ~n2999;
  assign n3182 = ~n3180 & ~n3181;
  assign n3183 = n2571 & n2628;
  assign n3184 = ~n2569 & n2645;
  assign n3185 = ~n3183 & ~n3184;
  assign n3186 = n2570 ^ n2569;
  assign n3187 = n2665 & ~n2670;
  assign n3188 = ~n2640 & n3187;
  assign n3189 = ~n3186 & ~n3188;
  assign n3190 = ~n2634 & ~n2661;
  assign n3191 = ~n2624 & n3190;
  assign n3192 = n2654 & n3191;
  assign n3193 = n2616 ^ n2593;
  assign n3194 = n3193 ^ n2572;
  assign n3195 = ~n2617 & ~n3194;
  assign n3196 = n2624 & n3195;
  assign n3197 = ~n2632 & ~n3196;
  assign n3198 = ~n3192 & ~n3197;
  assign n3199 = ~n3189 & ~n3198;
  assign n3200 = n3185 & n3199;
  assign n3201 = n3182 & n3200;
  assign n3202 = n2994 & n3201;
  assign n3203 = n2631 & n3202;
  assign n3204 = n3203 ^ x18;
  assign n3205 = n3204 ^ x180;
  assign n3206 = n3179 & n3205;
  assign n3207 = n1806 & n1815;
  assign n3208 = n1801 & n1824;
  assign n3209 = ~n3207 & ~n3208;
  assign n3210 = n1799 & n1820;
  assign n3211 = ~n1816 & n1834;
  assign n3212 = ~n3210 & ~n3211;
  assign n3213 = n3209 & n3212;
  assign n3214 = n1803 & n1841;
  assign n3215 = ~n1851 & n3060;
  assign n3216 = ~n1814 & n3215;
  assign n3217 = n1809 & ~n3216;
  assign n3218 = ~n1800 & n1832;
  assign n3219 = n1838 & ~n3218;
  assign n3220 = n1809 & n1849;
  assign n3221 = n1803 & ~n3060;
  assign n3222 = ~n3220 & ~n3221;
  assign n3223 = n1803 & n1814;
  assign n3224 = n1801 & n1850;
  assign n3225 = ~n1771 & ~n1806;
  assign n3226 = n1809 & ~n3225;
  assign n3227 = ~n3224 & ~n3226;
  assign n3228 = ~n3223 & n3227;
  assign n3229 = ~n3054 & n3228;
  assign n3230 = n3050 & n3229;
  assign n3231 = n3222 & n3230;
  assign n3232 = n3219 & n3231;
  assign n3233 = ~n3217 & n3232;
  assign n3234 = ~n3214 & n3233;
  assign n3235 = n3213 & n3234;
  assign n3236 = n1828 & n3235;
  assign n3237 = n3236 ^ x26;
  assign n3238 = n3237 ^ x179;
  assign n3239 = ~n1387 & n1566;
  assign n3240 = n1564 & n1572;
  assign n3241 = ~n1356 & n1596;
  assign n3242 = n1562 & ~n1612;
  assign n3243 = ~n1590 & n3242;
  assign n3244 = ~n1597 & n3243;
  assign n3245 = n1388 & ~n3244;
  assign n3246 = ~n3241 & ~n3245;
  assign n3247 = ~n1496 & n1553;
  assign n3248 = ~n1596 & ~n3247;
  assign n3249 = n1613 & n3248;
  assign n3250 = n1556 & ~n3249;
  assign n3251 = n1591 & ~n1603;
  assign n3252 = ~n1581 & n3251;
  assign n3253 = ~n1575 & ~n2696;
  assign n3254 = n1588 & n3253;
  assign n3255 = ~n3252 & ~n3254;
  assign n3256 = ~n1577 & ~n3255;
  assign n3257 = ~n1602 & ~n3256;
  assign n3258 = ~n3250 & ~n3257;
  assign n3259 = n3246 & n3258;
  assign n3260 = ~n3240 & n3259;
  assign n3261 = ~n3239 & n3260;
  assign n3262 = n1571 & n3261;
  assign n3263 = n2699 & n3262;
  assign n3264 = ~n1555 & n3263;
  assign n3265 = n3264 ^ x10;
  assign n3266 = n3265 ^ x181;
  assign n3267 = n3238 & ~n3266;
  assign n3268 = n3206 & n3267;
  assign n3269 = n3178 & n3268;
  assign n3270 = n3176 & n3177;
  assign n3271 = n3179 & ~n3205;
  assign n3272 = n3266 ^ n3238;
  assign n3273 = n3271 & n3272;
  assign n3274 = n3270 & n3273;
  assign n3275 = ~n3269 & ~n3274;
  assign n3276 = ~n3238 & n3266;
  assign n3277 = n3206 & n3276;
  assign n3278 = n3270 & n3277;
  assign n3279 = ~n3179 & ~n3205;
  assign n3280 = n3238 & n3266;
  assign n3281 = n3279 & n3280;
  assign n3282 = ~n3238 & ~n3266;
  assign n3283 = n3206 & n3282;
  assign n3284 = ~n3281 & ~n3283;
  assign n3285 = n3178 & ~n3284;
  assign n3286 = ~n3278 & ~n3285;
  assign n3287 = ~n3179 & n3267;
  assign n3288 = ~n3179 & n3205;
  assign n3289 = ~n3238 & n3288;
  assign n3290 = ~n3281 & ~n3289;
  assign n3291 = ~n3287 & n3290;
  assign n3292 = n3270 & ~n3291;
  assign n3293 = ~n3238 & n3279;
  assign n3294 = n3280 & n3288;
  assign n3295 = ~n3293 & ~n3294;
  assign n3296 = ~n3273 & n3295;
  assign n3297 = n3178 & ~n3296;
  assign n3298 = ~n3292 & ~n3297;
  assign n3299 = n3176 & ~n3177;
  assign n3300 = ~n3179 & n3282;
  assign n3301 = n3205 ^ n3179;
  assign n3302 = n3280 & n3301;
  assign n3303 = ~n3266 & n3279;
  assign n3304 = ~n3302 & ~n3303;
  assign n3305 = ~n3300 & n3304;
  assign n3306 = ~n3283 & n3305;
  assign n3307 = n3299 & n3306;
  assign n3308 = ~n3273 & n3307;
  assign n3309 = ~n3176 & ~n3177;
  assign n3310 = ~n3283 & ~n3293;
  assign n3311 = ~n3277 & n3305;
  assign n3312 = n3310 & n3311;
  assign n3313 = n3309 & ~n3312;
  assign n3314 = ~n3308 & ~n3313;
  assign n3315 = n3298 & n3314;
  assign n3316 = n3286 & n3315;
  assign n3317 = n3275 & n3316;
  assign n3318 = n3317 ^ n1050;
  assign n3319 = n3318 ^ x222;
  assign n3320 = n3141 & n3319;
  assign n3321 = n2621 & n2624;
  assign n3322 = ~n2997 & ~n3186;
  assign n3323 = ~n3321 & ~n3322;
  assign n3324 = ~n2569 & n2628;
  assign n3325 = ~n2619 & n3003;
  assign n3326 = n2662 & n3325;
  assign n3327 = ~n2651 & n3326;
  assign n3328 = n2632 & ~n3327;
  assign n3329 = ~n3324 & ~n3328;
  assign n3330 = ~n2645 & n2654;
  assign n3331 = ~n2621 & n3330;
  assign n3332 = n2639 & ~n3331;
  assign n3333 = n2672 & n3191;
  assign n3334 = ~n2640 & n2662;
  assign n3335 = ~n2643 & n3334;
  assign n3336 = ~n2571 & n3335;
  assign n3337 = ~n3333 & ~n3336;
  assign n3338 = ~n2569 & n3337;
  assign n3339 = ~n3332 & ~n3338;
  assign n3340 = n3329 & n3339;
  assign n3341 = n3323 & n3340;
  assign n3342 = n2659 & n3341;
  assign n3343 = n2649 & n3342;
  assign n3344 = n3343 ^ x40;
  assign n3345 = n3344 ^ x163;
  assign n3346 = ~n1816 & n1820;
  assign n3347 = n1801 & ~n1825;
  assign n3348 = ~n3346 & ~n3347;
  assign n3349 = ~n1811 & ~n1849;
  assign n3350 = n1815 & ~n3349;
  assign n3351 = ~n1814 & n3048;
  assign n3352 = n1809 & ~n3351;
  assign n3353 = ~n3350 & ~n3352;
  assign n3354 = n1816 & n1841;
  assign n3355 = n1803 & n1836;
  assign n3356 = ~n1829 & ~n1841;
  assign n3357 = ~n1814 & n3356;
  assign n3358 = n1801 & ~n3357;
  assign n3359 = ~n1851 & ~n3059;
  assign n3360 = n1815 & ~n3359;
  assign n3361 = ~n3358 & ~n3360;
  assign n3362 = ~n3355 & n3361;
  assign n3363 = n3047 & n3362;
  assign n3364 = n3222 & n3363;
  assign n3365 = n3219 & n3364;
  assign n3366 = ~n3354 & n3365;
  assign n3367 = n3353 & n3366;
  assign n3368 = n3348 & n3367;
  assign n3369 = n3053 & n3368;
  assign n3370 = n1808 & n3369;
  assign n3371 = n3370 ^ x48;
  assign n3372 = n3371 ^ x162;
  assign n3373 = ~n3345 & n3372;
  assign n3382 = n2008 & ~n2013;
  assign n3383 = n1931 & n2013;
  assign n3384 = ~n1999 & ~n3383;
  assign n3385 = ~n1932 & ~n3384;
  assign n3386 = ~n3382 & ~n3385;
  assign n3387 = n2018 & n2032;
  assign n3388 = n1998 & n2007;
  assign n3389 = ~n1996 & n2023;
  assign n3374 = ~n1931 & ~n2013;
  assign n3390 = ~n1967 & n3374;
  assign n3391 = ~n3389 & ~n3390;
  assign n3392 = ~n3388 & n3391;
  assign n3393 = n1932 & ~n3392;
  assign n3394 = ~n3387 & ~n3393;
  assign n3395 = n3386 & n3394;
  assign n3396 = ~n2022 & n3395;
  assign n3375 = n1932 & n3374;
  assign n3376 = n2023 & n2032;
  assign n3377 = ~n2026 & ~n2038;
  assign n3378 = ~n1932 & ~n3377;
  assign n3379 = ~n3376 & ~n3378;
  assign n3380 = ~n3375 & n3379;
  assign n3381 = ~n2005 & n3380;
  assign n3397 = n3396 ^ n3381;
  assign n3398 = ~n1900 & n3397;
  assign n3399 = n3398 ^ n3396;
  assign n3400 = ~n2022 & n3399;
  assign n3401 = n3400 ^ x56;
  assign n3402 = n3401 ^ x161;
  assign n3403 = n2566 ^ x164;
  assign n3404 = n3402 & ~n3403;
  assign n3405 = n3373 & n3404;
  assign n3406 = n2770 & n2798;
  assign n3407 = n2782 & n2797;
  assign n3408 = ~n3406 & ~n3407;
  assign n3409 = n2765 & n2800;
  assign n3410 = n2769 & n2782;
  assign n3411 = ~n3409 & ~n3410;
  assign n3412 = n2787 & n3159;
  assign n3413 = ~n2797 & n3156;
  assign n3414 = n2765 & ~n3413;
  assign n3415 = ~n2792 & n2810;
  assign n3416 = ~n2769 & n3415;
  assign n3417 = n2770 & ~n3416;
  assign n3418 = ~n3414 & ~n3417;
  assign n3419 = ~n3412 & n3418;
  assign n3420 = ~n2800 & ~n2807;
  assign n3421 = n3166 & n3420;
  assign n3422 = n2782 & ~n3421;
  assign n3423 = n2790 & ~n2804;
  assign n3424 = ~n3422 & ~n3423;
  assign n3425 = n3419 & n3424;
  assign n3426 = n3411 & n3425;
  assign n3427 = n3408 & n3426;
  assign n3428 = n3147 & n3427;
  assign n3429 = n3428 ^ x6;
  assign n3430 = n3429 ^ x160;
  assign n3431 = n2719 ^ x165;
  assign n3432 = n3430 & n3431;
  assign n3433 = n3345 & ~n3372;
  assign n3434 = n3404 & n3433;
  assign n3435 = n3432 & n3434;
  assign n3436 = ~n3430 & n3431;
  assign n3437 = n3345 & n3372;
  assign n3438 = ~n3402 & n3403;
  assign n3439 = n3437 & n3438;
  assign n3440 = n3436 & n3439;
  assign n3441 = ~n3430 & ~n3431;
  assign n3442 = n3434 & n3441;
  assign n3443 = ~n3440 & ~n3442;
  assign n3444 = n3373 & n3438;
  assign n3445 = ~n3402 & ~n3403;
  assign n3446 = n3433 & n3445;
  assign n3447 = ~n3444 & ~n3446;
  assign n3448 = n3436 & ~n3447;
  assign n3449 = n3443 & ~n3448;
  assign n3450 = ~n3345 & ~n3372;
  assign n3451 = n3438 & n3450;
  assign n3452 = n3436 & n3451;
  assign n3453 = n3430 & ~n3431;
  assign n3454 = n3446 & n3453;
  assign n3455 = ~n3452 & ~n3454;
  assign n3456 = n3402 & n3403;
  assign n3457 = n3437 & n3456;
  assign n3458 = n3436 & n3457;
  assign n3459 = n3373 & n3445;
  assign n3460 = ~n3444 & ~n3459;
  assign n3461 = n3432 & ~n3460;
  assign n3462 = ~n3458 & ~n3461;
  assign n3463 = ~n3439 & ~n3459;
  assign n3464 = n3453 & ~n3463;
  assign n3465 = n3431 ^ n3430;
  assign n3466 = n3437 & n3445;
  assign n3467 = ~n3451 & ~n3466;
  assign n3468 = ~n3465 & ~n3467;
  assign n3469 = n3433 & n3438;
  assign n3470 = ~n3431 & n3469;
  assign n3471 = n3402 & n3450;
  assign n3472 = ~n3403 & n3471;
  assign n3473 = ~n3457 & ~n3472;
  assign n3474 = n3432 & ~n3473;
  assign n3475 = ~n3470 & ~n3474;
  assign n3476 = ~n3468 & n3475;
  assign n3477 = ~n3464 & n3476;
  assign n3478 = n3433 & n3456;
  assign n3479 = n3445 & n3450;
  assign n3480 = ~n3478 & ~n3479;
  assign n3481 = n3436 & ~n3480;
  assign n3482 = n3373 & n3456;
  assign n3483 = n3404 & n3437;
  assign n3484 = ~n3482 & ~n3483;
  assign n3485 = n3453 ^ n3441;
  assign n3486 = ~n3403 & n3485;
  assign n3487 = n3486 ^ n3453;
  assign n3488 = n3471 & n3487;
  assign n3489 = n3484 & ~n3488;
  assign n3490 = ~n3431 & ~n3489;
  assign n3491 = ~n3481 & ~n3490;
  assign n3492 = n3477 & n3491;
  assign n3493 = n3462 & n3492;
  assign n3494 = n3455 & n3493;
  assign n3495 = n3449 & n3494;
  assign n3496 = ~n3435 & n3495;
  assign n3497 = ~n3405 & n3496;
  assign n3498 = n3497 ^ n1121;
  assign n3499 = n3498 ^ x221;
  assign n3500 = n3015 ^ x195;
  assign n3501 = n2050 ^ x190;
  assign n3502 = n3500 & ~n3501;
  assign n3503 = n1626 ^ x191;
  assign n3504 = n2989 ^ x194;
  assign n3505 = n3503 & ~n3504;
  assign n3506 = n2110 & n2141;
  assign n3507 = n2112 & n2130;
  assign n3508 = ~n2124 & n2510;
  assign n3509 = n2132 & ~n3508;
  assign n3510 = ~n3507 & ~n3509;
  assign n3511 = ~n3506 & n3510;
  assign n3512 = n2054 & n2159;
  assign n3513 = ~n2127 & n2141;
  assign n3514 = ~n3512 & ~n3513;
  assign n3515 = ~n2148 & n2167;
  assign n3516 = n2132 & ~n3515;
  assign n3517 = n2141 & n2143;
  assign n3518 = ~n2134 & n2169;
  assign n3519 = n2112 & ~n3518;
  assign n3520 = n2151 & n2510;
  assign n3521 = ~n2137 & ~n2150;
  assign n3522 = n2141 & ~n3521;
  assign n3523 = ~n2054 & ~n3522;
  assign n3524 = ~n3520 & ~n3523;
  assign n3525 = ~n3519 & ~n3524;
  assign n3526 = ~n3517 & n3525;
  assign n3527 = ~n3516 & n3526;
  assign n3528 = n3514 & n3527;
  assign n3529 = n3511 & n3528;
  assign n3530 = n2508 & n3529;
  assign n3531 = n2136 & n3530;
  assign n3532 = n2117 & n3531;
  assign n3533 = n3532 ^ x12;
  assign n3534 = n3533 ^ x193;
  assign n3535 = n2762 & n2770;
  assign n3536 = n2765 & ~n2808;
  assign n3537 = ~n3535 & ~n3536;
  assign n3538 = ~n2787 & n2791;
  assign n3539 = ~n2806 & n3154;
  assign n3540 = n2780 & n3539;
  assign n3541 = n2787 & ~n3540;
  assign n3542 = ~n2762 & ~n2786;
  assign n3543 = n2810 & n3542;
  assign n3544 = ~n2770 & n3543;
  assign n3545 = ~n2773 & ~n2782;
  assign n3546 = n2782 & ~n3542;
  assign n3547 = n3166 & ~n3546;
  assign n3548 = ~n3545 & ~n3547;
  assign n3549 = ~n3544 & n3548;
  assign n3550 = ~n2799 & ~n3549;
  assign n3551 = ~n2804 & ~n3550;
  assign n3552 = ~n3541 & ~n3551;
  assign n3553 = ~n3538 & n3552;
  assign n3554 = n3537 & n3553;
  assign n3555 = n3411 & n3554;
  assign n3556 = n3408 & n3555;
  assign n3557 = n3146 & n3556;
  assign n3558 = n3153 & n3557;
  assign n3559 = n3558 ^ x20;
  assign n3560 = n3559 ^ x192;
  assign n3561 = ~n3534 & n3560;
  assign n3562 = n3505 & n3561;
  assign n3563 = n3502 & n3562;
  assign n3564 = n3503 & n3504;
  assign n3565 = n3534 & n3560;
  assign n3566 = n3564 & n3565;
  assign n3567 = n3502 & n3566;
  assign n3568 = ~n3500 & n3501;
  assign n3569 = ~n3503 & n3504;
  assign n3570 = ~n3534 & ~n3560;
  assign n3571 = n3569 & n3570;
  assign n3572 = n3568 & n3571;
  assign n3573 = ~n3503 & ~n3504;
  assign n3574 = n3565 & n3573;
  assign n3575 = n3561 & n3569;
  assign n3576 = ~n3574 & ~n3575;
  assign n3577 = n3502 & ~n3576;
  assign n3578 = ~n3572 & ~n3577;
  assign n3579 = n3534 & ~n3560;
  assign n3580 = n3573 & n3579;
  assign n3581 = n3502 & n3580;
  assign n3582 = ~n3500 & ~n3501;
  assign n3583 = n3569 & n3579;
  assign n3584 = n3582 & n3583;
  assign n3585 = ~n3581 & ~n3584;
  assign n3586 = ~n3500 & n3574;
  assign n3587 = n3500 & n3501;
  assign n3588 = n3534 ^ n3504;
  assign n3589 = n3588 ^ n3560;
  assign n3590 = ~n3503 & ~n3560;
  assign n3591 = n3589 & n3590;
  assign n3592 = n3591 ^ n3589;
  assign n3593 = n3587 & n3592;
  assign n3594 = ~n3586 & ~n3593;
  assign n3595 = n3501 ^ n3500;
  assign n3596 = n3570 & n3573;
  assign n3597 = ~n3575 & ~n3596;
  assign n3598 = ~n3595 & ~n3597;
  assign n3599 = n3561 & n3564;
  assign n3600 = n3505 & n3570;
  assign n3601 = ~n3599 & ~n3600;
  assign n3602 = ~n3583 & n3601;
  assign n3603 = n3502 & ~n3602;
  assign n3604 = n3565 & n3569;
  assign n3605 = ~n3580 & ~n3604;
  assign n3606 = n3568 & ~n3605;
  assign n3607 = n3505 & n3579;
  assign n3608 = ~n3562 & ~n3566;
  assign n3609 = ~n3607 & n3608;
  assign n3610 = n3582 & ~n3609;
  assign n3611 = n3564 & n3570;
  assign n3612 = ~n3600 & ~n3611;
  assign n3613 = n3505 & n3565;
  assign n3614 = n3564 & n3579;
  assign n3615 = ~n3613 & ~n3614;
  assign n3616 = n3612 & n3615;
  assign n3617 = n3609 & ~n3614;
  assign n3618 = ~n3568 & n3617;
  assign n3619 = ~n3616 & ~n3618;
  assign n3620 = ~n3610 & ~n3619;
  assign n3621 = ~n3500 & ~n3620;
  assign n3622 = ~n3606 & ~n3621;
  assign n3623 = ~n3603 & n3622;
  assign n3624 = ~n3598 & n3623;
  assign n3625 = n3594 & n3624;
  assign n3626 = n3585 & n3625;
  assign n3627 = n3578 & n3626;
  assign n3628 = ~n3567 & n3627;
  assign n3629 = ~n3563 & n3628;
  assign n3630 = n3629 ^ n1276;
  assign n3631 = n3630 ^ x223;
  assign n3632 = ~n3499 & n3631;
  assign n3633 = n3320 & n3632;
  assign n3634 = n2936 & n3633;
  assign n3635 = ~n3141 & ~n3319;
  assign n3636 = ~n3499 & ~n3631;
  assign n3637 = n3635 & n3636;
  assign n3638 = n2936 & n3637;
  assign n3639 = ~n2496 & n2935;
  assign n3640 = n3499 & n3631;
  assign n3641 = n3320 & n3640;
  assign n3642 = n3635 & n3640;
  assign n3643 = ~n3641 & ~n3642;
  assign n3644 = n3639 & ~n3643;
  assign n3645 = ~n3638 & ~n3644;
  assign n3646 = ~n3634 & n3645;
  assign n3647 = n3141 & ~n3319;
  assign n3648 = n3632 & n3647;
  assign n3649 = n2936 & n3648;
  assign n3650 = n3499 & ~n3631;
  assign n3651 = n3635 & n3650;
  assign n3652 = n3639 & n3651;
  assign n3653 = ~n3649 & ~n3652;
  assign n3654 = n2496 & ~n2935;
  assign n3655 = n3632 & n3635;
  assign n3656 = n3654 & n3655;
  assign n3657 = ~n2496 & ~n2935;
  assign n3658 = n3320 & n3636;
  assign n3659 = n3657 & n3658;
  assign n3660 = ~n3656 & ~n3659;
  assign n3661 = n3653 & n3660;
  assign n3662 = ~n3141 & n3319;
  assign n3663 = n3632 & n3662;
  assign n3664 = ~n3639 & ~n3654;
  assign n3665 = n3663 & ~n3664;
  assign n3666 = n3636 & n3662;
  assign n3667 = n3664 & n3666;
  assign n3668 = n3320 & n3650;
  assign n3669 = n3657 & n3668;
  assign n3670 = ~n3655 & ~n3658;
  assign n3671 = n3639 & ~n3670;
  assign n3672 = n3650 & n3662;
  assign n3673 = n3647 & n3650;
  assign n3674 = ~n3672 & ~n3673;
  assign n3675 = n3654 & ~n3674;
  assign n3676 = ~n3671 & ~n3675;
  assign n3677 = n3639 & n3666;
  assign n3678 = n3636 & n3647;
  assign n3679 = n3639 & n3678;
  assign n3680 = n2936 & n3668;
  assign n3681 = ~n3679 & ~n3680;
  assign n3682 = ~n3677 & n3681;
  assign n3683 = ~n3643 & n3654;
  assign n3684 = n3640 & n3662;
  assign n3685 = n3640 & n3647;
  assign n3686 = ~n3684 & ~n3685;
  assign n3687 = ~n3651 & n3686;
  assign n3688 = n3664 & ~n3687;
  assign n3689 = ~n3633 & ~n3678;
  assign n3690 = ~n2935 & ~n3689;
  assign n3691 = ~n3688 & ~n3690;
  assign n3692 = ~n3683 & n3691;
  assign n3693 = n3682 & n3692;
  assign n3694 = n3676 & n3693;
  assign n3695 = ~n3669 & n3694;
  assign n3696 = ~n3667 & n3695;
  assign n3697 = ~n3665 & n3696;
  assign n3698 = n3661 & n3697;
  assign n3699 = n3646 & n3698;
  assign n3700 = n3699 ^ n2989;
  assign n3701 = n3700 ^ x292;
  assign n3702 = ~n1346 & n2442;
  assign n3703 = ~n2431 & ~n2457;
  assign n3704 = n2439 & ~n3703;
  assign n3705 = ~n3702 & ~n3704;
  assign n3706 = ~n1346 & n2440;
  assign n3707 = n1628 & ~n2448;
  assign n3708 = ~n3706 & ~n3707;
  assign n3709 = n2473 & ~n2478;
  assign n3710 = n2439 & ~n2460;
  assign n3711 = ~n3709 & ~n3710;
  assign n3712 = n3708 & n3711;
  assign n3713 = n2447 & n2455;
  assign n3714 = ~n2445 & ~n2474;
  assign n3715 = ~n2480 & n3714;
  assign n3716 = n2186 & ~n3715;
  assign n3717 = n2051 ^ n1869;
  assign n3718 = ~n2182 & n3717;
  assign n3719 = n2455 & n3718;
  assign n3720 = ~n2425 & n2448;
  assign n3721 = ~n2473 & n3720;
  assign n3722 = n2439 & ~n3721;
  assign n3723 = ~n3719 & ~n3722;
  assign n3724 = ~n2186 & ~n2463;
  assign n3725 = ~n2468 & ~n3724;
  assign n3726 = n2184 & ~n2422;
  assign n3727 = n2186 & n2425;
  assign n3728 = ~n2436 & ~n2458;
  assign n3729 = ~n1628 & ~n2425;
  assign n3730 = ~n3728 & ~n3729;
  assign n3731 = ~n3727 & ~n3730;
  assign n3732 = ~n3726 & n3731;
  assign n3733 = ~n2437 & ~n3732;
  assign n3734 = ~n3725 & ~n3733;
  assign n3735 = n3723 & n3734;
  assign n3736 = ~n3716 & n3735;
  assign n3737 = ~n3713 & n3736;
  assign n3738 = n3712 & n3737;
  assign n3739 = n3705 & n3738;
  assign n3740 = n3739 ^ n2240;
  assign n3741 = n3740 ^ x243;
  assign n3742 = n3077 ^ x202;
  assign n3743 = n3401 ^ x207;
  assign n3744 = n3742 & n3743;
  assign n3745 = ~n2120 & ~n2143;
  assign n3746 = ~n2158 & n3745;
  assign n3747 = n2132 & ~n3746;
  assign n3748 = ~n2130 & n2151;
  assign n3749 = n2141 & ~n3748;
  assign n3750 = n2141 & n2159;
  assign n3751 = n2112 & ~n3521;
  assign n3752 = ~n2115 & n2160;
  assign n3753 = ~n2148 & n3752;
  assign n3754 = n2054 & ~n3753;
  assign n3755 = ~n3751 & ~n3754;
  assign n3756 = ~n3750 & n3755;
  assign n3757 = ~n2163 & n3756;
  assign n3758 = ~n3749 & n3757;
  assign n3759 = ~n3747 & n3758;
  assign n3760 = n3511 & n3759;
  assign n3761 = n2507 & n3760;
  assign n3762 = n2504 & n3761;
  assign n3763 = n2129 & n3762;
  assign n3764 = n2501 & n3763;
  assign n3765 = n3764 ^ x14;
  assign n3766 = n3765 ^ x205;
  assign n3767 = n2964 ^ x203;
  assign n3768 = n3766 & ~n3767;
  assign n3769 = n3429 ^ x206;
  assign n3770 = ~n1286 & ~n2836;
  assign n3771 = n1288 & ~n2845;
  assign n3772 = ~n3770 & ~n3771;
  assign n3773 = n989 & n1292;
  assign n3774 = ~n1283 & n1329;
  assign n3775 = ~n1301 & n3774;
  assign n3776 = n1285 & ~n3775;
  assign n3777 = ~n3773 & ~n3776;
  assign n3778 = n1278 ^ n1051;
  assign n3779 = ~n1122 & n3778;
  assign n3780 = n1284 & n3779;
  assign n3781 = ~n1288 & ~n1306;
  assign n3782 = ~n989 & n2844;
  assign n3783 = ~n3781 & ~n3782;
  assign n3784 = ~n1295 & ~n3783;
  assign n3785 = ~n1290 & n3784;
  assign n3786 = n1286 & ~n3785;
  assign n3787 = ~n3780 & ~n3786;
  assign n3788 = n3777 & n3787;
  assign n3789 = n3772 & n3788;
  assign n3790 = n2834 & n3789;
  assign n3791 = ~n1280 & n3790;
  assign n3792 = ~n1323 & n3791;
  assign n3793 = n3792 ^ x22;
  assign n3794 = n3793 ^ x204;
  assign n3795 = ~n3769 & ~n3794;
  assign n3796 = n3768 & n3795;
  assign n3797 = n3744 & n3796;
  assign n3798 = ~n3742 & ~n3743;
  assign n3799 = n3769 & ~n3794;
  assign n3800 = n3768 & n3799;
  assign n3801 = n3798 & n3800;
  assign n3802 = ~n3797 & ~n3801;
  assign n3803 = ~n3742 & n3743;
  assign n3804 = n3766 & n3767;
  assign n3805 = ~n3769 & n3794;
  assign n3806 = n3804 & n3805;
  assign n3807 = ~n3766 & n3767;
  assign n3808 = n3769 & n3794;
  assign n3809 = n3807 & n3808;
  assign n3810 = n3795 & n3807;
  assign n3811 = ~n3809 & ~n3810;
  assign n3812 = ~n3806 & n3811;
  assign n3813 = n3803 & ~n3812;
  assign n3814 = n3799 & n3807;
  assign n3815 = n3744 & n3814;
  assign n3816 = n3742 & ~n3743;
  assign n3817 = ~n3811 & n3816;
  assign n3818 = ~n3815 & ~n3817;
  assign n3819 = n3743 ^ n3742;
  assign n3820 = n3768 & n3805;
  assign n3821 = ~n3819 & n3820;
  assign n3822 = ~n3766 & ~n3767;
  assign n3823 = n3808 & n3822;
  assign n3824 = n3795 & n3822;
  assign n3825 = ~n3823 & ~n3824;
  assign n3826 = n3816 & ~n3825;
  assign n3827 = ~n3821 & ~n3826;
  assign n3828 = n3795 & n3804;
  assign n3829 = n3816 & n3828;
  assign n3830 = n3804 & n3808;
  assign n3831 = n3799 & n3822;
  assign n3832 = ~n3828 & ~n3831;
  assign n3833 = ~n3830 & n3832;
  assign n3834 = ~n3820 & n3833;
  assign n3835 = ~n3823 & n3834;
  assign n3836 = n3803 & ~n3835;
  assign n3837 = ~n3829 & ~n3836;
  assign n3838 = n3768 & n3808;
  assign n3839 = n3805 & n3822;
  assign n3840 = n3799 & n3804;
  assign n3841 = ~n3839 & ~n3840;
  assign n3842 = ~n3838 & n3841;
  assign n3843 = n3742 & ~n3842;
  assign n3844 = n3805 & n3807;
  assign n3845 = ~n3824 & ~n3844;
  assign n3846 = ~n3819 & ~n3845;
  assign n3847 = ~n3814 & n3833;
  assign n3848 = n3798 & ~n3847;
  assign n3849 = ~n3846 & ~n3848;
  assign n3850 = ~n3843 & n3849;
  assign n3851 = n3837 & n3850;
  assign n3852 = n3827 & n3851;
  assign n3853 = n3818 & n3852;
  assign n3854 = ~n3813 & n3853;
  assign n3855 = n3802 & n3854;
  assign n3856 = n3855 ^ n2270;
  assign n3857 = n3856 ^ x239;
  assign n3858 = n2688 ^ x172;
  assign n3859 = n3237 ^ x177;
  assign n3860 = n3858 & ~n3859;
  assign n3861 = ~n3858 & n3859;
  assign n3862 = ~n3860 & ~n3861;
  assign n3863 = n2528 ^ x173;
  assign n3864 = ~n2022 & n3381;
  assign n3865 = n3864 ^ n3396;
  assign n3866 = n1900 & ~n3865;
  assign n3867 = n3866 ^ n3396;
  assign n3868 = n3867 ^ x50;
  assign n3869 = n3868 ^ x174;
  assign n3870 = n3863 & ~n3869;
  assign n3871 = n3175 ^ x176;
  assign n3872 = n2367 & n2382;
  assign n3873 = n2242 & n2377;
  assign n3874 = ~n3872 & ~n3873;
  assign n3875 = n2216 & n2406;
  assign n3876 = ~n2369 & n2396;
  assign n3877 = n2395 & ~n2539;
  assign n3878 = ~n2241 & n2405;
  assign n3879 = ~n2393 & n2402;
  assign n3880 = ~n2391 & n3879;
  assign n3881 = n2368 & ~n3880;
  assign n3882 = ~n3878 & ~n3881;
  assign n3883 = ~n3877 & n3882;
  assign n3884 = n2242 & n2406;
  assign n3885 = ~n2367 & ~n2393;
  assign n3886 = ~n2360 & n2394;
  assign n3887 = ~n3885 & ~n3886;
  assign n3888 = ~n2377 & ~n3887;
  assign n3889 = n2216 & ~n3888;
  assign n3890 = ~n3884 & ~n3889;
  assign n3891 = n3883 & n3890;
  assign n3892 = n2938 & n3891;
  assign n3893 = ~n2358 & n3892;
  assign n3894 = ~n3876 & n3893;
  assign n3895 = ~n3875 & n3894;
  assign n3896 = n3874 & n3895;
  assign n3897 = n2942 & n3896;
  assign n3898 = n2531 & n3897;
  assign n3899 = n3898 ^ x42;
  assign n3900 = n3899 ^ x175;
  assign n3901 = n3871 & ~n3900;
  assign n3902 = n3870 & n3901;
  assign n3903 = ~n3862 & n3902;
  assign n3904 = ~n3858 & ~n3859;
  assign n3905 = n3871 & n3900;
  assign n3906 = n3870 & n3905;
  assign n3907 = n3863 & n3869;
  assign n3908 = ~n3871 & n3900;
  assign n3909 = n3907 & n3908;
  assign n3910 = ~n3906 & ~n3909;
  assign n3911 = n3904 & ~n3910;
  assign n3912 = ~n3903 & ~n3911;
  assign n3913 = n3858 & n3859;
  assign n3914 = ~n3863 & n3869;
  assign n3915 = n3908 & n3914;
  assign n3916 = n3913 & n3915;
  assign n3917 = n3905 & n3907;
  assign n3918 = n3861 & n3917;
  assign n3919 = n3870 & n3908;
  assign n3920 = n3860 & n3919;
  assign n3921 = ~n3918 & ~n3920;
  assign n3922 = ~n3916 & n3921;
  assign n3923 = n3901 & n3907;
  assign n3924 = ~n3871 & ~n3900;
  assign n3925 = n3870 & n3924;
  assign n3926 = ~n3923 & ~n3925;
  assign n3927 = n3904 & ~n3926;
  assign n3928 = n3860 & n3917;
  assign n3929 = n3861 & n3919;
  assign n3930 = n3907 & n3924;
  assign n3931 = n3901 & n3914;
  assign n3932 = ~n3915 & ~n3931;
  assign n3933 = ~n3861 & n3932;
  assign n3934 = ~n3863 & ~n3869;
  assign n3935 = n3908 & n3934;
  assign n3936 = n3901 & n3934;
  assign n3937 = ~n3935 & ~n3936;
  assign n3938 = n3932 & n3937;
  assign n3939 = ~n3933 & ~n3938;
  assign n3940 = n3905 & n3914;
  assign n3941 = n3905 & n3934;
  assign n3942 = ~n3940 & ~n3941;
  assign n3943 = ~n3860 & n3938;
  assign n3944 = ~n3942 & ~n3943;
  assign n3945 = ~n3939 & ~n3944;
  assign n3946 = ~n3930 & n3945;
  assign n3947 = ~n3862 & ~n3946;
  assign n3948 = n3924 & n3934;
  assign n3949 = ~n3941 & ~n3948;
  assign n3950 = ~n3940 & n3949;
  assign n3951 = n3913 & ~n3950;
  assign n3952 = n3914 & n3924;
  assign n3953 = ~n3931 & n3949;
  assign n3954 = n3904 & ~n3953;
  assign n3955 = ~n3919 & n3926;
  assign n3956 = ~n3913 & n3953;
  assign n3957 = ~n3955 & ~n3956;
  assign n3958 = ~n3954 & ~n3957;
  assign n3959 = ~n3952 & n3958;
  assign n3960 = n3862 & ~n3959;
  assign n3961 = ~n3951 & ~n3960;
  assign n3962 = ~n3947 & n3961;
  assign n3963 = ~n3929 & n3962;
  assign n3964 = ~n3928 & n3963;
  assign n3965 = ~n3927 & n3964;
  assign n3966 = n3922 & n3965;
  assign n3967 = n3912 & n3966;
  assign n3968 = n3967 ^ n2321;
  assign n3969 = n3968 ^ x242;
  assign n3970 = ~n3857 & n3969;
  assign n3971 = ~n3114 & n3125;
  assign n3972 = ~n3105 & ~n3109;
  assign n3973 = n2990 & ~n3972;
  assign n3974 = n3041 & n3088;
  assign n3975 = ~n3087 & ~n3974;
  assign n3976 = n3097 & n3975;
  assign n3977 = n3045 & n3976;
  assign n3978 = n3977 ^ n3975;
  assign n3979 = n2991 & ~n3978;
  assign n3980 = n3127 & ~n3974;
  assign n3981 = ~n3112 & n3980;
  assign n3982 = ~n3080 & n3981;
  assign n3983 = n3095 & ~n3982;
  assign n3984 = ~n3979 & ~n3983;
  assign n3985 = ~n3112 & n3119;
  assign n3986 = n3086 & ~n3985;
  assign n3987 = n2990 ^ n2965;
  assign n3988 = ~n3081 & ~n3125;
  assign n3989 = n3083 & n3086;
  assign n3990 = ~n3101 & ~n3989;
  assign n3991 = ~n3094 & n3990;
  assign n3992 = ~n3089 & n3991;
  assign n3993 = ~n3988 & ~n3992;
  assign n3994 = n3987 & n3993;
  assign n3995 = ~n3986 & ~n3994;
  assign n3996 = n3984 & n3995;
  assign n3997 = n3092 & n3996;
  assign n3998 = ~n3973 & n3997;
  assign n3999 = ~n3971 & n3998;
  assign n4000 = n3108 & n3999;
  assign n4001 = ~n3096 & n4000;
  assign n4002 = n4001 ^ n2350;
  assign n4003 = n4002 ^ x240;
  assign n4004 = n3441 & n3451;
  assign n4005 = n3436 & n3483;
  assign n4006 = ~n4004 & ~n4005;
  assign n4007 = n3436 & n3482;
  assign n4008 = n3432 & n3439;
  assign n4009 = ~n3444 & ~n3457;
  assign n4010 = n3441 & ~n4009;
  assign n4011 = ~n4008 & ~n4010;
  assign n4012 = ~n4007 & n4011;
  assign n4013 = ~n3466 & ~n3469;
  assign n4014 = n3453 & ~n4013;
  assign n4015 = n3451 & n3453;
  assign n4016 = n3403 & n3471;
  assign n4017 = ~n3405 & ~n4016;
  assign n4018 = ~n3483 & n4017;
  assign n4019 = n3441 & ~n4018;
  assign n4020 = ~n4015 & ~n4019;
  assign n4021 = n3432 & n3466;
  assign n4022 = ~n3459 & n3473;
  assign n4023 = n3436 & ~n4022;
  assign n4024 = ~n4021 & ~n4023;
  assign n4025 = ~n3469 & ~n3479;
  assign n4026 = ~n3465 & ~n4025;
  assign n4027 = ~n3457 & ~n3459;
  assign n4028 = ~n3453 & n4027;
  assign n4029 = ~n3405 & ~n3478;
  assign n4030 = ~n3472 & n4029;
  assign n4031 = ~n3432 & n4030;
  assign n4032 = ~n4028 & ~n4031;
  assign n4033 = ~n3482 & ~n4032;
  assign n4034 = n3430 & ~n4033;
  assign n4035 = ~n4026 & ~n4034;
  assign n4036 = n4024 & n4035;
  assign n4037 = n4020 & n4036;
  assign n4038 = ~n4014 & n4037;
  assign n4039 = n3455 & n4038;
  assign n4040 = ~n3448 & n4039;
  assign n4041 = n4012 & n4040;
  assign n4042 = ~n3435 & n4041;
  assign n4043 = n4006 & n4042;
  assign n4044 = n4043 ^ n2294;
  assign n4045 = n4044 ^ x241;
  assign n4046 = n4003 & ~n4045;
  assign n4047 = n3970 & n4046;
  assign n4048 = ~n3741 & n4047;
  assign n4049 = n3271 & n3276;
  assign n4050 = n3266 ^ n3179;
  assign n4051 = ~n3301 & n4050;
  assign n4052 = ~n3272 & n4051;
  assign n4053 = n4052 ^ n3272;
  assign n4054 = ~n4049 & n4053;
  assign n4055 = ~n3268 & n4054;
  assign n4056 = n3309 & ~n4055;
  assign n4057 = n3238 & ~n4050;
  assign n4058 = n3205 & n4057;
  assign n4059 = ~n4049 & ~n4058;
  assign n4060 = n3276 & n3288;
  assign n4061 = n3179 & n3238;
  assign n4062 = n4061 ^ n3266;
  assign n4063 = ~n3205 & ~n4062;
  assign n4064 = ~n4060 & ~n4063;
  assign n4065 = n4059 & n4064;
  assign n4066 = n3299 & n4065;
  assign n4067 = ~n4056 & ~n4066;
  assign n4068 = n3310 & ~n4058;
  assign n4069 = n3270 & ~n4068;
  assign n4070 = n3178 & ~n4064;
  assign n4071 = ~n4069 & ~n4070;
  assign n4072 = n4067 & n4071;
  assign n4073 = n3286 & n4072;
  assign n4074 = n3275 & n4073;
  assign n4075 = n4074 ^ n2215;
  assign n4076 = n4075 ^ x238;
  assign n4077 = ~n3741 & ~n4076;
  assign n4078 = ~n4003 & ~n4045;
  assign n4079 = n3970 & n4078;
  assign n4080 = ~n3857 & ~n3969;
  assign n4081 = n4046 & n4080;
  assign n4082 = ~n4079 & ~n4081;
  assign n4083 = n4077 & ~n4082;
  assign n4084 = ~n4048 & ~n4083;
  assign n4085 = n3741 & n4076;
  assign n4086 = ~n4077 & ~n4085;
  assign n4087 = ~n4003 & n4045;
  assign n4088 = n4080 & n4087;
  assign n4089 = ~n4086 & n4088;
  assign n4090 = n3741 & ~n4076;
  assign n4091 = n4003 & n4090;
  assign n4092 = n3857 & n4091;
  assign n4093 = ~n4089 & ~n4092;
  assign n4094 = n4084 & n4093;
  assign n4095 = n4003 & n4045;
  assign n4096 = n3970 & n4095;
  assign n4097 = ~n4081 & ~n4096;
  assign n4098 = ~n4079 & n4097;
  assign n4099 = n4085 & ~n4098;
  assign n4100 = ~n3741 & n4076;
  assign n4101 = n4078 & n4080;
  assign n4102 = n4097 & ~n4101;
  assign n4103 = n4100 & ~n4102;
  assign n4104 = n3857 & ~n3969;
  assign n4105 = n4078 & n4104;
  assign n4106 = n3857 & n3969;
  assign n4107 = n4095 & n4106;
  assign n4108 = n4087 & n4104;
  assign n4109 = ~n4107 & ~n4108;
  assign n4110 = ~n4096 & n4109;
  assign n4111 = ~n4105 & n4110;
  assign n4112 = n4077 & ~n4111;
  assign n4113 = n4078 & n4106;
  assign n4114 = n4080 & n4095;
  assign n4115 = n3970 & n4087;
  assign n4116 = ~n4101 & ~n4115;
  assign n4117 = ~n4114 & n4116;
  assign n4118 = ~n4113 & n4117;
  assign n4119 = n4090 & ~n4118;
  assign n4120 = n4095 & n4104;
  assign n4121 = n4046 & n4106;
  assign n4122 = ~n4108 & ~n4121;
  assign n4123 = ~n4120 & n4122;
  assign n4124 = ~n4105 & n4123;
  assign n4125 = ~n4100 & n4124;
  assign n4126 = n4003 ^ n3969;
  assign n4127 = n3857 & n4126;
  assign n4128 = n4100 & n4127;
  assign n4129 = ~n4085 & ~n4128;
  assign n4130 = ~n4125 & ~n4129;
  assign n4131 = ~n4119 & ~n4130;
  assign n4132 = ~n4112 & n4131;
  assign n4133 = ~n4103 & n4132;
  assign n4134 = ~n4099 & n4133;
  assign n4135 = n4094 & n4134;
  assign n4136 = n4135 ^ n2964;
  assign n4137 = n4136 ^ x297;
  assign n4138 = n3701 & n4137;
  assign n4139 = n3277 & n3299;
  assign n4140 = n3268 & n3309;
  assign n4141 = ~n4139 & ~n4140;
  assign n4142 = n3178 & n3312;
  assign n4143 = n3270 & ~n3306;
  assign n4144 = ~n4142 & ~n4143;
  assign n4145 = ~n3291 & n3299;
  assign n4146 = ~n3179 & n3280;
  assign n4147 = n3310 & ~n4146;
  assign n4148 = n3309 & ~n4147;
  assign n4149 = ~n4145 & ~n4148;
  assign n4150 = n4144 & n4149;
  assign n4151 = n4141 & n4150;
  assign n4152 = ~n3273 & n4151;
  assign n4153 = n4152 ^ n1355;
  assign n4154 = n4153 ^ x255;
  assign n4155 = n2864 & n2886;
  assign n4156 = n2568 & n2908;
  assign n4157 = ~n4155 & ~n4156;
  assign n4158 = n2568 & n2919;
  assign n4159 = n2868 & n2870;
  assign n4160 = n2866 & n2898;
  assign n4161 = ~n4159 & ~n4160;
  assign n4162 = ~n4158 & n4161;
  assign n4163 = ~n2879 & ~n2915;
  assign n4164 = ~n2906 & ~n4163;
  assign n4165 = n2890 & n2910;
  assign n4166 = ~n2901 & n4165;
  assign n4167 = n2568 & ~n4166;
  assign n4168 = ~n2889 & n2911;
  assign n4169 = n2866 & ~n4168;
  assign n4170 = ~n4167 & ~n4169;
  assign n4171 = ~n4164 & n4170;
  assign n4172 = ~n2877 & ~n2907;
  assign n4173 = ~n2898 & n4172;
  assign n4174 = n2870 & ~n4173;
  assign n4175 = n2826 ^ n2689;
  assign n4176 = n4175 ^ n2883;
  assign n4177 = ~n2720 & ~n4176;
  assign n4178 = n4177 ^ n2883;
  assign n4179 = n2886 & n4178;
  assign n4180 = ~n4174 & ~n4179;
  assign n4181 = n4171 & n4180;
  assign n4182 = n2875 & n4181;
  assign n4183 = n4162 & n4182;
  assign n4184 = ~n2902 & n4183;
  assign n4185 = ~n2904 & n4184;
  assign n4186 = n4157 & n4185;
  assign n4187 = n4186 ^ n1386;
  assign n4188 = n4187 ^ x250;
  assign n4189 = n4154 & n4188;
  assign n4190 = n3083 & n3125;
  assign n4191 = n3086 & n3109;
  assign n4192 = ~n4190 & ~n4191;
  assign n4193 = n3097 & n3100;
  assign n4194 = n2990 & n4193;
  assign n4195 = n3101 & n3987;
  assign n4196 = ~n4194 & ~n4195;
  assign n4197 = ~n3087 & n3111;
  assign n4198 = n3125 & ~n4197;
  assign n4199 = n3086 & ~n3127;
  assign n4200 = ~n4198 & ~n4199;
  assign n4201 = n4196 & n4200;
  assign n4202 = n2991 & ~n3129;
  assign n4203 = n3095 & n3132;
  assign n4204 = ~n4202 & ~n4203;
  assign n4205 = n4201 & n4204;
  assign n4206 = ~n3099 & n4205;
  assign n4207 = n4192 & n4206;
  assign n4208 = n3092 & n4207;
  assign n4209 = n4208 ^ n1521;
  assign n4210 = n4209 ^ x254;
  assign n4211 = ~n3583 & ~n3596;
  assign n4212 = n3582 & ~n4211;
  assign n4213 = n3578 & ~n4212;
  assign n4214 = n3561 & n3573;
  assign n4215 = n3582 & n4214;
  assign n4216 = n3568 & ~n3597;
  assign n4217 = ~n4215 & ~n4216;
  assign n4218 = ~n3562 & ~n3574;
  assign n4219 = n3615 & n4218;
  assign n4220 = ~n3583 & n4219;
  assign n4221 = n3568 & ~n4220;
  assign n4222 = ~n3571 & n3601;
  assign n4223 = ~n3566 & n4222;
  assign n4224 = n3582 & ~n4223;
  assign n4225 = ~n4221 & ~n4224;
  assign n4226 = ~n3595 & n3607;
  assign n4227 = ~n3611 & ~n3613;
  assign n4228 = ~n3607 & n4227;
  assign n4229 = n4211 & n4228;
  assign n4230 = n3502 & ~n4229;
  assign n4231 = n3612 & ~n4214;
  assign n4232 = ~n3599 & ~n3614;
  assign n4233 = ~n3604 & n4232;
  assign n4234 = n4231 & n4233;
  assign n4235 = ~n3580 & n4234;
  assign n4236 = n3587 & ~n4235;
  assign n4237 = ~n4230 & ~n4236;
  assign n4238 = ~n4226 & n4237;
  assign n4239 = n4225 & n4238;
  assign n4240 = n4217 & n4239;
  assign n4241 = n4213 & n4240;
  assign n4242 = ~n3563 & n4241;
  assign n4243 = n4242 ^ n1551;
  assign n4244 = n4243 ^ x251;
  assign n4245 = n4210 & ~n4244;
  assign n4246 = n3861 & n3948;
  assign n4247 = n3860 & n3931;
  assign n4248 = ~n4246 & ~n4247;
  assign n4249 = n3913 & ~n3937;
  assign n4250 = n4248 & ~n4249;
  assign n4251 = ~n3906 & ~n3917;
  assign n4252 = ~n3925 & n4251;
  assign n4253 = n3860 & ~n4252;
  assign n4254 = n3860 & ~n3949;
  assign n4255 = n3926 & ~n3940;
  assign n4256 = n3913 & ~n4255;
  assign n4257 = ~n4254 & ~n4256;
  assign n4258 = n3910 & ~n3948;
  assign n4259 = n3862 & ~n4258;
  assign n4260 = ~n3902 & n3938;
  assign n4261 = n3904 & ~n4260;
  assign n4262 = ~n4259 & ~n4261;
  assign n4263 = n4257 & n4262;
  assign n4264 = ~n3862 & n3923;
  assign n4265 = n3937 & ~n3952;
  assign n4266 = ~n3919 & n4265;
  assign n4267 = ~n3940 & n4266;
  assign n4268 = n3861 & ~n4267;
  assign n4269 = ~n4264 & ~n4268;
  assign n4270 = n4263 & n4269;
  assign n4271 = n3921 & n4270;
  assign n4272 = ~n4253 & n4271;
  assign n4273 = n4250 & n4272;
  assign n4274 = n4273 ^ n1456;
  assign n4275 = n4274 ^ x252;
  assign n4276 = n3444 & n3453;
  assign n4277 = n3436 & ~n4017;
  assign n4278 = ~n4276 & ~n4277;
  assign n4279 = ~n3431 & n3434;
  assign n4280 = n3453 & ~n4018;
  assign n4281 = ~n4279 & ~n4280;
  assign n4282 = n3430 & n3472;
  assign n4283 = n3439 & ~n3465;
  assign n4284 = ~n4282 & ~n4283;
  assign n4285 = ~n3459 & ~n3479;
  assign n4286 = ~n3444 & n4285;
  assign n4287 = ~n3469 & n4286;
  assign n4288 = n3436 & ~n4287;
  assign n4289 = ~n3446 & ~n3482;
  assign n4290 = ~n3478 & n4289;
  assign n4291 = n3432 & ~n4290;
  assign n4292 = ~n3457 & n3484;
  assign n4293 = n4285 & n4292;
  assign n4294 = n3441 & ~n4293;
  assign n4295 = ~n4291 & ~n4294;
  assign n4296 = ~n4288 & n4295;
  assign n4297 = n4284 & n4296;
  assign n4298 = n4281 & n4297;
  assign n4299 = n3462 & n4298;
  assign n4300 = n4278 & n4299;
  assign n4301 = ~n4014 & n4300;
  assign n4302 = ~n3435 & n4301;
  assign n4303 = n4006 & n4302;
  assign n4304 = n4303 ^ n1495;
  assign n4305 = n4304 ^ x253;
  assign n4306 = n4275 & ~n4305;
  assign n4307 = n4245 & n4306;
  assign n4308 = ~n4210 & ~n4244;
  assign n4309 = ~n4275 & ~n4305;
  assign n4310 = n4308 & n4309;
  assign n4311 = ~n4307 & ~n4310;
  assign n4312 = n4189 & ~n4311;
  assign n4313 = n4154 & ~n4188;
  assign n4314 = ~n4210 & n4244;
  assign n4315 = n4306 & n4314;
  assign n4316 = n4313 & n4315;
  assign n4317 = ~n4154 & n4188;
  assign n4318 = ~n4275 & n4305;
  assign n4319 = n4245 & n4318;
  assign n4320 = n4275 & n4305;
  assign n4321 = n4245 & n4320;
  assign n4322 = ~n4319 & ~n4321;
  assign n4323 = n4317 & ~n4322;
  assign n4324 = ~n4316 & ~n4323;
  assign n4325 = n4210 & n4244;
  assign n4326 = n4320 & n4325;
  assign n4327 = n4318 & n4325;
  assign n4328 = n4314 & n4320;
  assign n4329 = ~n4327 & ~n4328;
  assign n4330 = ~n4326 & n4329;
  assign n4331 = n4313 & ~n4330;
  assign n4332 = n4245 & n4309;
  assign n4333 = n4306 & n4308;
  assign n4334 = ~n4332 & ~n4333;
  assign n4335 = n4317 & ~n4334;
  assign n4336 = ~n4331 & ~n4335;
  assign n4337 = n4308 & n4320;
  assign n4338 = ~n4332 & ~n4337;
  assign n4339 = n4189 & ~n4338;
  assign n4340 = ~n4154 & ~n4188;
  assign n4341 = n4308 & n4318;
  assign n4342 = ~n4321 & n4338;
  assign n4343 = ~n4341 & n4342;
  assign n4344 = n4340 & ~n4343;
  assign n4345 = n4309 & n4314;
  assign n4346 = n4317 & n4345;
  assign n4347 = n4314 & n4318;
  assign n4348 = ~n4326 & ~n4347;
  assign n4349 = n4317 & ~n4348;
  assign n4350 = ~n4346 & ~n4349;
  assign n4351 = n4189 & n4315;
  assign n4352 = n4307 & n4313;
  assign n4353 = ~n4351 & ~n4352;
  assign n4354 = n4306 & n4325;
  assign n4355 = ~n4345 & ~n4354;
  assign n4356 = n4340 & ~n4355;
  assign n4357 = n4317 & n4354;
  assign n4358 = ~n4327 & n4348;
  assign n4359 = n4189 & ~n4358;
  assign n4360 = ~n4357 & ~n4359;
  assign n4361 = n4309 & n4325;
  assign n4362 = ~n4347 & ~n4361;
  assign n4363 = n4340 & ~n4362;
  assign n4364 = ~n4310 & ~n4319;
  assign n4365 = ~n4333 & n4364;
  assign n4366 = n4313 & ~n4365;
  assign n4367 = ~n4363 & ~n4366;
  assign n4368 = n4360 & n4367;
  assign n4369 = ~n4356 & n4368;
  assign n4370 = n4353 & n4369;
  assign n4371 = n4350 & n4370;
  assign n4372 = ~n4344 & n4371;
  assign n4373 = ~n4339 & n4372;
  assign n4374 = n4336 & n4373;
  assign n4375 = n4324 & n4374;
  assign n4376 = ~n4312 & n4375;
  assign n4377 = n4376 ^ n3039;
  assign n4378 = n4377 ^ x295;
  assign n4379 = n3856 ^ x237;
  assign n4380 = n3861 & n3931;
  assign n4381 = n3860 & n3952;
  assign n4382 = ~n3925 & ~n3930;
  assign n4383 = n3913 & ~n4382;
  assign n4384 = ~n4381 & ~n4383;
  assign n4385 = ~n4380 & n4384;
  assign n4386 = ~n3862 & n3915;
  assign n4387 = ~n3929 & ~n4386;
  assign n4388 = ~n3935 & n3950;
  assign n4389 = n3904 & ~n4388;
  assign n4390 = ~n3902 & ~n3936;
  assign n4391 = n3860 & ~n4390;
  assign n4392 = n3926 & n4251;
  assign n4393 = n3861 & ~n4392;
  assign n4394 = ~n4391 & ~n4393;
  assign n4395 = ~n3902 & ~n3909;
  assign n4396 = ~n3930 & n4395;
  assign n4397 = ~n3923 & n4396;
  assign n4398 = n3904 & ~n4397;
  assign n4399 = n3942 & n4395;
  assign n4400 = ~n3935 & n4399;
  assign n4401 = ~n3952 & n4400;
  assign n4402 = n3913 & ~n4401;
  assign n4403 = ~n4398 & ~n4402;
  assign n4404 = n4394 & n4403;
  assign n4405 = ~n4253 & n4404;
  assign n4406 = ~n4389 & n4405;
  assign n4407 = n4387 & n4406;
  assign n4408 = n4385 & n4407;
  assign n4409 = n4248 & n4408;
  assign n4410 = n4409 ^ n1930;
  assign n4411 = n4410 ^ x232;
  assign n4412 = ~n4379 & n4411;
  assign n4413 = n4075 ^ x236;
  assign n4414 = n2870 & n2908;
  assign n4415 = ~n2865 & ~n4414;
  assign n4416 = n2568 & n2915;
  assign n4417 = n2870 & ~n2899;
  assign n4418 = ~n4416 & ~n4417;
  assign n4419 = ~n2872 & n4172;
  assign n4420 = n2866 & ~n4419;
  assign n4421 = ~n2868 & ~n2907;
  assign n4422 = n2886 & ~n4421;
  assign n4423 = ~n2864 & ~n2919;
  assign n4424 = ~n2901 & n4423;
  assign n4425 = n2870 & ~n4424;
  assign n4426 = ~n2889 & n2899;
  assign n4427 = n2568 & ~n4426;
  assign n4428 = ~n4425 & ~n4427;
  assign n4429 = n2886 & n2893;
  assign n4430 = ~n2879 & n2910;
  assign n4431 = ~n2884 & n4430;
  assign n4432 = n2866 & ~n4431;
  assign n4433 = ~n4429 & ~n4432;
  assign n4434 = n4428 & n4433;
  assign n4435 = ~n2902 & n4434;
  assign n4436 = ~n2904 & n4435;
  assign n4437 = n4157 & n4436;
  assign n4438 = ~n4422 & n4437;
  assign n4439 = ~n4420 & n4438;
  assign n4440 = n4418 & n4439;
  assign n4441 = n4415 & n4440;
  assign n4442 = n4162 & n4441;
  assign n4443 = n2892 & n4442;
  assign n4444 = n4443 ^ n2592;
  assign n4445 = n4444 ^ x234;
  assign n4446 = n4413 & n4445;
  assign n4447 = n3587 & ~n4211;
  assign n4448 = ~n3571 & ~n3613;
  assign n4449 = n3502 & ~n4448;
  assign n4450 = ~n4447 & ~n4449;
  assign n4451 = n3597 & ~n3614;
  assign n4452 = n3502 & ~n4451;
  assign n4453 = n4228 & n4233;
  assign n4454 = n3568 & ~n4453;
  assign n4455 = ~n4452 & ~n4454;
  assign n4456 = ~n3607 & n4218;
  assign n4457 = ~n3604 & n4456;
  assign n4458 = n3612 & n4457;
  assign n4459 = n3582 & ~n4458;
  assign n4460 = ~n3575 & n4228;
  assign n4461 = ~n3580 & n4460;
  assign n4462 = ~n3599 & n4461;
  assign n4463 = n3587 & ~n4462;
  assign n4464 = ~n4459 & ~n4463;
  assign n4465 = n4455 & n4464;
  assign n4466 = n3585 & n4465;
  assign n4467 = n4450 & n4466;
  assign n4468 = n4217 & n4467;
  assign n4469 = ~n3567 & n4468;
  assign n4470 = ~n3563 & n4469;
  assign n4471 = n4470 ^ n2615;
  assign n4472 = n4471 ^ x235;
  assign n4473 = n3453 & n3469;
  assign n4474 = n3430 & n3451;
  assign n4475 = ~n4473 & ~n4474;
  assign n4476 = ~n3431 & n3459;
  assign n4477 = n3432 & ~n4285;
  assign n4478 = ~n4476 & ~n4477;
  assign n4479 = n4475 & n4478;
  assign n4480 = n3434 & n3436;
  assign n4481 = ~n3466 & n4029;
  assign n4482 = n3441 & ~n4481;
  assign n4483 = n3473 & ~n3478;
  assign n4484 = ~n3483 & n4483;
  assign n4485 = ~n3453 & n4484;
  assign n4486 = n3432 & ~n4483;
  assign n4487 = n4292 & ~n4486;
  assign n4488 = ~n3472 & n4487;
  assign n4489 = ~n4485 & ~n4488;
  assign n4490 = n3430 & n4489;
  assign n4491 = ~n4482 & ~n4490;
  assign n4492 = ~n4480 & n4491;
  assign n4493 = n4479 & n4492;
  assign n4494 = n4278 & n4493;
  assign n4495 = n4012 & n4494;
  assign n4496 = n3449 & n4495;
  assign n4497 = n4006 & n4496;
  assign n4498 = n4497 ^ n1899;
  assign n4499 = n4498 ^ x233;
  assign n4500 = ~n4472 & ~n4499;
  assign n4501 = n4446 & n4500;
  assign n4502 = ~n4413 & ~n4445;
  assign n4503 = n4500 & n4502;
  assign n4504 = ~n4501 & ~n4503;
  assign n4505 = n4412 & ~n4504;
  assign n4506 = ~n4379 & ~n4411;
  assign n4507 = n4413 & ~n4445;
  assign n4508 = n4500 & n4507;
  assign n4509 = n4506 & n4508;
  assign n4510 = n4379 & n4411;
  assign n4511 = n4472 & ~n4499;
  assign n4512 = n4446 & n4511;
  assign n4513 = n4502 & n4511;
  assign n4514 = ~n4512 & ~n4513;
  assign n4515 = n4510 & ~n4514;
  assign n4516 = ~n4509 & ~n4515;
  assign n4517 = ~n4505 & n4516;
  assign n4518 = n4412 & n4512;
  assign n4519 = n4379 & ~n4411;
  assign n4520 = n4472 & n4499;
  assign n4521 = ~n4413 & n4445;
  assign n4522 = n4520 & n4521;
  assign n4523 = ~n4472 & n4499;
  assign n4524 = n4446 & n4523;
  assign n4525 = n4502 & n4523;
  assign n4526 = n4507 & n4523;
  assign n4527 = ~n4525 & ~n4526;
  assign n4528 = ~n4524 & n4527;
  assign n4529 = ~n4522 & n4528;
  assign n4530 = n4519 & ~n4529;
  assign n4531 = ~n4518 & ~n4530;
  assign n4532 = ~n4379 & n4513;
  assign n4533 = n4507 & n4511;
  assign n4534 = ~n4525 & ~n4533;
  assign n4535 = n4506 & ~n4534;
  assign n4536 = ~n4532 & ~n4535;
  assign n4537 = n4500 & n4521;
  assign n4538 = ~n4508 & ~n4537;
  assign n4539 = n4510 & ~n4538;
  assign n4540 = n4506 & n4526;
  assign n4541 = n4511 & n4521;
  assign n4542 = n4519 & n4541;
  assign n4543 = n4521 & n4523;
  assign n4544 = n4506 & n4543;
  assign n4545 = ~n4542 & ~n4544;
  assign n4546 = n4446 & n4520;
  assign n4547 = ~n4524 & ~n4546;
  assign n4548 = n4506 & ~n4547;
  assign n4549 = n4502 & n4520;
  assign n4550 = ~n4524 & ~n4549;
  assign n4551 = n4507 & n4520;
  assign n4552 = ~n4522 & ~n4551;
  assign n4553 = n4550 & n4552;
  assign n4554 = n4510 & ~n4553;
  assign n4555 = ~n4548 & ~n4554;
  assign n4556 = ~n4512 & ~n4537;
  assign n4557 = ~n4533 & n4556;
  assign n4558 = n4519 & ~n4557;
  assign n4559 = ~n4526 & n4552;
  assign n4560 = ~n4549 & n4559;
  assign n4561 = n4412 & ~n4560;
  assign n4562 = ~n4558 & ~n4561;
  assign n4563 = n4555 & n4562;
  assign n4564 = n4545 & n4563;
  assign n4565 = ~n4540 & n4564;
  assign n4566 = ~n4539 & n4565;
  assign n4567 = n4536 & n4566;
  assign n4568 = n4531 & n4567;
  assign n4569 = n4517 & n4568;
  assign n4570 = n4569 ^ n3015;
  assign n4571 = n4570 ^ x293;
  assign n4572 = n4378 & n4571;
  assign n4573 = n2934 ^ x227;
  assign n4574 = n3744 & n3844;
  assign n4575 = n3798 & ~n3811;
  assign n4576 = ~n4574 & ~n4575;
  assign n4577 = n3803 & n3820;
  assign n4578 = ~n3806 & ~n3809;
  assign n4579 = n3744 & ~n4578;
  assign n4580 = ~n4577 & ~n4579;
  assign n4581 = ~n3819 & n3828;
  assign n4582 = ~n3800 & ~n3839;
  assign n4583 = ~n3838 & n4582;
  assign n4584 = n3803 & ~n4583;
  assign n4585 = ~n4581 & ~n4584;
  assign n4586 = n3798 & n3814;
  assign n4588 = n3767 ^ n3766;
  assign n4589 = n4588 ^ n3794;
  assign n4587 = n3767 & n3799;
  assign n4590 = n4589 ^ n4587;
  assign n4591 = n3816 & n4590;
  assign n4592 = n3811 & ~n3830;
  assign n4593 = ~n3814 & n4592;
  assign n4594 = n3803 & ~n4593;
  assign n4595 = ~n3820 & n4583;
  assign n4596 = n3798 & ~n4595;
  assign n4597 = ~n3796 & ~n3831;
  assign n4598 = ~n3838 & n4597;
  assign n4599 = ~n3824 & n4598;
  assign n4600 = n3744 & ~n4599;
  assign n4601 = ~n4596 & ~n4600;
  assign n4602 = ~n4594 & n4601;
  assign n4603 = ~n4591 & n4602;
  assign n4604 = ~n4586 & n4603;
  assign n4605 = n4585 & n4604;
  assign n4606 = n4580 & n4605;
  assign n4607 = n4576 & n4606;
  assign n4608 = n4607 ^ n1966;
  assign n4609 = n4608 ^ x229;
  assign n4610 = n4410 ^ x230;
  assign n4611 = ~n4609 & ~n4610;
  assign n4612 = n3140 ^ x226;
  assign n4613 = n4498 ^ x231;
  assign n4614 = n4612 & ~n4613;
  assign n4615 = n4611 & n4614;
  assign n4616 = ~n4573 & n4615;
  assign n4617 = ~n4612 & ~n4613;
  assign n4618 = n2425 & n2439;
  assign n4619 = ~n2463 & ~n4618;
  assign n4620 = ~n2437 & n3726;
  assign n4621 = ~n2457 & n3728;
  assign n4622 = n2186 & ~n4621;
  assign n4623 = ~n4620 & ~n4622;
  assign n4624 = ~n2428 & ~n2459;
  assign n4625 = n1628 & ~n4624;
  assign n4626 = ~n2431 & n2484;
  assign n4627 = n2439 & ~n4626;
  assign n4628 = ~n2475 & ~n2478;
  assign n4629 = ~n2447 & ~n2473;
  assign n4630 = n2186 & ~n4629;
  assign n4631 = n2460 & ~n2466;
  assign n4632 = ~n2428 & n4631;
  assign n4633 = n2439 & ~n4632;
  assign n4634 = ~n4630 & ~n4633;
  assign n4635 = ~n4628 & n4634;
  assign n4636 = n1628 & ~n3721;
  assign n4637 = n2433 & n2484;
  assign n4638 = ~n2466 & n4637;
  assign n4639 = n2455 & ~n4638;
  assign n4640 = ~n4636 & ~n4639;
  assign n4641 = n4635 & n4640;
  assign n4642 = ~n4627 & n4641;
  assign n4643 = ~n4625 & n4642;
  assign n4644 = n4623 & n4643;
  assign n4645 = n4619 & n4644;
  assign n4646 = n4645 ^ n1995;
  assign n4647 = n4646 ^ x228;
  assign n4650 = n4609 & ~n4610;
  assign n4648 = ~n4609 & n4610;
  assign n4649 = n4573 & n4648;
  assign n4651 = n4650 ^ n4649;
  assign n4652 = ~n4647 & n4651;
  assign n4653 = n4652 ^ n4649;
  assign n4654 = n4617 & n4653;
  assign n4655 = ~n4616 & ~n4654;
  assign n4656 = n4612 & n4613;
  assign n4657 = ~n4573 & ~n4647;
  assign n4658 = n4610 ^ n4609;
  assign n4659 = ~n4657 & ~n4658;
  assign n4660 = n4647 ^ n4610;
  assign n4661 = n4658 & n4660;
  assign n4662 = ~n4573 & n4661;
  assign n4663 = ~n4659 & ~n4662;
  assign n4664 = n4656 & ~n4663;
  assign n4665 = n4573 & n4647;
  assign n4666 = n4611 & n4665;
  assign n4667 = n4609 & n4610;
  assign n4668 = n4647 & n4667;
  assign n4669 = ~n4662 & ~n4668;
  assign n4670 = ~n4666 & n4669;
  assign n4671 = n4617 & ~n4670;
  assign n4672 = ~n4664 & ~n4671;
  assign n4673 = ~n4612 & n4613;
  assign n4674 = ~n4573 & n4667;
  assign n4675 = ~n4657 & ~n4665;
  assign n4676 = n4650 & n4675;
  assign n4677 = ~n4674 & ~n4676;
  assign n4678 = n4573 & ~n4609;
  assign n4679 = n4678 ^ n4611;
  assign n4680 = n4647 & n4679;
  assign n4681 = n4680 ^ n4678;
  assign n4682 = n4677 & ~n4681;
  assign n4683 = n4673 & n4682;
  assign n4684 = ~n4573 & n4647;
  assign n4685 = ~n4650 & n4684;
  assign n4686 = n4573 & ~n4658;
  assign n4687 = ~n4647 & n4686;
  assign n4688 = n4650 & ~n4675;
  assign n4689 = ~n4687 & ~n4688;
  assign n4690 = ~n4685 & n4689;
  assign n4691 = n4614 & ~n4690;
  assign n4692 = ~n4683 & ~n4691;
  assign n4693 = n4672 & n4692;
  assign n4694 = n4655 & n4693;
  assign n4695 = n4694 ^ n3044;
  assign n4696 = n4695 ^ x294;
  assign n4697 = n3498 ^ x219;
  assign n4698 = n3587 & ~n4457;
  assign n4699 = n3502 & ~n4231;
  assign n4700 = ~n4698 & ~n4699;
  assign n4701 = ~n3500 & n3562;
  assign n4702 = ~n3595 & ~n3601;
  assign n4703 = ~n4701 & ~n4702;
  assign n4704 = ~n3604 & n3615;
  assign n4705 = n3582 & ~n4704;
  assign n4706 = ~n3566 & n4461;
  assign n4707 = n3568 & ~n4706;
  assign n4708 = ~n4705 & ~n4707;
  assign n4709 = n4703 & n4708;
  assign n4710 = n4700 & n4709;
  assign n4711 = n4450 & n4710;
  assign n4712 = n4213 & n4711;
  assign n4713 = ~n3567 & n4712;
  assign n4714 = n4713 ^ n1798;
  assign n4715 = n4714 ^ x214;
  assign n4716 = ~n4697 & n4715;
  assign n4717 = ~n3800 & ~n3814;
  assign n4718 = n3744 & ~n4717;
  assign n4719 = ~n3828 & ~n3840;
  assign n4720 = ~n3830 & n4719;
  assign n4721 = n4597 & n4720;
  assign n4722 = ~n3844 & n4721;
  assign n4723 = n3816 & ~n4722;
  assign n4724 = ~n4718 & ~n4723;
  assign n4725 = n3798 & n3823;
  assign n4726 = ~n3806 & ~n3830;
  assign n4727 = ~n3831 & n4726;
  assign n4728 = ~n3819 & ~n4727;
  assign n4729 = ~n3796 & ~n3823;
  assign n4730 = n3842 & n4729;
  assign n4731 = n3803 & ~n4730;
  assign n4732 = ~n4728 & ~n4731;
  assign n4733 = ~n4725 & n4732;
  assign n4734 = n4724 & n4733;
  assign n4735 = n3827 & n4734;
  assign n4736 = n4576 & n4735;
  assign n4737 = ~n3813 & n4736;
  assign n4738 = n3802 & n4737;
  assign n4739 = n4738 ^ n1735;
  assign n4740 = n4739 ^ x215;
  assign n4741 = n3861 & n3935;
  assign n4742 = n3860 & n3948;
  assign n4743 = ~n4741 & ~n4742;
  assign n4744 = n3862 & n3923;
  assign n4745 = ~n3917 & ~n3941;
  assign n4746 = n3913 & ~n4745;
  assign n4747 = ~n4744 & ~n4746;
  assign n4748 = n4743 & n4747;
  assign n4749 = n3910 & ~n3940;
  assign n4750 = ~n3862 & ~n4749;
  assign n4751 = n3904 & ~n4267;
  assign n4752 = ~n4750 & ~n4751;
  assign n4753 = n4748 & n4752;
  assign n4754 = n4385 & n4753;
  assign n4755 = n3912 & n4754;
  assign n4756 = n3922 & n4755;
  assign n4757 = n4250 & n4756;
  assign n4758 = n4757 ^ n1659;
  assign n4759 = n4758 ^ x216;
  assign n4760 = ~n4740 & ~n4759;
  assign n4761 = n2495 ^ x218;
  assign n4762 = n3109 & n3125;
  assign n4763 = ~n3105 & ~n3110;
  assign n4764 = ~n3098 & n4763;
  assign n4765 = n3095 & ~n4764;
  assign n4766 = ~n4762 & ~n4765;
  assign n4767 = n3086 & ~n3128;
  assign n4768 = ~n3080 & ~n3089;
  assign n4769 = n2990 & ~n4768;
  assign n4770 = ~n3094 & ~n3974;
  assign n4771 = n2991 & ~n4770;
  assign n4772 = n3095 & ~n3975;
  assign n4773 = ~n4771 & ~n4772;
  assign n4774 = ~n3118 & ~n4193;
  assign n4775 = ~n2991 & n4774;
  assign n4776 = n3987 & ~n4774;
  assign n4777 = n4763 & ~n4776;
  assign n4778 = ~n4775 & ~n4777;
  assign n4779 = ~n3112 & ~n4778;
  assign n4780 = ~n3095 & ~n4779;
  assign n4781 = n4773 & ~n4780;
  assign n4782 = n3103 & n4781;
  assign n4783 = ~n4769 & n4782;
  assign n4784 = ~n4767 & n4783;
  assign n4785 = n4766 & n4784;
  assign n4786 = n4192 & n4785;
  assign n4787 = ~n3989 & n4786;
  assign n4788 = ~n3096 & n4787;
  assign n4789 = n4788 ^ n1768;
  assign n4790 = n4789 ^ x217;
  assign n4791 = ~n4761 & ~n4790;
  assign n4792 = n4760 & n4791;
  assign n4793 = n4716 & n4792;
  assign n4794 = n4697 & n4715;
  assign n4795 = n4761 & n4790;
  assign n4796 = n4760 & n4795;
  assign n4797 = n4794 & n4796;
  assign n4798 = ~n4740 & n4759;
  assign n4799 = n4795 & n4798;
  assign n4800 = n4716 & n4799;
  assign n4801 = ~n4797 & ~n4800;
  assign n4802 = ~n4697 & ~n4715;
  assign n4803 = ~n4761 & n4790;
  assign n4804 = n4798 & n4803;
  assign n4805 = n4761 & ~n4790;
  assign n4806 = n4760 & n4805;
  assign n4807 = ~n4804 & ~n4806;
  assign n4808 = n4802 & ~n4807;
  assign n4809 = n4740 & n4759;
  assign n4810 = n4803 & n4809;
  assign n4811 = n4805 & n4809;
  assign n4812 = ~n4810 & ~n4811;
  assign n4813 = n4716 & ~n4812;
  assign n4814 = ~n4808 & ~n4813;
  assign n4815 = n4801 & n4814;
  assign n4816 = ~n4793 & n4815;
  assign n4817 = n4697 & ~n4715;
  assign n4818 = n4792 & n4817;
  assign n4819 = n4791 & n4809;
  assign n4820 = n4794 & n4819;
  assign n4821 = n4798 & n4805;
  assign n4822 = n4817 & n4821;
  assign n4823 = ~n4820 & ~n4822;
  assign n4824 = ~n4818 & n4823;
  assign n4825 = n4791 & n4798;
  assign n4826 = n4716 & n4825;
  assign n4827 = ~n4716 & ~n4817;
  assign n4828 = n4760 & n4803;
  assign n4829 = n4827 & n4828;
  assign n4830 = n4794 & n4806;
  assign n4831 = ~n4829 & ~n4830;
  assign n4832 = ~n4826 & n4831;
  assign n4833 = n4740 & ~n4759;
  assign n4834 = n4791 & n4833;
  assign n4835 = n4795 & n4809;
  assign n4836 = ~n4825 & ~n4835;
  assign n4837 = ~n4834 & n4836;
  assign n4838 = ~n4799 & n4837;
  assign n4839 = n4794 & ~n4838;
  assign n4840 = n4805 & n4833;
  assign n4841 = ~n4796 & ~n4819;
  assign n4842 = ~n4840 & n4841;
  assign n4843 = n4716 & ~n4842;
  assign n4844 = n4803 & n4833;
  assign n4845 = ~n4835 & ~n4844;
  assign n4846 = ~n4811 & n4845;
  assign n4847 = ~n4821 & n4846;
  assign n4848 = ~n4834 & n4847;
  assign n4849 = n4802 & ~n4848;
  assign n4850 = n4795 & n4833;
  assign n4851 = ~n4810 & ~n4840;
  assign n4852 = ~n4850 & n4851;
  assign n4853 = ~n4844 & n4852;
  assign n4854 = ~n4811 & n4853;
  assign n4855 = ~n4804 & n4854;
  assign n4856 = n4817 & ~n4855;
  assign n4857 = ~n4849 & ~n4856;
  assign n4858 = ~n4843 & n4857;
  assign n4859 = ~n4839 & n4858;
  assign n4860 = n4832 & n4859;
  assign n4861 = n4824 & n4860;
  assign n4862 = n4816 & n4861;
  assign n4863 = n4862 ^ n3077;
  assign n4864 = n4863 ^ x296;
  assign n4865 = n4696 & ~n4864;
  assign n4866 = n4572 & n4865;
  assign n4867 = n4696 & n4864;
  assign n4868 = ~n4378 & n4571;
  assign n4869 = n4867 & n4868;
  assign n4870 = ~n4866 & ~n4869;
  assign n4871 = n4138 & ~n4870;
  assign n4872 = ~n3701 & n4137;
  assign n4873 = n4865 & n4868;
  assign n4874 = ~n4696 & n4864;
  assign n4875 = n4868 & n4874;
  assign n4876 = ~n4873 & ~n4875;
  assign n4877 = n4872 & ~n4876;
  assign n4878 = ~n4871 & ~n4877;
  assign n4879 = n4378 & ~n4571;
  assign n4880 = n4865 & n4879;
  assign n4881 = n4872 & n4880;
  assign n4882 = ~n4378 & ~n4571;
  assign n4883 = n4865 & n4882;
  assign n4884 = n4138 & n4883;
  assign n4885 = ~n4881 & ~n4884;
  assign n4886 = n4874 & n4882;
  assign n4887 = n4138 & n4886;
  assign n4888 = ~n3701 & ~n4137;
  assign n4889 = n4572 & n4867;
  assign n4890 = ~n4696 & ~n4864;
  assign n4891 = n4572 & n4890;
  assign n4892 = ~n4889 & ~n4891;
  assign n4893 = n4888 & ~n4892;
  assign n4894 = n4868 & n4890;
  assign n4895 = ~n4138 & ~n4888;
  assign n4896 = n4894 & ~n4895;
  assign n4897 = ~n4893 & ~n4896;
  assign n4898 = ~n4869 & ~n4880;
  assign n4899 = n4888 & ~n4898;
  assign n4900 = n4874 & n4879;
  assign n4901 = ~n4891 & ~n4900;
  assign n4902 = ~n4880 & n4901;
  assign n4903 = n4138 & ~n4902;
  assign n4904 = ~n4899 & ~n4903;
  assign n4905 = n3701 & ~n4137;
  assign n4906 = n4867 & n4879;
  assign n4907 = ~n4875 & ~n4891;
  assign n4908 = ~n4906 & n4907;
  assign n4909 = ~n4883 & ~n4886;
  assign n4910 = ~n4900 & n4909;
  assign n4911 = n4908 & n4910;
  assign n4912 = n4898 & n4911;
  assign n4913 = n4905 & n4912;
  assign n4914 = ~n4866 & ~n4906;
  assign n4915 = n4872 & ~n4914;
  assign n4916 = n4867 & n4882;
  assign n4917 = n4879 & n4890;
  assign n4918 = ~n4916 & ~n4917;
  assign n4919 = ~n4886 & n4918;
  assign n4920 = ~n3701 & ~n4919;
  assign n4921 = ~n4915 & ~n4920;
  assign n4922 = ~n4913 & n4921;
  assign n4923 = n4904 & n4922;
  assign n4924 = n4897 & n4923;
  assign n4925 = ~n4887 & n4924;
  assign n4926 = n4885 & n4925;
  assign n4927 = n4878 & n4926;
  assign n4928 = n4927 ^ n3140;
  assign n4929 = n4928 ^ x322;
  assign n4930 = n4313 & ~n4348;
  assign n4931 = ~n4334 & n4340;
  assign n4932 = ~n4930 & ~n4931;
  assign n4933 = n4317 & n4341;
  assign n4934 = n4189 & ~n4329;
  assign n4935 = ~n4933 & ~n4934;
  assign n4936 = ~n4307 & ~n4337;
  assign n4937 = ~n4321 & n4936;
  assign n4938 = n4313 & ~n4937;
  assign n4939 = ~n4322 & n4340;
  assign n4940 = n4340 & ~n4348;
  assign n4941 = n4188 ^ n4154;
  assign n4942 = ~n4315 & ~n4354;
  assign n4943 = ~n4941 & ~n4942;
  assign n4944 = ~n4940 & ~n4943;
  assign n4945 = ~n4310 & ~n4361;
  assign n4946 = n4313 & ~n4945;
  assign n4947 = n4334 & n4364;
  assign n4948 = n4189 & ~n4947;
  assign n4949 = ~n4328 & n4945;
  assign n4950 = ~n4354 & n4949;
  assign n4951 = n4317 & ~n4950;
  assign n4952 = ~n4948 & ~n4951;
  assign n4953 = ~n4946 & n4952;
  assign n4954 = n4944 & n4953;
  assign n4955 = ~n4939 & n4954;
  assign n4956 = ~n4938 & n4955;
  assign n4957 = ~n4346 & n4956;
  assign n4958 = n4324 & n4957;
  assign n4959 = n4935 & n4958;
  assign n4960 = n4932 & n4959;
  assign n4961 = n4960 ^ n2719;
  assign n4962 = n4961 ^ x261;
  assign n4963 = n3825 & n4720;
  assign n4964 = n3798 & ~n4963;
  assign n4965 = ~n3744 & ~n3839;
  assign n4966 = ~n4583 & ~n4965;
  assign n4967 = ~n3819 & n4966;
  assign n4968 = ~n4964 & ~n4967;
  assign n4969 = ~n3800 & n3835;
  assign n4970 = n3816 & ~n4969;
  assign n4971 = n3810 & ~n3819;
  assign n4972 = n4578 & n4598;
  assign n4973 = ~n3844 & n4972;
  assign n4974 = ~n3814 & n4973;
  assign n4975 = n3803 & ~n4974;
  assign n4976 = ~n4971 & ~n4975;
  assign n4977 = ~n4970 & n4976;
  assign n4978 = n4968 & n4977;
  assign n4979 = n4580 & n4978;
  assign n4980 = n3818 & n4979;
  assign n4981 = n3802 & n4980;
  assign n4982 = n4981 ^ n2759;
  assign n4983 = n4982 ^ x247;
  assign n4984 = n3740 ^ x245;
  assign n4985 = ~n4983 & ~n4984;
  assign n4986 = ~n3273 & n4068;
  assign n4987 = n3299 & ~n4986;
  assign n4988 = n3284 & n4064;
  assign n4989 = n3309 & ~n4988;
  assign n4990 = ~n4987 & ~n4989;
  assign n4991 = n3178 & n4055;
  assign n4992 = n3270 & ~n4065;
  assign n4993 = ~n4991 & ~n4992;
  assign n4994 = n4990 & n4993;
  assign n4995 = n4141 & n4994;
  assign n4996 = n4995 ^ n2729;
  assign n4997 = n4996 ^ x246;
  assign n4998 = n4187 ^ x248;
  assign n4999 = ~n4997 & n4998;
  assign n5000 = n4985 & n4999;
  assign n5001 = n4983 & ~n4984;
  assign n5002 = n4997 & ~n4998;
  assign n5003 = n5001 & n5002;
  assign n5004 = ~n5000 & ~n5003;
  assign n5005 = n4243 ^ x249;
  assign n5006 = n3968 ^ x244;
  assign n5007 = n5005 & ~n5006;
  assign n5008 = ~n5004 & n5007;
  assign n5009 = n5005 & n5006;
  assign n5010 = ~n4983 & n4984;
  assign n5011 = n4997 & n4998;
  assign n5012 = n5010 & n5011;
  assign n5013 = n4983 & n4984;
  assign n5014 = n5002 & n5013;
  assign n5015 = ~n5012 & ~n5014;
  assign n5016 = n5009 & ~n5015;
  assign n5017 = n4999 & n5010;
  assign n5018 = n5002 & n5010;
  assign n5019 = ~n5017 & ~n5018;
  assign n5020 = n5007 & ~n5019;
  assign n5021 = ~n5016 & ~n5020;
  assign n5022 = ~n5008 & n5021;
  assign n5023 = n4999 & n5001;
  assign n5024 = n5007 & n5023;
  assign n5025 = ~n5005 & n5006;
  assign n5026 = n4998 ^ n4997;
  assign n5027 = n4985 & ~n5026;
  assign n5028 = n5004 & ~n5012;
  assign n5029 = n5013 & ~n5026;
  assign n5030 = n5028 & ~n5029;
  assign n5031 = ~n5027 & n5030;
  assign n5032 = ~n5018 & n5031;
  assign n5033 = n5025 & ~n5032;
  assign n5034 = ~n5024 & ~n5033;
  assign n5035 = ~n5005 & ~n5006;
  assign n5036 = n5001 & n5011;
  assign n5037 = ~n4997 & ~n4998;
  assign n5038 = n5013 & n5037;
  assign n5039 = ~n4984 & n5026;
  assign n5040 = ~n5038 & ~n5039;
  assign n5041 = ~n5012 & n5040;
  assign n5042 = ~n5017 & n5041;
  assign n5043 = ~n5036 & n5042;
  assign n5044 = n5035 & n5043;
  assign n5045 = ~n5027 & ~n5036;
  assign n5046 = n5009 & ~n5045;
  assign n5047 = n4985 & n5002;
  assign n5048 = ~n5007 & ~n5038;
  assign n5049 = n5029 & ~n5048;
  assign n5050 = ~n5047 & ~n5049;
  assign n5051 = ~n5017 & n5050;
  assign n5052 = n5005 & ~n5051;
  assign n5053 = ~n5046 & ~n5052;
  assign n5054 = ~n5044 & n5053;
  assign n5055 = n5034 & n5054;
  assign n5056 = n5022 & n5055;
  assign n5057 = n5056 ^ n3429;
  assign n5058 = n5057 ^ x256;
  assign n5059 = n4962 & n5058;
  assign n5060 = n4519 & ~n4550;
  assign n5061 = ~n4501 & ~n4533;
  assign n5062 = n4412 & ~n5061;
  assign n5063 = ~n5060 & ~n5062;
  assign n5064 = ~n4379 & n4541;
  assign n5065 = ~n4525 & ~n4543;
  assign n5066 = n4519 & ~n5065;
  assign n5067 = ~n5064 & ~n5066;
  assign n5068 = n4412 & n4513;
  assign n5069 = n4411 ^ n4379;
  assign n5070 = ~n4533 & ~n4537;
  assign n5071 = ~n5069 & ~n5070;
  assign n5072 = ~n4501 & ~n4512;
  assign n5073 = ~n4508 & n5072;
  assign n5074 = n4519 & ~n5073;
  assign n5075 = ~n4546 & ~n4549;
  assign n5076 = ~n4551 & n5075;
  assign n5077 = n4506 & ~n5076;
  assign n5078 = ~n5074 & ~n5077;
  assign n5079 = ~n4503 & ~n4512;
  assign n5080 = n4510 & ~n5079;
  assign n5081 = ~n4546 & n4559;
  assign n5082 = n4510 & ~n5081;
  assign n5083 = n4528 & ~n4551;
  assign n5084 = n4412 & ~n5083;
  assign n5085 = ~n5082 & ~n5084;
  assign n5086 = ~n5080 & n5085;
  assign n5087 = n5078 & n5086;
  assign n5088 = n4545 & n5087;
  assign n5089 = ~n5071 & n5088;
  assign n5090 = ~n5068 & n5089;
  assign n5091 = n5067 & n5090;
  assign n5092 = n5063 & n5091;
  assign n5093 = ~n4540 & n5092;
  assign n5094 = n5093 ^ n3344;
  assign n5095 = n5094 ^ x259;
  assign n5096 = n4090 & n4113;
  assign n5097 = n4047 & n4085;
  assign n5098 = ~n5096 & ~n5097;
  assign n5099 = ~n4047 & ~n4114;
  assign n5100 = n4077 & ~n5099;
  assign n5101 = ~n4079 & ~n4088;
  assign n5102 = n4085 & ~n5101;
  assign n5103 = ~n5100 & ~n5102;
  assign n5104 = n4085 & n4101;
  assign n5105 = n4077 & n4079;
  assign n5106 = ~n5104 & ~n5105;
  assign n5107 = ~n3741 & n4105;
  assign n5108 = n4097 & ~n4115;
  assign n5109 = n4086 & ~n5108;
  assign n5110 = ~n5107 & ~n5109;
  assign n5111 = n4003 & n4104;
  assign n5112 = ~n4105 & ~n5111;
  assign n5113 = ~n4088 & n5112;
  assign n5114 = n4090 & ~n5113;
  assign n5115 = n4046 & n4104;
  assign n5116 = ~n4113 & ~n5115;
  assign n5117 = n4109 & n5116;
  assign n5118 = n4100 & ~n5117;
  assign n5119 = n4087 & n4106;
  assign n5120 = ~n4085 & n4123;
  assign n5121 = n4122 & ~n5115;
  assign n5122 = ~n4077 & n5121;
  assign n5123 = ~n5120 & ~n5122;
  assign n5124 = ~n5119 & ~n5123;
  assign n5125 = ~n4086 & ~n5124;
  assign n5126 = ~n5118 & ~n5125;
  assign n5127 = ~n5114 & n5126;
  assign n5128 = n5110 & n5127;
  assign n5129 = n5106 & n5128;
  assign n5130 = n5103 & n5129;
  assign n5131 = n5098 & n5130;
  assign n5132 = n5131 ^ n2566;
  assign n5133 = n5132 ^ x260;
  assign n5134 = ~n5095 & n5133;
  assign n5135 = n4573 & n4650;
  assign n5136 = n4647 & n5135;
  assign n5137 = ~n4647 & n4649;
  assign n5138 = ~n4685 & ~n5137;
  assign n5139 = n4617 & ~n5138;
  assign n5140 = ~n5136 & ~n5139;
  assign n5141 = n4610 ^ n4573;
  assign n5142 = n4647 & ~n5141;
  assign n5143 = ~n4609 & n5142;
  assign n5144 = ~n4687 & ~n5143;
  assign n5145 = ~n4662 & n5144;
  assign n5146 = ~n5135 & n5145;
  assign n5147 = n4673 & ~n5146;
  assign n5148 = n5140 & ~n5147;
  assign n5149 = ~n4647 & n4667;
  assign n5150 = n4610 & ~n4675;
  assign n5151 = ~n5149 & ~n5150;
  assign n5152 = n4614 & ~n5151;
  assign n5153 = n4647 & ~n4658;
  assign n5154 = ~n4688 & ~n5153;
  assign n5155 = ~n4674 & n5154;
  assign n5156 = ~n5137 & n5155;
  assign n5157 = n4656 & ~n5156;
  assign n5158 = ~n5152 & ~n5157;
  assign n5159 = n5148 & n5158;
  assign n5160 = n4655 & n5159;
  assign n5161 = n5160 ^ n3401;
  assign n5162 = n5161 ^ x257;
  assign n5163 = n4794 & n4804;
  assign n5164 = n4716 & n4821;
  assign n5165 = ~n5163 & ~n5164;
  assign n5166 = n4799 & n4802;
  assign n5167 = n4817 & n4840;
  assign n5168 = ~n5166 & ~n5167;
  assign n5169 = n5165 & n5168;
  assign n5170 = n4792 & n4794;
  assign n5171 = n4817 & ~n4846;
  assign n5172 = ~n5170 & ~n5171;
  assign n5173 = n4716 & n4804;
  assign n5174 = n4806 & n4827;
  assign n5175 = ~n5173 & ~n5174;
  assign n5176 = ~n4828 & ~n4834;
  assign n5177 = n4802 & ~n5176;
  assign n5185 = ~n4840 & ~n4844;
  assign n5186 = ~n4819 & n5185;
  assign n5187 = n4716 & ~n5186;
  assign n5188 = ~n4804 & n5176;
  assign n5189 = ~n4806 & n5188;
  assign n5190 = ~n4817 & ~n4834;
  assign n5191 = n5186 & n5190;
  assign n5192 = ~n5189 & ~n5191;
  assign n5193 = ~n5187 & ~n5192;
  assign n5178 = ~n4794 & n4812;
  assign n5179 = ~n4802 & ~n4811;
  assign n5180 = ~n4812 & ~n5179;
  assign n5181 = ~n4835 & ~n5180;
  assign n5182 = ~n5178 & ~n5181;
  assign n5183 = ~n4850 & ~n5182;
  assign n5184 = ~n4819 & n5183;
  assign n5194 = n5193 ^ n5184;
  assign n5195 = n4827 & n5194;
  assign n5196 = n5195 ^ n5193;
  assign n5197 = ~n5177 & n5196;
  assign n5198 = n5175 & n5197;
  assign n5199 = n5172 & n5198;
  assign n5200 = n4801 & n5199;
  assign n5201 = ~n4793 & n5200;
  assign n5202 = n5169 & n5201;
  assign n5203 = n5202 ^ n3371;
  assign n5204 = n5203 ^ x258;
  assign n5205 = n5162 & n5204;
  assign n5206 = n5134 & n5205;
  assign n5207 = n5059 & n5206;
  assign n5208 = ~n4962 & n5058;
  assign n5209 = n5095 & n5133;
  assign n5210 = n5205 & n5209;
  assign n5211 = n5208 & n5210;
  assign n5212 = ~n5207 & ~n5211;
  assign n5213 = n4962 & ~n5058;
  assign n5214 = ~n5095 & ~n5133;
  assign n5215 = n5205 & n5214;
  assign n5216 = n5095 & ~n5133;
  assign n5217 = n5205 & n5216;
  assign n5218 = n5162 & ~n5204;
  assign n5219 = n5209 & n5218;
  assign n5220 = ~n5217 & ~n5219;
  assign n5221 = ~n5215 & n5220;
  assign n5222 = n5213 & ~n5221;
  assign n5223 = n5216 & n5218;
  assign n5224 = n5059 & n5223;
  assign n5225 = ~n5162 & ~n5204;
  assign n5226 = n5134 & n5225;
  assign n5227 = ~n5215 & ~n5226;
  assign n5228 = n5208 & ~n5227;
  assign n5229 = ~n5224 & ~n5228;
  assign n5230 = ~n5222 & n5229;
  assign n5231 = ~n4962 & ~n5058;
  assign n5232 = n5214 & n5218;
  assign n5233 = n5231 & n5232;
  assign n5234 = ~n5162 & n5204;
  assign n5235 = n5209 & n5234;
  assign n5236 = n5213 & n5235;
  assign n5237 = n5216 & n5234;
  assign n5238 = n5059 & n5237;
  assign n5239 = ~n5236 & ~n5238;
  assign n5240 = ~n5233 & n5239;
  assign n5241 = n5206 & n5231;
  assign n5242 = n5208 & n5223;
  assign n5243 = ~n5241 & ~n5242;
  assign n5244 = ~n5059 & ~n5231;
  assign n5245 = n5134 & n5218;
  assign n5246 = ~n5244 & n5245;
  assign n5247 = n5209 & n5225;
  assign n5248 = n5134 & n5234;
  assign n5249 = n5216 & n5225;
  assign n5250 = ~n5248 & ~n5249;
  assign n5251 = ~n5215 & n5250;
  assign n5252 = ~n5247 & n5251;
  assign n5253 = n5059 & ~n5252;
  assign n5254 = ~n5246 & ~n5253;
  assign n5255 = ~n5235 & ~n5237;
  assign n5256 = ~n5247 & n5255;
  assign n5257 = ~n5206 & n5256;
  assign n5258 = n5208 & ~n5257;
  assign n5259 = n5214 & n5225;
  assign n5260 = ~n5248 & ~n5259;
  assign n5261 = ~n5210 & ~n5232;
  assign n5262 = n5260 & n5261;
  assign n5263 = n5213 & ~n5262;
  assign n5264 = n5214 & n5234;
  assign n5265 = n5256 & ~n5264;
  assign n5266 = ~n5217 & n5265;
  assign n5267 = n5231 & ~n5266;
  assign n5268 = ~n5263 & ~n5267;
  assign n5269 = ~n5258 & n5268;
  assign n5270 = n5254 & n5269;
  assign n5271 = n5243 & n5270;
  assign n5272 = n5240 & n5271;
  assign n5273 = n5230 & n5272;
  assign n5274 = n5212 & n5273;
  assign n5275 = n5274 ^ n4498;
  assign n5276 = n5275 ^ x327;
  assign n5277 = ~n4929 & n5276;
  assign n5278 = n4657 & n4673;
  assign n5279 = n4650 & n5278;
  assign n5280 = n4611 & n4656;
  assign n5281 = ~n4573 & n5280;
  assign n5282 = ~n5279 & ~n5281;
  assign n5283 = n4614 & n4663;
  assign n5284 = ~n4647 & n5135;
  assign n5285 = ~n4609 & n4665;
  assign n5286 = ~n5284 & ~n5285;
  assign n5287 = n4669 & n5286;
  assign n5288 = n4673 & ~n5287;
  assign n5289 = ~n5283 & ~n5288;
  assign n5290 = n4617 & ~n4682;
  assign n5291 = n4656 & ~n4690;
  assign n5292 = ~n5290 & ~n5291;
  assign n5293 = n5289 & n5292;
  assign n5294 = n5282 & n5293;
  assign n5295 = n5294 ^ n2050;
  assign n5296 = n5295 ^ x284;
  assign n5297 = n4077 & n4113;
  assign n5298 = ~n4082 & ~n4086;
  assign n5299 = ~n5297 & ~n5298;
  assign n5300 = ~n3741 & n4115;
  assign n5301 = ~n4105 & ~n5119;
  assign n5302 = n4109 & n5301;
  assign n5303 = ~n4114 & n5302;
  assign n5304 = n4085 & ~n5303;
  assign n5305 = ~n5300 & ~n5304;
  assign n5306 = ~n4096 & ~n4101;
  assign n5307 = ~n4088 & n5306;
  assign n5308 = n4100 & ~n5307;
  assign n5309 = n4098 & n4123;
  assign n5310 = ~n4114 & n5309;
  assign n5311 = n4090 & ~n5310;
  assign n5312 = ~n4121 & n5112;
  assign n5313 = ~n4077 & n5312;
  assign n5314 = ~n4107 & n4123;
  assign n5315 = ~n4100 & n5314;
  assign n5316 = ~n5313 & ~n5315;
  assign n5317 = ~n3741 & n5316;
  assign n5318 = ~n5311 & ~n5317;
  assign n5319 = ~n5308 & n5318;
  assign n5320 = n5305 & n5319;
  assign n5321 = n5299 & n5320;
  assign n5322 = n5098 & n5321;
  assign n5323 = n5322 ^ n2421;
  assign n5324 = n5323 ^ x283;
  assign n5325 = n5296 & n5324;
  assign n5326 = n4794 & n4799;
  assign n5327 = n4817 & n4819;
  assign n5328 = ~n5326 & ~n5327;
  assign n5329 = n4794 & ~n4852;
  assign n5330 = n4841 & n4846;
  assign n5331 = ~n4825 & n5330;
  assign n5332 = n4802 & ~n5331;
  assign n5333 = ~n5329 & ~n5332;
  assign n5334 = ~n4806 & n4853;
  assign n5335 = n4716 & ~n5334;
  assign n5336 = ~n4850 & n5188;
  assign n5337 = ~n4799 & n5336;
  assign n5338 = n4817 & ~n5337;
  assign n5339 = ~n5335 & ~n5338;
  assign n5340 = n5333 & n5339;
  assign n5341 = n4823 & n5340;
  assign n5342 = n5328 & n5341;
  assign n5343 = n4832 & n5342;
  assign n5344 = ~n4793 & n5343;
  assign n5345 = n5169 & n5344;
  assign n5346 = n5345 ^ n1868;
  assign n5347 = n5346 ^ x282;
  assign n5348 = n4209 ^ x208;
  assign n5349 = n4739 ^ x213;
  assign n5350 = n5348 & ~n5349;
  assign n5351 = n4153 ^ x209;
  assign n5352 = ~n1346 & n2473;
  assign n5353 = ~n2437 & n2480;
  assign n5354 = ~n5352 & ~n5353;
  assign n5355 = n2427 & n2439;
  assign n5356 = ~n2440 & n2475;
  assign n5357 = n2186 & ~n5356;
  assign n5358 = ~n5355 & ~n5357;
  assign n5359 = n5354 & n5358;
  assign n5360 = n1628 & n2447;
  assign n5361 = ~n2425 & ~n2445;
  assign n5362 = n2455 & ~n5361;
  assign n5363 = ~n2431 & n2460;
  assign n5364 = ~n2473 & n5363;
  assign n5365 = n2186 & ~n5364;
  assign n5366 = ~n2440 & n3714;
  assign n5367 = n2439 & ~n5366;
  assign n5368 = ~n2455 & n4631;
  assign n5369 = ~n3726 & n4624;
  assign n5370 = ~n2431 & n5369;
  assign n5371 = ~n1628 & n5370;
  assign n5372 = ~n5368 & ~n5371;
  assign n5373 = ~n1346 & n5372;
  assign n5374 = ~n5367 & ~n5373;
  assign n5375 = ~n5365 & n5374;
  assign n5376 = n4619 & n5375;
  assign n5377 = ~n5362 & n5376;
  assign n5378 = ~n5360 & n5377;
  assign n5379 = n5359 & n5378;
  assign n5380 = n3705 & n5379;
  assign n5381 = n5380 ^ n2107;
  assign n5382 = n5381 ^ x211;
  assign n5383 = n5351 & ~n5382;
  assign n5384 = n4714 ^ x212;
  assign n5385 = n2886 & n2894;
  assign n5386 = n2870 & n2879;
  assign n5387 = ~n5385 & ~n5386;
  assign n5388 = ~n2866 & ~n2886;
  assign n5389 = n2884 & ~n5388;
  assign n5390 = ~n2868 & ~n2915;
  assign n5391 = n2568 & ~n5390;
  assign n5392 = ~n5389 & ~n5391;
  assign n5393 = ~n2906 & ~n2920;
  assign n5394 = n2870 & n2888;
  assign n5395 = n2568 & ~n2910;
  assign n5396 = ~n5394 & ~n5395;
  assign n5397 = n2886 & n2908;
  assign n5398 = n2872 & ~n5388;
  assign n5399 = n2866 & ~n5390;
  assign n5400 = ~n5398 & ~n5399;
  assign n5401 = ~n5397 & n5400;
  assign n5402 = n5396 & n5401;
  assign n5403 = n4415 & n5402;
  assign n5404 = n2881 & n5403;
  assign n5405 = ~n2891 & n5404;
  assign n5406 = n4161 & n5405;
  assign n5407 = ~n5393 & n5406;
  assign n5408 = n5392 & n5407;
  assign n5409 = n5387 & n5408;
  assign n5410 = n2905 & n5409;
  assign n5411 = n2918 & n5410;
  assign n5412 = n4157 & n5411;
  assign n5413 = n5412 ^ n2084;
  assign n5414 = n5413 ^ x210;
  assign n5415 = ~n5384 & n5414;
  assign n5416 = n5383 & n5415;
  assign n5417 = n5350 & n5416;
  assign n5418 = ~n5348 & ~n5349;
  assign n5419 = ~n5384 & ~n5414;
  assign n5420 = n5383 & n5419;
  assign n5421 = n5418 & n5420;
  assign n5422 = ~n5417 & ~n5421;
  assign n5423 = n5348 & n5349;
  assign n5424 = ~n5351 & n5382;
  assign n5425 = n5415 & n5424;
  assign n5426 = n5423 & n5425;
  assign n5427 = n5384 & ~n5414;
  assign n5428 = n5424 & n5427;
  assign n5429 = n5350 & n5428;
  assign n5430 = n5384 & n5414;
  assign n5431 = ~n5351 & ~n5382;
  assign n5432 = n5430 & n5431;
  assign n5433 = n5419 & n5424;
  assign n5434 = ~n5432 & ~n5433;
  assign n5435 = n5423 & ~n5434;
  assign n5436 = n5424 & n5430;
  assign n5437 = ~n5348 & n5436;
  assign n5438 = ~n5435 & ~n5437;
  assign n5439 = ~n5429 & n5438;
  assign n5440 = ~n5418 & ~n5423;
  assign n5441 = n5428 & ~n5440;
  assign n5442 = n5427 & n5431;
  assign n5443 = ~n5425 & ~n5442;
  assign n5444 = n5350 & ~n5443;
  assign n5445 = ~n5441 & ~n5444;
  assign n5446 = n5418 & n5425;
  assign n5447 = n5350 & n5436;
  assign n5448 = ~n5446 & ~n5447;
  assign n5449 = ~n5348 & n5349;
  assign n5450 = n5351 & n5382;
  assign n5451 = n5415 & n5450;
  assign n5452 = n5427 & n5450;
  assign n5453 = ~n5451 & ~n5452;
  assign n5454 = ~n5416 & n5453;
  assign n5455 = n5449 & ~n5454;
  assign n5456 = n5415 & n5431;
  assign n5457 = n5418 & n5456;
  assign n5458 = n5383 & n5430;
  assign n5459 = n5430 & n5450;
  assign n5460 = n5419 & n5450;
  assign n5461 = ~n5459 & ~n5460;
  assign n5462 = ~n5458 & n5461;
  assign n5463 = n5350 & ~n5462;
  assign n5464 = ~n5457 & ~n5463;
  assign n5465 = n5419 & n5431;
  assign n5466 = ~n5432 & ~n5465;
  assign n5467 = ~n5420 & n5466;
  assign n5468 = ~n5459 & n5467;
  assign n5469 = n5449 & ~n5468;
  assign n5470 = n5383 & n5427;
  assign n5471 = ~n5451 & ~n5458;
  assign n5472 = ~n5423 & n5471;
  assign n5473 = ~n5416 & ~n5458;
  assign n5474 = n5418 & n5451;
  assign n5475 = ~n5460 & ~n5474;
  assign n5476 = n5473 & n5475;
  assign n5477 = ~n5472 & ~n5476;
  assign n5478 = ~n5470 & ~n5477;
  assign n5479 = ~n5440 & ~n5478;
  assign n5480 = ~n5469 & ~n5479;
  assign n5481 = n5464 & n5480;
  assign n5482 = ~n5455 & n5481;
  assign n5483 = n5448 & n5482;
  assign n5484 = n5445 & n5483;
  assign n5485 = n5439 & n5484;
  assign n5486 = ~n5426 & n5485;
  assign n5487 = n5422 & n5486;
  assign n5488 = n5487 ^ n2181;
  assign n5489 = n5488 ^ x281;
  assign n5490 = ~n5347 & n5489;
  assign n5491 = n5325 & n5490;
  assign n5492 = n5347 & ~n5489;
  assign n5493 = n5325 & n5492;
  assign n5494 = ~n5491 & ~n5493;
  assign n5495 = n4317 & n4361;
  assign n5496 = n4313 & n4333;
  assign n5497 = ~n5495 & ~n5496;
  assign n5498 = n4341 & ~n4941;
  assign n5499 = n4322 & n4942;
  assign n5500 = ~n4345 & n5499;
  assign n5501 = n4313 & ~n5500;
  assign n5502 = ~n5498 & ~n5501;
  assign n5503 = n4317 & ~n4937;
  assign n5504 = ~n4319 & n4329;
  assign n5505 = n4340 & ~n5504;
  assign n5506 = ~n4333 & ~n4337;
  assign n5507 = ~n4361 & n5506;
  assign n5508 = n4189 & ~n5507;
  assign n5509 = ~n5505 & ~n5508;
  assign n5510 = ~n5503 & n5509;
  assign n5511 = n5502 & n5510;
  assign n5512 = ~n4356 & n5511;
  assign n5513 = n5497 & n5512;
  assign n5514 = n4935 & n5513;
  assign n5515 = n4350 & n5514;
  assign n5516 = n4932 & n5515;
  assign n5517 = ~n4312 & n5516;
  assign n5518 = n5517 ^ n1626;
  assign n5519 = n5518 ^ x285;
  assign n5520 = n3637 & n3654;
  assign n5521 = n2936 & n3641;
  assign n5522 = n3637 & n3639;
  assign n5523 = ~n5521 & ~n5522;
  assign n5524 = n3641 & n3654;
  assign n5525 = n3657 & n3673;
  assign n5526 = ~n5524 & ~n5525;
  assign n5527 = ~n2935 & n3685;
  assign n5528 = ~n3658 & ~n3663;
  assign n5529 = n3639 & ~n5528;
  assign n5530 = ~n5527 & ~n5529;
  assign n5531 = ~n3672 & ~n3684;
  assign n5532 = n3654 & ~n5531;
  assign n5533 = ~n3642 & n3686;
  assign n5534 = ~n3672 & n5533;
  assign n5535 = n3639 & ~n5534;
  assign n5536 = n3670 & ~n3678;
  assign n5537 = n3654 & ~n5536;
  assign n5538 = ~n5535 & ~n5537;
  assign n5539 = ~n5532 & n5538;
  assign n5540 = n2936 & n3673;
  assign n5541 = ~n3648 & ~n3663;
  assign n5542 = n3657 & ~n5541;
  assign n5543 = ~n2936 & n5541;
  assign n5544 = ~n3651 & ~n3655;
  assign n5545 = ~n5543 & ~n5544;
  assign n5546 = ~n5542 & ~n5545;
  assign n5547 = ~n3666 & n5546;
  assign n5548 = ~n3642 & n5547;
  assign n5549 = ~n3633 & n5548;
  assign n5550 = n3664 & ~n5549;
  assign n5551 = ~n5540 & ~n5550;
  assign n5552 = n5539 & n5551;
  assign n5553 = n5530 & n5552;
  assign n5554 = n3681 & n5553;
  assign n5555 = n5526 & n5554;
  assign n5556 = n5523 & n5555;
  assign n5557 = ~n5520 & n5556;
  assign n5558 = ~n3669 & n5557;
  assign n5559 = n5558 ^ n1345;
  assign n5560 = n5559 ^ x280;
  assign n5561 = n5519 & ~n5560;
  assign n5562 = ~n5494 & n5561;
  assign n5563 = ~n5296 & ~n5324;
  assign n5564 = n5492 & n5563;
  assign n5565 = ~n5519 & n5560;
  assign n5566 = n5564 & n5565;
  assign n5567 = n5347 & n5489;
  assign n5568 = n5325 & n5567;
  assign n5569 = n5519 & n5560;
  assign n5570 = n5568 & n5569;
  assign n5571 = n5490 & n5563;
  assign n5572 = ~n5519 & ~n5560;
  assign n5573 = n5571 & n5572;
  assign n5574 = n5561 & n5564;
  assign n5575 = ~n5573 & ~n5574;
  assign n5576 = ~n5570 & n5575;
  assign n5577 = ~n5296 & n5324;
  assign n5578 = n5490 & n5577;
  assign n5579 = n5572 & n5578;
  assign n5580 = n5296 & ~n5324;
  assign n5581 = ~n5347 & ~n5489;
  assign n5582 = n5580 & n5581;
  assign n5583 = n5577 & n5581;
  assign n5584 = ~n5582 & ~n5583;
  assign n5585 = n5561 & ~n5584;
  assign n5586 = ~n5579 & ~n5585;
  assign n5587 = n5492 & n5577;
  assign n5588 = n5325 & n5581;
  assign n5589 = ~n5564 & ~n5588;
  assign n5590 = ~n5587 & n5589;
  assign n5591 = n5569 & ~n5590;
  assign n5592 = n5492 & n5580;
  assign n5593 = ~n5560 & n5592;
  assign n5594 = n5563 & n5567;
  assign n5595 = n5490 & n5580;
  assign n5596 = ~n5594 & ~n5595;
  assign n5597 = ~n5583 & n5596;
  assign n5598 = ~n5571 & n5597;
  assign n5599 = n5569 & ~n5598;
  assign n5600 = ~n5593 & ~n5599;
  assign n5601 = ~n5569 & ~n5572;
  assign n5602 = n5567 & n5577;
  assign n5603 = ~n5595 & ~n5602;
  assign n5604 = ~n5493 & ~n5582;
  assign n5605 = n5565 & ~n5604;
  assign n5606 = n5603 & ~n5605;
  assign n5607 = n5601 & ~n5606;
  assign n5608 = n5567 & n5580;
  assign n5609 = ~n5602 & ~n5608;
  assign n5610 = ~n5578 & n5609;
  assign n5611 = ~n5491 & n5610;
  assign n5612 = n5565 & ~n5611;
  assign n5613 = n5563 & n5581;
  assign n5614 = ~n5587 & ~n5608;
  assign n5615 = ~n5613 & n5614;
  assign n5616 = ~n5588 & n5615;
  assign n5617 = ~n5568 & n5616;
  assign n5618 = n5572 & ~n5617;
  assign n5619 = ~n5612 & ~n5618;
  assign n5620 = ~n5607 & n5619;
  assign n5621 = n5600 & n5620;
  assign n5622 = ~n5591 & n5621;
  assign n5623 = n5586 & n5622;
  assign n5624 = n5576 & n5623;
  assign n5625 = ~n5566 & n5624;
  assign n5626 = ~n5562 & n5625;
  assign n5627 = n5626 ^ n4646;
  assign n5628 = n5627 ^ x324;
  assign n5629 = ~n4827 & n4828;
  assign n5630 = ~n4834 & ~n4850;
  assign n5631 = n4716 & ~n5630;
  assign n5632 = ~n5629 & ~n5631;
  assign n5633 = ~n4796 & n4845;
  assign n5634 = n4817 & ~n5633;
  assign n5635 = ~n5180 & n5185;
  assign n5636 = ~n4825 & n5635;
  assign n5637 = n4827 & ~n5636;
  assign n5638 = ~n5634 & ~n5637;
  assign n5639 = n5632 & n5638;
  assign n5640 = n5328 & n5639;
  assign n5641 = n4824 & n5640;
  assign n5642 = n4816 & n5641;
  assign n5643 = n5169 & n5642;
  assign n5644 = n5643 ^ n3237;
  assign n5645 = n5644 ^ x273;
  assign n5646 = n4506 & ~n4552;
  assign n5647 = ~n4503 & ~n4533;
  assign n5648 = n4519 & ~n5647;
  assign n5649 = ~n5646 & ~n5648;
  assign n5650 = n4543 & ~n5069;
  assign n5651 = ~n4541 & n4552;
  assign n5652 = ~n4508 & n5651;
  assign n5653 = n4519 & ~n5652;
  assign n5654 = ~n5650 & ~n5653;
  assign n5655 = n4506 & n4546;
  assign n5656 = n4527 & n4556;
  assign n5657 = n5075 & n5656;
  assign n5658 = n4412 & ~n5657;
  assign n5659 = ~n4525 & ~n4541;
  assign n5660 = ~n4501 & n5659;
  assign n5661 = n4504 & ~n4508;
  assign n5662 = ~n4506 & n5661;
  assign n5663 = ~n5069 & ~n5662;
  assign n5664 = ~n5660 & n5663;
  assign n5665 = ~n4526 & ~n5663;
  assign n5666 = ~n4551 & n5665;
  assign n5667 = n4510 & ~n5666;
  assign n5668 = ~n5664 & ~n5667;
  assign n5669 = ~n5658 & n5668;
  assign n5670 = ~n5655 & n5669;
  assign n5671 = n5654 & n5670;
  assign n5672 = n4516 & n5671;
  assign n5673 = n5649 & n5672;
  assign n5674 = n5063 & n5673;
  assign n5675 = n5674 ^ n2688;
  assign n5676 = n5675 ^ x268;
  assign n5677 = ~n5645 & n5676;
  assign n5678 = n5010 & n5037;
  assign n5679 = ~n5009 & ~n5035;
  assign n5680 = n5678 & ~n5679;
  assign n5681 = n4985 & n5011;
  assign n5682 = n5001 & n5037;
  assign n5683 = ~n5681 & ~n5682;
  assign n5684 = ~n5007 & ~n5035;
  assign n5685 = ~n5683 & ~n5684;
  assign n5686 = ~n5014 & ~n5036;
  assign n5687 = n5007 & ~n5686;
  assign n5688 = n5009 & ~n5040;
  assign n5689 = ~n5687 & ~n5688;
  assign n5690 = ~n5685 & n5689;
  assign n5691 = ~n5030 & n5035;
  assign n5692 = n5025 & n5043;
  assign n5693 = ~n5691 & ~n5692;
  assign n5694 = n5690 & n5693;
  assign n5695 = n5022 & n5694;
  assign n5696 = ~n5680 & n5695;
  assign n5697 = n5696 ^ n3175;
  assign n5698 = n5697 ^ x272;
  assign n5699 = n5423 & n5436;
  assign n5700 = ~n5426 & ~n5699;
  assign n5701 = ~n5436 & ~n5458;
  assign n5702 = n5449 & ~n5701;
  assign n5703 = ~n5452 & ~n5459;
  assign n5704 = n5350 & ~n5703;
  assign n5705 = ~n5420 & ~n5460;
  assign n5706 = ~n5458 & n5705;
  assign n5707 = n5423 & ~n5706;
  assign n5708 = ~n5704 & ~n5707;
  assign n5709 = ~n5428 & ~n5433;
  assign n5710 = ~n5470 & n5709;
  assign n5711 = n5449 & ~n5710;
  assign n5712 = ~n5416 & n5461;
  assign n5713 = ~n5442 & n5712;
  assign n5714 = n5418 & ~n5713;
  assign n5715 = ~n5711 & ~n5714;
  assign n5716 = n5708 & n5715;
  assign n5717 = n5349 ^ n5348;
  assign n5718 = n5466 ^ n5456;
  assign n5719 = n5717 & ~n5718;
  assign n5720 = n5719 ^ n5456;
  assign n5721 = n5716 & ~n5720;
  assign n5722 = ~n5702 & n5721;
  assign n5723 = n5700 & n5722;
  assign n5724 = n5445 & n5723;
  assign n5725 = n5422 & n5724;
  assign n5726 = ~n5451 & n5725;
  assign n5727 = n5726 ^ n2528;
  assign n5728 = n5727 ^ x269;
  assign n5729 = ~n5698 & n5728;
  assign n5730 = n4617 & n5146;
  assign n5731 = n4613 & n5136;
  assign n5732 = ~n4649 & ~n4685;
  assign n5733 = ~n5135 & n5732;
  assign n5734 = n4673 & ~n5733;
  assign n5735 = ~n5731 & ~n5734;
  assign n5736 = ~n5730 & n5735;
  assign n5737 = n4656 & ~n5151;
  assign n5738 = n4614 & n5156;
  assign n5739 = ~n5737 & ~n5738;
  assign n5740 = n5736 & n5739;
  assign n5741 = n5282 & n5740;
  assign n5742 = n5741 ^ n3868;
  assign n5743 = n5742 ^ x270;
  assign n5744 = ~n4096 & ~n4114;
  assign n5745 = n4085 & ~n5744;
  assign n5746 = ~n4120 & n5301;
  assign n5747 = n4086 & ~n5746;
  assign n5748 = ~n5745 & ~n5747;
  assign n5749 = ~n3741 & n4088;
  assign n5750 = n4082 & n4116;
  assign n5751 = ~n4121 & n5750;
  assign n5752 = n4090 & ~n5751;
  assign n5753 = ~n5749 & ~n5752;
  assign n5754 = n5748 & n5753;
  assign n5755 = n4077 & n4115;
  assign n5756 = n4098 & ~n4107;
  assign n5757 = n4100 & ~n5756;
  assign n5758 = ~n4107 & n5121;
  assign n5759 = ~n4085 & n5758;
  assign n5760 = ~n4107 & n4122;
  assign n5761 = n4077 & ~n5760;
  assign n5762 = n5116 & ~n5761;
  assign n5763 = n5301 & n5762;
  assign n5764 = ~n5759 & ~n5763;
  assign n5765 = ~n4086 & n5764;
  assign n5766 = ~n5757 & ~n5765;
  assign n5767 = ~n5755 & n5766;
  assign n5768 = n5754 & n5767;
  assign n5769 = n5103 & n5768;
  assign n5770 = n5769 ^ n3899;
  assign n5771 = n5770 ^ x271;
  assign n5772 = ~n5743 & ~n5771;
  assign n5773 = n5729 & n5772;
  assign n5774 = n5677 & n5773;
  assign n5775 = ~n5743 & n5771;
  assign n5776 = n5698 & n5775;
  assign n5777 = n5728 & n5776;
  assign n5778 = n5677 & n5777;
  assign n5779 = n5698 & n5743;
  assign n5780 = ~n5771 & n5779;
  assign n5781 = ~n5728 & n5780;
  assign n5782 = n5645 & ~n5676;
  assign n5783 = n5781 & n5782;
  assign n5784 = ~n5778 & ~n5783;
  assign n5785 = ~n5774 & n5784;
  assign n5786 = n5645 & n5676;
  assign n5787 = n5777 & n5786;
  assign n5788 = n5729 & n5771;
  assign n5789 = ~n5743 & n5788;
  assign n5790 = n5771 & n5779;
  assign n5791 = n5728 & n5790;
  assign n5792 = ~n5789 & ~n5791;
  assign n5793 = n5677 & ~n5792;
  assign n5794 = ~n5787 & ~n5793;
  assign n5795 = ~n5728 & n5771;
  assign n5796 = ~n5743 & n5795;
  assign n5797 = ~n5698 & n5796;
  assign n5798 = n5698 & n5772;
  assign n5799 = ~n5728 & n5798;
  assign n5800 = n5743 & ~n5771;
  assign n5801 = ~n5698 & n5800;
  assign n5802 = ~n5728 & n5801;
  assign n5803 = ~n5799 & ~n5802;
  assign n5804 = ~n5797 & n5803;
  assign n5805 = n5782 & ~n5804;
  assign n5806 = ~n5645 & ~n5676;
  assign n5807 = n5779 & n5795;
  assign n5808 = ~n5791 & ~n5807;
  assign n5809 = n5698 & n5796;
  assign n5810 = ~n5698 & n5772;
  assign n5811 = ~n5728 & n5810;
  assign n5812 = ~n5809 & ~n5811;
  assign n5813 = n5808 & n5812;
  assign n5814 = ~n5797 & n5813;
  assign n5815 = n5806 & ~n5814;
  assign n5816 = ~n5805 & ~n5815;
  assign n5817 = ~n5786 & ~n5806;
  assign n5818 = n5728 & n5798;
  assign n5819 = n5743 & n5788;
  assign n5820 = n5728 & n5780;
  assign n5821 = ~n5819 & ~n5820;
  assign n5822 = ~n5818 & n5821;
  assign n5823 = ~n5817 & ~n5822;
  assign n5824 = n5729 & ~n5800;
  assign n5825 = n5792 & ~n5824;
  assign n5826 = n5782 & ~n5825;
  assign n5827 = ~n5823 & ~n5826;
  assign n5828 = n5729 & n5800;
  assign n5829 = n5743 & n5795;
  assign n5830 = ~n5698 & n5829;
  assign n5831 = ~n5809 & ~n5830;
  assign n5832 = ~n5828 & n5831;
  assign n5833 = ~n5811 & n5832;
  assign n5834 = n5786 & ~n5833;
  assign n5835 = ~n5799 & ~n5830;
  assign n5836 = ~n5781 & n5835;
  assign n5837 = ~n5802 & n5836;
  assign n5838 = n5677 & ~n5837;
  assign n5839 = ~n5834 & ~n5838;
  assign n5840 = n5827 & n5839;
  assign n5841 = n5816 & n5840;
  assign n5842 = n5794 & n5841;
  assign n5843 = n5785 & n5842;
  assign n5844 = n5843 ^ n4410;
  assign n5845 = n5844 ^ x326;
  assign n5846 = n5161 ^ x303;
  assign n5847 = n4863 ^ x298;
  assign n5848 = n5846 & ~n5847;
  assign n5849 = ~n5442 & ~n5456;
  assign n5850 = n5350 & ~n5849;
  assign n5851 = n5418 & ~n5709;
  assign n5852 = ~n5850 & ~n5851;
  assign n5853 = ~n5433 & n5443;
  assign n5854 = n5449 & ~n5853;
  assign n5855 = n5453 & n5705;
  assign n5856 = n5350 & ~n5855;
  assign n5857 = ~n5854 & ~n5856;
  assign n5858 = ~n5432 & n5473;
  assign n5859 = ~n5459 & n5858;
  assign n5860 = n5418 & ~n5859;
  assign n5861 = n5461 & ~n5470;
  assign n5862 = n5467 & n5861;
  assign n5863 = n5423 & ~n5862;
  assign n5864 = ~n5860 & ~n5863;
  assign n5865 = n5857 & n5864;
  assign n5866 = ~n5702 & n5865;
  assign n5867 = ~n5455 & n5866;
  assign n5868 = n5448 & n5867;
  assign n5869 = n5700 & n5868;
  assign n5870 = n5852 & n5869;
  assign n5871 = n5422 & n5870;
  assign n5872 = n5871 ^ n3765;
  assign n5873 = n5872 ^ x301;
  assign n5874 = n5057 ^ x302;
  assign n5875 = n5873 & ~n5874;
  assign n5876 = n4136 ^ x299;
  assign n5877 = n3633 & n3657;
  assign n5878 = n2936 & ~n3670;
  assign n5879 = ~n5877 & ~n5878;
  assign n5880 = n2496 & n3648;
  assign n5881 = n3651 & n3664;
  assign n5882 = ~n5880 & ~n5881;
  assign n5883 = n3654 & n3666;
  assign n5884 = n3657 & n3678;
  assign n5885 = n3643 & ~n3673;
  assign n5886 = n3657 & ~n5885;
  assign n5887 = ~n3663 & ~n3668;
  assign n5888 = n2936 & ~n5887;
  assign n5889 = ~n5886 & ~n5888;
  assign n5890 = ~n3633 & ~n3685;
  assign n5891 = n3654 & ~n5890;
  assign n5892 = ~n3648 & n3674;
  assign n5893 = n3639 & ~n5892;
  assign n5894 = ~n5891 & ~n5893;
  assign n5895 = n5889 & n5894;
  assign n5896 = n3676 & n5895;
  assign n5897 = ~n3669 & n5896;
  assign n5898 = ~n5884 & n5897;
  assign n5899 = ~n5883 & n5898;
  assign n5900 = n5882 & n5899;
  assign n5901 = n3645 & n5900;
  assign n5902 = n5523 & n5901;
  assign n5903 = n5879 & n5902;
  assign n5904 = ~n5520 & n5903;
  assign n5905 = ~n3655 & n5904;
  assign n5906 = n5905 ^ n3793;
  assign n5907 = n5906 ^ x300;
  assign n5908 = ~n5876 & n5907;
  assign n5909 = n5875 & n5908;
  assign n5910 = ~n5873 & n5874;
  assign n5911 = n5908 & n5910;
  assign n5912 = ~n5909 & ~n5911;
  assign n5913 = n5848 & ~n5912;
  assign n5914 = ~n5846 & ~n5847;
  assign n5915 = n5873 & n5874;
  assign n5916 = n5876 & n5907;
  assign n5917 = n5915 & n5916;
  assign n5918 = n5876 & ~n5907;
  assign n5919 = n5875 & n5918;
  assign n5920 = ~n5917 & ~n5919;
  assign n5921 = n5914 & ~n5920;
  assign n5922 = ~n5913 & ~n5921;
  assign n5923 = ~n5873 & ~n5874;
  assign n5924 = n5916 & n5923;
  assign n5925 = n5847 & n5924;
  assign n5926 = n5908 & n5923;
  assign n5927 = ~n5876 & ~n5907;
  assign n5928 = n5910 & n5927;
  assign n5929 = ~n5926 & ~n5928;
  assign n5930 = n5848 & ~n5929;
  assign n5931 = ~n5925 & ~n5930;
  assign n5932 = n5915 & n5918;
  assign n5933 = n5914 & n5932;
  assign n5934 = ~n5846 & n5847;
  assign n5935 = n5910 & n5918;
  assign n5936 = n5910 & n5916;
  assign n5937 = ~n5919 & ~n5936;
  assign n5938 = ~n5935 & n5937;
  assign n5939 = n5934 & ~n5938;
  assign n5940 = ~n5933 & ~n5939;
  assign n5941 = n5931 & n5940;
  assign n5942 = n5847 ^ n5846;
  assign n5943 = n5918 & n5923;
  assign n5944 = ~n5942 & n5943;
  assign n5945 = n5846 & n5847;
  assign n5946 = n5875 & n5916;
  assign n5947 = ~n5917 & ~n5946;
  assign n5948 = n5945 & ~n5947;
  assign n5949 = n5914 & ~n5929;
  assign n5950 = n5908 & n5915;
  assign n5951 = n5934 & n5950;
  assign n5952 = n5848 & n5917;
  assign n5953 = ~n5951 & ~n5952;
  assign n5954 = ~n5912 & n5914;
  assign n5955 = n5923 & n5927;
  assign n5956 = ~n5909 & ~n5928;
  assign n5957 = ~n5955 & n5956;
  assign n5958 = n5934 & ~n5957;
  assign n5959 = ~n5954 & ~n5958;
  assign n5960 = ~n5932 & n5937;
  assign n5961 = n5848 & ~n5960;
  assign n5962 = n5915 & n5927;
  assign n5963 = n5875 & n5927;
  assign n5964 = ~n5911 & ~n5955;
  assign n5965 = ~n5963 & n5964;
  assign n5966 = ~n5962 & n5965;
  assign n5967 = n5945 & ~n5966;
  assign n5968 = ~n5961 & ~n5967;
  assign n5969 = n5959 & n5968;
  assign n5970 = n5953 & n5969;
  assign n5971 = ~n5949 & n5970;
  assign n5972 = ~n5948 & n5971;
  assign n5973 = ~n5944 & n5972;
  assign n5974 = n5941 & n5973;
  assign n5975 = n5922 & n5974;
  assign n5976 = n5975 ^ n4608;
  assign n5977 = n5976 ^ x325;
  assign n5978 = n5845 & n5977;
  assign n5979 = ~n5628 & n5978;
  assign n5980 = n5727 ^ x267;
  assign n5981 = n5132 ^ x262;
  assign n5982 = n5980 & ~n5981;
  assign n5983 = n3648 & ~n3664;
  assign n5984 = n2496 & ~n3674;
  assign n5985 = ~n5983 & ~n5984;
  assign n5986 = n3664 & n3685;
  assign n5987 = ~n3655 & ~n3672;
  assign n5988 = n3657 & ~n5987;
  assign n5989 = ~n5986 & ~n5988;
  assign n5990 = ~n3668 & ~n3684;
  assign n5991 = n3639 & ~n5990;
  assign n5992 = ~n3651 & n5528;
  assign n5993 = ~n2935 & ~n5992;
  assign n5994 = ~n5991 & ~n5993;
  assign n5995 = n5989 & n5994;
  assign n5996 = n5985 & n5995;
  assign n5997 = ~n5522 & n5996;
  assign n5998 = n5526 & n5997;
  assign n5999 = n5879 & n5998;
  assign n6000 = n3646 & n5999;
  assign n6001 = n3682 & n6000;
  assign n6002 = ~n5520 & n6001;
  assign n6003 = n6002 ^ n2861;
  assign n6004 = n6003 ^ x264;
  assign n6005 = n5675 ^ x266;
  assign n6006 = n4961 ^ x263;
  assign n6007 = n5007 & n5012;
  assign n6008 = n5007 & n5038;
  assign n6009 = n5017 & ~n5035;
  assign n6010 = ~n6008 & ~n6009;
  assign n6011 = ~n5015 & n5025;
  assign n6012 = ~n5007 & ~n5025;
  assign n6013 = n5003 & ~n6012;
  assign n6014 = n4985 & n5026;
  assign n6015 = n5035 & n6014;
  assign n6016 = n5013 & ~n5679;
  assign n6017 = n4999 & n6016;
  assign n6018 = ~n6015 & ~n6017;
  assign n6019 = n5009 & n5014;
  assign n6020 = ~n5018 & ~n5029;
  assign n6021 = ~n5036 & n6020;
  assign n6022 = n5035 & ~n6021;
  assign n6023 = ~n6019 & ~n6022;
  assign n6024 = ~n5023 & ~n5027;
  assign n6025 = ~n5009 & n6024;
  assign n6026 = n6012 & ~n6014;
  assign n6027 = ~n5036 & n6026;
  assign n6028 = ~n6025 & ~n6027;
  assign n6029 = ~n5682 & ~n6028;
  assign n6030 = ~n5035 & ~n6029;
  assign n6031 = n6023 & ~n6030;
  assign n6032 = n6018 & n6031;
  assign n6033 = ~n6013 & n6032;
  assign n6034 = ~n6011 & n6033;
  assign n6035 = n6010 & n6034;
  assign n6036 = ~n6007 & n6035;
  assign n6037 = ~n5680 & n6036;
  assign n6038 = n6037 ^ n2825;
  assign n6039 = n6038 ^ x265;
  assign n6040 = ~n6006 & ~n6039;
  assign n6041 = n6005 & n6040;
  assign n6042 = n6004 & n6041;
  assign n6043 = ~n6004 & ~n6005;
  assign n6044 = ~n6006 & n6043;
  assign n6045 = ~n6039 & n6044;
  assign n6046 = ~n6042 & ~n6045;
  assign n6047 = n5982 & ~n6046;
  assign n6048 = n5980 & n5981;
  assign n6049 = n6006 & ~n6039;
  assign n6050 = n6004 & ~n6005;
  assign n6051 = n6049 & n6050;
  assign n6052 = n6048 & n6051;
  assign n6053 = ~n5980 & ~n5981;
  assign n6054 = n6006 & n6039;
  assign n6055 = n6043 & n6054;
  assign n6056 = n6005 & n6049;
  assign n6057 = n6004 & n6056;
  assign n6058 = ~n6055 & ~n6057;
  assign n6059 = n6053 & ~n6058;
  assign n6060 = ~n6052 & ~n6059;
  assign n6061 = ~n6047 & n6060;
  assign n6062 = n5981 & n6057;
  assign n6063 = ~n6004 & n6056;
  assign n6064 = ~n6055 & ~n6063;
  assign n6065 = n6048 & ~n6064;
  assign n6066 = ~n6062 & ~n6065;
  assign n6067 = n6050 & n6054;
  assign n6068 = ~n6063 & ~n6067;
  assign n6069 = n6053 & ~n6068;
  assign n6070 = ~n6006 & n6039;
  assign n6071 = n6005 & n6070;
  assign n6072 = ~n6004 & n6071;
  assign n6073 = n6039 & n6044;
  assign n6074 = ~n6072 & ~n6073;
  assign n6075 = n5982 & ~n6074;
  assign n6076 = n6050 & n6070;
  assign n6077 = n6048 & n6076;
  assign n6078 = ~n5980 & n5981;
  assign n6079 = ~n6046 & n6078;
  assign n6080 = ~n6077 & ~n6079;
  assign n6081 = n6004 & n6071;
  assign n6082 = n6048 & n6081;
  assign n6083 = n6078 & n6081;
  assign n6084 = n5982 & ~n6064;
  assign n6085 = ~n6083 & ~n6084;
  assign n6086 = ~n6004 & n6041;
  assign n6087 = ~n6076 & ~n6086;
  assign n6088 = n6053 & ~n6087;
  assign n6089 = n6040 & n6050;
  assign n6090 = ~n6072 & ~n6089;
  assign n6091 = n6048 & ~n6090;
  assign n6092 = ~n6081 & ~n6089;
  assign n6093 = n6053 & ~n6092;
  assign n6094 = n6005 & n6054;
  assign n6095 = n6004 & n6094;
  assign n6096 = ~n6051 & ~n6095;
  assign n6097 = n5982 & ~n6096;
  assign n6098 = ~n6004 & n6094;
  assign n6099 = ~n6067 & ~n6098;
  assign n6100 = ~n6005 & n6049;
  assign n6101 = ~n6004 & n6100;
  assign n6102 = ~n6073 & ~n6101;
  assign n6103 = n6099 & n6102;
  assign n6104 = n6078 & ~n6103;
  assign n6105 = ~n6097 & ~n6104;
  assign n6106 = ~n6093 & n6105;
  assign n6107 = ~n6091 & n6106;
  assign n6108 = ~n6088 & n6107;
  assign n6109 = n6085 & n6108;
  assign n6110 = ~n6082 & n6109;
  assign n6111 = n6080 & n6110;
  assign n6112 = ~n6075 & n6111;
  assign n6113 = ~n6069 & n6112;
  assign n6114 = n6066 & n6113;
  assign n6115 = n6061 & n6114;
  assign n6116 = n6115 ^ n2934;
  assign n6117 = n6116 ^ x323;
  assign n6118 = n5977 & n6117;
  assign n6119 = n5628 & n6118;
  assign n6120 = ~n5845 & ~n5977;
  assign n6121 = ~n6117 & n6120;
  assign n6122 = ~n6119 & ~n6121;
  assign n6123 = ~n5979 & n6122;
  assign n6124 = n6117 ^ n5628;
  assign n6125 = ~n5977 & ~n6124;
  assign n6126 = n5845 & n6125;
  assign n6127 = n6123 & ~n6126;
  assign n6128 = n5277 & n6127;
  assign n6129 = ~n4929 & ~n5276;
  assign n6130 = ~n5628 & ~n5977;
  assign n6131 = ~n5845 & n6130;
  assign n6132 = n5979 & n6117;
  assign n6133 = ~n6131 & ~n6132;
  assign n6134 = n5628 & ~n5977;
  assign n6135 = n5845 & n6134;
  assign n6136 = ~n6117 & n6135;
  assign n6137 = n6133 & ~n6136;
  assign n6138 = n5977 & n6124;
  assign n6139 = ~n5845 & n6138;
  assign n6140 = n6137 & ~n6139;
  assign n6141 = ~n6126 & n6140;
  assign n6142 = n6129 & ~n6141;
  assign n6143 = ~n6128 & ~n6142;
  assign n6144 = n4929 & n5276;
  assign n6145 = n5977 ^ n5845;
  assign n6146 = n5628 & ~n6145;
  assign n6147 = n6117 & n6146;
  assign n6148 = n5845 ^ n5628;
  assign n6149 = n6134 & n6148;
  assign n6150 = n6149 ^ n6148;
  assign n6151 = ~n6117 & n6150;
  assign n6152 = ~n6131 & ~n6151;
  assign n6153 = ~n5979 & n6152;
  assign n6154 = ~n6147 & n6153;
  assign n6155 = n6144 & ~n6154;
  assign n6156 = n4929 & ~n5276;
  assign n6158 = ~n5628 & ~n6117;
  assign n6157 = n6130 ^ n6117;
  assign n6159 = n6158 ^ n6157;
  assign n6160 = n5845 & ~n6159;
  assign n6161 = n6160 ^ n6158;
  assign n6162 = ~n6147 & ~n6161;
  assign n6163 = n6156 & ~n6162;
  assign n6164 = ~n6155 & ~n6163;
  assign n6165 = n6143 & n6164;
  assign n6166 = n6165 ^ n4695;
  assign n6167 = n6166 ^ x390;
  assign n6168 = n5844 ^ x328;
  assign n6169 = n5848 & n5924;
  assign n6170 = n5953 & ~n6169;
  assign n6171 = n5945 & ~n5964;
  assign n6172 = ~n5926 & ~n5962;
  assign n6173 = n5848 & ~n6172;
  assign n6174 = ~n6171 & ~n6173;
  assign n6175 = n5926 & n5945;
  assign n6176 = ~n5912 & n5934;
  assign n6177 = ~n6175 & ~n6176;
  assign n6178 = ~n5848 & n5963;
  assign n6179 = ~n5932 & ~n5946;
  assign n6180 = ~n5936 & ~n5962;
  assign n6181 = n6179 & n6180;
  assign n6182 = ~n5943 & n6181;
  assign n6183 = n5914 & ~n6182;
  assign n6184 = n5937 & ~n5950;
  assign n6185 = ~n5943 & n6184;
  assign n6186 = n5848 & ~n6185;
  assign n6187 = ~n5909 & n6179;
  assign n6188 = n5945 & ~n6187;
  assign n6189 = ~n5934 & ~n5935;
  assign n6190 = ~n5935 & ~n5943;
  assign n6191 = n5920 & n6190;
  assign n6192 = ~n6189 & ~n6191;
  assign n6193 = ~n6188 & ~n6192;
  assign n6194 = n5847 & ~n6193;
  assign n6195 = ~n6186 & ~n6194;
  assign n6196 = ~n6183 & n6195;
  assign n6197 = ~n6178 & n6196;
  assign n6198 = n6177 & n6197;
  assign n6199 = n6174 & n6198;
  assign n6200 = ~n5949 & n6199;
  assign n6201 = n6170 & n6200;
  assign n6202 = n6201 ^ n3856;
  assign n6203 = n6202 ^ x333;
  assign n6204 = ~n6168 & ~n6203;
  assign n6205 = n5697 ^ x274;
  assign n6206 = n5488 ^ x279;
  assign n6207 = n6205 & ~n6206;
  assign n6208 = n4345 & ~n4941;
  assign n6209 = n4340 & ~n4358;
  assign n6210 = ~n6208 & ~n6209;
  assign n6211 = n4313 & ~n4338;
  assign n6212 = ~n4347 & n4942;
  assign n6213 = n4317 & ~n6212;
  assign n6214 = ~n6211 & ~n6213;
  assign n6215 = ~n4326 & ~n4328;
  assign n6216 = n4189 & ~n6215;
  assign n6217 = ~n4319 & ~n4341;
  assign n6218 = n4189 & ~n6217;
  assign n6219 = ~n4327 & ~n4354;
  assign n6220 = n4313 & ~n6219;
  assign n6221 = ~n6218 & ~n6220;
  assign n6222 = n4340 & ~n4936;
  assign n6223 = ~n4310 & n4342;
  assign n6224 = n4317 & ~n6223;
  assign n6225 = ~n6222 & ~n6224;
  assign n6226 = n6221 & n6225;
  assign n6227 = n4932 & n6226;
  assign n6228 = ~n4312 & n6227;
  assign n6229 = ~n6216 & n6228;
  assign n6230 = n6214 & n6229;
  assign n6231 = n6210 & n6230;
  assign n6232 = n5497 & n6231;
  assign n6233 = n4353 & n6232;
  assign n6234 = n6233 ^ n3265;
  assign n6235 = n6234 ^ x277;
  assign n6236 = ~n4379 & n4543;
  assign n6237 = ~n4513 & n4556;
  assign n6238 = n4506 & ~n6237;
  assign n6239 = ~n6236 & ~n6238;
  assign n6240 = n4529 & n5061;
  assign n6241 = n4510 & ~n6240;
  assign n6242 = n5076 & n5659;
  assign n6243 = n4412 & ~n6242;
  assign n6244 = n5075 & n5660;
  assign n6245 = ~n4537 & n6244;
  assign n6246 = n4519 & ~n6245;
  assign n6247 = ~n6243 & ~n6246;
  assign n6248 = ~n6241 & n6247;
  assign n6249 = n6239 & n6248;
  assign n6250 = n5649 & n6249;
  assign n6251 = n4517 & n6250;
  assign n6252 = ~n4540 & n6251;
  assign n6253 = n6252 ^ n3204;
  assign n6254 = n6253 ^ x276;
  assign n6255 = n5644 ^ x275;
  assign n6256 = n5559 ^ x278;
  assign n6257 = ~n6255 & ~n6256;
  assign n6258 = n6254 & n6257;
  assign n6259 = ~n6235 & n6258;
  assign n6260 = n6256 ^ n6235;
  assign n6261 = n6255 & ~n6260;
  assign n6262 = ~n6254 & n6261;
  assign n6263 = ~n6259 & ~n6262;
  assign n6264 = ~n6235 & ~n6256;
  assign n6265 = n6235 ^ x276;
  assign n6266 = n6265 ^ n6253;
  assign n6267 = n6264 & ~n6266;
  assign n6268 = n6267 ^ n6266;
  assign n6269 = ~n6255 & ~n6268;
  assign n6270 = n6254 & n6256;
  assign n6271 = n6235 & n6270;
  assign n6272 = n6255 & n6264;
  assign n6273 = n6254 & n6272;
  assign n6274 = ~n6271 & ~n6273;
  assign n6275 = ~n6269 & n6274;
  assign n6276 = n6263 & n6275;
  assign n6277 = n6207 & n6276;
  assign n6278 = ~n6205 & ~n6206;
  assign n6279 = n6235 & n6255;
  assign n6280 = ~n6256 & n6279;
  assign n6281 = ~n6254 & n6280;
  assign n6282 = n6235 & n6256;
  assign n6283 = ~n6255 & n6282;
  assign n6284 = ~n6235 & ~n6270;
  assign n6285 = n6255 & n6284;
  assign n6286 = ~n6258 & ~n6285;
  assign n6287 = ~n6283 & n6286;
  assign n6288 = ~n6281 & n6287;
  assign n6289 = n6278 & ~n6288;
  assign n6290 = ~n6277 & ~n6289;
  assign n6291 = n6205 & n6206;
  assign n6292 = ~n6255 & n6270;
  assign n6293 = n6254 & n6280;
  assign n6294 = ~n6292 & ~n6293;
  assign n6295 = ~n6254 & n6257;
  assign n6296 = n6263 & ~n6295;
  assign n6297 = n6294 & n6296;
  assign n6298 = n6291 & ~n6297;
  assign n6299 = ~n6205 & n6206;
  assign n6300 = n6255 & n6270;
  assign n6301 = n6235 & n6257;
  assign n6302 = n6275 & ~n6301;
  assign n6303 = ~n6300 & n6302;
  assign n6304 = ~n6281 & n6303;
  assign n6305 = n6299 & ~n6304;
  assign n6306 = ~n6298 & ~n6305;
  assign n6307 = n6290 & n6306;
  assign n6308 = n6307 ^ n4075;
  assign n6309 = n6308 ^ x332;
  assign n6310 = n5295 ^ x286;
  assign n6311 = n4570 ^ x291;
  assign n6312 = n6310 & n6311;
  assign n6313 = n5518 ^ x287;
  assign n6314 = ~n5035 & n5036;
  assign n6315 = n5678 & ~n5684;
  assign n6316 = ~n6314 & ~n6315;
  assign n6317 = ~n5023 & ~n5682;
  assign n6318 = n5007 & ~n6317;
  assign n6319 = ~n5003 & n5683;
  assign n6320 = n5025 & ~n6319;
  assign n6321 = n4985 & n5037;
  assign n6322 = n5004 & ~n6321;
  assign n6323 = ~n5018 & n6322;
  assign n6324 = n5009 & ~n6323;
  assign n6325 = ~n6320 & ~n6324;
  assign n6326 = n5015 & n6317;
  assign n6327 = n5035 & ~n6326;
  assign n6328 = ~n5011 & ~n5025;
  assign n6329 = ~n5678 & ~n6007;
  assign n6330 = ~n5029 & n6329;
  assign n6331 = ~n5017 & n6330;
  assign n6332 = ~n6328 & ~n6331;
  assign n6333 = ~n6012 & n6332;
  assign n6334 = ~n6327 & ~n6333;
  assign n6335 = n6325 & n6334;
  assign n6336 = n5021 & n6335;
  assign n6337 = n6018 & n6336;
  assign n6338 = ~n6318 & n6337;
  assign n6339 = n6316 & n6338;
  assign n6340 = n6339 ^ n3559;
  assign n6341 = n6340 ^ x288;
  assign n6342 = n6313 & ~n6341;
  assign n6343 = n3700 ^ x290;
  assign n6344 = n5423 & n5456;
  assign n6345 = n5461 & n5473;
  assign n6346 = ~n5425 & n6345;
  assign n6347 = ~n5428 & n6346;
  assign n6348 = n5449 & ~n6347;
  assign n6349 = ~n6344 & ~n6348;
  assign n6350 = n5465 & n5717;
  assign n6351 = ~n5451 & n5861;
  assign n6352 = n5350 & ~n6351;
  assign n6353 = ~n5420 & ~n5459;
  assign n6354 = ~n5458 & n6353;
  assign n6355 = ~n5418 & n6354;
  assign n6356 = n5453 & n5473;
  assign n6357 = ~n5423 & n6356;
  assign n6358 = ~n6355 & ~n6357;
  assign n6359 = ~n5442 & ~n6358;
  assign n6360 = ~n5440 & ~n6359;
  assign n6361 = ~n6352 & ~n6360;
  assign n6362 = ~n6350 & n6361;
  assign n6363 = n6349 & n6362;
  assign n6364 = n5852 & n6363;
  assign n6365 = n5439 & n6364;
  assign n6366 = ~n5426 & n6365;
  assign n6367 = n6366 ^ n3533;
  assign n6368 = n6367 ^ x289;
  assign n6369 = n6343 & ~n6368;
  assign n6370 = n6342 & n6369;
  assign n6371 = n6312 & n6370;
  assign n6372 = ~n6310 & ~n6311;
  assign n6373 = n6313 & n6341;
  assign n6374 = ~n6343 & ~n6368;
  assign n6375 = n6373 & n6374;
  assign n6376 = n6372 & n6375;
  assign n6377 = ~n6371 & ~n6376;
  assign n6378 = ~n6313 & n6341;
  assign n6379 = n6343 & n6368;
  assign n6380 = n6378 & n6379;
  assign n6381 = n6374 & n6378;
  assign n6382 = ~n6380 & ~n6381;
  assign n6383 = n6312 & ~n6382;
  assign n6384 = n6310 & ~n6311;
  assign n6385 = ~n6343 & n6368;
  assign n6386 = n6373 & n6385;
  assign n6387 = n6369 & n6373;
  assign n6388 = ~n6386 & ~n6387;
  assign n6389 = n6384 & ~n6388;
  assign n6390 = ~n6383 & ~n6389;
  assign n6391 = n6373 & n6379;
  assign n6392 = n6384 & n6391;
  assign n6393 = n6312 & ~n6388;
  assign n6394 = ~n6392 & ~n6393;
  assign n6395 = n6342 & n6385;
  assign n6396 = ~n6372 & n6395;
  assign n6397 = n6378 & n6385;
  assign n6398 = ~n6313 & ~n6341;
  assign n6399 = n6369 & n6398;
  assign n6400 = ~n6397 & ~n6399;
  assign n6401 = n6312 & ~n6400;
  assign n6402 = ~n6396 & ~n6401;
  assign n6403 = n6342 & n6374;
  assign n6404 = ~n6310 & n6403;
  assign n6405 = ~n6310 & n6311;
  assign n6406 = ~n6381 & ~n6399;
  assign n6407 = ~n6391 & ~n6397;
  assign n6408 = n6342 & n6379;
  assign n6409 = n6369 & n6378;
  assign n6410 = ~n6408 & ~n6409;
  assign n6411 = n6407 & n6410;
  assign n6412 = n6406 & n6411;
  assign n6413 = n6405 & ~n6412;
  assign n6414 = ~n6404 & ~n6413;
  assign n6415 = n6372 & ~n6388;
  assign n6416 = n6379 & n6398;
  assign n6417 = n6374 & n6398;
  assign n6418 = n6385 & n6398;
  assign n6419 = ~n6380 & ~n6418;
  assign n6420 = ~n6417 & n6419;
  assign n6421 = ~n6384 & n6420;
  assign n6422 = ~n6370 & n6406;
  assign n6423 = ~n6372 & n6422;
  assign n6424 = ~n6421 & ~n6423;
  assign n6425 = ~n6416 & ~n6424;
  assign n6426 = ~n6311 & ~n6425;
  assign n6427 = ~n6415 & ~n6426;
  assign n6428 = n6414 & n6427;
  assign n6429 = n6402 & n6428;
  assign n6430 = n6394 & n6429;
  assign n6431 = n6390 & n6430;
  assign n6432 = n6377 & n6431;
  assign n6433 = n6432 ^ n4471;
  assign n6434 = n6433 ^ x331;
  assign n6435 = ~n6309 & ~n6434;
  assign n6436 = n5275 ^ x329;
  assign n6437 = n6078 & n6089;
  assign n6438 = ~n6073 & ~n6086;
  assign n6439 = n6048 & ~n6438;
  assign n6440 = ~n6437 & ~n6439;
  assign n6441 = n5982 & n6076;
  assign n6442 = ~n6064 & n6078;
  assign n6443 = ~n6441 & ~n6442;
  assign n6444 = n6048 & n6063;
  assign n6445 = n6078 & n6086;
  assign n6446 = ~n6444 & ~n6445;
  assign n6447 = n5981 & ~n6099;
  assign n6448 = n6074 & n6096;
  assign n6449 = n6053 & ~n6448;
  assign n6450 = ~n6042 & ~n6073;
  assign n6451 = ~n6098 & n6450;
  assign n6452 = ~n6100 & n6451;
  assign n6453 = ~n6063 & n6452;
  assign n6454 = ~n6081 & n6453;
  assign n6455 = n5982 & ~n6454;
  assign n6456 = ~n6449 & ~n6455;
  assign n6457 = ~n6447 & n6456;
  assign n6458 = n6446 & n6457;
  assign n6459 = n6060 & n6458;
  assign n6460 = ~n6093 & n6459;
  assign n6461 = n6443 & n6460;
  assign n6462 = n6440 & n6461;
  assign n6463 = ~n6082 & n6462;
  assign n6464 = n6080 & n6463;
  assign n6465 = n6464 ^ n4444;
  assign n6466 = n6465 ^ x330;
  assign n6467 = n6436 & ~n6466;
  assign n6468 = n6435 & n6467;
  assign n6469 = n6204 & n6468;
  assign n6470 = ~n6168 & n6203;
  assign n6471 = ~n6436 & ~n6466;
  assign n6472 = n6435 & n6471;
  assign n6473 = n6470 & n6472;
  assign n6474 = ~n6469 & ~n6473;
  assign n6475 = n6168 & n6203;
  assign n6476 = n6309 & n6434;
  assign n6477 = n6436 & n6466;
  assign n6478 = n6476 & n6477;
  assign n6479 = ~n6309 & n6434;
  assign n6480 = n6467 & n6479;
  assign n6481 = ~n6478 & ~n6480;
  assign n6482 = n6475 & ~n6481;
  assign n6483 = n6168 & ~n6203;
  assign n6484 = n6471 & n6476;
  assign n6485 = ~n6480 & ~n6484;
  assign n6486 = n6483 & ~n6485;
  assign n6487 = ~n6436 & n6466;
  assign n6488 = n6435 & n6487;
  assign n6489 = n6475 & n6488;
  assign n6490 = n6467 & n6476;
  assign n6491 = n6204 & n6490;
  assign n6492 = n6477 & n6479;
  assign n6493 = n6309 & ~n6434;
  assign n6494 = n6477 & n6493;
  assign n6495 = ~n6492 & ~n6494;
  assign n6496 = n6483 & ~n6495;
  assign n6497 = ~n6491 & ~n6496;
  assign n6498 = ~n6489 & n6497;
  assign n6499 = n6471 & n6493;
  assign n6500 = ~n6478 & ~n6499;
  assign n6501 = ~n6472 & n6500;
  assign n6502 = ~n6490 & n6501;
  assign n6503 = n6483 & ~n6502;
  assign n6504 = n6435 & n6477;
  assign n6505 = n6467 & n6493;
  assign n6506 = ~n6504 & ~n6505;
  assign n6507 = n6476 & n6487;
  assign n6508 = n6487 & n6493;
  assign n6509 = n6471 & n6479;
  assign n6510 = ~n6508 & ~n6509;
  assign n6511 = ~n6507 & n6510;
  assign n6512 = n6506 & n6511;
  assign n6513 = ~n6472 & n6512;
  assign n6514 = n6204 & ~n6513;
  assign n6515 = ~n6503 & ~n6514;
  assign n6516 = n6479 & n6487;
  assign n6517 = ~n6508 & ~n6516;
  assign n6518 = ~n6499 & n6517;
  assign n6519 = ~n6490 & ~n6504;
  assign n6520 = n6518 & n6519;
  assign n6521 = n6475 & ~n6520;
  assign n6522 = ~n6478 & n6506;
  assign n6523 = ~n6484 & n6522;
  assign n6524 = ~n6468 & n6523;
  assign n6525 = n6517 & n6524;
  assign n6526 = n6470 & ~n6525;
  assign n6527 = ~n6521 & ~n6526;
  assign n6528 = n6515 & n6527;
  assign n6529 = n6498 & n6528;
  assign n6530 = ~n6486 & n6529;
  assign n6531 = ~n6482 & n6530;
  assign n6532 = n6474 & n6531;
  assign n6533 = n6532 ^ n4570;
  assign n6534 = n6533 ^ x389;
  assign n6535 = n6167 & ~n6534;
  assign n6536 = ~n6259 & ~n6293;
  assign n6537 = ~n6235 & ~n6254;
  assign n6538 = ~n6255 & n6537;
  assign n6539 = ~n6254 & n6282;
  assign n6540 = ~n6538 & ~n6539;
  assign n6541 = ~n6300 & n6540;
  assign n6542 = n6207 & ~n6541;
  assign n6543 = n6257 & n6537;
  assign n6544 = ~n6292 & ~n6543;
  assign n6545 = n6274 & ~n6283;
  assign n6546 = n6255 ^ n6235;
  assign n6547 = n6256 ^ n6255;
  assign n6548 = n6546 & ~n6547;
  assign n6549 = ~n6254 & n6548;
  assign n6550 = n6545 & ~n6549;
  assign n6551 = n6544 & n6550;
  assign n6552 = n6299 & n6551;
  assign n6553 = ~n6542 & ~n6552;
  assign n6554 = n6270 & ~n6279;
  assign n6555 = ~n6281 & ~n6549;
  assign n6556 = ~n6554 & n6555;
  assign n6557 = n6278 & ~n6556;
  assign n6558 = n6291 & ~n6550;
  assign n6559 = ~n6557 & ~n6558;
  assign n6560 = n6553 & n6559;
  assign n6561 = n6536 & n6560;
  assign n6562 = n6561 ^ n4153;
  assign n6563 = n6562 ^ x351;
  assign n6564 = n6053 & ~n6450;
  assign n6565 = ~n6051 & ~n6057;
  assign n6566 = n6068 & n6565;
  assign n6567 = ~n6045 & ~n6072;
  assign n6568 = ~n6081 & n6567;
  assign n6569 = n6566 & n6568;
  assign n6570 = n6078 & ~n6569;
  assign n6571 = ~n6048 & ~n6053;
  assign n6572 = ~n6095 & ~n6101;
  assign n6573 = ~n6571 & ~n6572;
  assign n6574 = n6058 & n6099;
  assign n6575 = ~n6063 & n6574;
  assign n6576 = ~n6076 & n6575;
  assign n6577 = n5982 & ~n6576;
  assign n6578 = ~n6573 & ~n6577;
  assign n6579 = ~n6570 & n6578;
  assign n6580 = ~n6564 & n6579;
  assign n6581 = ~n6091 & n6580;
  assign n6582 = ~n6088 & n6581;
  assign n6583 = n6061 & n6582;
  assign n6584 = n6440 & n6583;
  assign n6585 = ~n6082 & n6584;
  assign n6586 = n6585 ^ n4187;
  assign n6587 = n6586 ^ x346;
  assign n6588 = ~n6563 & ~n6587;
  assign n6589 = n6405 & ~n6419;
  assign n6590 = ~n6409 & ~n6418;
  assign n6591 = n6384 & ~n6590;
  assign n6592 = ~n6589 & ~n6591;
  assign n6593 = n6312 & n6417;
  assign n6594 = n6384 & n6395;
  assign n6595 = n6312 & n6416;
  assign n6596 = ~n6594 & ~n6595;
  assign n6597 = ~n6593 & n6596;
  assign n6598 = n6312 & n6375;
  assign n6599 = ~n6387 & ~n6395;
  assign n6600 = n6405 & ~n6599;
  assign n6601 = ~n6370 & n6382;
  assign n6602 = n6372 & ~n6601;
  assign n6603 = ~n6600 & ~n6602;
  assign n6604 = ~n6598 & n6603;
  assign n6605 = ~n6310 & n6386;
  assign n6606 = n6380 & n6384;
  assign n6607 = ~n6605 & ~n6606;
  assign n6608 = n6312 & ~n6407;
  assign n6609 = n6410 & ~n6417;
  assign n6610 = n6372 & ~n6609;
  assign n6611 = ~n6384 & ~n6405;
  assign n6612 = ~n6403 & n6406;
  assign n6613 = ~n6611 & ~n6612;
  assign n6614 = ~n6610 & ~n6613;
  assign n6615 = ~n6608 & n6614;
  assign n6616 = n6607 & n6615;
  assign n6617 = n6394 & n6616;
  assign n6618 = n6377 & n6617;
  assign n6619 = n6604 & n6618;
  assign n6620 = n6597 & n6619;
  assign n6621 = n6592 & n6620;
  assign n6622 = n6621 ^ n4243;
  assign n6623 = n6622 ^ x347;
  assign n6624 = ~n5777 & ~n5819;
  assign n6625 = n5782 & ~n6624;
  assign n6626 = n5781 & n5806;
  assign n6627 = ~n5802 & ~n5807;
  assign n6628 = n5786 & ~n6627;
  assign n6629 = ~n6626 & ~n6628;
  assign n6630 = ~n5817 & n5818;
  assign n6631 = n5782 & ~n5835;
  assign n6632 = ~n6630 & ~n6631;
  assign n6633 = n5777 & ~n5817;
  assign n6634 = ~n5773 & ~n5820;
  assign n6635 = n6627 & n6634;
  assign n6636 = n5782 & ~n6635;
  assign n6637 = n5821 & n5832;
  assign n6638 = n5806 & ~n6637;
  assign n6639 = ~n5797 & ~n5828;
  assign n6640 = n5835 & n6639;
  assign n6641 = n5786 & ~n6640;
  assign n6642 = ~n6638 & ~n6641;
  assign n6643 = ~n5791 & n6634;
  assign n6644 = ~n5830 & n6643;
  assign n6645 = n5812 & n6644;
  assign n6646 = n6627 & n6645;
  assign n6647 = n5677 & ~n6646;
  assign n6648 = n6642 & ~n6647;
  assign n6649 = ~n6636 & n6648;
  assign n6650 = ~n6633 & n6649;
  assign n6651 = n6632 & n6650;
  assign n6652 = n6629 & n6651;
  assign n6653 = ~n6625 & n6652;
  assign n6654 = n6653 ^ n4274;
  assign n6655 = n6654 ^ x348;
  assign n6656 = n6623 & ~n6655;
  assign n6657 = n4138 & n4906;
  assign n6658 = n4138 & ~n4907;
  assign n6659 = ~n4873 & n4892;
  assign n6660 = n4898 & n6659;
  assign n6661 = ~n4886 & n6660;
  assign n6662 = n4905 & ~n6661;
  assign n6663 = ~n6658 & ~n6662;
  assign n6664 = n4888 & n4912;
  assign n6665 = n4882 & n4890;
  assign n6666 = ~n4916 & ~n6665;
  assign n6667 = n3701 & ~n6666;
  assign n6668 = n4892 & n4910;
  assign n6669 = n4872 & ~n6668;
  assign n6670 = ~n6667 & ~n6669;
  assign n6671 = ~n6664 & n6670;
  assign n6672 = n6663 & n6671;
  assign n6673 = ~n6657 & n6672;
  assign n6674 = n4885 & n6673;
  assign n6675 = n4878 & n6674;
  assign n6676 = n6675 ^ n4209;
  assign n6677 = n6676 ^ x350;
  assign n6678 = n5208 & n5217;
  assign n6679 = n5243 & ~n6678;
  assign n6680 = n5208 & n5219;
  assign n6681 = n5213 & n5249;
  assign n6682 = ~n6680 & ~n6681;
  assign n6683 = n5059 & n5232;
  assign n6684 = n5240 & ~n6683;
  assign n6685 = n5206 & n5213;
  assign n6686 = n5059 & n5235;
  assign n6687 = ~n6685 & ~n6686;
  assign n6688 = ~n5245 & n5260;
  assign n6689 = n5059 & ~n6688;
  assign n6690 = n5231 & ~n5252;
  assign n6691 = ~n6689 & ~n6690;
  assign n6692 = n5210 & ~n5244;
  assign n6693 = n5213 & n5226;
  assign n6694 = ~n6692 & ~n6693;
  assign n6695 = ~n5232 & ~n5264;
  assign n6696 = ~n5235 & n6695;
  assign n6697 = n5208 & ~n6696;
  assign n6698 = ~n5058 & n5237;
  assign n6699 = ~n6697 & ~n6698;
  assign n6700 = n6694 & n6699;
  assign n6701 = n6691 & n6700;
  assign n6702 = n6687 & n6701;
  assign n6703 = n6684 & n6702;
  assign n6704 = n6682 & n6703;
  assign n6705 = n5230 & n6704;
  assign n6706 = n6679 & n6705;
  assign n6707 = n6706 ^ n4304;
  assign n6708 = n6707 ^ x349;
  assign n6709 = ~n6677 & ~n6708;
  assign n6710 = n6656 & n6709;
  assign n6711 = n6588 & n6710;
  assign n6712 = n6563 & ~n6587;
  assign n6713 = ~n6623 & ~n6655;
  assign n6714 = ~n6677 & n6708;
  assign n6715 = n6713 & n6714;
  assign n6716 = ~n6623 & n6655;
  assign n6717 = n6677 & n6708;
  assign n6718 = n6716 & n6717;
  assign n6719 = ~n6715 & ~n6718;
  assign n6720 = n6712 & ~n6719;
  assign n6721 = ~n6711 & ~n6720;
  assign n6722 = ~n6563 & n6587;
  assign n6723 = n6710 & n6722;
  assign n6724 = ~n6677 & n6716;
  assign n6725 = n6708 & n6724;
  assign n6726 = n6677 & ~n6708;
  assign n6727 = n6713 & n6726;
  assign n6728 = ~n6725 & ~n6727;
  assign n6729 = n6712 & ~n6728;
  assign n6730 = ~n6723 & ~n6729;
  assign n6731 = n6656 & n6714;
  assign n6732 = n6588 & n6731;
  assign n6733 = n6563 & n6587;
  assign n6734 = n6623 & n6655;
  assign n6735 = n6714 & n6734;
  assign n6736 = n6726 & n6734;
  assign n6737 = ~n6735 & ~n6736;
  assign n6738 = n6733 & ~n6737;
  assign n6739 = ~n6732 & ~n6738;
  assign n6740 = n6656 & n6726;
  assign n6741 = n6712 & n6740;
  assign n6742 = ~n6719 & n6733;
  assign n6743 = ~n6741 & ~n6742;
  assign n6744 = ~n6731 & ~n6736;
  assign n6745 = n6722 & ~n6744;
  assign n6746 = ~n6708 & n6724;
  assign n6747 = n6733 & n6746;
  assign n6748 = n6733 & n6740;
  assign n6749 = n6712 & ~n6737;
  assign n6750 = ~n6748 & ~n6749;
  assign n6751 = ~n6747 & n6750;
  assign n6752 = n6587 ^ n6563;
  assign n6753 = n6713 & n6717;
  assign n6754 = ~n6752 & n6753;
  assign n6755 = n6709 & n6734;
  assign n6756 = n6712 & n6755;
  assign n6757 = ~n6754 & ~n6756;
  assign n6758 = n6710 & n6733;
  assign n6759 = n6709 & n6713;
  assign n6760 = n6717 & n6734;
  assign n6761 = n6656 & n6717;
  assign n6762 = ~n6760 & ~n6761;
  assign n6763 = n6716 & n6726;
  assign n6764 = ~n6746 & ~n6763;
  assign n6765 = n6762 & n6764;
  assign n6766 = ~n6759 & n6765;
  assign n6767 = n6588 & ~n6766;
  assign n6768 = n6728 & ~n6753;
  assign n6769 = ~n6763 & n6768;
  assign n6770 = ~n6760 & n6769;
  assign n6771 = n6722 & ~n6770;
  assign n6772 = ~n6767 & ~n6771;
  assign n6773 = ~n6758 & n6772;
  assign n6774 = n6757 & n6773;
  assign n6775 = n6751 & n6774;
  assign n6776 = ~n6745 & n6775;
  assign n6777 = n6743 & n6776;
  assign n6778 = n6739 & n6777;
  assign n6779 = n6730 & n6778;
  assign n6780 = n6721 & n6779;
  assign n6781 = n6780 ^ n4377;
  assign n6782 = n6781 ^ x391;
  assign n6783 = n5934 & n5963;
  assign n6784 = n5847 & n5955;
  assign n6785 = ~n6783 & ~n6784;
  assign n6786 = n5914 & n5950;
  assign n6787 = ~n5929 & n5945;
  assign n6788 = ~n6786 & ~n6787;
  assign n6789 = n6785 & n6788;
  assign n6790 = ~n5848 & n5962;
  assign n6791 = ~n5919 & ~n5935;
  assign n6792 = n5848 & ~n6791;
  assign n6793 = ~n5924 & ~n5936;
  assign n6794 = ~n5942 & ~n6793;
  assign n6795 = ~n5950 & ~n5955;
  assign n6796 = n5848 & ~n6795;
  assign n6797 = ~n6794 & ~n6796;
  assign n6798 = n5945 & ~n6179;
  assign n6799 = ~n5946 & n6190;
  assign n6800 = ~n5936 & n6799;
  assign n6801 = n5934 & ~n6800;
  assign n6802 = ~n6798 & ~n6801;
  assign n6803 = n6797 & n6802;
  assign n6804 = n5922 & n6803;
  assign n6805 = ~n6792 & n6804;
  assign n6806 = ~n6790 & n6805;
  assign n6807 = n6789 & n6806;
  assign n6808 = ~n5949 & n6807;
  assign n6809 = n6170 & n6808;
  assign n6810 = n6809 ^ n4739;
  assign n6811 = n6810 ^ x311;
  assign n6812 = n5786 & n5802;
  assign n6813 = ~n5677 & ~n5806;
  assign n6814 = n5797 & ~n6813;
  assign n6815 = ~n6812 & ~n6814;
  assign n6816 = ~n5789 & ~n5818;
  assign n6817 = n5782 & ~n6816;
  assign n6818 = ~n5799 & n6627;
  assign n6819 = n5677 & ~n6818;
  assign n6820 = ~n6817 & ~n6819;
  assign n6821 = ~n5809 & n5835;
  assign n6822 = ~n5817 & ~n6821;
  assign n6823 = n5828 & ~n6813;
  assign n6824 = n5806 & ~n6643;
  assign n6825 = ~n6823 & ~n6824;
  assign n6826 = ~n5811 & n6627;
  assign n6827 = n5782 & ~n6826;
  assign n6828 = ~n5818 & n6643;
  assign n6829 = n5677 & ~n6634;
  assign n6830 = ~n5786 & ~n6829;
  assign n6831 = ~n6828 & ~n6830;
  assign n6832 = ~n6827 & ~n6831;
  assign n6833 = n6825 & n6832;
  assign n6834 = n5784 & n6833;
  assign n6835 = ~n6822 & n6834;
  assign n6836 = n6820 & n6835;
  assign n6837 = n6815 & n6836;
  assign n6838 = ~n6625 & n6837;
  assign n6839 = n6838 ^ n4758;
  assign n6840 = n6839 ^ x312;
  assign n6841 = ~n6811 & ~n6840;
  assign n6842 = n5493 & n5572;
  assign n6843 = ~n5566 & ~n6842;
  assign n6844 = n5561 & n5568;
  assign n6845 = n5572 & n5595;
  assign n6846 = ~n6844 & ~n6845;
  assign n6847 = ~n5601 & n5613;
  assign n6848 = n6846 & ~n6847;
  assign n6849 = n5561 & n5613;
  assign n6850 = n5565 & n5583;
  assign n6851 = n5569 & n5582;
  assign n6852 = ~n6850 & ~n6851;
  assign n6853 = ~n6849 & n6852;
  assign n6854 = n5564 & n5572;
  assign n6855 = ~n5587 & ~n5592;
  assign n6856 = ~n5571 & n6855;
  assign n6857 = n5603 & n6856;
  assign n6858 = ~n5491 & n6857;
  assign n6859 = n5565 & ~n6858;
  assign n6860 = ~n6854 & ~n6859;
  assign n6861 = ~n5578 & ~n5594;
  assign n6862 = n5561 & ~n6861;
  assign n6863 = ~n5571 & ~n5578;
  assign n6864 = ~n5608 & n6863;
  assign n6865 = ~n5572 & n6864;
  assign n6866 = n5569 & ~n6863;
  assign n6867 = n5609 & ~n6866;
  assign n6868 = ~n5568 & n6867;
  assign n6869 = ~n6865 & ~n6868;
  assign n6870 = ~n5601 & n6869;
  assign n6871 = ~n6862 & ~n6870;
  assign n6872 = n6860 & n6871;
  assign n6873 = ~n5591 & n6872;
  assign n6874 = n6853 & n6873;
  assign n6875 = n5586 & n6874;
  assign n6876 = n6848 & n6875;
  assign n6877 = n6843 & n6876;
  assign n6878 = ~n5562 & n6877;
  assign n6879 = n6878 ^ n2495;
  assign n6880 = n6879 ^ x314;
  assign n6881 = n4572 & n4874;
  assign n6882 = ~n4866 & ~n6881;
  assign n6883 = ~n4875 & n6882;
  assign n6884 = ~n4917 & n6883;
  assign n6885 = n4138 & ~n6884;
  assign n6886 = ~n4873 & ~n6881;
  assign n6887 = n4909 & n6886;
  assign n6888 = ~n4906 & n6887;
  assign n6889 = n4888 & ~n6888;
  assign n6890 = ~n6885 & ~n6889;
  assign n6891 = ~n4869 & n4907;
  assign n6892 = ~n4905 & n6891;
  assign n6893 = ~n4865 & ~n4872;
  assign n6894 = n4572 & ~n6893;
  assign n6895 = n4898 & ~n6894;
  assign n6896 = ~n4875 & n6895;
  assign n6897 = ~n6892 & ~n6896;
  assign n6898 = ~n6665 & ~n6897;
  assign n6899 = n4918 & n6898;
  assign n6900 = ~n4900 & n6899;
  assign n6901 = n4895 & ~n6900;
  assign n6902 = n6890 & ~n6901;
  assign n6903 = n4897 & n6902;
  assign n6904 = ~n4887 & n6903;
  assign n6905 = ~n6657 & n6904;
  assign n6906 = n4885 & n6905;
  assign n6907 = n6906 ^ n4789;
  assign n6908 = n6907 ^ x313;
  assign n6909 = ~n6880 & n6908;
  assign n6910 = n6841 & n6909;
  assign n6911 = ~n5237 & n5260;
  assign n6912 = n5208 & ~n6911;
  assign n6913 = ~n5247 & n6688;
  assign n6914 = n5213 & ~n6913;
  assign n6915 = ~n6912 & ~n6914;
  assign n6916 = ~n5247 & ~n5264;
  assign n6917 = ~n5244 & ~n6916;
  assign n6918 = ~n5210 & ~n5223;
  assign n6919 = ~n5215 & n6918;
  assign n6920 = ~n5226 & n6919;
  assign n6921 = n5231 & ~n6920;
  assign n6922 = ~n6917 & ~n6921;
  assign n6923 = n6915 & n6922;
  assign n6924 = n5229 & n6923;
  assign n6925 = n6687 & n6924;
  assign n6926 = n6684 & n6925;
  assign n6927 = n6682 & n6926;
  assign n6928 = n5212 & n6927;
  assign n6929 = ~n5217 & n6928;
  assign n6930 = n6929 ^ n3498;
  assign n6931 = n6930 ^ x315;
  assign n6932 = ~n6310 & n6375;
  assign n6933 = ~n6391 & ~n6395;
  assign n6934 = ~n6416 & n6933;
  assign n6935 = ~n6403 & n6934;
  assign n6936 = n6372 & ~n6935;
  assign n6937 = ~n6932 & ~n6936;
  assign n6938 = ~n6386 & ~n6418;
  assign n6939 = ~n6370 & n6938;
  assign n6940 = ~n6403 & n6939;
  assign n6941 = n6312 & ~n6940;
  assign n6942 = n6400 & ~n6403;
  assign n6943 = ~n6409 & n6942;
  assign n6944 = ~n6405 & n6943;
  assign n6945 = ~n6384 & ~n6399;
  assign n6946 = ~n6942 & ~n6945;
  assign n6947 = n6590 & ~n6946;
  assign n6948 = ~n6417 & n6947;
  assign n6949 = ~n6944 & ~n6948;
  assign n6950 = ~n6408 & ~n6949;
  assign n6951 = ~n6611 & ~n6950;
  assign n6952 = ~n6941 & ~n6951;
  assign n6953 = n6937 & n6952;
  assign n6954 = n6596 & n6953;
  assign n6955 = n6390 & n6954;
  assign n6956 = n6604 & n6955;
  assign n6957 = n6956 ^ n4714;
  assign n6958 = n6957 ^ x310;
  assign n6959 = n6931 & ~n6958;
  assign n6960 = n6910 & n6959;
  assign n6961 = n6931 & n6958;
  assign n6962 = ~n6880 & ~n6908;
  assign n6963 = n6841 & n6962;
  assign n6964 = n6961 & n6963;
  assign n6965 = ~n6960 & ~n6964;
  assign n6966 = n6880 & ~n6908;
  assign n6967 = n6841 & n6966;
  assign n6968 = n6959 & n6967;
  assign n6969 = ~n6811 & n6840;
  assign n6970 = n6962 & n6969;
  assign n6971 = n6961 & n6970;
  assign n6972 = n6811 & ~n6840;
  assign n6973 = n6909 & n6972;
  assign n6974 = n6959 & n6973;
  assign n6975 = n6909 & n6969;
  assign n6976 = ~n6931 & ~n6958;
  assign n6977 = ~n6961 & ~n6976;
  assign n6978 = n6975 & ~n6977;
  assign n6979 = ~n6974 & ~n6978;
  assign n6980 = n6880 & n6908;
  assign n6981 = n6969 & n6980;
  assign n6982 = ~n6931 & n6958;
  assign n6983 = n6981 & n6982;
  assign n6984 = n6966 & n6969;
  assign n6985 = ~n6977 & n6984;
  assign n6986 = ~n6983 & ~n6985;
  assign n6987 = n6962 & n6972;
  assign n6988 = n6811 & n6840;
  assign n6989 = n6966 & n6988;
  assign n6990 = ~n6987 & ~n6989;
  assign n6991 = n6976 & ~n6990;
  assign n6992 = n6962 & n6988;
  assign n6993 = n6966 & n6972;
  assign n6994 = ~n6992 & ~n6993;
  assign n6995 = ~n6989 & n6994;
  assign n6996 = n6959 & ~n6995;
  assign n6997 = n6841 & n6980;
  assign n6998 = ~n6970 & ~n6997;
  assign n6999 = ~n6963 & n6998;
  assign n7000 = n6982 & ~n6999;
  assign n7001 = ~n6996 & ~n7000;
  assign n7002 = n6961 & n6997;
  assign n7003 = ~n6910 & ~n6967;
  assign n7004 = n6976 & ~n7003;
  assign n7013 = n6980 & n6988;
  assign n7014 = ~n6961 & ~n6973;
  assign n7007 = n6972 & n6980;
  assign n7015 = n6973 & n6976;
  assign n7016 = ~n6987 & ~n7015;
  assign n7017 = ~n7007 & n7016;
  assign n7018 = ~n7014 & ~n7017;
  assign n7019 = ~n7013 & ~n7018;
  assign n7005 = n6909 & n6988;
  assign n7006 = n6959 & n6981;
  assign n7008 = ~n6993 & ~n7007;
  assign n7009 = ~n6973 & n7008;
  assign n7010 = n6982 & ~n7009;
  assign n7011 = ~n7006 & ~n7010;
  assign n7012 = ~n7005 & n7011;
  assign n7020 = n7019 ^ n7012;
  assign n7021 = n6977 & n7020;
  assign n7022 = n7021 ^ n7019;
  assign n7023 = ~n7004 & n7022;
  assign n7024 = ~n7002 & n7023;
  assign n7025 = n7001 & n7024;
  assign n7026 = ~n6991 & n7025;
  assign n7027 = n6986 & n7026;
  assign n7028 = n6979 & n7027;
  assign n7029 = ~n6971 & n7028;
  assign n7030 = ~n6968 & n7029;
  assign n7031 = n6965 & n7030;
  assign n7032 = n7031 ^ n4863;
  assign n7033 = n7032 ^ x392;
  assign n7034 = ~n6782 & n7033;
  assign n7035 = n6535 & n7034;
  assign n7036 = n6879 ^ x316;
  assign n7037 = n6116 ^ x321;
  assign n7038 = ~n7036 & n7037;
  assign n7039 = n4928 ^ x320;
  assign n7040 = ~n6311 & n6391;
  assign n7041 = n6375 & ~n6611;
  assign n7042 = ~n7040 & ~n7041;
  assign n7043 = n6372 & n6386;
  assign n7044 = n6312 & ~n6406;
  assign n7045 = ~n7043 & ~n7044;
  assign n7046 = n7042 & n7045;
  assign n7047 = n6370 & n6405;
  assign n7048 = n6384 & n6387;
  assign n7049 = ~n7047 & ~n7048;
  assign n7050 = ~n6403 & ~n6408;
  assign n7051 = ~n6310 & ~n7050;
  assign n7052 = ~n6400 & n6405;
  assign n7053 = n6406 & n6419;
  assign n7054 = n6372 & ~n7053;
  assign n7055 = ~n7052 & ~n7054;
  assign n7056 = ~n6397 & ~n6416;
  assign n7057 = n6384 & ~n7056;
  assign n7058 = n6388 & n7050;
  assign n7059 = n6312 & ~n7058;
  assign n7060 = ~n7057 & ~n7059;
  assign n7061 = n7055 & n7060;
  assign n7062 = n6592 & n7061;
  assign n7063 = ~n7051 & n7062;
  assign n7064 = n7049 & n7063;
  assign n7065 = n7046 & n7064;
  assign n7066 = n6597 & n7065;
  assign n7067 = n7066 ^ n3630;
  assign n7068 = n7067 ^ x319;
  assign n7069 = n7039 & ~n7068;
  assign n7070 = n6536 & n6550;
  assign n7071 = n6207 & n7070;
  assign n7072 = n6278 & ~n6551;
  assign n7073 = ~n7071 & ~n7072;
  assign n7074 = n6536 & n6541;
  assign n7075 = n6291 & ~n7074;
  assign n7076 = ~n6235 & n6300;
  assign n7077 = n6555 & ~n7076;
  assign n7078 = n6294 & n7077;
  assign n7079 = ~n6259 & n7078;
  assign n7080 = n6299 & ~n7079;
  assign n7081 = ~n7075 & ~n7080;
  assign n7082 = n7073 & n7081;
  assign n7083 = n7082 ^ n3318;
  assign n7084 = n7083 ^ x318;
  assign n7085 = n6930 ^ x317;
  assign n7086 = ~n7084 & ~n7085;
  assign n7087 = n7069 & n7086;
  assign n7088 = n7038 & n7087;
  assign n7089 = n7036 & n7037;
  assign n7090 = ~n7039 & ~n7068;
  assign n7091 = n7084 & n7085;
  assign n7092 = n7090 & n7091;
  assign n7093 = ~n7084 & n7085;
  assign n7094 = n7069 & n7093;
  assign n7095 = ~n7092 & ~n7094;
  assign n7096 = n7089 & ~n7095;
  assign n7097 = ~n7039 & n7068;
  assign n7098 = n7084 & ~n7085;
  assign n7099 = n7097 & n7098;
  assign n7100 = n7069 & n7098;
  assign n7101 = ~n7099 & ~n7100;
  assign n7102 = n7038 & ~n7101;
  assign n7103 = ~n7096 & ~n7102;
  assign n7104 = n7037 ^ n7036;
  assign n7105 = n7086 & n7097;
  assign n7106 = n7104 & n7105;
  assign n7107 = n7039 & n7068;
  assign n7108 = n7098 & n7107;
  assign n7109 = ~n7037 & n7108;
  assign n7110 = ~n7106 & ~n7109;
  assign n7111 = n7091 & n7097;
  assign n7112 = n7086 & n7090;
  assign n7113 = ~n7111 & ~n7112;
  assign n7114 = n7089 & ~n7113;
  assign n7115 = ~n7036 & ~n7037;
  assign n7116 = n7090 & n7098;
  assign n7117 = ~n7087 & ~n7112;
  assign n7118 = ~n7116 & n7117;
  assign n7119 = n7115 & ~n7118;
  assign n7120 = n7094 & n7115;
  assign n7121 = n7093 & n7107;
  assign n7122 = n7038 & n7121;
  assign n7123 = n7036 & ~n7037;
  assign n7124 = n7121 & n7123;
  assign n7125 = n7086 & n7107;
  assign n7126 = ~n7087 & ~n7125;
  assign n7127 = n7123 & ~n7126;
  assign n7128 = n7091 & n7107;
  assign n7129 = n7093 & n7097;
  assign n7130 = ~n7128 & ~n7129;
  assign n7131 = ~n7092 & n7130;
  assign n7132 = n7115 & ~n7131;
  assign n7133 = ~n7127 & ~n7132;
  assign n7134 = n7069 & n7091;
  assign n7135 = n7090 & n7093;
  assign n7136 = ~n7134 & ~n7135;
  assign n7137 = ~n7111 & n7136;
  assign n7138 = n7104 & ~n7137;
  assign n7139 = ~n7116 & ~n7125;
  assign n7140 = ~n7108 & n7139;
  assign n7141 = ~n7105 & n7140;
  assign n7142 = n7089 & ~n7141;
  assign n7143 = ~n7138 & ~n7142;
  assign n7144 = n7133 & n7143;
  assign n7145 = ~n7124 & n7144;
  assign n7146 = ~n7122 & n7145;
  assign n7147 = ~n7120 & n7146;
  assign n7148 = ~n7119 & n7147;
  assign n7149 = ~n7114 & n7148;
  assign n7150 = n7110 & n7149;
  assign n7151 = n7103 & n7150;
  assign n7152 = ~n7088 & n7151;
  assign n7153 = n7152 ^ n3700;
  assign n7154 = n7153 ^ x388;
  assign n7155 = n5565 & n5588;
  assign n7156 = n5569 & n5587;
  assign n7157 = ~n7155 & ~n7156;
  assign n7158 = ~n5560 & n5583;
  assign n7159 = n5588 & ~n5601;
  assign n7160 = ~n7158 & ~n7159;
  assign n7161 = ~n5582 & ~n5587;
  assign n7162 = n5565 & ~n7161;
  assign n7163 = ~n5491 & ~n5568;
  assign n7164 = n6861 & n7163;
  assign n7165 = ~n5592 & n7164;
  assign n7166 = n5569 & ~n7165;
  assign n7167 = ~n7162 & ~n7166;
  assign n7168 = ~n5493 & n5596;
  assign n7169 = n6856 & n7168;
  assign n7170 = n5561 & ~n7169;
  assign n7171 = n6863 & n7163;
  assign n7172 = n5565 & ~n7171;
  assign n7173 = ~n5594 & n5609;
  assign n7174 = ~n5571 & n7173;
  assign n7175 = n5572 & ~n7174;
  assign n7176 = ~n7172 & ~n7175;
  assign n7177 = ~n7170 & n7176;
  assign n7178 = n7167 & n7177;
  assign n7179 = n7160 & n7178;
  assign n7180 = n7157 & n7179;
  assign n7181 = n6848 & n7180;
  assign n7182 = ~n5566 & n7181;
  assign n7183 = n7182 ^ n3740;
  assign n7184 = n7183 ^ x339;
  assign n7185 = n6308 ^ x334;
  assign n7186 = n7184 & ~n7185;
  assign n7187 = n4869 & n4872;
  assign n7188 = ~n4894 & n4908;
  assign n7189 = n4918 & n7188;
  assign n7190 = n4905 & ~n7189;
  assign n7191 = ~n7187 & ~n7190;
  assign n7192 = ~n6665 & n6886;
  assign n7193 = n4138 & ~n7192;
  assign n7194 = n4910 & ~n4917;
  assign n7195 = n4888 & ~n7194;
  assign n7196 = ~n7193 & ~n7195;
  assign n7197 = n7191 & n7196;
  assign n7198 = n3701 & n4880;
  assign n7199 = n4889 & n4895;
  assign n7200 = n4870 & ~n6881;
  assign n7201 = ~n4872 & n7200;
  assign n7202 = ~n4900 & ~n4917;
  assign n7203 = ~n4906 & n7202;
  assign n7204 = ~n4888 & n7203;
  assign n7205 = ~n7201 & ~n7204;
  assign n7206 = ~n4894 & ~n7205;
  assign n7207 = ~n3701 & ~n7206;
  assign n7208 = ~n7199 & ~n7207;
  assign n7209 = ~n7198 & n7208;
  assign n7210 = n7197 & n7209;
  assign n7211 = ~n4887 & n7210;
  assign n7212 = ~n6657 & n7211;
  assign n7213 = n4878 & n7212;
  assign n7214 = n7213 ^ n4002;
  assign n7215 = n7214 ^ x336;
  assign n7216 = n6202 ^ x335;
  assign n7217 = n7215 & n7216;
  assign n7218 = n5782 & n5811;
  assign n7219 = n5799 & n5806;
  assign n7220 = n5782 & ~n6639;
  assign n7221 = n5821 & n5831;
  assign n7222 = ~n5781 & n7221;
  assign n7223 = ~n5797 & n7222;
  assign n7224 = n5677 & ~n7223;
  assign n7225 = n5792 & n5812;
  assign n7226 = ~n5828 & n7225;
  assign n7227 = ~n5817 & ~n7226;
  assign n7228 = ~n7224 & ~n7227;
  assign n7229 = ~n7220 & n7228;
  assign n7230 = ~n7219 & n7229;
  assign n7231 = ~n7218 & n7230;
  assign n7232 = n6632 & n7231;
  assign n7233 = n5785 & n7232;
  assign n7234 = n6629 & n7233;
  assign n7235 = ~n6625 & n7234;
  assign n7236 = n7235 ^ n3968;
  assign n7237 = n7236 ^ x338;
  assign n7238 = n5208 & n5245;
  assign n7239 = n5257 & n6919;
  assign n7240 = ~n5259 & n7239;
  assign n7241 = n5213 & ~n7240;
  assign n7242 = ~n7238 & ~n7241;
  assign n7243 = ~n5221 & n5231;
  assign n7244 = ~n5237 & n5261;
  assign n7245 = n5059 & ~n7244;
  assign n7246 = ~n5058 & ~n5231;
  assign n7247 = ~n5235 & ~n5249;
  assign n7248 = ~n5247 & n7247;
  assign n7249 = ~n5058 & n7248;
  assign n7250 = n5244 & ~n5259;
  assign n7251 = ~n5247 & n7250;
  assign n7252 = n4962 & n5250;
  assign n7253 = ~n7251 & ~n7252;
  assign n7254 = ~n5264 & ~n7253;
  assign n7255 = ~n7249 & ~n7254;
  assign n7256 = ~n5226 & ~n7255;
  assign n7257 = ~n7246 & ~n7256;
  assign n7258 = ~n7245 & ~n7257;
  assign n7259 = ~n7243 & n7258;
  assign n7260 = n7242 & n7259;
  assign n7261 = n6679 & n7260;
  assign n7262 = n5212 & n7261;
  assign n7263 = n7262 ^ n4044;
  assign n7264 = n7263 ^ x337;
  assign n7265 = n7237 & ~n7264;
  assign n7266 = n7217 & n7265;
  assign n7267 = n7186 & n7266;
  assign n7268 = n7215 & ~n7216;
  assign n7269 = n7237 & n7264;
  assign n7270 = n7268 & n7269;
  assign n7271 = n7186 & n7270;
  assign n7272 = ~n7184 & n7185;
  assign n7273 = ~n7215 & ~n7216;
  assign n7274 = n7269 & n7273;
  assign n7275 = ~n7237 & ~n7264;
  assign n7276 = n7273 & n7275;
  assign n7277 = ~n7274 & ~n7276;
  assign n7278 = n7272 & ~n7277;
  assign n7279 = ~n7271 & ~n7278;
  assign n7280 = ~n7215 & n7216;
  assign n7281 = n7275 & n7280;
  assign n7282 = ~n7266 & ~n7281;
  assign n7283 = n7272 & ~n7282;
  assign n7284 = ~n7184 & ~n7185;
  assign n7285 = n7269 & n7280;
  assign n7286 = n7284 & n7285;
  assign n7287 = ~n7237 & n7264;
  assign n7288 = n7273 & n7287;
  assign n7289 = n7186 & n7288;
  assign n7290 = ~n7286 & ~n7289;
  assign n7291 = n7184 & n7185;
  assign n7292 = n7280 & n7287;
  assign n7293 = n7265 & n7280;
  assign n7294 = ~n7292 & ~n7293;
  assign n7295 = n7291 & ~n7294;
  assign n7296 = ~n7284 & ~n7291;
  assign n7297 = n7268 & n7275;
  assign n7298 = n7296 & n7297;
  assign n7299 = n7272 & n7292;
  assign n7300 = n7186 & ~n7294;
  assign n7301 = ~n7299 & ~n7300;
  assign n7302 = n7217 & n7269;
  assign n7303 = n7265 & n7273;
  assign n7304 = ~n7302 & ~n7303;
  assign n7305 = n7272 & ~n7304;
  assign n7306 = ~n7281 & ~n7285;
  assign n7307 = n7186 & ~n7306;
  assign n7308 = ~n7305 & ~n7307;
  assign n7309 = n7217 & n7275;
  assign n7310 = n7217 & n7287;
  assign n7311 = n7284 & n7303;
  assign n7312 = n7268 & n7287;
  assign n7313 = n7265 & n7268;
  assign n7314 = ~n7312 & ~n7313;
  assign n7315 = ~n7311 & n7314;
  assign n7316 = n7277 & n7315;
  assign n7317 = ~n7310 & n7316;
  assign n7318 = ~n7309 & n7317;
  assign n7319 = ~n7296 & ~n7318;
  assign n7320 = n7308 & ~n7319;
  assign n7321 = n7301 & n7320;
  assign n7322 = ~n7298 & n7321;
  assign n7323 = ~n7295 & n7322;
  assign n7324 = n7290 & n7323;
  assign n7325 = ~n7283 & n7324;
  assign n7326 = n7279 & n7325;
  assign n7327 = ~n7267 & n7326;
  assign n7328 = n7327 ^ n4136;
  assign n7329 = n7328 ^ x393;
  assign n7330 = ~n7154 & ~n7329;
  assign n7331 = n7035 & n7330;
  assign n7332 = ~n7154 & n7329;
  assign n7333 = n6167 & n6534;
  assign n7334 = n7034 & n7333;
  assign n7335 = ~n6167 & n6534;
  assign n7336 = ~n6782 & ~n7033;
  assign n7337 = n7335 & n7336;
  assign n7338 = ~n7334 & ~n7337;
  assign n7339 = n7332 & ~n7338;
  assign n7340 = ~n7331 & ~n7339;
  assign n7341 = ~n6167 & ~n6534;
  assign n7342 = n7034 & n7341;
  assign n7343 = n7332 & n7342;
  assign n7344 = n6782 & n7033;
  assign n7345 = n7335 & n7344;
  assign n7346 = n6782 & ~n7033;
  assign n7347 = n7333 & n7346;
  assign n7348 = ~n7345 & ~n7347;
  assign n7349 = n7330 & ~n7348;
  assign n7350 = ~n7343 & ~n7349;
  assign n7351 = n7154 & n7329;
  assign n7352 = n7335 & n7346;
  assign n7353 = n7034 & n7335;
  assign n7354 = ~n7347 & ~n7353;
  assign n7355 = ~n7352 & n7354;
  assign n7356 = n7351 & ~n7355;
  assign n7357 = n7035 & n7351;
  assign n7358 = n6535 & n7346;
  assign n7359 = n7332 & n7358;
  assign n7360 = ~n7357 & ~n7359;
  assign n7361 = n7333 & n7336;
  assign n7362 = n7341 & n7346;
  assign n7363 = ~n7361 & ~n7362;
  assign n7364 = n7154 & ~n7329;
  assign n7365 = ~n7332 & ~n7364;
  assign n7366 = ~n7363 & n7365;
  assign n7367 = n6535 & n7344;
  assign n7368 = n7336 & n7341;
  assign n7369 = ~n7367 & ~n7368;
  assign n7370 = n7351 & ~n7369;
  assign n7371 = ~n7366 & ~n7370;
  assign n7372 = n7341 & n7344;
  assign n7373 = ~n7362 & ~n7372;
  assign n7374 = n7354 & n7373;
  assign n7375 = n7369 & n7374;
  assign n7376 = ~n7334 & n7375;
  assign n7377 = ~n7035 & n7376;
  assign n7378 = n7364 & n7377;
  assign n7379 = ~n7342 & ~n7358;
  assign n7380 = ~n7353 & n7379;
  assign n7381 = n7330 & ~n7380;
  assign n7382 = ~n7035 & ~n7352;
  assign n7383 = n7373 & n7382;
  assign n7384 = n7332 & ~n7383;
  assign n7385 = ~n7381 & ~n7384;
  assign n7386 = ~n7378 & n7385;
  assign n7387 = n7371 & n7386;
  assign n7388 = n7360 & n7387;
  assign n7389 = ~n7356 & n7388;
  assign n7390 = n7350 & n7389;
  assign n7391 = n7340 & n7390;
  assign n7392 = n7391 ^ n4928;
  assign n7393 = n7392 ^ x418;
  assign n7394 = n6622 ^ x345;
  assign n7395 = n7236 ^ x340;
  assign n7396 = n7394 & n7395;
  assign n7397 = n7183 ^ x341;
  assign n7398 = n6288 & n6299;
  assign n7399 = ~n6276 & n6291;
  assign n7400 = ~n7398 & ~n7399;
  assign n7401 = n6207 & ~n6297;
  assign n7402 = n6278 & ~n6304;
  assign n7403 = ~n7401 & ~n7402;
  assign n7404 = n7400 & n7403;
  assign n7405 = n7404 ^ n4996;
  assign n7406 = n7405 ^ x342;
  assign n7407 = n7397 & ~n7406;
  assign n7408 = ~n5848 & n5928;
  assign n7409 = n5934 & ~n6172;
  assign n7410 = ~n7408 & ~n7409;
  assign n7411 = n5909 & ~n5942;
  assign n7412 = n6184 & n6190;
  assign n7413 = ~n5963 & n7412;
  assign n7414 = n5914 & ~n7413;
  assign n7415 = ~n7411 & ~n7414;
  assign n7416 = n5964 & n6179;
  assign n7417 = n5848 & ~n7416;
  assign n7418 = n5907 ^ n5874;
  assign n7419 = n5876 & ~n7418;
  assign n7420 = ~n5945 & ~n7419;
  assign n7421 = n5920 & ~n5924;
  assign n7422 = ~n5932 & n7421;
  assign n7423 = ~n5934 & n7422;
  assign n7424 = ~n7420 & ~n7423;
  assign n7425 = n5847 & n7424;
  assign n7426 = ~n7417 & ~n7425;
  assign n7427 = n7415 & n7426;
  assign n7428 = n7410 & n7427;
  assign n7429 = n6174 & n7428;
  assign n7430 = n6170 & n7429;
  assign n7431 = n7430 ^ n4982;
  assign n7432 = n7431 ^ x343;
  assign n7433 = n6586 ^ x344;
  assign n7434 = ~n7432 & n7433;
  assign n7435 = n7407 & n7434;
  assign n7436 = n7396 & n7435;
  assign n7437 = n7432 & ~n7433;
  assign n7438 = n7407 & n7437;
  assign n7439 = n7396 & n7438;
  assign n7440 = n7394 & ~n7395;
  assign n7441 = n7432 & n7433;
  assign n7442 = n7407 & n7441;
  assign n7443 = n7440 & n7442;
  assign n7444 = ~n7394 & n7395;
  assign n7445 = n7397 & n7406;
  assign n7446 = n7437 & n7445;
  assign n7447 = ~n7442 & ~n7446;
  assign n7448 = n7444 & ~n7447;
  assign n7449 = ~n7443 & ~n7448;
  assign n7450 = ~n7439 & n7449;
  assign n7451 = ~n7397 & ~n7406;
  assign n7452 = n7441 & n7451;
  assign n7453 = ~n7432 & ~n7433;
  assign n7454 = n7451 & n7453;
  assign n7455 = ~n7452 & ~n7454;
  assign n7456 = n7396 & ~n7455;
  assign n7457 = ~n7397 & n7406;
  assign n7458 = n7441 & n7457;
  assign n7459 = ~n7454 & ~n7458;
  assign n7460 = n7440 & ~n7459;
  assign n7461 = ~n7456 & ~n7460;
  assign n7462 = n7435 & n7444;
  assign n7463 = ~n7440 & ~n7444;
  assign n7464 = n7407 & n7453;
  assign n7465 = n7434 & n7457;
  assign n7466 = n7437 & n7451;
  assign n7467 = ~n7465 & ~n7466;
  assign n7468 = ~n7464 & n7467;
  assign n7469 = ~n7463 & ~n7468;
  assign n7470 = ~n7462 & ~n7469;
  assign n7471 = n7461 & n7470;
  assign n7472 = n7434 & n7451;
  assign n7473 = n7453 & n7457;
  assign n7474 = ~n7472 & ~n7473;
  assign n7475 = n7395 & ~n7474;
  assign n7476 = n7434 & n7445;
  assign n7477 = ~n7446 & ~n7476;
  assign n7478 = n7394 & ~n7477;
  assign n7479 = ~n7475 & ~n7478;
  assign n7480 = ~n7394 & ~n7395;
  assign n7481 = ~n7435 & ~n7476;
  assign n7482 = ~n7446 & n7459;
  assign n7483 = n7481 & n7482;
  assign n7484 = n7467 & n7483;
  assign n7485 = ~n7452 & n7484;
  assign n7486 = n7480 & n7485;
  assign n7487 = n7479 & ~n7486;
  assign n7488 = n7471 & n7487;
  assign n7489 = n7450 & n7488;
  assign n7490 = ~n7436 & n7489;
  assign n7491 = n7490 ^ n5057;
  assign n7492 = n7491 ^ x352;
  assign n7493 = n6710 & n6712;
  assign n7494 = n6722 & n6759;
  assign n7495 = ~n7493 & ~n7494;
  assign n7496 = n6588 & n6760;
  assign n7497 = n6733 & n6755;
  assign n7498 = ~n7496 & ~n7497;
  assign n7499 = ~n6761 & n6764;
  assign n7500 = n6712 & ~n7499;
  assign n7501 = ~n6731 & ~n6755;
  assign n7502 = n6762 & n7501;
  assign n7503 = ~n6727 & n7502;
  assign n7504 = ~n6715 & n7503;
  assign n7505 = n6722 & ~n7504;
  assign n7506 = ~n7500 & ~n7505;
  assign n7507 = ~n6563 & n6763;
  assign n7508 = ~n6735 & ~n6760;
  assign n7509 = n6733 & ~n7508;
  assign n7510 = n6715 & n6733;
  assign n7511 = n6588 & ~n6737;
  assign n7512 = ~n6752 & ~n6768;
  assign n7513 = ~n7511 & ~n7512;
  assign n7514 = ~n7510 & n7513;
  assign n7515 = ~n7509 & n7514;
  assign n7516 = ~n7507 & n7515;
  assign n7517 = n7506 & n7516;
  assign n7518 = n7498 & n7517;
  assign n7519 = n6750 & n7518;
  assign n7520 = n7495 & n7519;
  assign n7521 = n6721 & n7520;
  assign n7522 = n7521 ^ n4961;
  assign n7523 = n7522 ^ x357;
  assign n7524 = ~n7492 & ~n7523;
  assign n7525 = n6959 & n6984;
  assign n7526 = n6963 & n6976;
  assign n7527 = ~n6967 & ~n7007;
  assign n7528 = n6961 & ~n7527;
  assign n7529 = ~n7526 & ~n7528;
  assign n7530 = ~n7525 & n7529;
  assign n7531 = n6976 & n7007;
  assign n7532 = ~n7015 & ~n7531;
  assign n7533 = n6959 & n7013;
  assign n7534 = ~n6989 & ~n7005;
  assign n7535 = n6982 & ~n7534;
  assign n7536 = ~n7533 & ~n7535;
  assign n7537 = n6959 & ~n7534;
  assign n7538 = ~n6910 & ~n6963;
  assign n7539 = ~n6981 & n7538;
  assign n7540 = n6982 & ~n7539;
  assign n7541 = ~n7537 & ~n7540;
  assign n7542 = n6982 & n7013;
  assign n7543 = n6961 & n6973;
  assign n7544 = n6959 & n6987;
  assign n7545 = ~n7543 & ~n7544;
  assign n7546 = ~n7542 & n7545;
  assign n7547 = n6959 & n6975;
  assign n7548 = n6982 & ~n7527;
  assign n7549 = ~n7547 & ~n7548;
  assign n7550 = ~n6987 & ~n6992;
  assign n7551 = ~n6981 & n7550;
  assign n7552 = n6961 & ~n7551;
  assign n7553 = n6994 & ~n7013;
  assign n7554 = ~n6984 & n7553;
  assign n7555 = n6976 & ~n7554;
  assign n7556 = ~n7552 & ~n7555;
  assign n7557 = n7549 & n7556;
  assign n7558 = n7546 & n7557;
  assign n7559 = n6979 & n7558;
  assign n7560 = n7541 & n7559;
  assign n7561 = n7536 & n7560;
  assign n7562 = n7532 & n7561;
  assign n7563 = ~n6971 & n7562;
  assign n7564 = ~n6968 & n7563;
  assign n7565 = n7530 & n7564;
  assign n7566 = n7565 ^ n5203;
  assign n7567 = n7566 ^ x354;
  assign n7568 = n6470 & n6505;
  assign n7569 = n6204 & n6480;
  assign n7570 = ~n7568 & ~n7569;
  assign n7571 = ~n6203 & n6505;
  assign n7572 = n6470 & ~n6519;
  assign n7573 = ~n7571 & ~n7572;
  assign n7574 = n6204 & ~n6501;
  assign n7575 = ~n6204 & ~n6475;
  assign n7576 = ~n6488 & ~n6507;
  assign n7577 = ~n7575 & ~n7576;
  assign n7578 = n6470 & n6494;
  assign n7579 = n6468 & n6483;
  assign n7580 = ~n7578 & ~n7579;
  assign n7581 = n6436 ^ n6309;
  assign n7582 = n6436 ^ n6434;
  assign n7583 = n7582 ^ n6466;
  assign n7584 = n7581 & n7583;
  assign n7585 = n6475 & n7584;
  assign n7586 = n6466 ^ n6309;
  assign n7587 = n6466 ^ n6436;
  assign n7588 = n7582 & ~n7587;
  assign n7589 = n7586 & n7588;
  assign n7590 = n7589 ^ n7586;
  assign n7591 = ~n6470 & ~n7590;
  assign n7592 = ~n6509 & n6518;
  assign n7593 = n6470 & ~n7592;
  assign n7594 = ~n6483 & ~n7593;
  assign n7595 = ~n7591 & ~n7594;
  assign n7596 = ~n7585 & ~n7595;
  assign n7597 = n7580 & n7596;
  assign n7598 = ~n7577 & n7597;
  assign n7599 = ~n7574 & n7598;
  assign n7600 = n7573 & n7599;
  assign n7601 = n6497 & n7600;
  assign n7602 = n7570 & n7601;
  assign n7603 = ~n6482 & n7602;
  assign n7604 = n7603 ^ n5094;
  assign n7605 = n7604 ^ x355;
  assign n7606 = ~n7567 & ~n7605;
  assign n7607 = n6117 & n6130;
  assign n7608 = n5845 & n7607;
  assign n7609 = n5978 & n6158;
  assign n7610 = ~n7608 & ~n7609;
  assign n7611 = n5628 & n5977;
  assign n7612 = ~n5845 & n7611;
  assign n7613 = n7612 ^ n6134;
  assign n7614 = ~n6117 & n7613;
  assign n7615 = n7614 ^ n7612;
  assign n7616 = n6133 & ~n7615;
  assign n7617 = n7610 & n7616;
  assign n7618 = n6144 & ~n7617;
  assign n7619 = ~n6126 & ~n6139;
  assign n7620 = ~n6147 & n7619;
  assign n7621 = n5277 & ~n7620;
  assign n7622 = ~n7618 & ~n7621;
  assign n7623 = ~n5845 & n6118;
  assign n7624 = n6158 ^ n6134;
  assign n7625 = ~n5845 & n7624;
  assign n7626 = n7625 ^ n6134;
  assign n7627 = ~n7623 & ~n7626;
  assign n7628 = n6129 & ~n7627;
  assign n7629 = n5978 & ~n6117;
  assign n7630 = n6120 & ~n6158;
  assign n7631 = ~n7629 & ~n7630;
  assign n7632 = ~n6139 & n7631;
  assign n7633 = n6156 & ~n7632;
  assign n7634 = ~n7628 & ~n7633;
  assign n7635 = n7622 & n7634;
  assign n7636 = n7610 & n7635;
  assign n7637 = n7636 ^ n5161;
  assign n7638 = n7637 ^ x353;
  assign n7639 = n7270 & n7272;
  assign n7640 = n7284 & n7313;
  assign n7641 = ~n7639 & ~n7640;
  assign n7642 = n7284 & n7288;
  assign n7643 = ~n7285 & ~n7310;
  assign n7644 = n7272 & ~n7643;
  assign n7645 = ~n7642 & ~n7644;
  assign n7646 = ~n7296 & n7303;
  assign n7647 = n7277 & ~n7292;
  assign n7648 = ~n7312 & n7647;
  assign n7649 = ~n7281 & n7648;
  assign n7650 = n7186 & ~n7649;
  assign n7651 = ~n7646 & ~n7650;
  assign n7652 = n7645 & n7651;
  assign n7653 = ~n7291 & n7309;
  assign n7654 = ~n7297 & n7314;
  assign n7655 = n7291 & ~n7654;
  assign n7656 = n7281 & n7291;
  assign n7657 = n7294 & ~n7656;
  assign n7658 = ~n7281 & ~n7293;
  assign n7659 = ~n7284 & n7658;
  assign n7660 = ~n7657 & ~n7659;
  assign n7661 = ~n7302 & ~n7660;
  assign n7662 = ~n7310 & n7661;
  assign n7663 = ~n7296 & ~n7662;
  assign n7664 = ~n7655 & ~n7663;
  assign n7665 = ~n7653 & n7664;
  assign n7666 = n7652 & n7665;
  assign n7667 = ~n7283 & n7666;
  assign n7668 = n7641 & n7667;
  assign n7669 = ~n7267 & n7668;
  assign n7670 = n7279 & n7669;
  assign n7671 = n7670 ^ n5132;
  assign n7672 = n7671 ^ x356;
  assign n7673 = ~n7638 & n7672;
  assign n7674 = n7606 & n7673;
  assign n7675 = n7524 & n7674;
  assign n7676 = n7492 & n7523;
  assign n7677 = n7567 & ~n7605;
  assign n7678 = ~n7638 & ~n7672;
  assign n7679 = n7677 & n7678;
  assign n7680 = n7676 & n7679;
  assign n7681 = ~n7675 & ~n7680;
  assign n7682 = n7638 & ~n7672;
  assign n7683 = n7606 & n7682;
  assign n7684 = n7676 & n7683;
  assign n7685 = ~n7567 & n7605;
  assign n7686 = n7638 & n7672;
  assign n7687 = n7685 & n7686;
  assign n7688 = n7676 & n7687;
  assign n7689 = n7682 & n7685;
  assign n7690 = n7524 & n7689;
  assign n7691 = ~n7688 & ~n7690;
  assign n7692 = n7492 & ~n7523;
  assign n7693 = n7567 & n7605;
  assign n7694 = n7682 & n7693;
  assign n7695 = n7692 & n7694;
  assign n7696 = ~n7492 & n7523;
  assign n7697 = n7606 & n7686;
  assign n7698 = n7677 & n7682;
  assign n7699 = ~n7697 & ~n7698;
  assign n7700 = n7696 & ~n7699;
  assign n7701 = ~n7695 & ~n7700;
  assign n7702 = n7691 & n7701;
  assign n7703 = n7673 & n7677;
  assign n7704 = n7696 & n7703;
  assign n7705 = n7686 & n7693;
  assign n7706 = n7524 & n7705;
  assign n7707 = ~n7704 & ~n7706;
  assign n7708 = n7673 & n7693;
  assign n7709 = n7606 & n7678;
  assign n7710 = ~n7708 & ~n7709;
  assign n7711 = n7676 & ~n7710;
  assign n7712 = n7677 & n7686;
  assign n7713 = ~n7683 & ~n7712;
  assign n7714 = n7692 & ~n7713;
  assign n7715 = ~n7711 & ~n7714;
  assign n7716 = n7707 & n7715;
  assign n7717 = n7676 & n7705;
  assign n7718 = n7692 & n7705;
  assign n7719 = ~n7674 & ~n7694;
  assign n7720 = n7676 & ~n7719;
  assign n7721 = ~n7718 & ~n7720;
  assign n7722 = ~n7687 & ~n7698;
  assign n7723 = n7524 & ~n7722;
  assign n7724 = n7678 & n7685;
  assign n7725 = ~n7708 & ~n7724;
  assign n7726 = ~n7712 & n7725;
  assign n7727 = ~n7694 & n7726;
  assign n7728 = ~n7689 & n7727;
  assign n7729 = n7696 & ~n7728;
  assign n7730 = n7678 & n7693;
  assign n7731 = ~n7679 & ~n7730;
  assign n7732 = ~n7692 & n7731;
  assign n7733 = n7673 & n7685;
  assign n7734 = ~n7679 & ~n7733;
  assign n7735 = ~n7524 & n7734;
  assign n7736 = ~n7674 & n7735;
  assign n7737 = ~n7732 & ~n7736;
  assign n7738 = ~n7703 & ~n7737;
  assign n7739 = ~n7523 & ~n7738;
  assign n7740 = ~n7729 & ~n7739;
  assign n7741 = ~n7723 & n7740;
  assign n7742 = n7721 & n7741;
  assign n7743 = ~n7717 & n7742;
  assign n7744 = n7716 & n7743;
  assign n7745 = n7702 & n7744;
  assign n7746 = ~n7684 & n7745;
  assign n7747 = n7681 & n7746;
  assign n7748 = n7747 ^ n5275;
  assign n7749 = n7748 ^ x423;
  assign n7750 = ~n7393 & n7749;
  assign n7751 = n7522 ^ x359;
  assign n7752 = n7115 & ~n7130;
  assign n7753 = n7089 & ~n7101;
  assign n7754 = ~n7752 & ~n7753;
  assign n7755 = n7038 & n7128;
  assign n7756 = ~n7122 & ~n7755;
  assign n7757 = n7089 & n7108;
  assign n7758 = n7123 & n7128;
  assign n7759 = ~n7757 & ~n7758;
  assign n7760 = ~n7129 & ~n7134;
  assign n7761 = n7104 & ~n7760;
  assign n7762 = ~n7099 & n7139;
  assign n7763 = n7038 & ~n7762;
  assign n7764 = n7089 & n7135;
  assign n7765 = ~n7117 & n7123;
  assign n7766 = ~n7764 & ~n7765;
  assign n7767 = ~n7037 & n7111;
  assign n7768 = n7123 & ~n7139;
  assign n7769 = ~n7767 & ~n7768;
  assign n7770 = ~n7105 & ~n7121;
  assign n7771 = n7089 & ~n7770;
  assign n7772 = ~n7112 & ~n7125;
  assign n7773 = n7101 & n7772;
  assign n7774 = n7115 & ~n7773;
  assign n7775 = ~n7771 & ~n7774;
  assign n7776 = n7769 & n7775;
  assign n7777 = n7766 & n7776;
  assign n7778 = ~n7763 & n7777;
  assign n7779 = ~n7761 & n7778;
  assign n7780 = n7759 & n7779;
  assign n7781 = ~n7096 & n7780;
  assign n7782 = n7756 & n7781;
  assign n7783 = n7754 & n7782;
  assign n7784 = ~n7120 & n7783;
  assign n7785 = ~n7088 & n7784;
  assign n7786 = n7785 ^ n6003;
  assign n7787 = n7786 ^ x360;
  assign n7788 = n7751 & n7787;
  assign n7789 = n7445 & n7453;
  assign n7790 = n7463 & n7789;
  assign n7791 = ~n7447 & n7480;
  assign n7792 = ~n7790 & ~n7791;
  assign n7793 = ~n7439 & n7792;
  assign n7794 = n7465 & n7480;
  assign n7795 = n7441 & n7445;
  assign n7796 = n7396 & n7795;
  assign n7797 = ~n7794 & ~n7796;
  assign n7798 = n7480 & n7795;
  assign n7799 = n7438 & n7444;
  assign n7800 = n7440 & n7446;
  assign n7801 = ~n7799 & ~n7800;
  assign n7802 = ~n7455 & n7463;
  assign n7803 = n7437 & n7457;
  assign n7804 = ~n7465 & ~n7803;
  assign n7805 = ~n7476 & n7804;
  assign n7806 = n7396 & ~n7805;
  assign n7807 = ~n7802 & ~n7806;
  assign n7808 = n7801 & n7807;
  assign n7809 = n7464 & n7480;
  assign n7810 = ~n7472 & ~n7803;
  assign n7811 = ~n7466 & n7810;
  assign n7812 = n7481 & n7811;
  assign n7813 = ~n7458 & n7812;
  assign n7814 = ~n7473 & n7813;
  assign n7815 = ~n7463 & ~n7814;
  assign n7816 = ~n7809 & ~n7815;
  assign n7817 = n7808 & n7816;
  assign n7818 = ~n7798 & n7817;
  assign n7819 = n7797 & n7818;
  assign n7820 = n7793 & n7819;
  assign n7821 = n7820 ^ n6038;
  assign n7822 = n7821 ^ x361;
  assign n7823 = n6204 & n6494;
  assign n7824 = ~n6499 & ~n6509;
  assign n7825 = n6475 & ~n7824;
  assign n7826 = ~n7823 & ~n7825;
  assign n7827 = ~n6507 & n6518;
  assign n7828 = n6204 & ~n7827;
  assign n7829 = n6506 & n7576;
  assign n7830 = n6483 & ~n7829;
  assign n7831 = ~n7828 & ~n7830;
  assign n7832 = n6475 & ~n6524;
  assign n7833 = ~n6484 & ~n6492;
  assign n7834 = n6511 & n7833;
  assign n7835 = ~n6490 & n7834;
  assign n7836 = n6470 & ~n7835;
  assign n7837 = ~n7832 & ~n7836;
  assign n7838 = n7831 & n7837;
  assign n7839 = n7570 & n7838;
  assign n7840 = n6498 & n7839;
  assign n7841 = n7826 & n7840;
  assign n7842 = ~n6486 & n7841;
  assign n7843 = n6474 & n7842;
  assign n7844 = n7843 ^ n5675;
  assign n7845 = n7844 ^ x362;
  assign n7846 = ~n7822 & n7845;
  assign n7847 = n7788 & n7846;
  assign n7848 = n7751 & ~n7787;
  assign n7849 = n7822 & ~n7845;
  assign n7850 = n7848 & n7849;
  assign n7851 = ~n7847 & ~n7850;
  assign n7852 = n6562 ^ x305;
  assign n7853 = n5569 & n5602;
  assign n7854 = n6863 & n7168;
  assign n7855 = n5565 & ~n7854;
  assign n7856 = ~n7853 & ~n7855;
  assign n7857 = n5572 & ~n5611;
  assign n7858 = n5596 & n5614;
  assign n7859 = n5561 & ~n7858;
  assign n7860 = ~n5583 & ~n5592;
  assign n7861 = ~n5601 & ~n7860;
  assign n7862 = ~n7859 & ~n7861;
  assign n7863 = ~n7857 & n7862;
  assign n7864 = n7856 & n7863;
  assign n7865 = n7157 & n7864;
  assign n7866 = n6853 & n7865;
  assign n7867 = n5576 & n7866;
  assign n7868 = n6843 & n7867;
  assign n7869 = ~n6866 & n7868;
  assign n7870 = ~n5562 & n7869;
  assign n7871 = n7870 ^ n5381;
  assign n7872 = n7871 ^ x307;
  assign n7873 = n7852 & ~n7872;
  assign n7874 = n6078 & n6100;
  assign n7875 = ~n6086 & n6102;
  assign n7876 = n5982 & ~n7875;
  assign n7877 = ~n7874 & ~n7876;
  assign n7878 = n6053 & ~n6099;
  assign n7879 = ~n6565 & ~n6571;
  assign n7880 = n6048 & n6094;
  assign n7881 = ~n6057 & ~n6095;
  assign n7882 = n5982 & ~n7881;
  assign n7883 = ~n7880 & ~n7882;
  assign n7884 = n6076 & n6078;
  assign n7885 = ~n6086 & n6567;
  assign n7886 = ~n6053 & n7885;
  assign n7887 = ~n6048 & ~n6081;
  assign n7888 = n7875 & n7887;
  assign n7889 = ~n7886 & ~n7888;
  assign n7890 = ~n6571 & n7889;
  assign n7891 = ~n7884 & ~n7890;
  assign n7892 = n7883 & n7891;
  assign n7893 = n6085 & n7892;
  assign n7894 = n6080 & n7893;
  assign n7895 = ~n7879 & n7894;
  assign n7896 = ~n7878 & n7895;
  assign n7897 = n7877 & n7896;
  assign n7898 = n6443 & n7897;
  assign n7899 = n7898 ^ n5413;
  assign n7900 = n7899 ^ x306;
  assign n7901 = n6957 ^ x308;
  assign n7902 = n7900 & ~n7901;
  assign n7903 = n7873 & n7902;
  assign n7904 = n6676 ^ x304;
  assign n7905 = n6810 ^ x309;
  assign n7906 = ~n7904 & n7905;
  assign n7907 = n7852 & n7872;
  assign n7908 = n7900 & n7901;
  assign n7909 = n7907 & n7908;
  assign n7910 = n7906 & n7909;
  assign n7911 = ~n7904 & ~n7905;
  assign n7912 = ~n7852 & ~n7872;
  assign n7913 = ~n7900 & n7901;
  assign n7914 = n7912 & n7913;
  assign n7915 = n7911 & n7914;
  assign n7916 = n7904 & ~n7905;
  assign n7917 = ~n7852 & n7872;
  assign n7918 = n7913 & n7917;
  assign n7919 = n7916 & n7918;
  assign n7920 = ~n7915 & ~n7919;
  assign n7921 = ~n7910 & n7920;
  assign n7922 = n7904 & n7905;
  assign n7923 = ~n7900 & ~n7901;
  assign n7924 = n7907 & n7923;
  assign n7925 = n7922 & n7924;
  assign n7926 = n7873 & n7923;
  assign n7927 = n7922 & n7926;
  assign n7928 = n7909 & n7922;
  assign n7929 = n7908 & n7912;
  assign n7930 = n7906 & n7929;
  assign n7931 = ~n7928 & ~n7930;
  assign n7932 = n7907 & n7913;
  assign n7933 = n7906 & n7932;
  assign n7934 = ~n7911 & ~n7922;
  assign n7935 = n7902 & n7917;
  assign n7936 = ~n7934 & n7935;
  assign n7937 = ~n7933 & ~n7936;
  assign n7938 = n7902 & n7912;
  assign n7939 = ~n7929 & ~n7938;
  assign n7940 = ~n7914 & n7939;
  assign n7941 = n7922 & ~n7940;
  assign n7942 = n7908 & n7917;
  assign n7943 = n7917 & n7923;
  assign n7944 = ~n7942 & ~n7943;
  assign n7945 = n7873 & n7913;
  assign n7946 = n7873 & n7908;
  assign n7947 = n7902 & n7907;
  assign n7948 = ~n7946 & ~n7947;
  assign n7949 = ~n7945 & n7948;
  assign n7950 = n7944 & n7949;
  assign n7951 = ~n7938 & n7950;
  assign n7952 = n7916 & ~n7951;
  assign n7953 = n7912 & n7923;
  assign n7954 = ~n7914 & ~n7953;
  assign n7955 = n7944 & n7954;
  assign n7956 = n7906 & ~n7955;
  assign n7957 = ~n7926 & n7948;
  assign n7958 = ~n7918 & n7957;
  assign n7959 = ~n7924 & n7958;
  assign n7960 = n7911 & ~n7959;
  assign n7961 = ~n7956 & ~n7960;
  assign n7962 = ~n7952 & n7961;
  assign n7963 = ~n7941 & n7962;
  assign n7964 = n7937 & n7963;
  assign n7965 = n7931 & n7964;
  assign n7966 = ~n7927 & n7965;
  assign n7967 = ~n7925 & n7966;
  assign n7968 = n7921 & n7967;
  assign n7969 = ~n7903 & n7968;
  assign n7970 = n7969 ^ n5727;
  assign n7971 = n7970 ^ x363;
  assign n7972 = n7671 ^ x358;
  assign n7973 = ~n7971 & ~n7972;
  assign n7974 = ~n7851 & n7973;
  assign n7975 = ~n7751 & n7787;
  assign n7976 = n7846 & n7975;
  assign n7977 = ~n7751 & ~n7787;
  assign n7978 = n7849 & n7977;
  assign n7979 = ~n7976 & ~n7978;
  assign n7980 = n7971 & ~n7972;
  assign n7981 = ~n7979 & n7980;
  assign n7982 = ~n7822 & ~n7845;
  assign n7983 = n7977 & n7982;
  assign n7984 = ~n7971 & n7972;
  assign n7985 = n7983 & n7984;
  assign n7986 = n7788 & n7849;
  assign n7987 = n7980 & n7986;
  assign n7988 = n7822 & n7845;
  assign n7989 = n7975 & n7988;
  assign n7990 = n7984 & n7989;
  assign n7991 = n7848 & n7988;
  assign n7992 = n7971 & n7972;
  assign n7993 = n7991 & n7992;
  assign n7994 = ~n7990 & ~n7993;
  assign n7995 = ~n7987 & n7994;
  assign n7996 = ~n7985 & n7995;
  assign n7997 = n7847 & n7971;
  assign n7998 = n7850 & n7972;
  assign n7999 = ~n7997 & ~n7998;
  assign n8000 = n7977 & n7988;
  assign n8001 = ~n7845 & n7975;
  assign n8002 = ~n7822 & n8001;
  assign n8003 = ~n8000 & ~n8002;
  assign n8004 = n7992 & ~n8003;
  assign n8005 = n7822 & n8001;
  assign n8006 = n7846 & n7848;
  assign n8007 = ~n8000 & ~n8006;
  assign n8008 = ~n8005 & n8007;
  assign n8009 = n7973 & ~n8008;
  assign n8010 = ~n8004 & ~n8009;
  assign n8011 = n7846 & n7977;
  assign n8012 = ~n7983 & ~n8011;
  assign n8013 = ~n7986 & n8012;
  assign n8014 = n7972 ^ n7971;
  assign n8015 = ~n8013 & ~n8014;
  assign n8016 = n7848 & n7982;
  assign n8017 = ~n7991 & ~n8016;
  assign n8018 = ~n7989 & ~n8002;
  assign n8019 = n8017 & n8018;
  assign n8020 = n7980 & ~n8019;
  assign n8021 = n7788 & n7988;
  assign n8022 = ~n7976 & ~n8021;
  assign n8023 = n7788 & n7982;
  assign n8024 = ~n8006 & ~n8023;
  assign n8025 = n8022 & n8024;
  assign n8026 = ~n7978 & n8025;
  assign n8027 = n7984 & ~n8026;
  assign n8028 = ~n8020 & ~n8027;
  assign n8029 = ~n8015 & n8028;
  assign n8030 = n8010 & n8029;
  assign n8031 = n7999 & n8030;
  assign n8032 = n7996 & n8031;
  assign n8033 = ~n7981 & n8032;
  assign n8034 = ~n7974 & n8033;
  assign n8035 = n8034 ^ n6116;
  assign n8036 = n8035 ^ x419;
  assign n8037 = n6959 & n7007;
  assign n8038 = n6982 & ~n6994;
  assign n8039 = ~n8037 & ~n8038;
  assign n8040 = ~n6970 & ~n6981;
  assign n8041 = n6959 & ~n8040;
  assign n8042 = ~n6975 & ~n6993;
  assign n8043 = n6976 & ~n8042;
  assign n8044 = ~n8041 & ~n8043;
  assign n8045 = ~n6973 & ~n6984;
  assign n8046 = n6982 & ~n8045;
  assign n8047 = ~n6971 & n7534;
  assign n8048 = ~n6967 & n8047;
  assign n8049 = ~n6997 & n8048;
  assign n8050 = ~n6977 & ~n8049;
  assign n8051 = ~n8046 & ~n8050;
  assign n8052 = n8044 & n8051;
  assign n8053 = n7546 & n8052;
  assign n8054 = n8039 & n8053;
  assign n8055 = n7541 & n8054;
  assign n8056 = ~n7015 & n8055;
  assign n8057 = n6965 & n8056;
  assign n8058 = n7530 & n8057;
  assign n8059 = n8058 ^ n5644;
  assign n8060 = n8059 ^ x369;
  assign n8061 = n7844 ^ x364;
  assign n8062 = n8060 & n8061;
  assign n8063 = n7396 & ~n7482;
  assign n8064 = n7444 & n7485;
  assign n8065 = ~n8063 & ~n8064;
  assign n8066 = n7435 & n7480;
  assign n8067 = ~n7395 & ~n7810;
  assign n8068 = ~n8066 & ~n8067;
  assign n8069 = ~n7394 & ~n7480;
  assign n8070 = ~n7467 & ~n8069;
  assign n8071 = ~n7464 & ~n7476;
  assign n8072 = ~n7452 & n8071;
  assign n8073 = ~n7438 & n8072;
  assign n8074 = n7440 & ~n8073;
  assign n8075 = ~n8070 & ~n8074;
  assign n8076 = n8068 & n8075;
  assign n8077 = n8065 & n8076;
  assign n8078 = n7793 & n8077;
  assign n8079 = ~n7436 & n8078;
  assign n8080 = n8079 ^ n5697;
  assign n8081 = n8080 ^ x368;
  assign n8082 = n7970 ^ x365;
  assign n8083 = n8081 & ~n8082;
  assign n8084 = n6156 & n7617;
  assign n8085 = n6129 & n7620;
  assign n8086 = n7610 & n8085;
  assign n8087 = ~n8084 & ~n8086;
  assign n8088 = n7610 & n7627;
  assign n8089 = n5277 & ~n8088;
  assign n8090 = ~n7608 & n7632;
  assign n8091 = n6144 & ~n8090;
  assign n8092 = ~n8089 & ~n8091;
  assign n8093 = n8087 & n8092;
  assign n8094 = n8093 ^ n5742;
  assign n8095 = n8094 ^ x366;
  assign n8096 = n7270 & n7284;
  assign n8097 = n7291 & n7313;
  assign n8098 = ~n8096 & ~n8097;
  assign n8099 = ~n7288 & ~n7312;
  assign n8100 = ~n7296 & ~n8099;
  assign n8101 = ~n7302 & ~n7309;
  assign n8102 = ~n7285 & n8101;
  assign n8103 = n7272 & ~n8102;
  assign n8104 = ~n8100 & ~n8103;
  assign n8105 = ~n7274 & n8101;
  assign n8106 = ~n7266 & n8105;
  assign n8107 = n7291 & ~n8106;
  assign n8108 = ~n7303 & n7643;
  assign n8109 = n7658 & n8108;
  assign n8110 = n7284 & ~n8109;
  assign n8111 = n7272 & ~n7314;
  assign n8112 = ~n7276 & n8101;
  assign n8113 = ~n7297 & n8112;
  assign n8114 = ~n7313 & n8113;
  assign n8115 = n7186 & ~n8114;
  assign n8116 = ~n8111 & ~n8115;
  assign n8117 = ~n8110 & n8116;
  assign n8118 = ~n8107 & n8117;
  assign n8119 = n8104 & n8118;
  assign n8120 = n8098 & n8119;
  assign n8121 = ~n7656 & n8120;
  assign n8122 = n7301 & n8121;
  assign n8123 = n7279 & n8122;
  assign n8124 = n8123 ^ n5770;
  assign n8125 = n8124 ^ x367;
  assign n8126 = ~n8095 & n8125;
  assign n8127 = n8083 & n8126;
  assign n8128 = n8062 & n8127;
  assign n8129 = ~n8060 & ~n8061;
  assign n8130 = n8081 & n8082;
  assign n8131 = n8095 & ~n8125;
  assign n8132 = n8130 & n8131;
  assign n8133 = n8129 & n8132;
  assign n8134 = ~n8128 & ~n8133;
  assign n8135 = ~n8081 & ~n8082;
  assign n8136 = n8126 & n8135;
  assign n8137 = n8062 & n8136;
  assign n8138 = ~n8095 & ~n8125;
  assign n8139 = n8130 & n8138;
  assign n8140 = n8129 & n8139;
  assign n8141 = ~n8137 & ~n8140;
  assign n8142 = ~n8081 & n8082;
  assign n8143 = n8095 & n8142;
  assign n8144 = n8129 & n8143;
  assign n8145 = n8060 & ~n8061;
  assign n8146 = n8132 & n8145;
  assign n8147 = ~n8144 & ~n8146;
  assign n8148 = ~n8060 & n8061;
  assign n8149 = n8139 & n8148;
  assign n8150 = n8095 & n8125;
  assign n8151 = n8083 & n8150;
  assign n8152 = n8131 & n8135;
  assign n8153 = ~n8151 & ~n8152;
  assign n8154 = n8062 & ~n8153;
  assign n8155 = ~n8149 & ~n8154;
  assign n8156 = n8061 ^ n8060;
  assign n8157 = n8130 & n8150;
  assign n8158 = n8126 & n8130;
  assign n8159 = n8138 & n8142;
  assign n8160 = ~n8158 & ~n8159;
  assign n8161 = ~n8157 & n8160;
  assign n8162 = n8156 & ~n8161;
  assign n8163 = ~n8139 & ~n8159;
  assign n8164 = ~n8143 & n8163;
  assign n8165 = n8062 & ~n8164;
  assign n8166 = ~n8127 & ~n8136;
  assign n8167 = n8135 & n8138;
  assign n8168 = ~n8151 & ~n8167;
  assign n8169 = n8166 & n8168;
  assign n8170 = n8129 & ~n8169;
  assign n8171 = ~n8165 & ~n8170;
  assign n8172 = n8135 & n8150;
  assign n8173 = n8083 & n8131;
  assign n8174 = ~n8172 & ~n8173;
  assign n8175 = n8126 & n8142;
  assign n8176 = ~n8167 & ~n8175;
  assign n8177 = n8174 & n8176;
  assign n8178 = n8145 & ~n8177;
  assign n8179 = n8083 & n8138;
  assign n8180 = n8174 & ~n8179;
  assign n8181 = ~n8152 & n8180;
  assign n8182 = n8148 & ~n8181;
  assign n8183 = ~n8178 & ~n8182;
  assign n8184 = n8171 & n8183;
  assign n8185 = ~n8162 & n8184;
  assign n8186 = n8155 & n8185;
  assign n8187 = n8147 & n8186;
  assign n8188 = n8141 & n8187;
  assign n8189 = n8134 & n8188;
  assign n8190 = n8189 ^ n5844;
  assign n8191 = n8190 ^ x422;
  assign n8192 = n7637 ^ x399;
  assign n8193 = n7032 ^ x394;
  assign n8194 = ~n8192 & ~n8193;
  assign n8195 = n7491 ^ x398;
  assign n8196 = n7922 & n7938;
  assign n8197 = ~n7945 & ~n7947;
  assign n8198 = ~n7903 & n8197;
  assign n8199 = n7906 & ~n8198;
  assign n8200 = ~n8196 & ~n8199;
  assign n8201 = n7904 & n7929;
  assign n8202 = n7922 & n7943;
  assign n8203 = ~n8201 & ~n8202;
  assign n8204 = ~n7934 & n7942;
  assign n8205 = ~n7926 & n8198;
  assign n8206 = ~n7935 & n8205;
  assign n8207 = ~n7924 & n8206;
  assign n8208 = n7916 & ~n8207;
  assign n8209 = ~n8204 & ~n8208;
  assign n8210 = ~n7938 & ~n7953;
  assign n8211 = n7911 & ~n8210;
  assign n8212 = ~n7918 & ~n7953;
  assign n8213 = n7939 & n8212;
  assign n8214 = n7906 & ~n8213;
  assign n8215 = ~n7932 & ~n7946;
  assign n8216 = ~n7911 & n8215;
  assign n8217 = ~n7909 & ~n7924;
  assign n8218 = ~n7922 & n8217;
  assign n8219 = n7948 & n8218;
  assign n8220 = ~n8216 & ~n8219;
  assign n8221 = ~n7934 & n8220;
  assign n8222 = ~n8214 & ~n8221;
  assign n8223 = ~n8211 & n8222;
  assign n8224 = n8209 & n8223;
  assign n8225 = n8203 & n8224;
  assign n8226 = n8200 & n8225;
  assign n8227 = ~n7927 & n8226;
  assign n8228 = ~n7925 & n8227;
  assign n8229 = n7921 & n8228;
  assign n8230 = n8229 ^ n5872;
  assign n8231 = n8230 ^ x397;
  assign n8232 = n8195 & n8231;
  assign n8233 = n7094 & n7104;
  assign n8234 = ~n7087 & ~n7134;
  assign n8235 = n7115 & ~n8234;
  assign n8236 = ~n8233 & ~n8235;
  assign n8237 = n7089 & ~n7130;
  assign n8238 = n7037 & ~n7139;
  assign n8239 = ~n8237 & ~n8238;
  assign n8240 = n8236 & n8239;
  assign n8241 = n7038 & ~n7113;
  assign n8242 = ~n7092 & ~n7128;
  assign n8243 = n7123 & ~n8242;
  assign n8244 = ~n7105 & ~n7116;
  assign n8245 = n7101 & n8244;
  assign n8246 = ~n7123 & n8245;
  assign n8247 = ~n7108 & ~n7116;
  assign n8248 = ~n7111 & n8247;
  assign n8249 = ~n7087 & n8248;
  assign n8250 = ~n7115 & n8249;
  assign n8251 = ~n8246 & ~n8250;
  assign n8252 = ~n8243 & ~n8251;
  assign n8253 = ~n8241 & n8252;
  assign n8254 = n8240 & n8253;
  assign n8255 = n7103 & n8254;
  assign n8256 = n7754 & n8255;
  assign n8257 = ~n7124 & n8256;
  assign n8258 = ~n7122 & n8257;
  assign n8259 = n8258 ^ n5906;
  assign n8260 = n8259 ^ x396;
  assign n8261 = n7328 ^ x395;
  assign n8262 = ~n8260 & ~n8261;
  assign n8263 = n8232 & n8262;
  assign n8264 = n8194 & n8263;
  assign n8265 = n8192 & n8193;
  assign n8266 = ~n8195 & n8231;
  assign n8267 = n8262 & n8266;
  assign n8268 = n8260 & ~n8261;
  assign n8269 = n8232 & n8268;
  assign n8270 = ~n8267 & ~n8269;
  assign n8271 = n8265 & ~n8270;
  assign n8272 = ~n8264 & ~n8271;
  assign n8273 = ~n8195 & ~n8231;
  assign n8274 = n8260 & n8261;
  assign n8275 = n8273 & n8274;
  assign n8276 = n8265 & n8275;
  assign n8277 = ~n8260 & n8261;
  assign n8278 = n8266 & n8277;
  assign n8279 = n8194 & n8278;
  assign n8280 = n8266 & n8268;
  assign n8281 = n8194 & n8280;
  assign n8282 = ~n8192 & n8193;
  assign n8283 = n8232 & n8277;
  assign n8284 = n8232 & n8274;
  assign n8285 = ~n8283 & ~n8284;
  assign n8286 = n8282 & ~n8285;
  assign n8287 = n8192 & ~n8193;
  assign n8288 = n8268 & n8273;
  assign n8289 = ~n8269 & ~n8288;
  assign n8290 = n8287 & ~n8289;
  assign n8291 = ~n8286 & ~n8290;
  assign n8292 = n8273 & n8277;
  assign n8293 = n8282 & n8292;
  assign n8294 = n8266 & n8274;
  assign n8295 = n8193 & n8294;
  assign n8296 = ~n8293 & ~n8295;
  assign n8297 = ~n8263 & ~n8280;
  assign n8298 = n8287 & ~n8297;
  assign n8299 = n8195 & ~n8231;
  assign n8300 = n8262 & n8299;
  assign n8301 = n8262 & n8273;
  assign n8302 = n8274 & n8299;
  assign n8303 = ~n8278 & ~n8302;
  assign n8304 = ~n8301 & n8303;
  assign n8305 = ~n8300 & n8304;
  assign n8306 = n8265 & ~n8305;
  assign n8307 = ~n8298 & ~n8306;
  assign n8308 = n8277 & n8299;
  assign n8309 = ~n8292 & ~n8302;
  assign n8310 = n8289 & n8309;
  assign n8311 = ~n8308 & n8310;
  assign n8312 = n8194 & ~n8311;
  assign n8313 = ~n8284 & n8309;
  assign n8314 = ~n8308 & n8313;
  assign n8315 = n8287 & ~n8314;
  assign n8316 = n8260 ^ n8231;
  assign n8317 = ~n8261 & n8316;
  assign n8318 = n8282 & n8317;
  assign n8319 = ~n8315 & ~n8318;
  assign n8320 = ~n8312 & n8319;
  assign n8321 = n8307 & n8320;
  assign n8322 = n8296 & n8321;
  assign n8323 = n8291 & n8322;
  assign n8324 = ~n8281 & n8323;
  assign n8325 = ~n8279 & n8324;
  assign n8326 = ~n8276 & n8325;
  assign n8327 = n8272 & n8326;
  assign n8328 = n8327 ^ n5976;
  assign n8329 = n8328 ^ x421;
  assign n8330 = n8191 & ~n8329;
  assign n8331 = n8036 & n8330;
  assign n8547 = ~n8191 & n8329;
  assign n8332 = n6712 & n6760;
  assign n8333 = n6722 & ~n6764;
  assign n8334 = ~n8332 & ~n8333;
  assign n8335 = ~n6752 & n6759;
  assign n8336 = n6724 & ~n6768;
  assign n8337 = n6733 & n8336;
  assign n8338 = ~n8335 & ~n8337;
  assign n8339 = n6718 & n6722;
  assign n8340 = ~n6731 & ~n6763;
  assign n8341 = n6712 & ~n8340;
  assign n8342 = ~n8339 & ~n8341;
  assign n8343 = n6587 & n6761;
  assign n8344 = n6768 & n7501;
  assign n8345 = ~n6740 & n8344;
  assign n8346 = n6588 & ~n8345;
  assign n8347 = ~n8343 & ~n8346;
  assign n8348 = n8342 & n8347;
  assign n8349 = n8338 & n8348;
  assign n8350 = ~n6742 & n8349;
  assign n8351 = n7498 & n8350;
  assign n8352 = n8334 & n8351;
  assign n8353 = n6751 & n8352;
  assign n8354 = n7495 & n8353;
  assign n8355 = ~n6745 & n8354;
  assign n8356 = n6730 & n8355;
  assign n8357 = n8356 ^ n5518;
  assign n8358 = n8357 ^ x381;
  assign n8359 = n7092 & n7104;
  assign n8360 = n7038 & n7094;
  assign n8361 = ~n7129 & ~n7135;
  assign n8362 = n7115 & ~n8361;
  assign n8363 = n7760 & n7772;
  assign n8364 = ~n7099 & n8363;
  assign n8365 = ~n7092 & n8364;
  assign n8366 = n7089 & ~n8365;
  assign n8367 = ~n8362 & ~n8366;
  assign n8368 = ~n7037 & n7134;
  assign n8369 = ~n7100 & ~n7105;
  assign n8370 = n7123 & ~n8369;
  assign n8371 = ~n7111 & n8244;
  assign n8372 = n7038 & ~n8371;
  assign n8373 = ~n7099 & n7140;
  assign n8374 = n7115 & ~n8373;
  assign n8375 = ~n8372 & ~n8374;
  assign n8376 = ~n8370 & n8375;
  assign n8377 = ~n8368 & n8376;
  assign n8378 = n8367 & n8377;
  assign n8379 = n7766 & n8378;
  assign n8380 = ~n7088 & n8379;
  assign n8381 = ~n8360 & n8380;
  assign n8382 = ~n8359 & n8381;
  assign n8383 = n7759 & n8382;
  assign n8384 = n7756 & n8383;
  assign n8385 = ~n7120 & n8384;
  assign n8386 = ~n7124 & n8385;
  assign n8387 = n8386 ^ n5559;
  assign n8388 = n8387 ^ x376;
  assign n8389 = n8358 & n8388;
  assign n8390 = n6154 & n6156;
  assign n8391 = ~n6127 & n6129;
  assign n8392 = ~n8390 & ~n8391;
  assign n8393 = n5277 & ~n6141;
  assign n8394 = n6144 & ~n6162;
  assign n8395 = ~n8393 & ~n8394;
  assign n8396 = n8392 & n8395;
  assign n8397 = n8396 ^ n5295;
  assign n8398 = n8397 ^ x380;
  assign n8399 = n6976 & ~n6998;
  assign n8400 = ~n6910 & ~n6997;
  assign n8401 = ~n6975 & n8400;
  assign n8402 = n6982 & ~n8401;
  assign n8403 = ~n8399 & ~n8402;
  assign n8404 = ~n6992 & ~n7005;
  assign n8405 = ~n6963 & n8404;
  assign n8406 = n6959 & ~n8405;
  assign n8407 = n6994 & ~n7005;
  assign n8408 = ~n6975 & n8407;
  assign n8409 = n6961 & ~n8408;
  assign n8410 = ~n8406 & ~n8409;
  assign n8411 = n8403 & n8410;
  assign n8412 = ~n6991 & n8411;
  assign n8413 = n6986 & n8412;
  assign n8414 = n8039 & n8413;
  assign n8415 = n7536 & n8414;
  assign n8416 = n7532 & n8415;
  assign n8417 = ~n6968 & n8416;
  assign n8418 = n6965 & n8417;
  assign n8419 = n7530 & n8418;
  assign n8420 = n8419 ^ n5346;
  assign n8421 = n8420 ^ x378;
  assign n8422 = ~n8398 & ~n8421;
  assign n8423 = n7944 & ~n7946;
  assign n8424 = ~n7924 & n8423;
  assign n8425 = n7906 & ~n8424;
  assign n8426 = n7940 & n7957;
  assign n8427 = ~n7909 & n8426;
  assign n8428 = n7916 & ~n8427;
  assign n8429 = ~n8425 & ~n8428;
  assign n8430 = ~n7935 & n7939;
  assign n8431 = n7911 & ~n8430;
  assign n8432 = ~n7942 & n7954;
  assign n8433 = n7922 & ~n8432;
  assign n8434 = ~n7911 & ~n7947;
  assign n8435 = ~n7903 & n8218;
  assign n8436 = ~n8434 & ~n8435;
  assign n8437 = ~n7932 & ~n8436;
  assign n8438 = ~n7934 & ~n8437;
  assign n8439 = ~n8433 & ~n8438;
  assign n8440 = ~n8431 & n8439;
  assign n8441 = n8429 & n8440;
  assign n8442 = n7920 & n8441;
  assign n8443 = n7931 & n8442;
  assign n8444 = n8200 & n8443;
  assign n8445 = ~n7927 & n8444;
  assign n8446 = n8445 ^ n5488;
  assign n8447 = n8446 ^ x377;
  assign n8448 = n7266 & n7284;
  assign n8449 = n7186 & n7310;
  assign n8450 = n7276 & ~n7296;
  assign n8451 = ~n7274 & ~n7297;
  assign n8452 = ~n7312 & n8451;
  assign n8453 = n7272 & ~n8452;
  assign n8454 = ~n8450 & ~n8453;
  assign n8455 = n8101 & n8108;
  assign n8456 = ~n7288 & n8455;
  assign n8457 = n7291 & ~n8456;
  assign n8458 = n7277 & ~n7313;
  assign n8459 = ~n7288 & n8458;
  assign n8460 = n7186 & ~n8459;
  assign n8461 = ~n8457 & ~n8460;
  assign n8462 = n7284 & ~n7643;
  assign n8463 = ~n7281 & ~n7309;
  assign n8464 = n7272 & ~n8463;
  assign n8465 = ~n8462 & ~n8464;
  assign n8466 = n7294 & n8465;
  assign n8467 = ~n7184 & ~n8466;
  assign n8468 = n8461 & ~n8467;
  assign n8469 = n8454 & n8468;
  assign n8470 = ~n8449 & n8469;
  assign n8471 = ~n8448 & n8470;
  assign n8472 = ~n7300 & n8471;
  assign n8473 = n7641 & n8472;
  assign n8474 = n8098 & n8473;
  assign n8475 = ~n7267 & n8474;
  assign n8476 = n8475 ^ n5323;
  assign n8477 = n8476 ^ x379;
  assign n8478 = ~n8447 & ~n8477;
  assign n8479 = n8422 & n8478;
  assign n8480 = n8389 & n8479;
  assign n8481 = n8358 & ~n8388;
  assign n8482 = ~n8398 & n8421;
  assign n8483 = n8447 & n8477;
  assign n8484 = n8482 & n8483;
  assign n8485 = n8398 & n8421;
  assign n8486 = n8447 & ~n8477;
  assign n8487 = n8485 & n8486;
  assign n8488 = ~n8484 & ~n8487;
  assign n8489 = n8481 & ~n8488;
  assign n8490 = ~n8480 & ~n8489;
  assign n8491 = ~n8358 & n8388;
  assign n8492 = n8422 & n8486;
  assign n8493 = ~n8487 & ~n8492;
  assign n8494 = n8491 & ~n8493;
  assign n8495 = n8483 & n8485;
  assign n8496 = ~n8358 & n8495;
  assign n8497 = n8422 & n8483;
  assign n8498 = n8491 & n8497;
  assign n8499 = ~n8496 & ~n8498;
  assign n8500 = n8398 & ~n8421;
  assign n8501 = n8483 & n8500;
  assign n8502 = ~n8497 & ~n8501;
  assign n8503 = n8481 & ~n8502;
  assign n8504 = ~n8447 & n8477;
  assign n8505 = n8485 & n8504;
  assign n8506 = n8389 & n8505;
  assign n8507 = n8422 & n8504;
  assign n8508 = n8491 & n8507;
  assign n8509 = n8478 & n8500;
  assign n8510 = n8481 & n8509;
  assign n8511 = ~n8508 & ~n8510;
  assign n8512 = ~n8358 & ~n8388;
  assign n8513 = n8486 & n8500;
  assign n8514 = ~n8492 & ~n8513;
  assign n8515 = n8512 & ~n8514;
  assign n8516 = ~n8447 & n8482;
  assign n8517 = ~n8479 & ~n8516;
  assign n8518 = ~n8491 & n8517;
  assign n8519 = ~n8477 & n8516;
  assign n8520 = ~n8505 & ~n8519;
  assign n8521 = ~n8509 & n8520;
  assign n8522 = n8491 & ~n8521;
  assign n8523 = ~n8481 & ~n8522;
  assign n8524 = ~n8518 & ~n8523;
  assign n8525 = n8477 & n8516;
  assign n8526 = n8478 & n8485;
  assign n8527 = ~n8525 & ~n8526;
  assign n8528 = n8482 & n8486;
  assign n8529 = n8500 & n8504;
  assign n8530 = ~n8501 & ~n8513;
  assign n8531 = ~n8529 & n8530;
  assign n8532 = ~n8528 & n8531;
  assign n8533 = n8527 & n8532;
  assign n8534 = n8388 ^ n8358;
  assign n8535 = ~n8533 & ~n8534;
  assign n8536 = ~n8524 & ~n8535;
  assign n8537 = ~n8515 & n8536;
  assign n8538 = n8511 & n8537;
  assign n8539 = ~n8506 & n8538;
  assign n8540 = ~n8503 & n8539;
  assign n8541 = n8499 & n8540;
  assign n8542 = ~n8494 & n8541;
  assign n8543 = n8490 & n8542;
  assign n8544 = n8543 ^ n5627;
  assign n8545 = n8544 ^ x420;
  assign n8546 = ~n8036 & n8545;
  assign n8548 = n8547 ^ n8546;
  assign n8549 = ~n8331 & ~n8548;
  assign n8550 = n7750 & ~n8549;
  assign n8551 = n7393 & n7749;
  assign n8552 = ~n8191 & ~n8329;
  assign n8553 = n8036 & n8545;
  assign n8554 = ~n8552 & n8553;
  assign n8555 = n8191 & n8329;
  assign n8556 = ~n8545 & n8555;
  assign n8557 = ~n8554 & ~n8556;
  assign n8558 = ~n8036 & n8552;
  assign n8559 = ~n8036 & ~n8545;
  assign n8560 = ~n8329 & n8559;
  assign n8561 = ~n8558 & ~n8560;
  assign n8562 = n8557 & n8561;
  assign n8563 = n8551 & ~n8562;
  assign n8564 = ~n8550 & ~n8563;
  assign n8565 = n7393 & ~n7749;
  assign n8566 = n8329 & n8559;
  assign n8567 = n8329 ^ n8191;
  assign n8568 = n8545 & ~n8567;
  assign n8569 = ~n8566 & ~n8568;
  assign n8570 = ~n8545 & n8552;
  assign n8571 = n8570 ^ n8545;
  assign n8572 = n8571 ^ n8329;
  assign n8573 = n8036 & ~n8572;
  assign n8574 = n8569 & ~n8573;
  assign n8575 = n8565 & n8574;
  assign n8576 = ~n7393 & ~n7749;
  assign n8577 = n8329 & ~n8545;
  assign n8578 = n8036 & n8577;
  assign n8579 = ~n8553 & ~n8559;
  assign n8580 = ~n8191 & n8579;
  assign n8581 = ~n8578 & ~n8580;
  assign n8582 = n8545 & n8547;
  assign n8583 = n8330 & ~n8579;
  assign n8584 = ~n8582 & ~n8583;
  assign n8585 = n8581 & n8584;
  assign n8586 = n8576 & n8585;
  assign n8587 = ~n8575 & ~n8586;
  assign n8588 = n8564 & n8587;
  assign n8589 = n8588 ^ n8094;
  assign n8590 = n8589 ^ x462;
  assign n8591 = n8136 & n8145;
  assign n8592 = n8129 & n8173;
  assign n8593 = n8127 & n8148;
  assign n8594 = n8156 & n8157;
  assign n8595 = ~n8593 & ~n8594;
  assign n8596 = ~n8592 & n8595;
  assign n8597 = n8129 & n8167;
  assign n8598 = n8125 & n8143;
  assign n8599 = ~n8158 & ~n8598;
  assign n8600 = n8129 & ~n8599;
  assign n8601 = ~n8132 & ~n8159;
  assign n8602 = n8062 & ~n8601;
  assign n8603 = ~n8600 & ~n8602;
  assign n8604 = ~n8597 & n8603;
  assign n8605 = n8062 & n8172;
  assign n8606 = n8134 & ~n8605;
  assign n8607 = n8125 ^ n8095;
  assign n8608 = n8142 & n8607;
  assign n8609 = ~n8139 & ~n8608;
  assign n8610 = n8156 & ~n8609;
  assign n8611 = ~n8127 & ~n8159;
  assign n8612 = ~n8152 & n8611;
  assign n8613 = n8129 & ~n8612;
  assign n8614 = ~n8610 & ~n8613;
  assign n8615 = n8145 & ~n8180;
  assign n8616 = ~n8152 & ~n8175;
  assign n8617 = n8168 & n8616;
  assign n8618 = n8062 & ~n8617;
  assign n8619 = ~n8151 & n8174;
  assign n8620 = n8148 & ~n8619;
  assign n8621 = ~n8618 & ~n8620;
  assign n8622 = ~n8615 & n8621;
  assign n8623 = n8614 & n8622;
  assign n8624 = n8606 & n8623;
  assign n8625 = n8604 & n8624;
  assign n8626 = n8596 & n8625;
  assign n8627 = ~n8591 & n8626;
  assign n8628 = n8627 ^ n7236;
  assign n8629 = n8628 ^ x436;
  assign n8630 = n8397 ^ x382;
  assign n8631 = n6533 ^ x387;
  assign n8632 = ~n8630 & ~n8631;
  assign n8633 = n8357 ^ x383;
  assign n8634 = n7911 & n7929;
  assign n8635 = n7904 & n7935;
  assign n8636 = ~n8634 & ~n8635;
  assign n8637 = n7906 & ~n7957;
  assign n8638 = n7922 & n7942;
  assign n8639 = n7914 & n7916;
  assign n8640 = n7906 & ~n7940;
  assign n8641 = ~n8639 & ~n8640;
  assign n8642 = n7905 ^ n7904;
  assign n8643 = ~n7909 & n8212;
  assign n8644 = n8643 ^ n7943;
  assign n8645 = ~n8642 & ~n8644;
  assign n8646 = n8645 ^ n7943;
  assign n8647 = n8641 & ~n8646;
  assign n8648 = n7911 & ~n8198;
  assign n8649 = ~n7926 & ~n7932;
  assign n8650 = ~n7903 & n8649;
  assign n8651 = n7916 & ~n8650;
  assign n8652 = ~n8196 & ~n8651;
  assign n8653 = ~n7946 & n8652;
  assign n8654 = n7904 & ~n8653;
  assign n8655 = ~n8648 & ~n8654;
  assign n8656 = n8647 & n8655;
  assign n8657 = ~n7925 & n8656;
  assign n8658 = ~n8638 & n8657;
  assign n8659 = ~n8637 & n8658;
  assign n8660 = n8636 & n8659;
  assign n8661 = n7921 & n8660;
  assign n8662 = n8661 ^ n6367;
  assign n8663 = n8662 ^ x385;
  assign n8664 = ~n8633 & n8663;
  assign n8665 = n7153 ^ x386;
  assign n8666 = n7440 & ~n7481;
  assign n8667 = n7459 & ~n7803;
  assign n8668 = n7480 & ~n8667;
  assign n8669 = ~n8666 & ~n8668;
  assign n8670 = n7394 & n7464;
  assign n8671 = ~n7476 & ~n7789;
  assign n8672 = n7444 & ~n8671;
  assign n8678 = ~n7435 & ~n7438;
  assign n8679 = ~n7440 & n8678;
  assign n8680 = ~n7458 & ~n7803;
  assign n8681 = ~n7452 & n8680;
  assign n8682 = ~n7480 & n8681;
  assign n8683 = ~n8679 & ~n8682;
  assign n8684 = ~n7789 & ~n8683;
  assign n8673 = ~n7396 & n7811;
  assign n8674 = n7467 & ~n7473;
  assign n8675 = ~n7444 & n8674;
  assign n8676 = ~n8673 & ~n8675;
  assign n8677 = ~n7452 & ~n8676;
  assign n8685 = n8684 ^ n8677;
  assign n8686 = n7395 & n8685;
  assign n8687 = n8686 ^ n8684;
  assign n8688 = ~n7798 & n8687;
  assign n8689 = ~n8672 & n8688;
  assign n8690 = ~n8670 & n8689;
  assign n8691 = n8669 & n8690;
  assign n8692 = n7797 & n8691;
  assign n8693 = n7450 & n8692;
  assign n8694 = ~n7436 & n8693;
  assign n8695 = n8694 ^ n6340;
  assign n8696 = n8695 ^ x384;
  assign n8697 = n8665 & ~n8696;
  assign n8698 = n8664 & n8697;
  assign n8699 = ~n8633 & ~n8663;
  assign n8700 = ~n8665 & ~n8696;
  assign n8701 = n8699 & n8700;
  assign n8702 = ~n8698 & ~n8701;
  assign n8703 = n8632 & ~n8702;
  assign n8704 = n8630 & n8631;
  assign n8705 = ~n8665 & n8696;
  assign n8706 = n8699 & n8705;
  assign n8707 = n8633 & n8663;
  assign n8708 = n8700 & n8707;
  assign n8709 = n8633 & ~n8663;
  assign n8710 = n8697 & n8709;
  assign n8711 = ~n8708 & ~n8710;
  assign n8712 = ~n8706 & n8711;
  assign n8713 = n8704 & ~n8712;
  assign n8714 = n8631 ^ n8630;
  assign n8715 = n8664 & n8705;
  assign n8716 = n8714 & n8715;
  assign n8717 = ~n8630 & n8631;
  assign n8718 = n8665 & n8696;
  assign n8719 = n8699 & n8718;
  assign n8720 = ~n8698 & ~n8719;
  assign n8721 = n8717 & ~n8720;
  assign n8722 = ~n8716 & ~n8721;
  assign n8723 = n8664 & n8718;
  assign n8724 = n8704 & n8723;
  assign n8725 = n8630 & ~n8631;
  assign n8726 = n8705 & n8709;
  assign n8727 = n8725 & n8726;
  assign n8728 = ~n8724 & ~n8727;
  assign n8729 = n8664 & n8700;
  assign n8730 = n8704 & n8729;
  assign n8731 = n8701 & n8714;
  assign n8732 = n8700 & n8709;
  assign n8733 = ~n8706 & ~n8732;
  assign n8734 = n8632 & ~n8733;
  assign n8735 = ~n8731 & ~n8734;
  assign n8736 = ~n8730 & n8735;
  assign n8737 = n8697 & n8699;
  assign n8738 = n8632 & n8737;
  assign n8739 = ~n8719 & ~n8737;
  assign n8740 = n8705 & n8707;
  assign n8741 = n8697 & n8707;
  assign n8742 = ~n8740 & ~n8741;
  assign n8743 = n8739 & n8742;
  assign n8744 = ~n8698 & n8743;
  assign n8745 = n8725 & ~n8744;
  assign n8746 = n8707 & n8718;
  assign n8747 = n8709 & n8718;
  assign n8748 = ~n8746 & ~n8747;
  assign n8749 = ~n8708 & n8748;
  assign n8750 = n8632 & ~n8749;
  assign n8751 = ~n8732 & ~n8747;
  assign n8752 = ~n8741 & n8751;
  assign n8753 = n8704 & ~n8752;
  assign n8754 = n8711 & ~n8740;
  assign n8755 = ~n8726 & n8754;
  assign n8756 = n8717 & ~n8755;
  assign n8757 = ~n8753 & ~n8756;
  assign n8758 = ~n8750 & n8757;
  assign n8759 = ~n8745 & n8758;
  assign n8760 = ~n8738 & n8759;
  assign n8761 = n8736 & n8760;
  assign n8762 = n8728 & n8761;
  assign n8763 = n8722 & n8762;
  assign n8764 = ~n8713 & n8763;
  assign n8765 = ~n8703 & n8764;
  assign n8766 = n8765 ^ n6622;
  assign n8767 = n8766 ^ x441;
  assign n8768 = ~n8629 & ~n8767;
  assign n8769 = n7984 & n7986;
  assign n8770 = n7996 & ~n8769;
  assign n8771 = ~n7851 & n7980;
  assign n8772 = n8005 & ~n8014;
  assign n8773 = ~n8771 & ~n8772;
  assign n8774 = ~n7978 & ~n8011;
  assign n8775 = ~n7972 & ~n8774;
  assign n8776 = n7983 & n7992;
  assign n8777 = ~n8775 & ~n8776;
  assign n8778 = ~n7850 & ~n7991;
  assign n8779 = ~n8006 & n8778;
  assign n8780 = n7984 & ~n8779;
  assign n8781 = ~n7989 & n8024;
  assign n8782 = n7980 & ~n8781;
  assign n8783 = ~n8780 & ~n8782;
  assign n8784 = n7972 & ~n8003;
  assign n8785 = ~n8016 & n8022;
  assign n8786 = ~n8014 & ~n8785;
  assign n8787 = ~n8784 & ~n8786;
  assign n8788 = n8783 & n8787;
  assign n8789 = n8777 & n8788;
  assign n8790 = n8773 & n8789;
  assign n8791 = n8770 & n8790;
  assign n8792 = ~n7974 & n8791;
  assign n8793 = n8792 ^ n6586;
  assign n8794 = n8793 ^ x440;
  assign n8795 = n8268 & n8299;
  assign n8796 = n8194 & n8795;
  assign n8797 = n8282 & n8795;
  assign n8798 = ~n8294 & ~n8302;
  assign n8799 = n8287 & ~n8798;
  assign n8800 = ~n8797 & ~n8799;
  assign n8801 = ~n8796 & n8800;
  assign n8802 = n8193 ^ n8192;
  assign n8803 = n8260 & ~n8802;
  assign n8804 = ~n8261 & n8803;
  assign n8805 = n8273 & n8804;
  assign n8806 = ~n8275 & ~n8308;
  assign n8807 = n8287 & ~n8806;
  assign n8808 = n8194 & n8284;
  assign n8809 = ~n8280 & ~n8300;
  assign n8810 = n8287 & ~n8809;
  assign n8811 = ~n8808 & ~n8810;
  assign n8812 = n8278 & n8282;
  assign n8813 = n8265 & n8308;
  assign n8814 = ~n8812 & ~n8813;
  assign n8815 = n8193 & n8263;
  assign n8816 = ~n8283 & ~n8292;
  assign n8817 = ~n8301 & n8816;
  assign n8818 = n8194 & ~n8817;
  assign n8819 = ~n8815 & ~n8818;
  assign n8820 = ~n8270 & n8287;
  assign n8821 = ~n8294 & n8309;
  assign n8822 = n8265 & ~n8821;
  assign n8823 = n8313 & n8809;
  assign n8824 = n8282 & ~n8823;
  assign n8825 = ~n8822 & ~n8824;
  assign n8826 = ~n8820 & n8825;
  assign n8827 = n8819 & n8826;
  assign n8828 = n8814 & n8827;
  assign n8829 = n8811 & n8828;
  assign n8830 = ~n8279 & n8829;
  assign n8831 = ~n8807 & n8830;
  assign n8832 = ~n8805 & n8831;
  assign n8833 = n8801 & n8832;
  assign n8834 = n8272 & n8833;
  assign n8835 = n8834 ^ n7431;
  assign n8836 = n8835 ^ x439;
  assign n8837 = n8794 & ~n8836;
  assign n8838 = n8080 ^ x370;
  assign n8839 = n8446 ^ x375;
  assign n8840 = n8838 & n8839;
  assign n8841 = n8059 ^ x371;
  assign n8842 = n8387 ^ x374;
  assign n8843 = ~n6563 & n6753;
  assign n8844 = n6655 & n6726;
  assign n8845 = n8844 ^ n6716;
  assign n8846 = ~n6753 & ~n8845;
  assign n8847 = ~n6710 & n8846;
  assign n8848 = n6712 & ~n8847;
  assign n8849 = ~n8843 & ~n8848;
  assign n8850 = n6715 & n6722;
  assign n8851 = ~n6727 & ~n6759;
  assign n8852 = n6733 & ~n8851;
  assign n8853 = n6733 & ~n7501;
  assign n8854 = ~n6735 & n6762;
  assign n8855 = ~n6710 & n8854;
  assign n8856 = n6722 & ~n8855;
  assign n8857 = ~n6740 & ~n8845;
  assign n8858 = n6588 & ~n8857;
  assign n8859 = ~n8856 & ~n8858;
  assign n8860 = ~n8853 & n8859;
  assign n8861 = n6739 & n8860;
  assign n8862 = ~n8852 & n8861;
  assign n8863 = ~n8850 & n8862;
  assign n8864 = n8849 & n8863;
  assign n8865 = ~n6711 & n8864;
  assign n8866 = n8334 & n8865;
  assign n8867 = n6743 & n8866;
  assign n8868 = n8867 ^ n6234;
  assign n8869 = n8868 ^ x373;
  assign n8904 = ~n8842 & n8869;
  assign n8871 = n6470 & ~n6481;
  assign n8872 = n6483 & ~n6519;
  assign n8873 = ~n8871 & ~n8872;
  assign n8874 = ~n6507 & ~n6516;
  assign n8875 = n6475 & ~n8874;
  assign n8876 = ~n6436 & n6493;
  assign n8877 = ~n6507 & ~n8876;
  assign n8878 = ~n6483 & n8877;
  assign n8879 = n6434 ^ n6309;
  assign n8880 = n8879 ^ n6466;
  assign n8881 = ~n6436 & ~n8880;
  assign n8882 = n6483 & n8881;
  assign n8883 = ~n6470 & ~n8882;
  assign n8884 = ~n8878 & ~n8883;
  assign n8885 = ~n8875 & ~n8884;
  assign n8886 = ~n6203 & n6492;
  assign n8887 = ~n6488 & ~n6494;
  assign n8888 = ~n6468 & n8887;
  assign n8889 = ~n6204 & n8888;
  assign n8890 = ~n6509 & n7576;
  assign n8891 = ~n6475 & n8890;
  assign n8892 = ~n8889 & ~n8891;
  assign n8893 = ~n6480 & ~n8892;
  assign n8894 = ~n7575 & ~n8893;
  assign n8895 = ~n8886 & ~n8894;
  assign n8896 = n8885 & n8895;
  assign n8897 = n8873 & n8896;
  assign n8898 = n7573 & n8897;
  assign n8899 = n7826 & n8898;
  assign n8900 = n6474 & n8899;
  assign n8901 = n8900 ^ n6253;
  assign n8902 = n8901 ^ x372;
  assign n8870 = n8869 ^ n8842;
  assign n8903 = n8902 ^ n8870;
  assign n8905 = n8904 ^ n8903;
  assign n8906 = ~n8841 & n8905;
  assign n8907 = n8906 ^ n8870;
  assign n8908 = n8840 & ~n8907;
  assign n8909 = ~n8838 & ~n8839;
  assign n8910 = n8842 & ~n8869;
  assign n8911 = n8902 & n8910;
  assign n8912 = ~n8841 & ~n8902;
  assign n8913 = ~n8869 & n8912;
  assign n8914 = ~n8911 & ~n8913;
  assign n8915 = ~n8841 & n8902;
  assign n8916 = n8904 & n8915;
  assign n8917 = n8841 & ~n8910;
  assign n8918 = ~n8902 & n8917;
  assign n8919 = ~n8916 & ~n8918;
  assign n8920 = n8914 & n8919;
  assign n8921 = n8909 & ~n8920;
  assign n8922 = ~n8908 & ~n8921;
  assign n8923 = n8838 & ~n8839;
  assign n8924 = n8841 & n8902;
  assign n8925 = ~n8842 & ~n8869;
  assign n8926 = n8924 & n8925;
  assign n8927 = n8842 & n8915;
  assign n8928 = n8842 & n8869;
  assign n8929 = n8902 & n8928;
  assign n8930 = ~n8927 & ~n8929;
  assign n8931 = ~n8926 & n8930;
  assign n8932 = n8910 ^ n8841;
  assign n8933 = n8931 & ~n8932;
  assign n8934 = ~n8902 & n8933;
  assign n8935 = n8934 ^ n8931;
  assign n8936 = n8923 & ~n8935;
  assign n8937 = ~n8838 & n8839;
  assign n8938 = n8869 & n8924;
  assign n8939 = ~n8841 & n8925;
  assign n8940 = ~n8938 & ~n8939;
  assign n8941 = n8841 & n8928;
  assign n8942 = ~n8912 & ~n8924;
  assign n8943 = n8842 & ~n8942;
  assign n8944 = ~n8941 & ~n8943;
  assign n8945 = n8940 & n8944;
  assign n8946 = n8937 & n8945;
  assign n8947 = ~n8936 & ~n8946;
  assign n8948 = n8922 & n8947;
  assign n8949 = n8948 ^ n7405;
  assign n8950 = n8949 ^ x438;
  assign n8951 = n8481 & n8507;
  assign n8952 = n8389 & ~n8488;
  assign n8953 = ~n8951 & ~n8952;
  assign n8954 = ~n8495 & ~n8528;
  assign n8955 = n8491 & ~n8954;
  assign n8956 = n8484 & n8491;
  assign n8957 = ~n8388 & ~n8514;
  assign n8958 = ~n8956 & ~n8957;
  assign n8959 = n8487 & n8512;
  assign n8960 = n8481 & ~n8520;
  assign n8961 = ~n8959 & ~n8960;
  assign n8962 = n8502 & ~n8526;
  assign n8963 = n8520 & n8962;
  assign n8964 = n8389 & ~n8963;
  assign n8965 = ~n8491 & ~n8529;
  assign n8966 = ~n8516 & n8965;
  assign n8967 = ~n8479 & ~n8501;
  assign n8968 = ~n8512 & n8967;
  assign n8969 = ~n8966 & ~n8968;
  assign n8970 = ~n8509 & ~n8969;
  assign n8971 = ~n8497 & n8970;
  assign n8972 = ~n8358 & ~n8971;
  assign n8973 = ~n8964 & ~n8972;
  assign n8974 = n8961 & n8973;
  assign n8975 = n8958 & n8974;
  assign n8976 = ~n8955 & n8975;
  assign n8977 = n8490 & n8976;
  assign n8978 = n8953 & n8977;
  assign n8979 = n8511 & n8978;
  assign n8980 = n8979 ^ n7183;
  assign n8981 = n8980 ^ x437;
  assign n8982 = n8950 & n8981;
  assign n8983 = n8837 & n8982;
  assign n8984 = n8768 & n8983;
  assign n8985 = ~n8629 & n8767;
  assign n8986 = ~n8794 & n8836;
  assign n8987 = ~n8950 & ~n8981;
  assign n8988 = n8986 & n8987;
  assign n8989 = n8985 & n8988;
  assign n8990 = n8629 & n8767;
  assign n8991 = n8950 & ~n8981;
  assign n8992 = n8986 & n8991;
  assign n8993 = n8837 & n8987;
  assign n8994 = ~n8992 & ~n8993;
  assign n8995 = n8990 & ~n8994;
  assign n8996 = ~n8989 & ~n8995;
  assign n8997 = ~n8984 & n8996;
  assign n8998 = n8982 & n8986;
  assign n8999 = n8990 & n8998;
  assign n9000 = ~n8794 & ~n8836;
  assign n9001 = n8990 & n8991;
  assign n9002 = n9000 & n9001;
  assign n9003 = ~n8999 & ~n9002;
  assign n9004 = n8982 & n9000;
  assign n9005 = ~n8950 & n8981;
  assign n9006 = n8837 & n9005;
  assign n9007 = ~n9004 & ~n9006;
  assign n9008 = n8985 & ~n9007;
  assign n9009 = n9003 & ~n9008;
  assign n9010 = n8629 & ~n8767;
  assign n9011 = ~n8985 & ~n9010;
  assign n9012 = n9000 & n9005;
  assign n9013 = n9011 & n9012;
  assign n9014 = ~n8629 & ~n8994;
  assign n9015 = ~n9013 & ~n9014;
  assign n9016 = n8794 & n8991;
  assign n9017 = ~n8998 & ~n9016;
  assign n9018 = n8985 & ~n9017;
  assign n9019 = n8986 & n9005;
  assign n9020 = n8794 & n8836;
  assign n9021 = n8982 & n9020;
  assign n9022 = ~n9019 & ~n9021;
  assign n9023 = n8837 & n8991;
  assign n9024 = ~n8988 & ~n9023;
  assign n9025 = n9022 & n9024;
  assign n9026 = n8768 & ~n9025;
  assign n9027 = ~n9018 & ~n9026;
  assign n9028 = n9015 & n9027;
  assign n9029 = n8987 & n9020;
  assign n9030 = ~n8983 & ~n9019;
  assign n9031 = ~n9029 & n9030;
  assign n9032 = n8990 & ~n9031;
  assign n9033 = n8991 & n9020;
  assign n9034 = n8991 & n9000;
  assign n9035 = ~n8993 & ~n9034;
  assign n9036 = ~n9033 & n9035;
  assign n9037 = ~n8992 & ~n9029;
  assign n9038 = ~n8983 & n9037;
  assign n9039 = ~n9006 & n9038;
  assign n9040 = n9036 & n9039;
  assign n9041 = ~n9019 & n9040;
  assign n9042 = n9010 & n9041;
  assign n9043 = ~n9032 & ~n9042;
  assign n9044 = n9028 & n9043;
  assign n9045 = n9009 & n9044;
  assign n9046 = n8997 & n9045;
  assign n9047 = n9046 ^ n8080;
  assign n9048 = n9047 ^ x464;
  assign n9049 = n8590 & ~n9048;
  assign n9050 = n8840 & ~n8935;
  assign n9051 = ~n8920 & n8937;
  assign n9052 = ~n9050 & ~n9051;
  assign n9053 = n8907 & n8923;
  assign n9054 = n8909 & ~n8945;
  assign n9055 = ~n9053 & ~n9054;
  assign n9056 = n9052 & n9055;
  assign n9057 = n9056 ^ n6308;
  assign n9058 = n9057 ^ x430;
  assign n9059 = n8980 ^ x435;
  assign n9060 = n9058 & n9059;
  assign n9061 = n8628 ^ x434;
  assign n9062 = ~n7358 & n7369;
  assign n9063 = n7330 & ~n9062;
  assign n9064 = n7348 & ~n7361;
  assign n9065 = ~n7334 & n9064;
  assign n9066 = n7364 & ~n9065;
  assign n9067 = ~n9063 & ~n9066;
  assign n9068 = n7333 & n7344;
  assign n9069 = ~n7337 & ~n9068;
  assign n9070 = ~n7352 & ~n7353;
  assign n9071 = n9069 & n9070;
  assign n9072 = n7351 & ~n9071;
  assign n9073 = n7364 & ~n7379;
  assign n9074 = n7360 & ~n9073;
  assign n9075 = n6535 & n7336;
  assign n9076 = n7351 & n9075;
  assign n9077 = ~n7351 & ~n7364;
  assign n9078 = ~n7373 & ~n9077;
  assign n9079 = ~n9076 & ~n9078;
  assign n9080 = ~n7361 & ~n9068;
  assign n9081 = n9070 & n9080;
  assign n9082 = n7330 & ~n9081;
  assign n9083 = ~n7351 & ~n7361;
  assign n9084 = ~n7345 & n9083;
  assign n9085 = ~n7372 & n9084;
  assign n9086 = ~n7367 & n9085;
  assign n9087 = ~n7353 & n9086;
  assign n9088 = n7332 & ~n9087;
  assign n9089 = ~n9082 & ~n9088;
  assign n9090 = n9079 & n9089;
  assign n9091 = n9074 & n9090;
  assign n9092 = ~n9072 & n9091;
  assign n9093 = n9067 & n9092;
  assign n9094 = n7340 & n9093;
  assign n9095 = n9094 ^ n7214;
  assign n9096 = n9095 ^ x432;
  assign n9097 = ~n9061 & ~n9096;
  assign n9098 = n7676 & n7712;
  assign n9099 = n7524 & n7694;
  assign n9100 = ~n9098 & ~n9099;
  assign n9101 = ~n7674 & ~n7724;
  assign n9102 = n7696 & ~n9101;
  assign n9103 = ~n7717 & ~n9102;
  assign n9104 = n7638 & n7693;
  assign n9105 = n7696 & n9104;
  assign n9106 = n7676 & n7689;
  assign n9107 = ~n9105 & ~n9106;
  assign n9108 = ~n7679 & n7713;
  assign n9109 = n7696 & ~n9108;
  assign n9110 = ~n7730 & ~n7733;
  assign n9111 = n7722 & n9101;
  assign n9112 = n9110 & n9111;
  assign n9113 = n7692 & ~n9112;
  assign n9114 = ~n9109 & ~n9113;
  assign n9115 = n7676 & ~n9110;
  assign n9116 = n7699 & ~n7703;
  assign n9117 = ~n7709 & n9116;
  assign n9118 = ~n7733 & n9117;
  assign n9119 = n7524 & ~n9118;
  assign n9120 = ~n9115 & ~n9119;
  assign n9121 = n9114 & n9120;
  assign n9122 = n7716 & n9121;
  assign n9123 = n9107 & n9122;
  assign n9124 = n9103 & n9123;
  assign n9125 = n9100 & n9124;
  assign n9126 = n7681 & n9125;
  assign n9127 = n9126 ^ n7263;
  assign n9128 = n9127 ^ x433;
  assign n9129 = n8287 & n8292;
  assign n9130 = n8265 & n8280;
  assign n9131 = ~n9129 & ~n9130;
  assign n9132 = n8265 & n8288;
  assign n9133 = ~n8278 & ~n8795;
  assign n9134 = n8287 & ~n9133;
  assign n9135 = ~n9132 & ~n9134;
  assign n9136 = n8193 & n8283;
  assign n9137 = ~n8275 & ~n8300;
  assign n9138 = n8194 & ~n9137;
  assign n9139 = n8308 & ~n8802;
  assign n9140 = ~n8287 & n8301;
  assign n9141 = ~n9139 & ~n9140;
  assign n9142 = n8284 & n8287;
  assign n9143 = n8282 & ~n8310;
  assign n9144 = ~n9142 & ~n9143;
  assign n9145 = n9141 & n9144;
  assign n9146 = ~n9138 & n9145;
  assign n9147 = ~n9136 & n9146;
  assign n9148 = n9135 & n9147;
  assign n9149 = ~n8812 & n9148;
  assign n9150 = n8800 & n9149;
  assign n9151 = n9131 & n9150;
  assign n9152 = n8811 & n9151;
  assign n9153 = ~n8281 & n9152;
  assign n9154 = ~n8279 & n9153;
  assign n9155 = ~n8276 & n9154;
  assign n9156 = n8272 & n9155;
  assign n9157 = n9156 ^ n6202;
  assign n9158 = n9157 ^ x431;
  assign n9159 = n9128 & ~n9158;
  assign n9160 = n9097 & n9159;
  assign n9161 = n9061 & ~n9096;
  assign n9162 = ~n9128 & ~n9158;
  assign n9163 = n9161 & n9162;
  assign n9164 = ~n9160 & ~n9163;
  assign n9165 = n9060 & ~n9164;
  assign n9166 = ~n9058 & n9059;
  assign n9167 = ~n9061 & n9096;
  assign n9168 = n9162 & n9167;
  assign n9169 = ~n9163 & ~n9168;
  assign n9170 = n9166 & ~n9169;
  assign n9171 = ~n9128 & n9158;
  assign n9172 = n9097 & n9171;
  assign n9173 = n9128 & n9158;
  assign n9174 = n9161 & n9173;
  assign n9175 = ~n9172 & ~n9174;
  assign n9176 = n9060 & ~n9175;
  assign n9177 = n9058 & ~n9059;
  assign n9178 = n9061 & n9096;
  assign n9179 = n9159 & n9178;
  assign n9180 = ~n9160 & ~n9179;
  assign n9181 = n9177 & ~n9180;
  assign n9182 = ~n9176 & ~n9181;
  assign n9183 = ~n9170 & n9182;
  assign n9184 = n9173 & n9178;
  assign n9185 = ~n9059 & n9184;
  assign n9186 = n9161 & n9171;
  assign n9187 = n9060 & n9186;
  assign n9188 = ~n9185 & ~n9187;
  assign n9189 = ~n9058 & ~n9059;
  assign n9190 = n9171 & n9178;
  assign n9191 = n9097 & n9173;
  assign n9192 = ~n9190 & ~n9191;
  assign n9193 = n9189 & ~n9192;
  assign n9194 = ~n9166 & ~n9177;
  assign n9195 = n9167 & n9173;
  assign n9196 = ~n9172 & ~n9195;
  assign n9197 = ~n9174 & n9196;
  assign n9198 = ~n9194 & ~n9197;
  assign n9199 = ~n9193 & ~n9198;
  assign n9200 = n9188 & n9199;
  assign n9201 = ~n9169 & n9177;
  assign n9202 = n9159 & n9161;
  assign n9203 = n9097 & n9162;
  assign n9204 = ~n9202 & ~n9203;
  assign n9205 = ~n9190 & n9204;
  assign n9206 = n9166 & ~n9205;
  assign n9207 = ~n9201 & ~n9206;
  assign n9208 = n9167 & n9171;
  assign n9209 = n9159 & n9167;
  assign n9210 = ~n9179 & ~n9209;
  assign n9211 = ~n9189 & n9210;
  assign n9212 = ~n9160 & ~n9202;
  assign n9213 = n9060 & n9179;
  assign n9214 = n9162 & n9178;
  assign n9215 = ~n9209 & ~n9214;
  assign n9216 = ~n9213 & n9215;
  assign n9217 = n9212 & n9216;
  assign n9218 = ~n9211 & ~n9217;
  assign n9219 = n9194 & ~n9218;
  assign n9220 = ~n9208 & n9219;
  assign n9221 = n9220 ^ n9194;
  assign n9222 = n9207 & ~n9221;
  assign n9223 = n9200 & n9222;
  assign n9224 = n9183 & n9223;
  assign n9225 = ~n9165 & n9224;
  assign n9226 = n9225 ^ n8124;
  assign n9227 = n9226 ^ x463;
  assign n9228 = ~n7368 & ~n7372;
  assign n9229 = n7351 & ~n9228;
  assign n9230 = n7362 & ~n7365;
  assign n9231 = ~n9229 & ~n9230;
  assign n9232 = n7334 & n7351;
  assign n9233 = ~n7342 & ~n9075;
  assign n9234 = ~n9077 & ~n9233;
  assign n9235 = ~n9232 & ~n9234;
  assign n9236 = ~n7337 & ~n7353;
  assign n9237 = n7364 & ~n9236;
  assign n9238 = ~n7035 & n7348;
  assign n9239 = ~n7365 & ~n9238;
  assign n9240 = ~n9237 & ~n9239;
  assign n9241 = n9235 & n9240;
  assign n9242 = n7332 & ~n7369;
  assign n9243 = n7330 & n7377;
  assign n9244 = ~n9242 & ~n9243;
  assign n9245 = n9241 & n9244;
  assign n9246 = ~n7339 & n9245;
  assign n9247 = ~n7356 & n9246;
  assign n9248 = n9231 & n9247;
  assign n9249 = n9248 ^ n6676;
  assign n9250 = n9249 ^ x400;
  assign n9251 = n8282 & n8301;
  assign n9252 = n8283 & n8287;
  assign n9253 = n8275 & n8282;
  assign n9254 = n8193 & n8267;
  assign n9255 = ~n9253 & ~n9254;
  assign n9256 = n8265 & n8284;
  assign n9257 = n8194 & ~n8313;
  assign n9258 = ~n9256 & ~n9257;
  assign n9259 = n9255 & n9258;
  assign n9260 = ~n8287 & n8300;
  assign n9261 = ~n8263 & ~n8294;
  assign n9262 = ~n8802 & ~n9261;
  assign n9263 = ~n8267 & ~n8795;
  assign n9264 = n8287 & ~n9263;
  assign n9265 = ~n9262 & ~n9264;
  assign n9266 = ~n9260 & n9265;
  assign n9267 = n9259 & n9266;
  assign n9268 = n8814 & n9267;
  assign n9269 = n8291 & n9268;
  assign n9270 = ~n8276 & n9269;
  assign n9271 = ~n9252 & n9270;
  assign n9272 = ~n9251 & n9271;
  assign n9273 = n9131 & n9272;
  assign n9274 = n8801 & n9273;
  assign n9275 = ~n8281 & n9274;
  assign n9276 = n9275 ^ n6810;
  assign n9277 = n9276 ^ x405;
  assign n9278 = ~n9250 & n9277;
  assign n9279 = n7978 & n7984;
  assign n9280 = n7973 & n7983;
  assign n9281 = ~n9279 & ~n9280;
  assign n9282 = n7972 & n8011;
  assign n9283 = ~n8005 & n8022;
  assign n9284 = ~n8011 & n9283;
  assign n9285 = n7980 & ~n9284;
  assign n9286 = ~n9282 & ~n9285;
  assign n9287 = n7971 & n8016;
  assign n9288 = n8018 & ~n8023;
  assign n9289 = ~n7850 & n9288;
  assign n9290 = n7992 & ~n9289;
  assign n9291 = ~n7991 & ~n8021;
  assign n9292 = ~n7847 & n9291;
  assign n9293 = n7984 & ~n9292;
  assign n9294 = n8025 & n8778;
  assign n9295 = n7973 & ~n9294;
  assign n9296 = ~n9293 & ~n9295;
  assign n9297 = ~n9290 & n9296;
  assign n9298 = ~n9287 & n9297;
  assign n9299 = n9286 & n9298;
  assign n9300 = n9281 & n9299;
  assign n9301 = n8773 & n9300;
  assign n9302 = n8770 & n9301;
  assign n9303 = n9302 ^ n7899;
  assign n9304 = n9303 ^ x402;
  assign n9305 = ~n8702 & n8704;
  assign n9306 = ~n8711 & n8725;
  assign n9307 = ~n8723 & ~n8726;
  assign n9308 = n8632 & ~n9307;
  assign n9309 = ~n9306 & ~n9308;
  assign n9310 = ~n9305 & n9309;
  assign n9311 = n8725 & n8729;
  assign n9312 = n8739 & ~n8746;
  assign n9313 = ~n8740 & n9312;
  assign n9314 = n8714 & ~n9313;
  assign n9315 = ~n9311 & ~n9314;
  assign n9316 = n8704 & n8715;
  assign n9317 = ~n8696 & n8709;
  assign n9318 = ~n8706 & ~n9317;
  assign n9319 = ~n8715 & n9318;
  assign n9320 = n8717 & ~n9319;
  assign n9321 = ~n8714 & ~n8751;
  assign n9322 = ~n8708 & ~n8726;
  assign n9323 = n8704 & ~n9322;
  assign n9324 = n8632 & ~n8742;
  assign n9325 = ~n9323 & ~n9324;
  assign n9326 = ~n9321 & n9325;
  assign n9327 = ~n9320 & n9326;
  assign n9328 = ~n9316 & n9327;
  assign n9329 = n9315 & n9328;
  assign n9330 = n8728 & n9329;
  assign n9331 = n9310 & n9330;
  assign n9332 = ~n8703 & n9331;
  assign n9333 = n9332 ^ n6957;
  assign n9334 = n9333 ^ x404;
  assign n9335 = n9304 & n9334;
  assign n9336 = ~n8902 & n8910;
  assign n9337 = n8841 & n9336;
  assign n9338 = n8910 & n8915;
  assign n9339 = n8841 & n8904;
  assign n9340 = n8910 ^ n8902;
  assign n9341 = ~n8932 & ~n9340;
  assign n9342 = ~n9339 & n9341;
  assign n9343 = n9342 ^ n9339;
  assign n9344 = ~n9338 & ~n9343;
  assign n9345 = n8909 & ~n9344;
  assign n9346 = ~n8841 & n8928;
  assign n9347 = n8902 & n8925;
  assign n9348 = ~n8842 & n8942;
  assign n9349 = ~n9347 & ~n9348;
  assign n9350 = ~n9346 & n9349;
  assign n9351 = n8923 & ~n9350;
  assign n9352 = ~n9345 & ~n9351;
  assign n9353 = n8904 & n8924;
  assign n9354 = ~n8870 & ~n8902;
  assign n9355 = ~n8869 & n8942;
  assign n9356 = ~n9354 & ~n9355;
  assign n9357 = ~n9353 & n9356;
  assign n9358 = n8840 & ~n9357;
  assign n9359 = ~n8869 & n8924;
  assign n9360 = n8904 & n8942;
  assign n9361 = ~n9359 & ~n9360;
  assign n9362 = ~n9336 & n9361;
  assign n9363 = ~n8943 & n9362;
  assign n9364 = n8937 & ~n9363;
  assign n9365 = ~n9358 & ~n9364;
  assign n9366 = n9352 & n9365;
  assign n9367 = ~n9337 & n9366;
  assign n9368 = n9367 ^ n6562;
  assign n9369 = n9368 ^ x401;
  assign n9370 = n8389 & n8507;
  assign n9371 = ~n8955 & ~n9370;
  assign n9372 = ~n8492 & ~n8497;
  assign n9373 = ~n8388 & ~n9372;
  assign n9374 = n8491 & ~n8514;
  assign n9375 = ~n9373 & ~n9374;
  assign n9376 = ~n8487 & ~n8528;
  assign n9377 = n8481 & ~n9376;
  assign n9378 = ~n8519 & n8527;
  assign n9379 = n8389 & ~n9378;
  assign n9380 = ~n9377 & ~n9379;
  assign n9381 = ~n8484 & ~n8501;
  assign n9382 = n8512 & ~n9381;
  assign n9383 = ~n8479 & ~n8526;
  assign n9384 = ~n8505 & n9383;
  assign n9385 = ~n8497 & n9384;
  assign n9386 = n8491 & ~n9385;
  assign n9387 = ~n8479 & n8520;
  assign n9388 = n8965 & n9387;
  assign n9389 = n8481 & ~n9388;
  assign n9390 = ~n8509 & n8527;
  assign n9391 = ~n8479 & n9390;
  assign n9392 = n8512 & ~n9391;
  assign n9393 = ~n8495 & n8530;
  assign n9394 = ~n8484 & n9393;
  assign n9395 = n8389 & ~n9394;
  assign n9396 = ~n9392 & ~n9395;
  assign n9397 = ~n9389 & n9396;
  assign n9398 = ~n9386 & n9397;
  assign n9399 = ~n9382 & n9398;
  assign n9400 = n9380 & n9399;
  assign n9401 = n9375 & n9400;
  assign n9402 = n9371 & n9401;
  assign n9403 = n9402 ^ n7871;
  assign n9404 = n9403 ^ x403;
  assign n9405 = n9369 & ~n9404;
  assign n9406 = n9335 & n9405;
  assign n9407 = n9278 & n9406;
  assign n9408 = ~n9369 & n9404;
  assign n9409 = n9335 & n9408;
  assign n9410 = n9278 & n9409;
  assign n9411 = n9250 & ~n9277;
  assign n9412 = ~n9304 & n9334;
  assign n9413 = ~n9369 & ~n9404;
  assign n9414 = n9412 & n9413;
  assign n9415 = n9411 & n9414;
  assign n9416 = ~n9410 & ~n9415;
  assign n9417 = n9405 & n9412;
  assign n9418 = n9278 & n9417;
  assign n9419 = ~n9250 & ~n9277;
  assign n9420 = n9408 & n9412;
  assign n9421 = ~n9304 & ~n9334;
  assign n9422 = n9405 & n9421;
  assign n9423 = n9304 & ~n9334;
  assign n9424 = n9413 & n9423;
  assign n9425 = ~n9414 & ~n9424;
  assign n9426 = ~n9422 & n9425;
  assign n9427 = ~n9420 & n9426;
  assign n9428 = n9419 & ~n9427;
  assign n9429 = n9369 & n9404;
  assign n9430 = n9423 & n9429;
  assign n9431 = n9405 & n9423;
  assign n9432 = n9419 & n9431;
  assign n9433 = n9250 & n9277;
  assign n9434 = n9408 & n9423;
  assign n9435 = ~n9420 & ~n9434;
  assign n9436 = ~n9409 & n9435;
  assign n9437 = ~n9424 & n9436;
  assign n9438 = n9433 & ~n9437;
  assign n9439 = n9421 & n9429;
  assign n9440 = ~n9406 & ~n9422;
  assign n9441 = ~n9439 & n9440;
  assign n9442 = n9433 & ~n9441;
  assign n9443 = n9408 & n9421;
  assign n9444 = n9413 & n9421;
  assign n9445 = n9335 & n9413;
  assign n9446 = ~n9444 & ~n9445;
  assign n9447 = ~n9443 & n9446;
  assign n9448 = ~n9420 & n9447;
  assign n9449 = n9278 & ~n9448;
  assign n9450 = ~n9442 & ~n9449;
  assign n9451 = ~n9438 & n9450;
  assign n9452 = n9335 & n9429;
  assign n9453 = ~n9439 & ~n9452;
  assign n9454 = n9419 & ~n9453;
  assign n9455 = n9412 & n9429;
  assign n9456 = n9446 & ~n9452;
  assign n9457 = ~n9455 & n9456;
  assign n9458 = ~n9431 & n9457;
  assign n9459 = ~n9434 & n9458;
  assign n9460 = n9411 & ~n9459;
  assign n9461 = ~n9454 & ~n9460;
  assign n9462 = n9451 & n9461;
  assign n9463 = ~n9432 & n9462;
  assign n9464 = ~n9430 & n9463;
  assign n9465 = ~n9428 & n9464;
  assign n9466 = ~n9418 & n9465;
  assign n9467 = n9416 & n9466;
  assign n9468 = ~n9407 & n9467;
  assign n9469 = n9468 ^ n7970;
  assign n9470 = n9469 ^ x461;
  assign n9471 = ~n9227 & ~n9470;
  assign n9472 = n9049 & n9471;
  assign n9473 = n8590 & n9048;
  assign n9474 = n9227 & ~n9470;
  assign n9475 = n9473 & n9474;
  assign n9476 = ~n9472 & ~n9475;
  assign n9477 = n9333 ^ x406;
  assign n9478 = n7676 & n7703;
  assign n9479 = n7681 & ~n9478;
  assign n9480 = ~n7687 & ~n7705;
  assign n9481 = ~n7703 & n9480;
  assign n9482 = n7696 & ~n9481;
  assign n9483 = ~n7689 & n9110;
  assign n9484 = n7524 & ~n9483;
  assign n9485 = ~n9482 & ~n9484;
  assign n9486 = ~n7674 & ~n7730;
  assign n9487 = n7676 & ~n9486;
  assign n9488 = n7696 & ~n7710;
  assign n9489 = ~n7694 & n7713;
  assign n9490 = n7524 & ~n9489;
  assign n9491 = ~n7697 & n7727;
  assign n9492 = n7734 & n9491;
  assign n9493 = n7692 & ~n9492;
  assign n9494 = ~n9490 & ~n9493;
  assign n9495 = ~n9488 & n9494;
  assign n9496 = ~n9106 & n9495;
  assign n9497 = n9103 & n9496;
  assign n9498 = ~n7684 & n9497;
  assign n9499 = ~n7698 & n9498;
  assign n9500 = ~n9487 & n9499;
  assign n9501 = n9485 & n9500;
  assign n9502 = n9479 & n9501;
  assign n9503 = n9502 ^ n6930;
  assign n9504 = n9503 ^ x411;
  assign n9505 = n9477 & n9504;
  assign n9506 = n7351 & n7358;
  assign n9507 = n7330 & ~n9069;
  assign n9508 = ~n9506 & ~n9507;
  assign n9515 = ~n7035 & n9083;
  assign n9516 = n7382 & n9080;
  assign n9517 = ~n7334 & n9516;
  assign n9518 = ~n9515 & ~n9517;
  assign n9519 = n9228 & ~n9518;
  assign n9509 = n7364 & ~n9070;
  assign n9510 = n7332 & ~n7354;
  assign n9511 = ~n9509 & ~n9510;
  assign n9512 = ~n7367 & n9511;
  assign n9513 = ~n9075 & n9512;
  assign n9514 = ~n7334 & n9513;
  assign n9520 = n9519 ^ n9514;
  assign n9521 = ~n7365 & n9520;
  assign n9522 = n9521 ^ n9519;
  assign n9523 = n9508 & n9522;
  assign n9524 = n9231 & n9523;
  assign n9525 = n7350 & n9524;
  assign n9526 = n9074 & n9525;
  assign n9527 = n9526 ^ n6907;
  assign n9528 = n9527 ^ x409;
  assign n9529 = n9276 ^ x407;
  assign n9530 = n9528 & ~n9529;
  assign n9531 = n8148 & n8152;
  assign n9532 = n8095 ^ n8082;
  assign n9533 = n8095 ^ n8081;
  assign n9534 = n9533 ^ n8125;
  assign n9535 = ~n9532 & n9534;
  assign n9536 = n8062 & n9535;
  assign n9537 = n8145 & n8157;
  assign n9538 = n8148 & n8175;
  assign n9539 = ~n9537 & ~n9538;
  assign n9540 = n9533 ^ n8082;
  assign n9541 = n8125 ^ n8082;
  assign n9542 = ~n9532 & n9541;
  assign n9543 = ~n9540 & n9542;
  assign n9544 = n9543 ^ n9540;
  assign n9545 = n8156 & ~n9544;
  assign n9546 = ~n8136 & ~n8179;
  assign n9547 = n8616 & n9546;
  assign n9548 = ~n8151 & n9547;
  assign n9549 = n8129 & ~n9548;
  assign n9550 = ~n9545 & ~n9549;
  assign n9551 = n9539 & n9550;
  assign n9552 = ~n9536 & n9551;
  assign n9553 = ~n9531 & n9552;
  assign n9554 = n8606 & n9553;
  assign n9555 = n8603 & n9554;
  assign n9556 = ~n8591 & n9555;
  assign n9557 = n9556 ^ n6839;
  assign n9558 = n9557 ^ x408;
  assign n9559 = n8512 & ~n9387;
  assign n9560 = n8389 & ~n8514;
  assign n9561 = ~n9559 & ~n9560;
  assign n9562 = n8481 & n8529;
  assign n9563 = ~n8388 & n8525;
  assign n9564 = ~n8501 & n8527;
  assign n9565 = n8491 & ~n9564;
  assign n9566 = ~n8529 & n9383;
  assign n9567 = n8389 & ~n9566;
  assign n9568 = ~n9565 & ~n9567;
  assign n9569 = n8502 & ~n8513;
  assign n9570 = ~n8528 & n9569;
  assign n9571 = n8512 & ~n9570;
  assign n9572 = ~n8519 & n9372;
  assign n9573 = ~n8495 & n9572;
  assign n9574 = n8481 & ~n9573;
  assign n9575 = ~n9571 & ~n9574;
  assign n9576 = n9568 & n9575;
  assign n9577 = n9371 & n9576;
  assign n9578 = ~n8494 & n9577;
  assign n9579 = ~n9563 & n9578;
  assign n9580 = ~n9562 & n9579;
  assign n9581 = n9561 & n9580;
  assign n9582 = n8953 & n9581;
  assign n9583 = n8511 & n9582;
  assign n9584 = n9583 ^ n6879;
  assign n9585 = n9584 ^ x410;
  assign n9586 = n9558 & ~n9585;
  assign n9587 = n9530 & n9586;
  assign n9588 = n9505 & n9587;
  assign n9589 = n9477 & ~n9504;
  assign n9590 = ~n9528 & ~n9529;
  assign n9591 = n9558 & n9585;
  assign n9592 = n9590 & n9591;
  assign n9593 = ~n9558 & ~n9585;
  assign n9594 = n9590 & n9593;
  assign n9595 = ~n9592 & ~n9594;
  assign n9596 = n9589 & ~n9595;
  assign n9597 = ~n9588 & ~n9596;
  assign n9598 = ~n9528 & n9529;
  assign n9599 = n9591 & n9598;
  assign n9600 = n9530 & n9591;
  assign n9601 = ~n9599 & ~n9600;
  assign n9602 = n9589 & ~n9601;
  assign n9603 = ~n9477 & ~n9504;
  assign n9604 = n9600 & n9603;
  assign n9605 = n9528 & n9529;
  assign n9606 = ~n9558 & n9585;
  assign n9607 = n9605 & n9606;
  assign n9608 = n9586 & n9605;
  assign n9609 = ~n9607 & ~n9608;
  assign n9610 = n9589 & ~n9609;
  assign n9611 = ~n9604 & ~n9610;
  assign n9612 = n9587 & n9603;
  assign n9613 = ~n9477 & n9504;
  assign n9614 = n9594 & n9613;
  assign n9615 = n9530 & n9606;
  assign n9616 = n9586 & n9590;
  assign n9617 = ~n9615 & ~n9616;
  assign n9618 = n9505 & ~n9617;
  assign n9619 = ~n9614 & ~n9618;
  assign n9620 = ~n9612 & n9619;
  assign n9621 = n9586 & n9598;
  assign n9622 = n9505 & n9621;
  assign n9623 = n9598 & n9606;
  assign n9624 = n9613 & n9623;
  assign n9625 = ~n9622 & ~n9624;
  assign n9626 = n9505 & n9600;
  assign n9627 = n9590 & n9606;
  assign n9628 = n9603 & n9627;
  assign n9629 = ~n9626 & ~n9628;
  assign n9630 = n9530 & n9593;
  assign n9631 = ~n9592 & ~n9630;
  assign n9632 = n9613 & ~n9631;
  assign n9633 = n9599 & n9603;
  assign n9634 = n9603 & n9608;
  assign n9635 = ~n9633 & ~n9634;
  assign n9636 = n9504 ^ n9477;
  assign n9637 = n9623 & ~n9636;
  assign n9638 = n9593 & n9598;
  assign n9639 = ~n9630 & ~n9638;
  assign n9640 = n9589 & ~n9639;
  assign n9641 = ~n9637 & ~n9640;
  assign n9642 = n9593 & n9605;
  assign n9643 = ~n9477 & n9642;
  assign n9644 = ~n9599 & ~n9642;
  assign n9645 = n9505 & ~n9644;
  assign n9646 = ~n9643 & ~n9645;
  assign n9647 = n9641 & n9646;
  assign n9648 = n9603 & n9616;
  assign n9649 = n9591 & n9605;
  assign n9650 = ~n9621 & ~n9649;
  assign n9651 = ~n9615 & n9650;
  assign n9652 = n9613 & ~n9651;
  assign n9653 = ~n9648 & ~n9652;
  assign n9654 = n9647 & n9653;
  assign n9655 = n9635 & n9654;
  assign n9656 = ~n9632 & n9655;
  assign n9657 = n9629 & n9656;
  assign n9658 = n9625 & n9657;
  assign n9659 = n9620 & n9658;
  assign n9660 = n9611 & n9659;
  assign n9661 = ~n9602 & n9660;
  assign n9662 = n9597 & n9661;
  assign n9663 = n9662 ^ n8059;
  assign n9664 = n9663 ^ x465;
  assign n9665 = n8190 ^ x424;
  assign n9666 = n9157 ^ x429;
  assign n9667 = n9665 & n9666;
  assign n9668 = n9057 ^ x428;
  assign n9669 = n7984 & n8000;
  assign n9670 = n7976 & ~n8014;
  assign n9671 = ~n9669 & ~n9670;
  assign n9672 = n8003 & n8017;
  assign n9673 = n7973 & ~n9672;
  assign n9674 = ~n8023 & n9291;
  assign n9675 = n7980 & ~n9674;
  assign n9676 = ~n9673 & ~n9675;
  assign n9677 = n7971 & ~n8012;
  assign n9678 = n7847 & n7984;
  assign n9679 = n8024 & ~n9678;
  assign n9680 = ~n8005 & n9679;
  assign n9681 = ~n7986 & n9680;
  assign n9682 = n7972 & ~n9681;
  assign n9683 = ~n9677 & ~n9682;
  assign n9684 = n9676 & n9683;
  assign n9685 = n9671 & n9684;
  assign n9686 = n7995 & n9685;
  assign n9687 = n9281 & n9686;
  assign n9688 = ~n7981 & n9687;
  assign n9689 = ~n7974 & n9688;
  assign n9690 = n9689 ^ n6465;
  assign n9691 = n9690 ^ x426;
  assign n9692 = n9668 & n9691;
  assign n9693 = ~n8726 & ~n8746;
  assign n9694 = n8717 & ~n9693;
  assign n9695 = n8725 & ~n8742;
  assign n9696 = ~n9694 & ~n9695;
  assign n9697 = n8632 & n8715;
  assign n9698 = n8723 & n8725;
  assign n9699 = ~n9697 & ~n9698;
  assign n9700 = n8704 & n8740;
  assign n9701 = n8632 & n8698;
  assign n9702 = ~n9700 & ~n9701;
  assign n9703 = ~n8711 & ~n8714;
  assign n9704 = ~n8719 & ~n8747;
  assign n9705 = n8630 & ~n9704;
  assign n9706 = ~n8729 & n8743;
  assign n9707 = n8717 & ~n9706;
  assign n9708 = ~n9705 & ~n9707;
  assign n9709 = ~n9703 & n9708;
  assign n9710 = n9702 & n9709;
  assign n9711 = n8736 & n9710;
  assign n9712 = n9699 & n9711;
  assign n9713 = n9310 & n9712;
  assign n9714 = n9696 & n9713;
  assign n9715 = n9714 ^ n6433;
  assign n9716 = n9715 ^ x427;
  assign n9717 = n7748 ^ x425;
  assign n9718 = n9716 & ~n9717;
  assign n9719 = n9692 & n9718;
  assign n9720 = n9667 & n9719;
  assign n9721 = ~n9665 & ~n9666;
  assign n9722 = ~n9668 & n9691;
  assign n9723 = n9716 & n9717;
  assign n9724 = n9722 & n9723;
  assign n9725 = n9721 & n9724;
  assign n9726 = ~n9665 & n9666;
  assign n9727 = ~n9668 & ~n9691;
  assign n9728 = ~n9716 & ~n9717;
  assign n9729 = n9727 & n9728;
  assign n9730 = n9726 & n9729;
  assign n9731 = n9665 & ~n9666;
  assign n9732 = n9723 & n9727;
  assign n9733 = n9692 & n9723;
  assign n9734 = ~n9732 & ~n9733;
  assign n9735 = n9731 & ~n9734;
  assign n9736 = ~n9730 & ~n9735;
  assign n9737 = ~n9725 & n9736;
  assign n9738 = ~n9716 & n9717;
  assign n9739 = n9727 & n9738;
  assign n9740 = n9731 & n9739;
  assign n9741 = ~n9667 & ~n9721;
  assign n9742 = n9722 & n9738;
  assign n9743 = n9668 & ~n9691;
  assign n9744 = n9723 & n9743;
  assign n9745 = ~n9742 & ~n9744;
  assign n9746 = ~n9741 & ~n9745;
  assign n9747 = ~n9740 & ~n9746;
  assign n9748 = n9721 & n9733;
  assign n9749 = n9718 & n9743;
  assign n9750 = n9728 & n9743;
  assign n9751 = n9718 & n9722;
  assign n9752 = ~n9750 & ~n9751;
  assign n9753 = ~n9749 & n9752;
  assign n9754 = n9726 & ~n9753;
  assign n9755 = n9738 & n9743;
  assign n9756 = n9665 & n9755;
  assign n9757 = n9692 & n9728;
  assign n9758 = n9722 & n9728;
  assign n9759 = ~n9749 & ~n9758;
  assign n9760 = ~n9757 & n9759;
  assign n9761 = ~n9719 & n9760;
  assign n9762 = n9731 & ~n9761;
  assign n9763 = ~n9756 & ~n9762;
  assign n9764 = n9692 & n9738;
  assign n9765 = ~n9732 & ~n9744;
  assign n9766 = ~n9724 & n9765;
  assign n9767 = ~n9764 & n9766;
  assign n9768 = n9726 & ~n9767;
  assign n9769 = n9718 & n9727;
  assign n9770 = ~n9757 & ~n9769;
  assign n9771 = ~n9729 & n9770;
  assign n9772 = ~n9721 & n9771;
  assign n9773 = ~n9739 & ~n9751;
  assign n9774 = ~n9757 & n9773;
  assign n9775 = ~n9667 & n9774;
  assign n9776 = ~n9772 & ~n9775;
  assign n9777 = ~n9750 & ~n9776;
  assign n9778 = ~n9741 & ~n9777;
  assign n9779 = ~n9768 & ~n9778;
  assign n9780 = n9763 & n9779;
  assign n9781 = ~n9754 & n9780;
  assign n9782 = ~n9748 & n9781;
  assign n9783 = n9747 & n9782;
  assign n9784 = n9737 & n9783;
  assign n9785 = ~n9720 & n9784;
  assign n9786 = n9785 ^ n7844;
  assign n9787 = n9786 ^ x460;
  assign n9788 = n9664 & n9787;
  assign n9789 = ~n9476 & n9788;
  assign n9790 = ~n8590 & n9048;
  assign n9791 = n9227 & n9470;
  assign n9792 = n9790 & n9791;
  assign n9793 = n9049 & n9791;
  assign n9794 = ~n9792 & ~n9793;
  assign n9795 = n9664 & ~n9787;
  assign n9796 = ~n9794 & n9795;
  assign n9797 = ~n9789 & ~n9796;
  assign n9798 = ~n8590 & ~n9048;
  assign n9799 = n9471 & n9798;
  assign n9800 = n9474 & n9790;
  assign n9801 = ~n9799 & ~n9800;
  assign n9802 = n9787 ^ n9664;
  assign n9803 = ~n9801 & ~n9802;
  assign n9804 = n9471 & n9473;
  assign n9805 = ~n9664 & n9804;
  assign n9806 = n9471 & n9790;
  assign n9807 = ~n9664 & ~n9787;
  assign n9808 = n9806 & n9807;
  assign n9809 = ~n9805 & ~n9808;
  assign n9810 = ~n9227 & n9470;
  assign n9811 = n9790 & n9810;
  assign n9812 = n9049 & n9810;
  assign n9813 = ~n9811 & ~n9812;
  assign n9814 = n9048 ^ n8590;
  assign n9815 = n9791 & ~n9814;
  assign n9816 = n9813 & ~n9815;
  assign n9817 = ~n9802 & ~n9816;
  assign n9818 = n9049 & n9474;
  assign n9819 = ~n9806 & ~n9818;
  assign n9820 = ~n9799 & n9819;
  assign n9821 = ~n9804 & n9820;
  assign n9822 = n9795 & ~n9821;
  assign n9823 = ~n9817 & ~n9822;
  assign n9824 = n9474 & n9798;
  assign n9825 = ~n9812 & ~n9824;
  assign n9826 = n9795 & ~n9825;
  assign n9827 = ~n9664 & n9787;
  assign n9828 = n9814 ^ n9227;
  assign n9829 = n9471 & ~n9828;
  assign n9830 = n9829 ^ n9828;
  assign n9831 = ~n9824 & n9830;
  assign n9832 = n9827 & ~n9831;
  assign n9833 = ~n9826 & ~n9832;
  assign n9834 = n9823 & n9833;
  assign n9835 = n9809 & n9834;
  assign n9836 = ~n9803 & n9835;
  assign n9837 = n9797 & n9836;
  assign n9838 = n9837 ^ n8628;
  assign n9839 = n9838 ^ x532;
  assign n9840 = n8035 ^ x417;
  assign n9841 = n9584 ^ x412;
  assign n9842 = n9840 & n9841;
  assign n9843 = n8717 & ~n8751;
  assign n9844 = ~n8719 & n9693;
  assign n9845 = ~n8714 & ~n9844;
  assign n9846 = ~n9843 & ~n9845;
  assign n9847 = n8714 & n8729;
  assign n9848 = ~n8701 & ~n8723;
  assign n9849 = n8704 & ~n9848;
  assign n9850 = ~n9847 & ~n9849;
  assign n9851 = ~n8737 & ~n9317;
  assign n9852 = n8725 & ~n9851;
  assign n9853 = ~n8708 & ~n8741;
  assign n9854 = n8632 & ~n9853;
  assign n9855 = ~n9852 & ~n9854;
  assign n9856 = n9850 & n9855;
  assign n9857 = n9846 & n9856;
  assign n9858 = n8722 & n9857;
  assign n9859 = n9699 & n9858;
  assign n9860 = ~n8713 & n9859;
  assign n9861 = n9696 & n9860;
  assign n9862 = ~n8703 & n9861;
  assign n9863 = n9862 ^ n7067;
  assign n9864 = n9863 ^ x415;
  assign n9865 = n7392 ^ x416;
  assign n9866 = ~n9864 & ~n9865;
  assign n9867 = n8923 & n9357;
  assign n9868 = n8909 & n9363;
  assign n9869 = ~n9867 & ~n9868;
  assign n9870 = n8910 & n8942;
  assign n9871 = ~n9343 & ~n9870;
  assign n9872 = n8937 & ~n9871;
  assign n9873 = ~n9337 & n9350;
  assign n9874 = n8840 & ~n9873;
  assign n9875 = ~n9872 & ~n9874;
  assign n9876 = n9869 & n9875;
  assign n9877 = n9876 ^ n7083;
  assign n9878 = n9877 ^ x414;
  assign n9879 = n9503 ^ x413;
  assign n9880 = ~n9878 & n9879;
  assign n9881 = n9866 & n9880;
  assign n9882 = n9842 & n9881;
  assign n9883 = ~n9864 & n9865;
  assign n9884 = n9878 & n9879;
  assign n9885 = n9883 & n9884;
  assign n9886 = ~n9840 & ~n9841;
  assign n9887 = ~n9842 & ~n9886;
  assign n9888 = n9885 & ~n9887;
  assign n9889 = ~n9882 & ~n9888;
  assign n9890 = n9864 & n9865;
  assign n9891 = n9880 & n9890;
  assign n9892 = n9886 & n9891;
  assign n9893 = n9840 & ~n9841;
  assign n9894 = n9878 & ~n9879;
  assign n9895 = n9866 & n9894;
  assign n9896 = n9893 & n9895;
  assign n9897 = ~n9892 & ~n9896;
  assign n9898 = n9884 & n9890;
  assign n9899 = n9893 & n9898;
  assign n9900 = n9864 & ~n9865;
  assign n9901 = n9880 & n9900;
  assign n9902 = n9893 & n9901;
  assign n9903 = ~n9899 & ~n9902;
  assign n9904 = ~n9878 & ~n9879;
  assign n9905 = n9866 & n9904;
  assign n9906 = n9890 & n9904;
  assign n9907 = ~n9905 & ~n9906;
  assign n9908 = n9842 & ~n9907;
  assign n9909 = n9903 & ~n9908;
  assign n9910 = n9884 & n9900;
  assign n9911 = ~n9891 & ~n9910;
  assign n9912 = n9842 & ~n9911;
  assign n9913 = n9890 & n9894;
  assign n9914 = ~n9895 & ~n9913;
  assign n9915 = ~n9887 & ~n9914;
  assign n9916 = ~n9912 & ~n9915;
  assign n9917 = ~n9840 & n9841;
  assign n9918 = n9880 & n9883;
  assign n9919 = ~n9901 & ~n9918;
  assign n9920 = n9866 & n9884;
  assign n9921 = ~n9898 & ~n9920;
  assign n9922 = n9919 & n9921;
  assign n9923 = n9917 & ~n9922;
  assign n9924 = n9883 & n9904;
  assign n9925 = n9900 & n9904;
  assign n9926 = ~n9924 & ~n9925;
  assign n9927 = n9883 & n9894;
  assign n9928 = ~n9881 & ~n9927;
  assign n9929 = n9926 & n9928;
  assign n9930 = n9893 & ~n9929;
  assign n9931 = ~n9923 & ~n9930;
  assign n9932 = n9894 & n9900;
  assign n9933 = n9887 & n9932;
  assign n9934 = ~n9913 & n9926;
  assign n9935 = n9917 & ~n9934;
  assign n9936 = ~n9910 & n9928;
  assign n9937 = ~n9924 & n9936;
  assign n9938 = n9886 & ~n9937;
  assign n9939 = ~n9935 & ~n9938;
  assign n9940 = ~n9933 & n9939;
  assign n9941 = n9931 & n9940;
  assign n9942 = n9916 & n9941;
  assign n9943 = n9909 & n9942;
  assign n9944 = n9897 & n9943;
  assign n9945 = n9889 & n9944;
  assign n9946 = n9945 ^ n7153;
  assign n9947 = n9946 ^ x482;
  assign n9948 = ~n9409 & ~n9420;
  assign n9949 = n9419 & ~n9948;
  assign n9950 = n9278 & n9431;
  assign n9951 = ~n9443 & ~n9445;
  assign n9952 = n9433 & ~n9951;
  assign n9953 = ~n9950 & ~n9952;
  assign n9954 = n9250 & ~n9425;
  assign n9955 = ~n9417 & ~n9430;
  assign n9956 = n9453 & n9955;
  assign n9957 = n9411 & ~n9956;
  assign n9958 = ~n9954 & ~n9957;
  assign n9959 = n9436 & ~n9444;
  assign n9960 = n9278 & ~n9959;
  assign n9961 = n9278 & ~n9453;
  assign n9962 = ~n9430 & ~n9455;
  assign n9963 = ~n9414 & ~n9443;
  assign n9964 = n9962 & n9963;
  assign n9965 = ~n9406 & n9964;
  assign n9966 = n9419 & ~n9965;
  assign n9967 = ~n9961 & ~n9966;
  assign n9968 = ~n9420 & ~n9444;
  assign n9969 = n9411 & ~n9968;
  assign n9970 = n9440 & ~n9452;
  assign n9971 = ~n9434 & n9970;
  assign n9972 = n9433 & ~n9971;
  assign n9973 = ~n9969 & ~n9972;
  assign n9974 = n9967 & n9973;
  assign n9975 = ~n9960 & n9974;
  assign n9976 = n9958 & n9975;
  assign n9977 = n9953 & n9976;
  assign n9978 = ~n9949 & n9977;
  assign n9979 = ~n9432 & n9978;
  assign n9980 = ~n9407 & n9979;
  assign n9981 = n9980 ^ n8662;
  assign n9982 = n9981 ^ x481;
  assign n9983 = n8793 ^ x442;
  assign n9984 = n9368 ^ x447;
  assign n9985 = n9983 & n9984;
  assign n9986 = n9249 ^ x446;
  assign n9987 = n8766 ^ x443;
  assign n9988 = n8132 & n8156;
  assign n9989 = n8062 & ~n8599;
  assign n9990 = ~n9988 & ~n9989;
  assign n9991 = ~n8172 & n9546;
  assign n9992 = n8129 & ~n9991;
  assign n9993 = n8168 & ~n8179;
  assign n9994 = n8060 & ~n9993;
  assign n9995 = ~n9992 & ~n9994;
  assign n9996 = n8145 & ~n8616;
  assign n9997 = n8160 & n8176;
  assign n9998 = ~n8173 & n9997;
  assign n9999 = n8148 & ~n9998;
  assign n10000 = ~n9996 & ~n9999;
  assign n10001 = n9995 & n10000;
  assign n10002 = n9990 & n10001;
  assign n10003 = n8141 & n10002;
  assign n10004 = n8604 & n10003;
  assign n10005 = n8596 & n10004;
  assign n10006 = ~n8591 & n10005;
  assign n10007 = n10006 ^ n6654;
  assign n10008 = n10007 ^ x444;
  assign n10009 = n7676 & ~n7725;
  assign n10010 = n7710 & ~n7712;
  assign n10011 = ~n7679 & n10010;
  assign n10012 = n7524 & ~n10011;
  assign n10013 = ~n10009 & ~n10012;
  assign n10014 = ~n7709 & n7734;
  assign n10015 = n7696 & ~n10014;
  assign n10016 = n9116 & n9483;
  assign n10017 = ~n7683 & n10016;
  assign n10018 = n7692 & ~n10017;
  assign n10019 = ~n10015 & ~n10018;
  assign n10020 = n10013 & n10019;
  assign n10021 = n7707 & n10020;
  assign n10022 = n9479 & n10021;
  assign n10023 = n9107 & n10022;
  assign n10024 = n9100 & n10023;
  assign n10025 = n7702 & n10024;
  assign n10026 = ~n7684 & n10025;
  assign n10027 = n10026 ^ n6707;
  assign n10028 = n10027 ^ x445;
  assign n10029 = n10008 & n10028;
  assign n10030 = n9987 & n10029;
  assign n10031 = ~n9986 & n10030;
  assign n10032 = n9985 & n10031;
  assign n10033 = n9983 & ~n9984;
  assign n10034 = n9986 & n9987;
  assign n10035 = ~n10008 & n10034;
  assign n10036 = ~n10028 & n10035;
  assign n10037 = n10033 & n10036;
  assign n10038 = ~n9983 & ~n9984;
  assign n10039 = ~n9987 & ~n10028;
  assign n10040 = n10008 & n10039;
  assign n10041 = ~n9986 & n10040;
  assign n10042 = ~n10008 & n10039;
  assign n10043 = n9986 & n10042;
  assign n10044 = ~n10041 & ~n10043;
  assign n10045 = n10038 & ~n10044;
  assign n10046 = ~n10037 & ~n10045;
  assign n10047 = ~n9986 & ~n10008;
  assign n10048 = n9987 & n10047;
  assign n10049 = n10028 & n10048;
  assign n10050 = n10029 & n10034;
  assign n10051 = ~n10049 & ~n10050;
  assign n10052 = n10033 & ~n10051;
  assign n10053 = n10039 & n10047;
  assign n10054 = n9986 & n10040;
  assign n10055 = ~n10053 & ~n10054;
  assign n10056 = n9985 & ~n10055;
  assign n10057 = ~n10052 & ~n10056;
  assign n10058 = ~n10028 & n10048;
  assign n10059 = n10033 & n10058;
  assign n10060 = ~n9983 & n9984;
  assign n10061 = n9987 & n10008;
  assign n10062 = ~n10028 & n10061;
  assign n10063 = ~n9986 & n10062;
  assign n10064 = ~n10050 & ~n10063;
  assign n10065 = n10060 & ~n10064;
  assign n10066 = ~n10059 & ~n10065;
  assign n10067 = n10008 & n10034;
  assign n10068 = ~n10028 & n10067;
  assign n10069 = ~n10058 & ~n10068;
  assign n10070 = n10038 & ~n10069;
  assign n10071 = ~n9987 & ~n10008;
  assign n10072 = n10028 & n10071;
  assign n10073 = n9986 & n10072;
  assign n10074 = ~n10041 & ~n10073;
  assign n10075 = n10060 & ~n10074;
  assign n10076 = ~n10070 & ~n10075;
  assign n10077 = n10066 & n10076;
  assign n10078 = ~n9987 & n10047;
  assign n10079 = n10028 & n10078;
  assign n10080 = n9985 & n10079;
  assign n10081 = n10060 & n10068;
  assign n10082 = ~n10080 & ~n10081;
  assign n10083 = ~n9984 & n10079;
  assign n10084 = n10028 & n10035;
  assign n10085 = ~n10031 & ~n10084;
  assign n10086 = ~n10073 & n10085;
  assign n10087 = n10038 & ~n10086;
  assign n10088 = ~n9987 & n10029;
  assign n10089 = n9986 & n10088;
  assign n10090 = n10060 & ~n10089;
  assign n10091 = ~n10048 & n10090;
  assign n10092 = n10091 ^ n10060;
  assign n10093 = ~n10087 & ~n10092;
  assign n10094 = ~n10083 & n10093;
  assign n10095 = n10054 & ~n10088;
  assign n10096 = n10095 ^ n10088;
  assign n10097 = n10033 & n10096;
  assign n10098 = n9987 ^ n9986;
  assign n10099 = n10008 ^ n9987;
  assign n10100 = ~n10098 & n10099;
  assign n10101 = n9985 & n10100;
  assign n10102 = ~n10097 & ~n10101;
  assign n10103 = n10094 & n10102;
  assign n10104 = n10082 & n10103;
  assign n10105 = n10077 & n10104;
  assign n10106 = n10057 & n10105;
  assign n10107 = n10046 & n10106;
  assign n10108 = ~n10032 & n10107;
  assign n10109 = n10108 ^ n8357;
  assign n10110 = n10109 ^ x479;
  assign n10111 = ~n9982 & n10110;
  assign n10112 = n9001 & n9020;
  assign n10113 = n8985 & n9029;
  assign n10114 = n8987 & n9000;
  assign n10115 = n8990 & n10114;
  assign n10116 = ~n10113 & ~n10115;
  assign n10117 = ~n10112 & n10116;
  assign n10118 = n9005 & n9020;
  assign n10119 = ~n8998 & ~n10118;
  assign n10120 = n9011 & ~n10119;
  assign n10121 = ~n8992 & n9024;
  assign n10122 = n9010 & ~n10121;
  assign n10123 = ~n10120 & ~n10122;
  assign n10124 = ~n8629 & n9012;
  assign n10125 = ~n9029 & n9035;
  assign n10126 = ~n8988 & n10125;
  assign n10127 = n8768 & ~n10126;
  assign n10128 = ~n10124 & ~n10127;
  assign n10129 = n10123 & n10128;
  assign n10130 = ~n8983 & ~n9004;
  assign n10131 = n8990 & ~n10130;
  assign n10132 = ~n8983 & ~n9021;
  assign n10133 = ~n9010 & n10132;
  assign n10134 = ~n9012 & n9022;
  assign n10135 = ~n9006 & n10134;
  assign n10136 = ~n8985 & n10135;
  assign n10137 = ~n10133 & ~n10136;
  assign n10138 = ~n9033 & ~n10137;
  assign n10139 = ~n9011 & ~n10138;
  assign n10140 = ~n10131 & ~n10139;
  assign n10141 = n10129 & n10140;
  assign n10142 = ~n9008 & n10141;
  assign n10143 = n8997 & n10142;
  assign n10144 = n10117 & n10143;
  assign n10145 = n10144 ^ n8695;
  assign n10146 = n10145 ^ x480;
  assign n10147 = n10111 & n10146;
  assign n10148 = ~n9947 & n10147;
  assign n10149 = ~n8329 & n8546;
  assign n10150 = ~n8570 & ~n10149;
  assign n10151 = n8545 ^ n8191;
  assign n10152 = n10151 ^ n8036;
  assign n10153 = ~n8329 & n10151;
  assign n10154 = ~n10152 & n10153;
  assign n10155 = n10154 ^ n10152;
  assign n10156 = n10150 & n10155;
  assign n10157 = n8551 & ~n10156;
  assign n10158 = ~n8036 & ~n8572;
  assign n10159 = n8036 & n8555;
  assign n10160 = n8552 & ~n8559;
  assign n10161 = ~n10159 & ~n10160;
  assign n10162 = ~n10158 & n10161;
  assign n10163 = n8565 & n10162;
  assign n10164 = ~n10157 & ~n10163;
  assign n10165 = ~n8036 & n8555;
  assign n10166 = n8329 & n8546;
  assign n10167 = ~n10165 & ~n10166;
  assign n10168 = n8545 & n8552;
  assign n10169 = ~n8545 & ~n8555;
  assign n10170 = n8036 & n10169;
  assign n10171 = ~n10168 & ~n10170;
  assign n10172 = n10167 & n10171;
  assign n10173 = n8576 & ~n10172;
  assign n10174 = n8329 & ~n10151;
  assign n10175 = ~n8329 & n8553;
  assign n10176 = ~n10158 & ~n10175;
  assign n10177 = ~n10174 & n10176;
  assign n10178 = n7750 & ~n10177;
  assign n10179 = ~n10173 & ~n10178;
  assign n10180 = n10164 & n10179;
  assign n10181 = n10180 ^ n8397;
  assign n10182 = n10181 ^ x478;
  assign n10183 = n9729 & n9731;
  assign n10184 = ~n9720 & ~n10183;
  assign n10185 = ~n9739 & ~n9764;
  assign n10186 = n9726 & ~n10185;
  assign n10187 = n9731 & ~n9770;
  assign n10188 = ~n10186 & ~n10187;
  assign n10189 = n9719 & n9731;
  assign n10190 = n9667 & n9758;
  assign n10191 = ~n10189 & ~n10190;
  assign n10192 = ~n9724 & ~n9755;
  assign n10193 = n9726 & ~n10192;
  assign n10194 = ~n9755 & n9766;
  assign n10195 = n9731 & ~n10194;
  assign n10196 = n9667 & n9724;
  assign n10197 = ~n9726 & ~n10196;
  assign n10198 = ~n9751 & ~n10196;
  assign n10199 = ~n9719 & n10198;
  assign n10200 = n9759 & n10199;
  assign n10201 = ~n10197 & ~n10200;
  assign n10202 = ~n10195 & ~n10201;
  assign n10203 = ~n10193 & n10202;
  assign n10204 = ~n9739 & ~n9749;
  assign n10205 = n9721 & ~n10204;
  assign n10206 = ~n9750 & ~n9769;
  assign n10207 = ~n9721 & n9765;
  assign n10208 = ~n9733 & ~n9742;
  assign n10209 = ~n9755 & n10208;
  assign n10210 = ~n9667 & n10209;
  assign n10211 = ~n10207 & ~n10210;
  assign n10212 = n10206 & ~n10211;
  assign n10213 = ~n9764 & n10212;
  assign n10214 = ~n9741 & ~n10213;
  assign n10215 = ~n10205 & ~n10214;
  assign n10216 = n10203 & n10215;
  assign n10217 = n10191 & n10216;
  assign n10218 = n10188 & n10217;
  assign n10219 = n10184 & n10218;
  assign n10220 = n10219 ^ n6533;
  assign n10221 = n10220 ^ x483;
  assign n10222 = ~n10182 & ~n10221;
  assign n10223 = n10148 & n10222;
  assign n10224 = n10182 & n10221;
  assign n10225 = n9982 & ~n10110;
  assign n10226 = n9947 & ~n10146;
  assign n10227 = n10225 & n10226;
  assign n10228 = n10224 & n10227;
  assign n10229 = ~n10223 & ~n10228;
  assign n10230 = n10111 & n10226;
  assign n10231 = n10222 & n10230;
  assign n10232 = ~n10182 & n10221;
  assign n10233 = n9982 & n10110;
  assign n10234 = ~n9947 & ~n10146;
  assign n10235 = n10233 & n10234;
  assign n10236 = n10232 & n10235;
  assign n10237 = ~n10231 & ~n10236;
  assign n10238 = n9947 & n10146;
  assign n10239 = n10225 & n10238;
  assign n10240 = ~n9982 & ~n10110;
  assign n10241 = n10234 & n10240;
  assign n10242 = ~n10239 & ~n10241;
  assign n10243 = n10222 & ~n10242;
  assign n10244 = n9947 & n10147;
  assign n10245 = ~n9947 & n10146;
  assign n10246 = n10233 & n10245;
  assign n10247 = ~n10244 & ~n10246;
  assign n10248 = n10221 & ~n10247;
  assign n10249 = n10225 & n10245;
  assign n10250 = n10233 & n10238;
  assign n10251 = ~n10148 & ~n10230;
  assign n10252 = ~n10250 & n10251;
  assign n10253 = ~n10241 & n10252;
  assign n10254 = ~n10249 & n10253;
  assign n10255 = n10224 & ~n10254;
  assign n10256 = ~n10248 & ~n10255;
  assign n10257 = n10182 & ~n10221;
  assign n10258 = n10111 & n10234;
  assign n10259 = ~n10235 & ~n10250;
  assign n10260 = ~n10258 & n10259;
  assign n10261 = n10238 & n10240;
  assign n10262 = n10225 & n10234;
  assign n10263 = ~n10261 & ~n10262;
  assign n10264 = n10240 & n10245;
  assign n10265 = n10226 & n10240;
  assign n10266 = ~n10264 & ~n10265;
  assign n10267 = ~n10239 & n10266;
  assign n10268 = n10263 & n10267;
  assign n10269 = n10260 & n10268;
  assign n10270 = n10257 & ~n10269;
  assign n10271 = n10226 & n10233;
  assign n10272 = ~n10246 & ~n10271;
  assign n10273 = ~n10261 & n10272;
  assign n10274 = ~n10264 & n10273;
  assign n10275 = n10222 & ~n10274;
  assign n10276 = ~n10239 & ~n10262;
  assign n10277 = ~n10258 & n10276;
  assign n10278 = n10266 & n10277;
  assign n10279 = n10232 & ~n10278;
  assign n10280 = ~n10275 & ~n10279;
  assign n10281 = ~n10270 & n10280;
  assign n10282 = n10256 & n10281;
  assign n10283 = ~n10243 & n10282;
  assign n10284 = n10237 & n10283;
  assign n10285 = n10229 & n10284;
  assign n10286 = n10285 ^ n8766;
  assign n10287 = n10286 ^ x537;
  assign n10288 = n9839 & n10287;
  assign n10289 = n9047 ^ x466;
  assign n10290 = n9250 & ~n9435;
  assign n10291 = n9423 ^ n9405;
  assign n10292 = n9419 & n10291;
  assign n10293 = ~n10290 & ~n10292;
  assign n10294 = n9409 & n9411;
  assign n10295 = n9456 & n9962;
  assign n10296 = ~n9422 & n10295;
  assign n10297 = n9278 & ~n10296;
  assign n10298 = ~n9433 & n9453;
  assign n10299 = ~n9417 & ~n9439;
  assign n10300 = ~n9411 & n10299;
  assign n10301 = ~n10298 & ~n10300;
  assign n10302 = ~n9406 & ~n10301;
  assign n10303 = ~n9431 & n10302;
  assign n10304 = n9250 & ~n10303;
  assign n10305 = ~n10297 & ~n10304;
  assign n10306 = ~n10294 & n10305;
  assign n10307 = n10293 & n10306;
  assign n10308 = n9953 & n10307;
  assign n10309 = ~n9949 & n10308;
  assign n10310 = n9416 & n10309;
  assign n10311 = n10310 ^ n8446;
  assign n10312 = n10311 ^ x471;
  assign n10313 = ~n10289 & n10312;
  assign n10314 = n9842 & n9925;
  assign n10315 = n9886 & n9913;
  assign n10316 = ~n10314 & ~n10315;
  assign n10317 = n9893 & n9924;
  assign n10318 = n9917 & ~n9921;
  assign n10319 = ~n10317 & ~n10318;
  assign n10320 = ~n9898 & ~n9913;
  assign n10321 = n9842 & ~n10320;
  assign n10322 = ~n9906 & ~n9932;
  assign n10323 = n9886 & ~n10322;
  assign n10324 = ~n10321 & ~n10323;
  assign n10325 = ~n9911 & n9917;
  assign n10326 = ~n9895 & n9919;
  assign n10327 = ~n9887 & ~n10326;
  assign n10328 = ~n9905 & ~n9927;
  assign n10329 = n9926 & n10328;
  assign n10330 = n9917 & ~n10329;
  assign n10331 = ~n9927 & ~n9932;
  assign n10332 = ~n9905 & n9911;
  assign n10333 = ~n9920 & n10332;
  assign n10334 = n10331 & n10333;
  assign n10335 = n9893 & ~n10334;
  assign n10336 = ~n10330 & ~n10335;
  assign n10337 = ~n9902 & n10336;
  assign n10338 = ~n10327 & n10337;
  assign n10339 = ~n10325 & n10338;
  assign n10340 = n10324 & n10339;
  assign n10341 = ~n9892 & n10340;
  assign n10342 = n10319 & n10341;
  assign n10343 = n9889 & n10342;
  assign n10344 = n10316 & n10343;
  assign n10345 = n10344 ^ n8387;
  assign n10346 = n10345 ^ x470;
  assign n10347 = n9663 ^ x467;
  assign n10348 = n9985 & n10073;
  assign n10349 = n10044 & ~n10054;
  assign n10350 = n10038 & ~n10349;
  assign n10351 = ~n10348 & ~n10350;
  assign n10352 = ~n9986 & n10088;
  assign n10353 = ~n9984 & n10352;
  assign n10354 = n10051 & ~n10084;
  assign n10355 = n10060 & ~n10354;
  assign n10356 = n9985 & n10063;
  assign n10357 = ~n10036 & ~n10049;
  assign n10358 = ~n10042 & n10357;
  assign n10359 = ~n10063 & n10358;
  assign n10360 = ~n10089 & n10359;
  assign n10361 = ~n10068 & n10360;
  assign n10362 = n10033 & ~n10361;
  assign n10363 = n10349 & ~n10352;
  assign n10364 = n10060 & ~n10363;
  assign n10365 = n9984 ^ n9983;
  assign n10366 = ~n10032 & n10354;
  assign n10367 = ~n10031 & ~n10050;
  assign n10368 = ~n10038 & n10367;
  assign n10369 = ~n10366 & ~n10368;
  assign n10370 = ~n10058 & ~n10369;
  assign n10371 = ~n10365 & ~n10370;
  assign n10372 = ~n10364 & ~n10371;
  assign n10373 = ~n10362 & n10372;
  assign n10374 = ~n10356 & n10373;
  assign n10375 = ~n10355 & n10374;
  assign n10376 = ~n10353 & n10375;
  assign n10377 = n10351 & n10376;
  assign n10378 = n10082 & n10377;
  assign n10379 = ~n10056 & n10378;
  assign n10380 = n10379 ^ n8868;
  assign n10381 = n10380 ^ x469;
  assign n10382 = ~n10347 & n10381;
  assign n10383 = n10346 & n10382;
  assign n10384 = n9770 & n10185;
  assign n10385 = ~n9749 & n10384;
  assign n10386 = n9667 & ~n10385;
  assign n10387 = n9716 ^ n9691;
  assign n10388 = n10387 ^ n9668;
  assign n10389 = ~n9717 & n10388;
  assign n10390 = n9721 & n10389;
  assign n10391 = ~n10386 & ~n10390;
  assign n10392 = n9731 & ~n9774;
  assign n10393 = ~n9741 & n9755;
  assign n10394 = ~n9666 & ~n9745;
  assign n10395 = ~n10393 & ~n10394;
  assign n10396 = n9734 & n9774;
  assign n10397 = n9759 & n10396;
  assign n10398 = n9726 & ~n10397;
  assign n10399 = n10395 & ~n10398;
  assign n10400 = ~n10392 & n10399;
  assign n10401 = n10391 & n10400;
  assign n10402 = n9737 & n10401;
  assign n10403 = n10184 & n10402;
  assign n10404 = ~n10196 & n10403;
  assign n10405 = n10404 ^ n8901;
  assign n10406 = n10405 ^ x468;
  assign n10407 = n10346 & n10406;
  assign n10408 = n10347 & ~n10381;
  assign n10409 = ~n10407 & n10408;
  assign n10410 = ~n10383 & ~n10409;
  assign n10412 = ~n10346 & ~n10406;
  assign n10411 = ~n10346 & n10406;
  assign n10413 = n10412 ^ n10411;
  assign n10414 = ~n10347 & n10413;
  assign n10415 = n10414 ^ n10412;
  assign n10416 = n10410 & ~n10415;
  assign n10417 = n10313 & n10416;
  assign n10418 = n10289 & n10312;
  assign n10419 = n10347 & n10381;
  assign n10420 = n10411 & n10419;
  assign n10421 = n10381 ^ n10346;
  assign n10422 = ~n10406 & ~n10421;
  assign n10423 = ~n10347 & n10422;
  assign n10424 = n10346 & n10408;
  assign n10425 = n10406 ^ n10381;
  assign n10426 = n10406 ^ n10346;
  assign n10427 = n10425 & ~n10426;
  assign n10428 = ~n10424 & n10427;
  assign n10429 = n10428 ^ n10424;
  assign n10430 = ~n10423 & ~n10429;
  assign n10431 = ~n10420 & n10430;
  assign n10432 = n10418 & n10431;
  assign n10433 = ~n10417 & ~n10432;
  assign n10434 = n10289 & ~n10312;
  assign n10435 = ~n10347 & n10407;
  assign n10436 = n10412 & ~n10419;
  assign n10437 = ~n10435 & ~n10436;
  assign n10438 = n10346 & ~n10406;
  assign n10439 = n10419 & n10438;
  assign n10440 = ~n10347 & ~n10381;
  assign n10441 = ~n10346 & n10440;
  assign n10442 = ~n10439 & ~n10441;
  assign n10443 = n10437 & n10442;
  assign n10444 = ~n10420 & n10443;
  assign n10445 = n10434 & ~n10444;
  assign n10446 = ~n10289 & ~n10312;
  assign n10447 = n10406 & n10408;
  assign n10448 = n10438 & n10440;
  assign n10449 = n10347 & n10411;
  assign n10450 = n10449 ^ n10346;
  assign n10451 = ~n10407 & n10450;
  assign n10452 = n10381 & ~n10451;
  assign n10453 = ~n10448 & ~n10452;
  assign n10454 = ~n10447 & n10453;
  assign n10455 = n10446 & ~n10454;
  assign n10456 = ~n10445 & ~n10455;
  assign n10457 = n10433 & n10456;
  assign n10458 = n10457 ^ n8949;
  assign n10459 = n10458 ^ x534;
  assign n10460 = ~n8549 & n8576;
  assign n10461 = n8551 & ~n8574;
  assign n10462 = ~n10460 & ~n10461;
  assign n10463 = n7750 & ~n8585;
  assign n10464 = n8547 & n8553;
  assign n10465 = n8191 & ~n8579;
  assign n10466 = ~n10159 & ~n10465;
  assign n10467 = ~n8558 & n10466;
  assign n10468 = n8565 & ~n10467;
  assign n10469 = ~n10464 & ~n10468;
  assign n10470 = ~n10463 & n10469;
  assign n10471 = n10462 & n10470;
  assign n10472 = n10471 ^ n7637;
  assign n10473 = n10472 ^ x495;
  assign n10474 = n9589 & n9621;
  assign n10475 = ~n9587 & n9644;
  assign n10476 = n9613 & ~n10475;
  assign n10477 = ~n10474 & ~n10476;
  assign n10478 = n9603 & n9642;
  assign n10479 = n9625 & ~n10478;
  assign n10480 = n9630 & ~n9636;
  assign n10481 = n9505 & n9627;
  assign n10482 = ~n10480 & ~n10481;
  assign n10483 = ~n9477 & n9592;
  assign n10484 = ~n9609 & n9613;
  assign n10485 = ~n10483 & ~n10484;
  assign n10486 = ~n9638 & ~n9649;
  assign n10487 = ~n9636 & ~n10486;
  assign n10488 = ~n9608 & n9617;
  assign n10489 = ~n9594 & n10488;
  assign n10490 = ~n9623 & n10489;
  assign n10491 = n9589 & ~n10490;
  assign n10492 = ~n10487 & ~n10491;
  assign n10493 = n10485 & n10492;
  assign n10494 = n9629 & n10493;
  assign n10495 = n10482 & n10494;
  assign n10496 = n9620 & n10495;
  assign n10497 = n10479 & n10496;
  assign n10498 = ~n9602 & n10497;
  assign n10499 = n10477 & n10498;
  assign n10500 = ~n9633 & n10499;
  assign n10501 = n10500 ^ n7032;
  assign n10502 = n10501 ^ x490;
  assign n10503 = n10473 & n10502;
  assign n10504 = ~n9431 & n9962;
  assign n10505 = n9278 & ~n10504;
  assign n10506 = n9411 & ~n9426;
  assign n10507 = ~n10505 & ~n10506;
  assign n10508 = n9250 & n9409;
  assign n10509 = n9435 & n9951;
  assign n10510 = n9419 & ~n10509;
  assign n10511 = ~n10508 & ~n10510;
  assign n10512 = ~n9434 & n9446;
  assign n10513 = n9433 & ~n10512;
  assign n10514 = ~n9439 & n10504;
  assign n10515 = n9411 & ~n10514;
  assign n10516 = ~n9417 & ~n9422;
  assign n10517 = n9453 & n10516;
  assign n10518 = n9433 & ~n10517;
  assign n10519 = ~n10515 & ~n10518;
  assign n10520 = n9419 & ~n9970;
  assign n10521 = ~n9409 & n9963;
  assign n10522 = ~n9434 & n10521;
  assign n10523 = n9278 & ~n10522;
  assign n10524 = ~n10520 & ~n10523;
  assign n10525 = n10519 & n10524;
  assign n10526 = ~n9432 & n10525;
  assign n10527 = ~n10513 & n10526;
  assign n10528 = n10511 & n10527;
  assign n10529 = n10507 & n10528;
  assign n10530 = ~n9407 & n10529;
  assign n10531 = n10530 ^ n8230;
  assign n10532 = n10531 ^ x493;
  assign n10533 = n9163 & n9189;
  assign n10534 = ~n9168 & ~n9179;
  assign n10535 = n9177 & ~n10534;
  assign n10536 = ~n10533 & ~n10535;
  assign n10537 = n9160 & n9189;
  assign n10538 = n9168 & n9194;
  assign n10539 = ~n10537 & ~n10538;
  assign n10540 = ~n9059 & n9214;
  assign n10541 = n9177 & n9203;
  assign n10542 = ~n10540 & ~n10541;
  assign n10543 = n9192 & n9196;
  assign n10544 = n9060 & ~n10543;
  assign n10545 = ~n9184 & ~n9191;
  assign n10546 = ~n9179 & n10545;
  assign n10547 = ~n9172 & n10546;
  assign n10548 = n9189 & ~n10547;
  assign n10549 = ~n10544 & ~n10548;
  assign n10550 = n9096 ^ n9061;
  assign n10551 = n9158 & n10550;
  assign n10552 = ~n9166 & ~n10551;
  assign n10553 = n9204 & ~n9209;
  assign n10554 = ~n9186 & n10553;
  assign n10555 = ~n9177 & n10554;
  assign n10556 = ~n10552 & ~n10555;
  assign n10557 = ~n9194 & n10556;
  assign n10558 = n10549 & ~n10557;
  assign n10559 = n9158 & n9166;
  assign n10560 = n9096 & n10559;
  assign n10561 = n10558 & ~n10560;
  assign n10562 = n10542 & n10561;
  assign n10563 = n10539 & n10562;
  assign n10564 = ~n9213 & n10563;
  assign n10565 = n10536 & n10564;
  assign n10566 = ~n9165 & n10565;
  assign n10567 = n10566 ^ n7328;
  assign n10568 = n10567 ^ x491;
  assign n10591 = n9881 & n9886;
  assign n10592 = n9887 & ~n9907;
  assign n10593 = ~n10591 & ~n10592;
  assign n10594 = ~n9887 & n9898;
  assign n10595 = n9842 & ~n10331;
  assign n10596 = ~n10594 & ~n10595;
  assign n10597 = ~n9918 & ~n9920;
  assign n10598 = ~n9925 & n10597;
  assign n10599 = n9887 & ~n10598;
  assign n10600 = ~n9891 & n9914;
  assign n10601 = n9917 & ~n10600;
  assign n10602 = ~n10599 & ~n10601;
  assign n10603 = n9893 & n9927;
  assign n10604 = n9919 & n9926;
  assign n10605 = n9886 & ~n10604;
  assign n10606 = ~n10603 & ~n10605;
  assign n10607 = n10602 & n10606;
  assign n10608 = n10596 & n10607;
  assign n10609 = n10593 & n10608;
  assign n10610 = n9909 & n10609;
  assign n10611 = n9889 & n10610;
  assign n10612 = n10316 & n10611;
  assign n10613 = n10612 ^ n8259;
  assign n10614 = n10613 ^ x492;
  assign n10569 = n8990 & n9006;
  assign n10570 = n8985 & n8992;
  assign n10571 = ~n10569 & ~n10570;
  assign n10572 = ~n9011 & ~n9022;
  assign n10573 = n8990 & ~n9030;
  assign n10574 = ~n10572 & ~n10573;
  assign n10575 = n8837 & n9001;
  assign n10576 = ~n9023 & ~n10114;
  assign n10577 = n10130 & n10576;
  assign n10578 = n8994 & n10577;
  assign n10579 = n9010 & ~n10578;
  assign n10580 = ~n10575 & ~n10579;
  assign n10581 = n8985 & ~n9035;
  assign n10582 = n8768 & n9041;
  assign n10583 = ~n10581 & ~n10582;
  assign n10584 = n10580 & n10583;
  assign n10585 = n10574 & n10584;
  assign n10586 = n10571 & n10585;
  assign n10587 = n9009 & n10586;
  assign n10588 = n10117 & n10587;
  assign n10589 = n10588 ^ n7491;
  assign n10590 = n10589 ^ x494;
  assign n10615 = n10614 ^ n10590;
  assign n10616 = ~n10568 & ~n10615;
  assign n10617 = ~n10532 & n10616;
  assign n10618 = n10503 & n10617;
  assign n10619 = ~n10473 & ~n10502;
  assign n10620 = ~n10590 & ~n10614;
  assign n10621 = ~n10568 & n10620;
  assign n10622 = n10532 & n10621;
  assign n10623 = n10619 & n10622;
  assign n10624 = n10502 ^ n10473;
  assign n10625 = n10614 ^ n10532;
  assign n10626 = n10615 & ~n10625;
  assign n10627 = ~n10568 & n10626;
  assign n10628 = ~n10624 & n10627;
  assign n10629 = ~n10623 & ~n10628;
  assign n10630 = ~n10473 & n10502;
  assign n10631 = n10590 & ~n10614;
  assign n10632 = ~n10568 & n10631;
  assign n10633 = ~n10532 & n10632;
  assign n10634 = ~n10568 & n10614;
  assign n10635 = ~n10590 & n10634;
  assign n10636 = ~n10532 & n10635;
  assign n10637 = ~n10633 & ~n10636;
  assign n10638 = n10630 & ~n10637;
  assign n10639 = n10473 & ~n10502;
  assign n10640 = ~n10532 & n10568;
  assign n10641 = n10614 & n10640;
  assign n10642 = ~n10590 & n10641;
  assign n10643 = n10532 & n10568;
  assign n10644 = n10614 & n10643;
  assign n10645 = n10590 & n10644;
  assign n10646 = ~n10642 & ~n10645;
  assign n10647 = n10631 & n10643;
  assign n10648 = ~n10590 & n10644;
  assign n10649 = ~n10647 & ~n10648;
  assign n10650 = n10646 & n10649;
  assign n10651 = n10639 & ~n10650;
  assign n10652 = n10620 & n10643;
  assign n10653 = n10630 & n10652;
  assign n10654 = n10620 & n10640;
  assign n10655 = n10630 & n10654;
  assign n10656 = n10590 & n10641;
  assign n10657 = n10619 & n10656;
  assign n10658 = ~n10655 & ~n10657;
  assign n10659 = ~n10645 & ~n10656;
  assign n10660 = n10630 & ~n10659;
  assign n10661 = n10631 & n10640;
  assign n10662 = ~n10652 & ~n10654;
  assign n10663 = ~n10661 & n10662;
  assign n10664 = n10619 & ~n10663;
  assign n10665 = ~n10660 & ~n10664;
  assign n10666 = n10646 & ~n10652;
  assign n10667 = ~n10647 & n10666;
  assign n10668 = n10503 & ~n10667;
  assign n10669 = n10532 & n10632;
  assign n10670 = ~n10617 & ~n10636;
  assign n10671 = ~n10669 & n10670;
  assign n10672 = n10639 & ~n10671;
  assign n10673 = ~n10668 & ~n10672;
  assign n10674 = n10665 & n10673;
  assign n10675 = n10658 & n10674;
  assign n10676 = ~n10653 & n10675;
  assign n10677 = ~n10651 & n10676;
  assign n10678 = ~n10638 & n10677;
  assign n10679 = n10629 & n10678;
  assign n10680 = n10590 & n10634;
  assign n10681 = n10532 & n10680;
  assign n10682 = n10630 & n10669;
  assign n10683 = n10681 & ~n10682;
  assign n10684 = ~n10473 & n10683;
  assign n10685 = n10684 ^ n10682;
  assign n10686 = n10679 & ~n10685;
  assign n10687 = ~n10618 & n10686;
  assign n10688 = n10687 ^ n8835;
  assign n10689 = n10688 ^ x535;
  assign n10690 = ~n10459 & ~n10689;
  assign n10691 = n10109 ^ x477;
  assign n10692 = n10345 ^ x472;
  assign n10693 = n10691 & n10692;
  assign n10694 = ~n9190 & ~n9195;
  assign n10695 = ~n9059 & ~n10694;
  assign n10696 = ~n9172 & n9204;
  assign n10697 = ~n9208 & n10696;
  assign n10698 = n9177 & ~n10697;
  assign n10699 = ~n10695 & ~n10698;
  assign n10700 = n9194 & ~n10545;
  assign n10701 = n9192 & ~n9195;
  assign n10702 = n9210 & n10701;
  assign n10703 = ~n9186 & n10702;
  assign n10704 = n9166 & ~n10703;
  assign n10705 = ~n10700 & ~n10704;
  assign n10706 = ~n9186 & ~n9202;
  assign n10707 = ~n9060 & n10706;
  assign n10708 = ~n9189 & n9215;
  assign n10709 = ~n10707 & ~n10708;
  assign n10710 = n9169 & ~n10709;
  assign n10711 = n9194 & ~n10710;
  assign n10712 = n10705 & ~n10711;
  assign n10713 = n10699 & n10712;
  assign n10714 = n9183 & n10713;
  assign n10715 = n10714 ^ n8476;
  assign n10716 = n10715 ^ x475;
  assign n10717 = n10311 ^ x473;
  assign n10718 = n10716 & ~n10717;
  assign n10719 = n10181 ^ x476;
  assign n10720 = ~n9623 & ~n9642;
  assign n10721 = n9589 & ~n10720;
  assign n10722 = n9609 & ~n9623;
  assign n10723 = ~n9600 & n10722;
  assign n10724 = n9505 & ~n10723;
  assign n10725 = ~n9587 & ~n9638;
  assign n10726 = ~n9600 & n10725;
  assign n10727 = ~n9607 & n10726;
  assign n10728 = ~n9621 & n10727;
  assign n10729 = n9613 & ~n10728;
  assign n10730 = ~n9616 & ~n9627;
  assign n10731 = n9589 & ~n10730;
  assign n10732 = n9617 & n9650;
  assign n10733 = n9603 & ~n10732;
  assign n10734 = ~n10731 & ~n10733;
  assign n10735 = ~n10729 & n10734;
  assign n10736 = ~n10724 & n10735;
  assign n10737 = ~n10721 & n10736;
  assign n10738 = ~n9632 & n10737;
  assign n10739 = n10482 & n10738;
  assign n10740 = n9611 & n10739;
  assign n10741 = n10479 & n10740;
  assign n10742 = ~n9633 & n10741;
  assign n10743 = n9597 & n10742;
  assign n10744 = n10743 ^ n8420;
  assign n10745 = n10744 ^ x474;
  assign n10746 = ~n10719 & n10745;
  assign n10747 = n10718 & n10746;
  assign n10748 = n10693 & n10747;
  assign n10749 = ~n10691 & n10692;
  assign n10750 = ~n10716 & n10717;
  assign n10751 = ~n10719 & ~n10745;
  assign n10752 = n10750 & n10751;
  assign n10753 = n10749 & n10752;
  assign n10754 = ~n10691 & ~n10692;
  assign n10755 = n10719 & n10745;
  assign n10756 = n10750 & n10755;
  assign n10757 = n10716 & n10717;
  assign n10758 = n10746 & n10757;
  assign n10759 = ~n10756 & ~n10758;
  assign n10760 = n10754 & ~n10759;
  assign n10761 = ~n10753 & ~n10760;
  assign n10762 = n10752 & n10754;
  assign n10763 = n10691 & ~n10692;
  assign n10764 = n10718 & n10755;
  assign n10765 = ~n10716 & ~n10717;
  assign n10766 = n10755 & n10765;
  assign n10767 = n10718 & n10751;
  assign n10768 = ~n10766 & ~n10767;
  assign n10769 = ~n10764 & n10768;
  assign n10770 = n10763 & ~n10769;
  assign n10771 = ~n10762 & ~n10770;
  assign n10772 = n10746 & n10750;
  assign n10773 = ~n10693 & ~n10754;
  assign n10774 = n10772 & ~n10773;
  assign n10775 = n10719 & ~n10745;
  assign n10776 = n10718 & n10775;
  assign n10777 = n10751 & n10765;
  assign n10778 = ~n10776 & ~n10777;
  assign n10779 = ~n10766 & n10778;
  assign n10780 = n10693 & ~n10779;
  assign n10781 = ~n10774 & ~n10780;
  assign n10782 = n10757 & n10775;
  assign n10783 = n10755 & n10757;
  assign n10784 = n10751 & n10757;
  assign n10785 = ~n10783 & ~n10784;
  assign n10786 = ~n10782 & n10785;
  assign n10787 = n10692 & ~n10786;
  assign n10788 = n10750 & n10775;
  assign n10789 = ~n10772 & ~n10788;
  assign n10790 = ~n10783 & n10789;
  assign n10791 = ~n10752 & n10790;
  assign n10792 = ~n10747 & n10791;
  assign n10793 = n10763 & ~n10792;
  assign n10794 = n10746 & n10765;
  assign n10795 = n10765 & n10775;
  assign n10796 = ~n10794 & ~n10795;
  assign n10797 = ~n10776 & n10796;
  assign n10798 = ~n10754 & n10797;
  assign n10799 = ~n10747 & n10798;
  assign n10800 = ~n10767 & n10778;
  assign n10801 = ~n10788 & n10800;
  assign n10802 = ~n10749 & n10801;
  assign n10803 = ~n10799 & ~n10802;
  assign n10804 = ~n10691 & n10803;
  assign n10805 = ~n10793 & ~n10804;
  assign n10806 = ~n10787 & n10805;
  assign n10807 = n10781 & n10806;
  assign n10808 = n10771 & n10807;
  assign n10809 = n10761 & n10808;
  assign n10810 = ~n10748 & n10809;
  assign n10811 = n10810 ^ n8980;
  assign n10812 = n10811 ^ x533;
  assign n10813 = n9469 ^ x459;
  assign n10814 = n9177 & n9202;
  assign n10815 = n9189 & n9209;
  assign n10816 = ~n10814 & ~n10815;
  assign n10817 = ~n9059 & n9172;
  assign n10818 = n9194 & n9214;
  assign n10819 = n9060 & n9203;
  assign n10820 = n9177 & ~n10545;
  assign n10821 = ~n10819 & ~n10820;
  assign n10822 = ~n9186 & ~n9208;
  assign n10823 = ~n9194 & ~n10822;
  assign n10824 = n9212 & n10534;
  assign n10825 = n9196 & n10824;
  assign n10826 = n9166 & ~n10825;
  assign n10827 = n9192 & ~n9208;
  assign n10828 = ~n9189 & n10827;
  assign n10829 = ~n9060 & n10701;
  assign n10830 = ~n10828 & ~n10829;
  assign n10831 = ~n9174 & ~n10830;
  assign n10832 = n9194 & ~n10831;
  assign n10833 = ~n10826 & ~n10832;
  assign n10834 = ~n10823 & n10833;
  assign n10835 = n10821 & n10834;
  assign n10836 = ~n10818 & n10835;
  assign n10837 = ~n10817 & n10836;
  assign n10838 = n10816 & n10837;
  assign n10839 = n10536 & n10838;
  assign n10840 = ~n9165 & n10839;
  assign n10841 = n10840 ^ n7671;
  assign n10842 = n10841 ^ x454;
  assign n10843 = n10813 & ~n10842;
  assign n10844 = ~n8988 & n10576;
  assign n10845 = ~n9011 & ~n10844;
  assign n10846 = ~n9012 & n9036;
  assign n10847 = n9011 & ~n10846;
  assign n10848 = ~n9004 & ~n10118;
  assign n10849 = n9022 & n10848;
  assign n10850 = n8768 & ~n10849;
  assign n10851 = ~n9006 & n9031;
  assign n10852 = n8985 & ~n10851;
  assign n10853 = ~n10850 & ~n10852;
  assign n10854 = ~n10847 & n10853;
  assign n10855 = ~n10845 & n10854;
  assign n10856 = ~n8988 & n10119;
  assign n10857 = n8990 & ~n10856;
  assign n10858 = ~n8998 & n9039;
  assign n10859 = n9010 & ~n10858;
  assign n10860 = ~n10857 & ~n10859;
  assign n10861 = n10855 & n10860;
  assign n10862 = n10571 & n10861;
  assign n10863 = n10862 ^ n7821;
  assign n10864 = n10863 ^ x457;
  assign n10865 = n10033 & n10068;
  assign n10866 = n9985 & n10084;
  assign n10867 = ~n9984 & n10089;
  assign n10868 = ~n10866 & ~n10867;
  assign n10869 = ~n10865 & n10868;
  assign n10870 = n10068 & ~n10365;
  assign n10871 = n10031 & n10033;
  assign n10872 = n10051 & ~n10063;
  assign n10873 = n10038 & ~n10872;
  assign n10874 = ~n10042 & n10074;
  assign n10875 = n9985 & ~n10874;
  assign n10876 = ~n10873 & ~n10875;
  assign n10877 = ~n10053 & ~n10096;
  assign n10878 = n10357 & n10877;
  assign n10879 = n10060 & ~n10878;
  assign n10880 = n10033 & n10078;
  assign n10881 = ~n10073 & ~n10880;
  assign n10882 = ~n9984 & ~n10881;
  assign n10883 = ~n10879 & ~n10882;
  assign n10884 = n10876 & n10883;
  assign n10885 = ~n10871 & n10884;
  assign n10886 = ~n10870 & n10885;
  assign n10887 = n10046 & n10886;
  assign n10888 = n10869 & n10887;
  assign n10889 = n10066 & n10888;
  assign n10890 = ~n10032 & n10889;
  assign n10891 = ~n10356 & n10890;
  assign n10892 = n10891 ^ n7522;
  assign n10893 = n10892 ^ x455;
  assign n10894 = ~n10864 & ~n10893;
  assign n10895 = ~n9885 & ~n9891;
  assign n10896 = n9842 & ~n10895;
  assign n10897 = ~n9918 & n10331;
  assign n10898 = ~n9881 & n10897;
  assign n10899 = n9917 & ~n10898;
  assign n10900 = ~n10896 & ~n10899;
  assign n10901 = ~n9885 & ~n9910;
  assign n10902 = n9893 & ~n10901;
  assign n10903 = ~n9913 & n10328;
  assign n10904 = ~n9886 & n10903;
  assign n10905 = ~n9925 & n10331;
  assign n10906 = ~n9842 & n10905;
  assign n10907 = ~n10904 & ~n10906;
  assign n10908 = n10597 & ~n10907;
  assign n10909 = ~n9887 & ~n10908;
  assign n10910 = ~n10902 & ~n10909;
  assign n10911 = n10900 & n10910;
  assign n10912 = n9903 & n10911;
  assign n10913 = n10593 & n10912;
  assign n10914 = n10319 & n10913;
  assign n10915 = n9897 & n10914;
  assign n10916 = n10316 & n10915;
  assign n10917 = n10916 ^ n7786;
  assign n10918 = n10917 ^ x456;
  assign n10919 = n9786 ^ x458;
  assign n10920 = n10918 & n10919;
  assign n10921 = n10894 & n10920;
  assign n10922 = ~n10918 & ~n10919;
  assign n10923 = n10894 & n10922;
  assign n10924 = ~n10921 & ~n10923;
  assign n10925 = n10843 & ~n10924;
  assign n10926 = ~n10813 & ~n10842;
  assign n10927 = ~n10864 & n10893;
  assign n10928 = n10920 & n10927;
  assign n10929 = n10864 & n10893;
  assign n10930 = n10922 & n10929;
  assign n10931 = ~n10928 & ~n10930;
  assign n10932 = n10926 & ~n10931;
  assign n10933 = ~n10925 & ~n10932;
  assign n10934 = n10918 & ~n10919;
  assign n10935 = n10927 & n10934;
  assign n10936 = n10842 & n10935;
  assign n10937 = ~n10813 & n10842;
  assign n10938 = ~n10918 & n10919;
  assign n10939 = n10927 & n10938;
  assign n10940 = n10929 & n10934;
  assign n10941 = ~n10939 & ~n10940;
  assign n10942 = ~n10928 & n10941;
  assign n10943 = n10937 & ~n10942;
  assign n10944 = ~n10936 & ~n10943;
  assign n10945 = n10813 & n10842;
  assign n10946 = n10864 & ~n10893;
  assign n10947 = n10920 & n10946;
  assign n10948 = n10945 & n10947;
  assign n10949 = n10934 & n10946;
  assign n10950 = ~n10939 & ~n10949;
  assign n10951 = n10843 & ~n10950;
  assign n10952 = n10842 ^ n10813;
  assign n10953 = n10920 & n10929;
  assign n10954 = n10922 & n10927;
  assign n10955 = ~n10953 & ~n10954;
  assign n10956 = ~n10952 & ~n10955;
  assign n10957 = n10929 & n10938;
  assign n10958 = n10931 & ~n10940;
  assign n10959 = ~n10957 & n10958;
  assign n10960 = n10843 & ~n10959;
  assign n10961 = n10894 & n10938;
  assign n10962 = n10922 & n10946;
  assign n10963 = ~n10961 & ~n10962;
  assign n10964 = ~n10949 & n10963;
  assign n10965 = ~n10921 & n10964;
  assign n10966 = n10926 & ~n10965;
  assign n10967 = ~n10960 & ~n10966;
  assign n10968 = ~n10956 & n10967;
  assign n10969 = n10938 & n10946;
  assign n10970 = n10894 & n10934;
  assign n10971 = ~n10969 & ~n10970;
  assign n10972 = n10945 & ~n10963;
  assign n10973 = ~n10923 & ~n10947;
  assign n10974 = n10937 & ~n10973;
  assign n10975 = ~n10972 & ~n10974;
  assign n10976 = n10971 & n10975;
  assign n10977 = n10842 & ~n10976;
  assign n10978 = n10968 & ~n10977;
  assign n10979 = ~n10951 & n10978;
  assign n10980 = ~n10948 & n10979;
  assign n10981 = n10944 & n10980;
  assign n10982 = n10933 & n10981;
  assign n10983 = n10982 ^ n8793;
  assign n10984 = n10983 ^ x536;
  assign n10985 = n10812 & n10984;
  assign n10986 = n10690 & n10985;
  assign n10987 = ~n10459 & n10689;
  assign n10988 = n10812 & ~n10984;
  assign n10989 = n10987 & n10988;
  assign n10990 = ~n10986 & ~n10989;
  assign n10991 = n10288 & ~n10990;
  assign n10992 = ~n9839 & n10287;
  assign n10993 = n10459 & ~n10689;
  assign n10994 = n10985 & n10993;
  assign n10995 = n10690 & n10988;
  assign n10996 = ~n10994 & ~n10995;
  assign n10997 = n10992 & ~n10996;
  assign n10998 = ~n10991 & ~n10997;
  assign n10999 = ~n10812 & n10984;
  assign n11000 = n10993 & n10999;
  assign n11001 = ~n10812 & ~n10984;
  assign n11002 = n10987 & n11001;
  assign n11003 = ~n11000 & ~n11002;
  assign n11004 = n10288 & ~n11003;
  assign n11005 = n10987 & n10999;
  assign n11006 = n10992 & n11005;
  assign n11007 = ~n9839 & ~n10287;
  assign n11008 = n10988 & n10993;
  assign n11009 = ~n10986 & ~n11008;
  assign n11010 = n11007 & ~n11009;
  assign n11011 = ~n11006 & ~n11010;
  assign n11012 = ~n11004 & n11011;
  assign n11013 = n10989 & n10992;
  assign n11014 = n10985 & n10987;
  assign n11015 = n10459 & n10689;
  assign n11016 = n10988 & n11015;
  assign n11017 = ~n11014 & ~n11016;
  assign n11018 = n11007 & ~n11017;
  assign n11019 = ~n11013 & ~n11018;
  assign n11020 = n9839 & ~n10287;
  assign n11021 = n10999 & n11015;
  assign n11022 = n10812 ^ n10459;
  assign n11023 = n10812 ^ n10689;
  assign n11024 = n11023 ^ n10984;
  assign n11025 = ~n11022 & ~n11024;
  assign n11026 = ~n11021 & ~n11025;
  assign n11027 = n11003 & n11026;
  assign n11028 = ~n10986 & n11027;
  assign n11029 = n11020 & n11028;
  assign n11030 = n10690 & n10999;
  assign n11031 = n11001 & n11015;
  assign n11032 = ~n11030 & ~n11031;
  assign n11033 = n11003 & n11032;
  assign n11034 = ~n9839 & ~n11033;
  assign n11035 = n10690 & n11001;
  assign n11036 = ~n11021 & ~n11035;
  assign n11037 = ~n11016 & n11036;
  assign n11038 = ~n11008 & n11037;
  assign n11039 = n10288 & ~n11038;
  assign n11040 = ~n11034 & ~n11039;
  assign n11041 = ~n11029 & n11040;
  assign n11042 = n11019 & n11041;
  assign n11043 = n11012 & n11042;
  assign n11044 = n10998 & n11043;
  assign n11045 = n11044 ^ n9047;
  assign n11046 = n11045 ^ x562;
  assign n11047 = n9946 ^ x484;
  assign n11048 = n10567 ^ x489;
  assign n11049 = n11047 & n11048;
  assign n11050 = n8565 & ~n10156;
  assign n11051 = n8551 & ~n10162;
  assign n11052 = ~n11050 & ~n11051;
  assign n11053 = n7750 & n10172;
  assign n11054 = n8576 & ~n10177;
  assign n11055 = ~n11053 & ~n11054;
  assign n11056 = n11052 & n11055;
  assign n11057 = n11056 ^ n6166;
  assign n11058 = n11057 ^ x486;
  assign n11059 = n10501 ^ x488;
  assign n11060 = n11058 & n11059;
  assign n11061 = n10352 & ~n10365;
  assign n11062 = n10043 & ~n10060;
  assign n11063 = ~n11061 & ~n11062;
  assign n11064 = n9985 & ~n10051;
  assign n11065 = n10033 & ~n10074;
  assign n11066 = ~n11064 & ~n11065;
  assign n11067 = ~n10079 & n10357;
  assign n11068 = n10038 & ~n11067;
  assign n11069 = n10055 & n10085;
  assign n11070 = n10060 & ~n11069;
  assign n11071 = ~n11068 & ~n11070;
  assign n11072 = n11066 & n11071;
  assign n11073 = n11063 & n11072;
  assign n11074 = n10869 & n11073;
  assign n11075 = n10077 & n11074;
  assign n11076 = n10057 & n11075;
  assign n11077 = ~n10356 & n11076;
  assign n11078 = n11077 ^ n6781;
  assign n11079 = n11078 ^ x487;
  assign n11080 = n10220 ^ x485;
  assign n11081 = ~n11079 & n11080;
  assign n11082 = n11060 & n11081;
  assign n11083 = n11058 & ~n11059;
  assign n11084 = n11079 & n11080;
  assign n11085 = n11083 & n11084;
  assign n11086 = ~n11082 & ~n11085;
  assign n11087 = n11049 & ~n11086;
  assign n11088 = ~n11047 & n11048;
  assign n11089 = ~n11058 & n11059;
  assign n11090 = n11081 & n11089;
  assign n11091 = n11081 & n11083;
  assign n11092 = ~n11090 & ~n11091;
  assign n11093 = n11088 & ~n11092;
  assign n11094 = ~n11087 & ~n11093;
  assign n11095 = ~n11058 & ~n11059;
  assign n11096 = n11084 & n11095;
  assign n11097 = n11049 & n11096;
  assign n11098 = n11079 & ~n11080;
  assign n11099 = n11083 & n11098;
  assign n11100 = ~n11079 & ~n11080;
  assign n11101 = n11089 & n11100;
  assign n11102 = ~n11099 & ~n11101;
  assign n11103 = n11088 & ~n11102;
  assign n11104 = ~n11097 & ~n11103;
  assign n11105 = n11060 & n11098;
  assign n11106 = n11083 & n11100;
  assign n11107 = ~n11105 & ~n11106;
  assign n11108 = n11049 & ~n11107;
  assign n11109 = n11049 & n11090;
  assign n11110 = n11089 & n11098;
  assign n11111 = ~n11106 & ~n11110;
  assign n11112 = n11088 & ~n11111;
  assign n11113 = ~n11109 & ~n11112;
  assign n11114 = n11095 & n11100;
  assign n11115 = n11060 & n11100;
  assign n11116 = ~n11114 & ~n11115;
  assign n11117 = n11047 & ~n11116;
  assign n11118 = n11047 & ~n11048;
  assign n11119 = ~n11082 & ~n11091;
  assign n11120 = n11102 & n11119;
  assign n11121 = n11118 & ~n11120;
  assign n11122 = ~n11117 & ~n11121;
  assign n11123 = n11113 & n11122;
  assign n11124 = ~n11088 & ~n11118;
  assign n11125 = n11060 & n11084;
  assign n11126 = ~n11096 & ~n11125;
  assign n11127 = ~n11124 & ~n11126;
  assign n11128 = ~n11047 & ~n11048;
  assign n11129 = n11079 ^ n11059;
  assign n11130 = n11129 ^ n11080;
  assign n11131 = n11080 ^ n11058;
  assign n11132 = ~n11059 & ~n11131;
  assign n11133 = ~n11130 & n11132;
  assign n11134 = n11133 ^ n11130;
  assign n11135 = n11102 & n11134;
  assign n11136 = n11128 & n11135;
  assign n11137 = ~n11127 & ~n11136;
  assign n11138 = n11123 & n11137;
  assign n11139 = ~n11108 & n11138;
  assign n11140 = n11104 & n11139;
  assign n11141 = n11094 & n11140;
  assign n11142 = n11141 ^ n9249;
  assign n11143 = n11142 ^ x496;
  assign n11144 = n10619 & ~n10637;
  assign n11145 = n10666 & ~n10681;
  assign n11146 = n10639 & ~n11145;
  assign n11147 = n10658 & ~n11146;
  assign n11148 = n10622 & n10630;
  assign n11149 = n10503 & ~n10649;
  assign n11150 = ~n11148 & ~n11149;
  assign n11151 = n10590 ^ n10532;
  assign n11152 = n10634 & n11151;
  assign n11153 = n10639 & n11152;
  assign n11154 = ~n10656 & ~n10661;
  assign n11155 = n10630 & ~n11154;
  assign n11156 = ~n11153 & ~n11155;
  assign n11157 = n10630 & n10648;
  assign n11158 = ~n10532 & n10621;
  assign n11159 = ~n10619 & n11158;
  assign n11160 = ~n11157 & ~n11159;
  assign n11161 = n10639 & n10661;
  assign n11162 = ~n10624 & n10669;
  assign n11163 = ~n11161 & ~n11162;
  assign n11164 = n10619 & ~n10666;
  assign n11165 = n10637 & ~n10641;
  assign n11166 = n10503 & n11165;
  assign n11167 = n11166 ^ n10503;
  assign n11168 = ~n11164 & ~n11167;
  assign n11169 = n11163 & n11168;
  assign n11170 = n11160 & n11169;
  assign n11171 = n11156 & n11170;
  assign n11172 = n11150 & n11171;
  assign n11173 = ~n10685 & n11172;
  assign n11174 = n11147 & n11173;
  assign n11175 = ~n11144 & n11174;
  assign n11176 = n11175 ^ n9276;
  assign n11177 = n11176 ^ x501;
  assign n11178 = n11143 & n11177;
  assign n11179 = n10381 ^ n10347;
  assign n11180 = n10438 & ~n11179;
  assign n11181 = n10422 ^ n10407;
  assign n11182 = ~n10347 & n11181;
  assign n11183 = n11182 ^ n10407;
  assign n11184 = ~n11180 & ~n11183;
  assign n11185 = n10434 & ~n11184;
  assign n11186 = n10382 & n10407;
  assign n11187 = ~n10429 & ~n11186;
  assign n11188 = n10446 & ~n11187;
  assign n11189 = ~n11185 & ~n11188;
  assign n11190 = ~n10381 & n10407;
  assign n11191 = n10382 & n10413;
  assign n11192 = n11191 ^ n10412;
  assign n11193 = ~n11190 & ~n11192;
  assign n11194 = ~n11180 & n11193;
  assign n11195 = n10418 & n11194;
  assign n11196 = n10407 & n10408;
  assign n11197 = ~n10415 & ~n11196;
  assign n11198 = ~n11180 & n11197;
  assign n11199 = ~n10420 & n11198;
  assign n11200 = n10313 & ~n11199;
  assign n11201 = ~n11195 & ~n11200;
  assign n11202 = n11189 & n11201;
  assign n11203 = n10411 & ~n11179;
  assign n11204 = n11202 & ~n11203;
  assign n11205 = n11204 ^ n9368;
  assign n11206 = n11205 ^ x497;
  assign n11207 = ~n10776 & ~n10794;
  assign n11208 = ~n10767 & n11207;
  assign n11209 = n10749 & ~n11208;
  assign n11210 = ~n10691 & n10764;
  assign n11211 = ~n10758 & ~n10795;
  assign n11212 = n10785 & n11211;
  assign n11213 = ~n10752 & n11212;
  assign n11214 = n10693 & ~n11213;
  assign n11215 = n10759 & ~n10784;
  assign n11216 = ~n10782 & n11215;
  assign n11217 = n10754 & ~n11216;
  assign n11218 = ~n10752 & ~n10784;
  assign n11219 = n10789 & n11218;
  assign n11220 = n10749 & ~n11219;
  assign n11221 = ~n11217 & ~n11220;
  assign n11222 = ~n11214 & n11221;
  assign n11223 = ~n10768 & ~n10773;
  assign n11224 = ~n10764 & ~n10777;
  assign n11225 = ~n10794 & n11224;
  assign n11226 = n10789 & n11225;
  assign n11227 = ~n10782 & n11226;
  assign n11228 = ~n10756 & n11227;
  assign n11229 = ~n10747 & n11228;
  assign n11230 = n10763 & ~n11229;
  assign n11231 = ~n11223 & ~n11230;
  assign n11232 = n11222 & n11231;
  assign n11233 = ~n11210 & n11232;
  assign n11234 = ~n11209 & n11233;
  assign n11235 = ~n10762 & n11234;
  assign n11236 = ~n10748 & n11235;
  assign n11237 = n11236 ^ n9403;
  assign n11238 = n11237 ^ x499;
  assign n11239 = n11206 & n11238;
  assign n11240 = n10232 & n10271;
  assign n11241 = n10222 & ~n10259;
  assign n11242 = ~n10244 & n10272;
  assign n11243 = ~n10235 & n11242;
  assign n11244 = n10257 & ~n11243;
  assign n11245 = n10263 & ~n10265;
  assign n11246 = ~n10241 & n11245;
  assign n11247 = ~n10147 & n11246;
  assign n11248 = n10232 & ~n11247;
  assign n11249 = n10251 & n10277;
  assign n11250 = ~n10246 & n11249;
  assign n11251 = ~n10264 & n11250;
  assign n11252 = n10224 & ~n11251;
  assign n11253 = ~n10239 & ~n10264;
  assign n11254 = ~n10227 & n11253;
  assign n11255 = ~n10257 & n11254;
  assign n11256 = ~n10261 & ~n10265;
  assign n11257 = ~n10249 & n11256;
  assign n11258 = ~n10222 & n11257;
  assign n11259 = ~n11255 & ~n11258;
  assign n11260 = ~n10258 & ~n11259;
  assign n11261 = ~n10221 & ~n11260;
  assign n11262 = ~n11252 & ~n11261;
  assign n11263 = ~n11248 & n11262;
  assign n11264 = ~n11244 & n11263;
  assign n11265 = ~n11241 & n11264;
  assign n11266 = n10237 & n11265;
  assign n11267 = n10229 & n11266;
  assign n11268 = ~n11240 & n11267;
  assign n11269 = n11268 ^ n9333;
  assign n11270 = n11269 ^ x500;
  assign n11271 = ~n10947 & ~n10962;
  assign n11272 = n10926 & ~n11271;
  assign n11273 = n10843 & n10939;
  assign n11274 = ~n10924 & n10937;
  assign n11275 = ~n11273 & ~n11274;
  assign n11276 = ~n11272 & n11275;
  assign n11277 = n10843 & n10953;
  assign n11278 = n10945 & n10969;
  assign n11279 = ~n11277 & ~n11278;
  assign n11280 = n10926 & n10954;
  assign n11281 = ~n10947 & ~n10949;
  assign n11282 = n10937 & ~n11281;
  assign n11283 = ~n11280 & ~n11282;
  assign n11284 = ~n10923 & ~n10949;
  assign n11285 = n10945 & ~n11284;
  assign n11286 = ~n10930 & ~n10935;
  assign n11287 = ~n10843 & n11286;
  assign n11288 = ~n10939 & n11287;
  assign n11289 = ~n10937 & n10964;
  assign n11290 = ~n11288 & ~n11289;
  assign n11291 = ~n10954 & ~n11290;
  assign n11292 = n10952 & ~n11291;
  assign n11293 = ~n11285 & ~n11292;
  assign n11294 = n10843 & ~n10931;
  assign n11295 = ~n10935 & ~n10957;
  assign n11296 = n10926 & n10940;
  assign n11297 = ~n10940 & ~n10945;
  assign n11298 = n10953 & ~n11297;
  assign n11299 = ~n11296 & ~n11298;
  assign n11300 = n11295 & n11299;
  assign n11301 = ~n10928 & n11300;
  assign n11302 = ~n10961 & n11301;
  assign n11303 = ~n10952 & ~n11302;
  assign n11304 = ~n11294 & ~n11303;
  assign n11305 = n11293 & n11304;
  assign n11306 = n11283 & n11305;
  assign n11307 = n11279 & n11306;
  assign n11308 = n11276 & n11307;
  assign n11309 = n11308 ^ n9303;
  assign n11310 = n11309 ^ x498;
  assign n11311 = n11270 & n11310;
  assign n11312 = n11239 & n11311;
  assign n11313 = n11178 & n11312;
  assign n11314 = n11143 & ~n11177;
  assign n11315 = n11206 & n11311;
  assign n11316 = ~n11238 & n11315;
  assign n11317 = n11314 & n11316;
  assign n11318 = ~n11313 & ~n11317;
  assign n11319 = n11206 & ~n11270;
  assign n11320 = ~n11238 & ~n11310;
  assign n11321 = n11319 & n11320;
  assign n11322 = n11314 & n11321;
  assign n11323 = n11178 & n11321;
  assign n11324 = ~n11143 & n11177;
  assign n11325 = ~n11206 & ~n11270;
  assign n11326 = n11238 & n11325;
  assign n11327 = ~n11310 & n11326;
  assign n11328 = ~n11206 & n11311;
  assign n11329 = n11238 & n11328;
  assign n11330 = ~n11327 & ~n11329;
  assign n11331 = n11324 & ~n11330;
  assign n11332 = ~n11323 & ~n11331;
  assign n11333 = ~n11238 & n11325;
  assign n11334 = n11310 & n11333;
  assign n11335 = ~n11329 & ~n11334;
  assign n11336 = n11178 & ~n11335;
  assign n11337 = ~n11143 & ~n11177;
  assign n11338 = ~n11206 & n11270;
  assign n11339 = n11320 & n11338;
  assign n11340 = ~n11334 & ~n11339;
  assign n11341 = n11337 & ~n11340;
  assign n11342 = ~n11336 & ~n11341;
  assign n11343 = ~n11238 & n11319;
  assign n11344 = n11310 & n11343;
  assign n11345 = n11270 ^ n11238;
  assign n11346 = n11310 ^ n11270;
  assign n11347 = n11345 & n11346;
  assign n11348 = n11206 & n11347;
  assign n11349 = ~n11344 & ~n11348;
  assign n11350 = n11324 & ~n11349;
  assign n11351 = n11239 & ~n11270;
  assign n11352 = ~n11310 & n11351;
  assign n11353 = n11337 & n11352;
  assign n11354 = ~n11238 & n11328;
  assign n11355 = n11324 & n11354;
  assign n11356 = ~n11353 & ~n11355;
  assign n11357 = ~n11177 & n11312;
  assign n11358 = n11310 & n11326;
  assign n11359 = ~n11344 & ~n11358;
  assign n11360 = ~n11354 & n11359;
  assign n11361 = n11337 & ~n11360;
  assign n11362 = ~n11357 & ~n11361;
  assign n11363 = ~n11178 & ~n11337;
  assign n11364 = n11239 & n11270;
  assign n11365 = ~n11310 & n11364;
  assign n11366 = ~n11363 & n11365;
  assign n11367 = ~n11316 & ~n11352;
  assign n11368 = n11324 & ~n11367;
  assign n11369 = n11310 & n11351;
  assign n11370 = n11320 & n11325;
  assign n11371 = ~n11339 & ~n11370;
  assign n11372 = ~n11314 & n11371;
  assign n11373 = n11238 & n11338;
  assign n11374 = ~n11310 & n11373;
  assign n11375 = ~n11178 & ~n11354;
  assign n11376 = n11340 & n11375;
  assign n11377 = ~n11374 & n11376;
  assign n11378 = ~n11372 & ~n11377;
  assign n11379 = ~n11369 & ~n11378;
  assign n11380 = n11143 & ~n11379;
  assign n11381 = ~n11368 & ~n11380;
  assign n11382 = ~n11366 & n11381;
  assign n11383 = n11362 & n11382;
  assign n11384 = n11356 & n11383;
  assign n11385 = ~n11350 & n11384;
  assign n11386 = n11342 & n11385;
  assign n11387 = n11332 & n11386;
  assign n11388 = ~n11322 & n11387;
  assign n11389 = n11318 & n11388;
  assign n11390 = n11389 ^ n10311;
  assign n11391 = n11390 ^ x567;
  assign n11392 = n11046 & ~n11391;
  assign n11857 = n9807 & n9824;
  assign n11858 = ~n9812 & ~n9818;
  assign n11859 = n9788 & ~n11858;
  assign n11860 = n9798 & n9810;
  assign n11861 = ~n9815 & ~n11860;
  assign n11862 = ~n9793 & n11861;
  assign n11863 = n9795 & ~n11862;
  assign n11864 = ~n11859 & ~n11863;
  assign n11865 = ~n9472 & ~n9804;
  assign n11866 = n9819 & n11865;
  assign n11867 = n9827 & ~n11866;
  assign n11868 = n9475 & n9807;
  assign n11408 = n9048 & n9810;
  assign n11409 = n9794 & ~n11408;
  assign n11869 = n9788 & ~n11409;
  assign n11412 = n9473 & n9791;
  assign n11870 = ~n9793 & ~n11408;
  assign n11871 = ~n11412 & n11870;
  assign n11872 = n9807 & ~n11871;
  assign n11873 = ~n11869 & ~n11872;
  assign n11874 = ~n9792 & n11861;
  assign n11875 = n9827 & ~n11874;
  assign n11876 = ~n9806 & ~n9824;
  assign n11877 = n11865 & n11876;
  assign n11878 = n9795 & ~n11877;
  assign n11879 = ~n11875 & ~n11878;
  assign n11880 = n11873 & n11879;
  assign n11881 = ~n11868 & n11880;
  assign n11882 = ~n11867 & n11881;
  assign n11883 = n11864 & n11882;
  assign n11884 = ~n9803 & n11883;
  assign n11885 = ~n11857 & n11884;
  assign n11886 = n11885 ^ n8190;
  assign n11887 = n11886 ^ x520;
  assign n11888 = n10639 & n10656;
  assign n11889 = n10619 & ~n10649;
  assign n11890 = ~n11888 & ~n11889;
  assign n11891 = n10622 & ~n10624;
  assign n11892 = n10473 & n10636;
  assign n11893 = n10630 & n10681;
  assign n11894 = ~n10645 & ~n11152;
  assign n11895 = ~n10661 & n11894;
  assign n11896 = n10630 & ~n11895;
  assign n11897 = ~n10654 & ~n10669;
  assign n11898 = ~n10502 & ~n11897;
  assign n11899 = n10532 & n10635;
  assign n11900 = ~n10661 & ~n11899;
  assign n11901 = n10503 & ~n11900;
  assign n11902 = ~n11898 & ~n11901;
  assign n11903 = ~n11896 & n11902;
  assign n11904 = n11150 & n11903;
  assign n11905 = ~n11893 & n11904;
  assign n11906 = ~n11892 & n11905;
  assign n11907 = ~n11891 & n11906;
  assign n11908 = n11890 & n11907;
  assign n11909 = n11147 & n11908;
  assign n11910 = ~n10653 & n11909;
  assign n11911 = ~n10618 & n11910;
  assign n11912 = ~n11144 & n11911;
  assign n11913 = n11912 ^ n9157;
  assign n11914 = n11913 ^ x525;
  assign n11915 = n11887 & ~n11914;
  assign n11916 = ~n10416 & n10446;
  assign n11917 = ~n10431 & n10434;
  assign n11918 = ~n11916 & ~n11917;
  assign n11919 = n10418 & ~n10444;
  assign n11920 = n10313 & ~n10454;
  assign n11921 = ~n11919 & ~n11920;
  assign n11922 = n11918 & n11921;
  assign n11923 = n11922 ^ n9057;
  assign n11924 = n11923 ^ x524;
  assign n11925 = ~n10961 & ~n10970;
  assign n11926 = n10937 & ~n11925;
  assign n11927 = ~n10954 & n11295;
  assign n11928 = n10843 & ~n11927;
  assign n11929 = ~n11926 & ~n11928;
  assign n11930 = n10926 & ~n10971;
  assign n11931 = n10963 & n11281;
  assign n11932 = n10945 & ~n11931;
  assign n11933 = n10941 & n11295;
  assign n11934 = n10945 & ~n11933;
  assign n11778 = n10931 & ~n10935;
  assign n11935 = ~n10953 & n11778;
  assign n11936 = n10926 & ~n11935;
  assign n11937 = ~n11934 & ~n11936;
  assign n11938 = ~n10930 & n10941;
  assign n11939 = ~n10957 & n11938;
  assign n11940 = n10937 & ~n11939;
  assign n11941 = ~n10921 & n11281;
  assign n11942 = ~n10962 & n11941;
  assign n11943 = n10843 & ~n11942;
  assign n11944 = ~n11940 & ~n11943;
  assign n11945 = n11937 & n11944;
  assign n11946 = ~n11932 & n11945;
  assign n11947 = ~n11930 & n11946;
  assign n11948 = n11929 & n11947;
  assign n11949 = n11276 & n11948;
  assign n11950 = n11949 ^ n9690;
  assign n11951 = n11950 ^ x522;
  assign n11952 = ~n11924 & n11951;
  assign n11702 = n10227 & n10257;
  assign n11703 = n10224 & ~n10247;
  assign n11704 = ~n11702 & ~n11703;
  assign n11953 = n10221 & n10249;
  assign n11954 = n10230 & n10257;
  assign n11955 = ~n11953 & ~n11954;
  assign n11956 = n10232 & n10261;
  assign n11957 = ~n10235 & n10267;
  assign n11958 = ~n10230 & n11957;
  assign n11959 = n10224 & ~n11958;
  assign n11960 = ~n11956 & ~n11959;
  assign n11961 = n11955 & n11960;
  assign n11962 = ~n10232 & ~n10257;
  assign n11963 = ~n10266 & ~n11962;
  assign n11964 = ~n10227 & ~n10262;
  assign n11965 = n10222 & ~n11964;
  assign n11966 = ~n10258 & n11962;
  assign n11967 = n10182 & n10259;
  assign n11968 = ~n11966 & ~n11967;
  assign n11969 = ~n10260 & n11968;
  assign n11970 = n10247 & ~n11969;
  assign n11971 = n10221 & ~n10260;
  assign n11972 = ~n10182 & n11971;
  assign n11973 = n11972 ^ n10221;
  assign n11974 = ~n11970 & ~n11973;
  assign n11975 = ~n11965 & ~n11974;
  assign n11976 = ~n11963 & n11975;
  assign n11977 = n11961 & n11976;
  assign n11978 = ~n10243 & n11977;
  assign n11979 = ~n10223 & n11978;
  assign n11980 = n11704 & n11979;
  assign n11981 = ~n11240 & n11980;
  assign n11982 = n11981 ^ n9715;
  assign n11983 = n11982 ^ x523;
  assign n11431 = n9721 & n9755;
  assign n11432 = n9731 & n9749;
  assign n11433 = ~n11431 & ~n11432;
  assign n11434 = ~n9741 & ~n9759;
  assign n11435 = n9667 & n9729;
  assign n11436 = ~n9666 & n9751;
  assign n11437 = n9731 & ~n10185;
  assign n11438 = ~n11436 & ~n11437;
  assign n11439 = n9734 & n9745;
  assign n11440 = n9721 & ~n11439;
  assign n11441 = ~n9744 & ~n9755;
  assign n11442 = n9665 & ~n11441;
  assign n11443 = ~n11440 & ~n11442;
  assign n11444 = n11438 & n11443;
  assign n11445 = n9667 & n9733;
  assign n11446 = ~n9732 & ~n9742;
  assign n11447 = n9726 & ~n11446;
  assign n11448 = ~n9757 & n10199;
  assign n11449 = ~n9750 & n11448;
  assign n11450 = ~n10197 & ~n11449;
  assign n11451 = ~n11447 & ~n11450;
  assign n11452 = ~n11445 & n11451;
  assign n11453 = n11444 & n11452;
  assign n11454 = ~n11435 & n11453;
  assign n11455 = ~n11434 & n11454;
  assign n11456 = n11433 & n11455;
  assign n11457 = n10188 & n11456;
  assign n11458 = ~n9720 & n11457;
  assign n11459 = n11458 ^ n7604;
  assign n11460 = n11459 ^ x451;
  assign n11461 = n10841 ^ x452;
  assign n11498 = ~n11460 & n11461;
  assign n11463 = n10472 ^ x449;
  assign n11464 = ~n9600 & ~n9621;
  assign n11465 = n9603 & ~n11464;
  assign n11466 = ~n9627 & n9639;
  assign n11467 = ~n9477 & ~n11466;
  assign n11468 = ~n11465 & ~n11467;
  assign n11469 = n9589 & ~n10726;
  assign n11470 = ~n9623 & ~n9649;
  assign n11471 = n9613 & ~n11470;
  assign n11472 = n9607 & ~n9636;
  assign n11473 = n9558 ^ n9529;
  assign n11474 = n9528 & ~n9585;
  assign n11475 = ~n11473 & n11474;
  assign n11476 = n11475 ^ n11473;
  assign n11477 = n9505 & ~n11476;
  assign n11478 = ~n11472 & ~n11477;
  assign n11479 = ~n11471 & n11478;
  assign n11480 = ~n11469 & n11479;
  assign n11481 = n11468 & n11480;
  assign n11482 = n9635 & n11481;
  assign n11483 = ~n10721 & n11482;
  assign n11484 = n10477 & n11483;
  assign n11485 = n9597 & n11484;
  assign n11486 = n11485 ^ n7566;
  assign n11487 = n11486 ^ x450;
  assign n11509 = ~n11463 & ~n11487;
  assign n11510 = n11498 & n11509;
  assign n11490 = n10589 ^ x448;
  assign n11491 = n10892 ^ x453;
  assign n11523 = n11490 & ~n11491;
  assign n11646 = n11510 & n11523;
  assign n11494 = ~n11490 & ~n11491;
  assign n11462 = n11460 & n11461;
  assign n11545 = n11462 & n11509;
  assign n11647 = n11494 & n11545;
  assign n11648 = ~n11646 & ~n11647;
  assign n11488 = ~n11463 & n11487;
  assign n11489 = n11462 & n11488;
  assign n11524 = n11489 & n11523;
  assign n11492 = ~n11490 & n11491;
  assign n11504 = n11463 & ~n11487;
  assign n11525 = n11462 & n11504;
  assign n11495 = n11463 & n11487;
  assign n11507 = n11460 & ~n11461;
  assign n11526 = n11495 & n11507;
  assign n11527 = ~n11525 & ~n11526;
  assign n11528 = n11492 & ~n11527;
  assign n11529 = ~n11524 & ~n11528;
  assign n11503 = n11490 & n11491;
  assign n11530 = n11488 & n11498;
  assign n11531 = n11503 & n11530;
  assign n11496 = ~n11460 & ~n11461;
  assign n11497 = n11495 & n11496;
  assign n11532 = n11492 & n11497;
  assign n11533 = ~n11531 & ~n11532;
  assign n11984 = n11489 & n11494;
  assign n11985 = n11533 & ~n11984;
  assign n11519 = n11462 & n11495;
  assign n11986 = n11492 & n11519;
  assign n11987 = n11490 & n11545;
  assign n11988 = ~n11986 & ~n11987;
  assign n11511 = n11507 & n11509;
  assign n11989 = n11503 & n11511;
  assign n11535 = n11488 & n11496;
  assign n11990 = n11494 & n11535;
  assign n11991 = ~n11989 & ~n11990;
  assign n11508 = n11488 & n11507;
  assign n11518 = ~n11494 & ~n11503;
  assign n11992 = n11518 & ~n11523;
  assign n11993 = n11508 & ~n11992;
  assign n11493 = n11489 & n11492;
  assign n11516 = n11504 & n11507;
  assign n11499 = n11495 & n11498;
  assign n11505 = n11498 & n11504;
  assign n11653 = ~n11499 & ~n11505;
  assign n11994 = ~n11497 & ~n11523;
  assign n11995 = n11653 & n11994;
  assign n11996 = ~n11516 & n11995;
  assign n11656 = ~n11516 & ~n11519;
  assign n11997 = ~n11499 & n11656;
  assign n11998 = ~n11497 & n11997;
  assign n11999 = n11523 & ~n11998;
  assign n12000 = ~n11503 & ~n11999;
  assign n12001 = ~n11996 & ~n12000;
  assign n11520 = n11496 & n11504;
  assign n12002 = ~n11492 & ~n11520;
  assign n11542 = n11496 & n11509;
  assign n11650 = ~n11530 & ~n11542;
  assign n12003 = ~n11520 & n11650;
  assign n12004 = ~n12002 & ~n12003;
  assign n12005 = ~n11526 & n11653;
  assign n12006 = ~n11494 & n12003;
  assign n12007 = ~n12005 & ~n12006;
  assign n12008 = ~n12004 & ~n12007;
  assign n12009 = ~n11490 & ~n12008;
  assign n12010 = ~n12001 & ~n12009;
  assign n12011 = ~n11493 & n12010;
  assign n12012 = ~n11993 & n12011;
  assign n12013 = n11991 & n12012;
  assign n12014 = n11988 & n12013;
  assign n12015 = n11985 & n12014;
  assign n12016 = n11529 & n12015;
  assign n12017 = n11648 & n12016;
  assign n12018 = n12017 ^ n7748;
  assign n12019 = n12018 ^ x521;
  assign n12020 = ~n11983 & n12019;
  assign n12021 = n11952 & n12020;
  assign n12022 = n11915 & n12021;
  assign n12023 = n11887 & n11914;
  assign n12024 = ~n11983 & ~n12019;
  assign n12025 = n11952 & n12024;
  assign n12026 = n12023 & n12025;
  assign n12027 = ~n11887 & n11914;
  assign n12028 = n11924 & n11951;
  assign n12029 = n12024 & n12028;
  assign n12030 = n12027 & n12029;
  assign n12031 = n11924 & ~n11951;
  assign n12032 = n11983 & ~n12019;
  assign n12033 = n12031 & n12032;
  assign n12034 = n11915 & n12033;
  assign n12035 = ~n12030 & ~n12034;
  assign n12036 = ~n12026 & n12035;
  assign n12037 = ~n12022 & n12036;
  assign n12038 = n11983 & n12019;
  assign n12039 = n12031 & n12038;
  assign n12040 = n12020 & n12031;
  assign n12041 = n11952 & n12038;
  assign n12042 = ~n12040 & ~n12041;
  assign n12043 = ~n12039 & n12042;
  assign n12044 = n11915 & ~n12043;
  assign n12045 = n11952 & n12032;
  assign n12046 = ~n11924 & ~n11951;
  assign n12047 = n12024 & n12046;
  assign n12048 = ~n12045 & ~n12047;
  assign n12049 = ~n12029 & n12048;
  assign n12050 = n11915 & ~n12049;
  assign n12051 = n12028 & n12032;
  assign n12052 = n12024 & n12031;
  assign n12053 = ~n12047 & ~n12052;
  assign n12054 = n12038 ^ n12020;
  assign n12055 = n11951 & n12054;
  assign n12056 = ~n11924 & n12055;
  assign n12057 = n12056 ^ n12038;
  assign n12058 = n12053 & ~n12057;
  assign n12059 = ~n12051 & n12058;
  assign n12060 = n12027 & ~n12059;
  assign n12061 = ~n12050 & ~n12060;
  assign n12062 = ~n11887 & ~n11914;
  assign n12063 = n12032 & n12046;
  assign n12064 = n12038 & n12046;
  assign n12065 = ~n12025 & ~n12051;
  assign n12066 = ~n12064 & n12065;
  assign n12067 = ~n12063 & n12066;
  assign n12068 = n12062 & ~n12067;
  assign n12069 = n12020 & n12046;
  assign n12070 = n12020 & n12028;
  assign n12071 = n12042 & ~n12070;
  assign n12072 = ~n12069 & n12071;
  assign n12073 = n12062 & ~n12072;
  assign n12074 = ~n12051 & ~n12063;
  assign n12075 = ~n12045 & ~n12052;
  assign n12076 = ~n12070 & n12075;
  assign n12077 = ~n12069 & n12076;
  assign n12078 = n12074 & n12077;
  assign n12079 = ~n12064 & n12078;
  assign n12080 = n12023 & ~n12079;
  assign n12081 = ~n12073 & ~n12080;
  assign n12082 = ~n12068 & n12081;
  assign n12083 = n12061 & n12082;
  assign n12084 = ~n12044 & n12083;
  assign n12085 = n12037 & n12084;
  assign n12086 = n12085 ^ n10405;
  assign n12087 = n12086 ^ x564;
  assign n11393 = n11205 ^ x543;
  assign n11394 = n10983 ^ x538;
  assign n11395 = ~n11393 & n11394;
  assign n11396 = n9788 & ~n9819;
  assign n11397 = n9810 & ~n9814;
  assign n11398 = n9795 & n11397;
  assign n11399 = ~n11396 & ~n11398;
  assign n11400 = n9476 & ~n9799;
  assign n11401 = n9827 & ~n11400;
  assign n11402 = ~n9800 & ~n9812;
  assign n11403 = ~n9804 & n11402;
  assign n11404 = n9807 & ~n11403;
  assign n11405 = ~n9792 & n9813;
  assign n11406 = ~n9824 & n11405;
  assign n11407 = n9788 & ~n11406;
  assign n11410 = n9807 & ~n11409;
  assign n11411 = ~n11407 & ~n11410;
  assign n11413 = ~n9800 & ~n11397;
  assign n11414 = ~n11412 & n11413;
  assign n11415 = n9827 & ~n11414;
  assign n11416 = n9476 & n9819;
  assign n11417 = n9795 & ~n11416;
  assign n11418 = ~n11415 & ~n11417;
  assign n11419 = n11411 & n11418;
  assign n11420 = ~n11404 & n11419;
  assign n11421 = ~n11401 & n11420;
  assign n11422 = n11399 & n11421;
  assign n11423 = n9797 & n11422;
  assign n11424 = ~n9818 & n11423;
  assign n11425 = n11424 ^ n10007;
  assign n11426 = n11425 ^ x540;
  assign n11427 = n10286 ^ x539;
  assign n11428 = n11142 ^ x542;
  assign n11429 = n11427 & n11428;
  assign n11430 = n11426 & n11429;
  assign n11500 = ~n11497 & ~n11499;
  assign n11501 = n11494 & ~n11500;
  assign n11502 = ~n11493 & ~n11501;
  assign n11506 = n11503 & n11505;
  assign n11512 = ~n11510 & ~n11511;
  assign n11513 = ~n11508 & n11512;
  assign n11514 = n11492 & ~n11513;
  assign n11515 = ~n11506 & ~n11514;
  assign n11517 = n11490 & n11516;
  assign n11521 = ~n11519 & ~n11520;
  assign n11522 = ~n11518 & ~n11521;
  assign n11534 = n11492 & n11499;
  assign n11536 = ~n11520 & ~n11535;
  assign n11537 = ~n11497 & ~n11510;
  assign n11538 = n11536 & n11537;
  assign n11539 = n11527 & n11538;
  assign n11540 = n11523 & ~n11539;
  assign n11541 = ~n11534 & ~n11540;
  assign n11543 = ~n11489 & ~n11542;
  assign n11544 = ~n11494 & n11543;
  assign n11546 = ~n11511 & ~n11530;
  assign n11547 = ~n11545 & n11546;
  assign n11548 = ~n11503 & n11547;
  assign n11549 = ~n11544 & ~n11548;
  assign n11550 = ~n11508 & ~n11549;
  assign n11551 = ~n11518 & ~n11550;
  assign n11552 = n11541 & ~n11551;
  assign n11553 = n11533 & n11552;
  assign n11554 = n11529 & n11553;
  assign n11555 = ~n11522 & n11554;
  assign n11556 = ~n11517 & n11555;
  assign n11557 = n11515 & n11556;
  assign n11558 = n11502 & n11557;
  assign n11559 = n11558 ^ n10027;
  assign n11560 = n11559 ^ x541;
  assign n11561 = n11430 & n11560;
  assign n11562 = n11395 & n11561;
  assign n11563 = n11393 & ~n11394;
  assign n11564 = n11426 & ~n11427;
  assign n11565 = n11428 & n11564;
  assign n11566 = n11560 & n11565;
  assign n11567 = n11563 & n11566;
  assign n11568 = ~n11562 & ~n11567;
  assign n11569 = ~n11426 & n11429;
  assign n11570 = n11560 & n11569;
  assign n11571 = n11395 & n11570;
  assign n11572 = n11426 & ~n11560;
  assign n11573 = ~n11427 & n11572;
  assign n11574 = ~n11428 & n11573;
  assign n11575 = n11563 & n11574;
  assign n11576 = ~n11571 & ~n11575;
  assign n11577 = n11568 & n11576;
  assign n11578 = ~n11393 & ~n11394;
  assign n11579 = ~n11560 & n11569;
  assign n11580 = n11578 & n11579;
  assign n11581 = ~n11428 & n11560;
  assign n11582 = n11427 & n11581;
  assign n11583 = n11426 & n11582;
  assign n11584 = n11394 & n11583;
  assign n11585 = ~n11580 & ~n11584;
  assign n11586 = ~n11426 & ~n11427;
  assign n11587 = n11428 & n11586;
  assign n11588 = n11560 & n11587;
  assign n11589 = n11564 & n11581;
  assign n11590 = ~n11588 & ~n11589;
  assign n11591 = n11563 & ~n11590;
  assign n11592 = n11393 & n11394;
  assign n11593 = n11427 & n11572;
  assign n11594 = ~n11428 & n11593;
  assign n11595 = n11592 & n11594;
  assign n11596 = n11581 & n11586;
  assign n11597 = ~n11566 & ~n11596;
  assign n11598 = n11592 & ~n11597;
  assign n11599 = n11394 ^ n11393;
  assign n11600 = ~n11426 & n11582;
  assign n11601 = n11429 & n11572;
  assign n11602 = ~n11600 & ~n11601;
  assign n11603 = ~n11599 & ~n11602;
  assign n11604 = n11560 ^ n11426;
  assign n11605 = ~n11427 & n11604;
  assign n11606 = n11395 & n11605;
  assign n11607 = ~n11603 & ~n11606;
  assign n11608 = ~n11426 & n11427;
  assign n11609 = ~n11428 & n11608;
  assign n11610 = ~n11560 & n11609;
  assign n11611 = ~n11393 & n11610;
  assign n11612 = ~n11566 & ~n11574;
  assign n11613 = n11590 & n11612;
  assign n11614 = n11578 & ~n11613;
  assign n11615 = ~n11560 & n11587;
  assign n11616 = ~n11428 & n11586;
  assign n11617 = ~n11560 & n11616;
  assign n11618 = ~n11615 & ~n11617;
  assign n11619 = n11592 & ~n11618;
  assign n11620 = ~n11601 & ~n11610;
  assign n11621 = ~n11561 & n11620;
  assign n11622 = ~n11579 & n11621;
  assign n11623 = n11563 & ~n11622;
  assign n11624 = ~n11619 & ~n11623;
  assign n11625 = ~n11614 & n11624;
  assign n11626 = ~n11611 & n11625;
  assign n11627 = n11607 & n11626;
  assign n11628 = ~n11598 & n11627;
  assign n11629 = ~n11595 & n11628;
  assign n11630 = ~n11591 & n11629;
  assign n11631 = n11585 & n11630;
  assign n11632 = n11577 & n11631;
  assign n11633 = n11632 ^ n10380;
  assign n11634 = n11633 ^ x565;
  assign n11635 = n10312 & n11203;
  assign n11636 = n10446 & n11199;
  assign n11637 = ~n11635 & ~n11636;
  assign n11638 = n10313 & ~n11187;
  assign n11639 = n10434 & ~n11194;
  assign n11640 = n10418 & ~n11184;
  assign n11641 = ~n11639 & ~n11640;
  assign n11642 = ~n11638 & n11641;
  assign n11643 = n11637 & n11642;
  assign n11644 = n11643 ^ n9877;
  assign n11645 = n11644 ^ x510;
  assign n11649 = n11490 & n11508;
  assign n11651 = n11523 & ~n11650;
  assign n11652 = ~n11649 & ~n11651;
  assign n11654 = n11492 & ~n11653;
  assign n11655 = ~n11518 & ~n11536;
  assign n11657 = n11537 & n11656;
  assign n11658 = n11494 & ~n11657;
  assign n11659 = ~n11542 & ~n11545;
  assign n11660 = n11546 & n11659;
  assign n11661 = n11492 & ~n11660;
  assign n11662 = ~n11658 & ~n11661;
  assign n11663 = ~n11519 & ~n11525;
  assign n11664 = ~n11497 & n11663;
  assign n11665 = n11523 & ~n11664;
  assign n11666 = ~n11516 & ~n11545;
  assign n11667 = ~n11489 & n11666;
  assign n11668 = ~n11499 & n11667;
  assign n11669 = n11503 & ~n11668;
  assign n11670 = ~n11665 & ~n11669;
  assign n11671 = n11662 & n11670;
  assign n11672 = ~n11655 & n11671;
  assign n11673 = ~n11654 & n11672;
  assign n11674 = n11652 & n11673;
  assign n11675 = ~n11493 & n11674;
  assign n11676 = n11648 & n11675;
  assign n11677 = ~n11526 & n11676;
  assign n11678 = n11677 ^ n9503;
  assign n11679 = n11678 ^ x509;
  assign n11680 = ~n11645 & n11679;
  assign n11681 = ~n11082 & n11126;
  assign n11682 = n11128 & ~n11681;
  assign n11683 = ~n11085 & ~n11105;
  assign n11684 = n11088 & ~n11683;
  assign n11685 = ~n11682 & ~n11684;
  assign n11686 = n11049 & ~n11111;
  assign n11687 = n11081 & n11095;
  assign n11688 = n11102 & ~n11687;
  assign n11689 = n11124 & ~n11688;
  assign n11690 = ~n11686 & ~n11689;
  assign n11691 = n11685 & n11690;
  assign n11692 = n11095 & n11098;
  assign n11693 = ~n11115 & ~n11692;
  assign n11694 = ~n11047 & ~n11693;
  assign n11695 = n11118 & n11135;
  assign n11696 = ~n11694 & ~n11695;
  assign n11697 = n11691 & n11696;
  assign n11698 = n11104 & n11697;
  assign n11699 = n11094 & n11698;
  assign n11700 = n11699 ^ n7392;
  assign n11701 = n11700 ^ x512;
  assign n11705 = ~n10249 & n10263;
  assign n11706 = n10257 & ~n11705;
  assign n11707 = n10266 & n10276;
  assign n11708 = n10222 & ~n11707;
  assign n11709 = ~n11706 & ~n11708;
  assign n11710 = ~n10265 & n10276;
  assign n11711 = ~n10249 & n11710;
  assign n11712 = n10232 & ~n11711;
  assign n11713 = ~n10258 & ~n10271;
  assign n11714 = n10224 & ~n11713;
  assign n11715 = ~n10147 & n10259;
  assign n11716 = n10257 & ~n11715;
  assign n11717 = ~n10241 & n10266;
  assign n11718 = ~n10227 & n11717;
  assign n11719 = n10224 & ~n11718;
  assign n11720 = ~n11716 & ~n11719;
  assign n11721 = ~n10222 & n10251;
  assign n11722 = ~n10250 & n10272;
  assign n11723 = ~n10232 & n11722;
  assign n11724 = ~n11721 & ~n11723;
  assign n11725 = ~n10258 & ~n11724;
  assign n11726 = ~n10182 & ~n11725;
  assign n11727 = n11720 & ~n11726;
  assign n11728 = ~n11240 & n11727;
  assign n11729 = ~n11714 & n11728;
  assign n11730 = ~n11712 & n11729;
  assign n11731 = n11709 & n11730;
  assign n11732 = n11704 & n11731;
  assign n11733 = n11732 ^ n9863;
  assign n11734 = n11733 ^ x511;
  assign n11735 = n11701 & n11734;
  assign n11736 = n11680 & n11735;
  assign n11737 = ~n10758 & ~n10782;
  assign n11738 = ~n10788 & n11737;
  assign n11739 = n10749 & ~n11738;
  assign n11740 = ~n10795 & n11224;
  assign n11741 = ~n10767 & n11740;
  assign n11742 = n10763 & ~n11741;
  assign n11743 = n10754 & ~n10785;
  assign n11744 = ~n10756 & n11218;
  assign n11745 = n10693 & ~n11744;
  assign n11746 = ~n10772 & n10786;
  assign n11747 = n10763 & ~n11746;
  assign n11748 = ~n11745 & ~n11747;
  assign n11749 = ~n11743 & n11748;
  assign n11750 = n10768 & ~n10794;
  assign n11751 = ~n10747 & n11750;
  assign n11752 = n10749 & ~n11751;
  assign n11753 = ~n10777 & n10798;
  assign n11754 = ~n10788 & n11225;
  assign n11755 = ~n10693 & n11754;
  assign n11756 = ~n11753 & ~n11755;
  assign n11757 = ~n10773 & n11756;
  assign n11758 = ~n11752 & ~n11757;
  assign n11759 = n11749 & n11758;
  assign n11760 = ~n11742 & n11759;
  assign n11761 = ~n11739 & n11760;
  assign n11762 = n10761 & n11761;
  assign n11763 = ~n10748 & n11762;
  assign n11764 = n11763 ^ n9584;
  assign n11765 = n11764 ^ x508;
  assign n11766 = n10941 & ~n10961;
  assign n11767 = n10926 & ~n11766;
  assign n11768 = ~n10969 & n11286;
  assign n11769 = ~n10962 & n11768;
  assign n11770 = n10843 & ~n11769;
  assign n11771 = ~n11767 & ~n11770;
  assign n11772 = n10937 & ~n11271;
  assign n11773 = ~n10970 & n11281;
  assign n11774 = ~n10952 & ~n11773;
  assign n11775 = ~n10928 & n11297;
  assign n11776 = ~n10957 & n11775;
  assign n11777 = ~n10954 & n11776;
  assign n11779 = ~n10939 & n11778;
  assign n11780 = ~n10937 & n11779;
  assign n11781 = ~n11777 & ~n11780;
  assign n11782 = n10842 & n11781;
  assign n11783 = ~n11774 & ~n11782;
  assign n11784 = ~n11772 & n11783;
  assign n11785 = n11771 & n11784;
  assign n11786 = n11279 & n11785;
  assign n11787 = n10933 & n11786;
  assign n11788 = n11275 & n11787;
  assign n11789 = n11788 ^ n8035;
  assign n11790 = n11789 ^ x513;
  assign n11791 = ~n11765 & n11790;
  assign n11792 = n11736 & n11791;
  assign n11793 = n11765 & n11790;
  assign n11794 = ~n11645 & ~n11679;
  assign n11795 = n11735 & n11794;
  assign n11796 = n11793 & n11795;
  assign n11797 = ~n11792 & ~n11796;
  assign n11798 = n11765 & ~n11790;
  assign n11799 = n11736 & n11798;
  assign n11800 = ~n11701 & ~n11734;
  assign n11801 = n11794 & n11800;
  assign n11802 = n11645 & ~n11679;
  assign n11803 = n11735 & n11802;
  assign n11804 = ~n11801 & ~n11803;
  assign n11805 = n11793 & ~n11804;
  assign n11806 = ~n11799 & ~n11805;
  assign n11807 = ~n11701 & n11734;
  assign n11808 = n11802 & n11807;
  assign n11809 = n11793 & n11808;
  assign n11810 = n11645 & n11679;
  assign n11811 = n11735 & n11810;
  assign n11812 = ~n11791 & ~n11798;
  assign n11813 = n11811 & ~n11812;
  assign n11814 = ~n11809 & ~n11813;
  assign n11815 = n11800 & n11810;
  assign n11816 = n11701 & ~n11734;
  assign n11817 = n11680 & n11816;
  assign n11818 = ~n11815 & ~n11817;
  assign n11819 = n11791 & ~n11818;
  assign n11820 = n11810 & n11816;
  assign n11821 = ~n11815 & ~n11820;
  assign n11822 = n11798 & ~n11821;
  assign n11823 = n11800 & n11802;
  assign n11824 = ~n11765 & ~n11790;
  assign n11825 = n11823 & n11824;
  assign n11826 = ~n11795 & ~n11803;
  assign n11827 = n11680 & ~n11701;
  assign n11828 = ~n11820 & ~n11827;
  assign n11829 = n11826 & n11828;
  assign n11830 = ~n11817 & n11829;
  assign n11831 = ~n11808 & n11830;
  assign n11832 = n11824 & ~n11831;
  assign n11833 = n11802 & n11816;
  assign n11834 = n11794 & n11816;
  assign n11835 = n11794 & n11807;
  assign n11836 = ~n11834 & ~n11835;
  assign n11837 = ~n11833 & n11836;
  assign n11838 = ~n11801 & n11837;
  assign n11839 = n11798 & ~n11838;
  assign n11840 = ~n11815 & n11828;
  assign n11841 = n11793 & ~n11840;
  assign n11842 = n11807 & n11810;
  assign n11843 = ~n11823 & n11836;
  assign n11844 = ~n11842 & n11843;
  assign n11845 = n11791 & ~n11844;
  assign n11846 = ~n11841 & ~n11845;
  assign n11847 = ~n11839 & n11846;
  assign n11848 = ~n11832 & n11847;
  assign n11849 = ~n11825 & n11848;
  assign n11850 = ~n11822 & n11849;
  assign n11851 = ~n11819 & n11850;
  assign n11852 = n11814 & n11851;
  assign n11853 = n11806 & n11852;
  assign n11854 = n11797 & n11853;
  assign n11855 = n11854 ^ n10345;
  assign n11856 = n11855 ^ x566;
  assign n12227 = n11634 & n11856;
  assign n12228 = n12087 & n12227;
  assign n12089 = n11678 ^ x507;
  assign n12090 = n11269 ^ x502;
  assign n12091 = n12089 & ~n12090;
  assign n12092 = n11764 ^ x506;
  assign n12093 = n11084 & n11089;
  assign n12094 = n11049 & n12093;
  assign n12095 = ~n11101 & ~n11106;
  assign n12096 = n11128 & ~n12095;
  assign n12097 = ~n12094 & ~n12096;
  assign n12098 = n11047 & n11085;
  assign n12099 = n11124 & n11687;
  assign n12100 = ~n12098 & ~n12099;
  assign n12101 = n11105 & n11128;
  assign n12102 = n11088 & n11096;
  assign n12103 = ~n11091 & ~n12093;
  assign n12104 = n11126 & n12103;
  assign n12105 = n11128 & ~n12104;
  assign n12106 = ~n11101 & ~n11692;
  assign n12107 = n11049 & ~n12106;
  assign n12108 = ~n12105 & ~n12107;
  assign n12109 = ~n11082 & ~n11090;
  assign n12110 = ~n11099 & n11693;
  assign n12111 = n12109 & n12110;
  assign n12112 = ~n11110 & n12111;
  assign n12113 = ~n11114 & n12112;
  assign n12114 = ~n11124 & ~n12113;
  assign n12115 = n12108 & ~n12114;
  assign n12116 = ~n11108 & n12115;
  assign n12117 = ~n12102 & n12116;
  assign n12118 = ~n12101 & n12117;
  assign n12119 = n12100 & n12118;
  assign n12120 = ~n11109 & n12119;
  assign n12121 = n12097 & n12120;
  assign n12122 = n12121 ^ n9527;
  assign n12123 = n12122 ^ x505;
  assign n12124 = ~n12092 & ~n12123;
  assign n12125 = n11176 ^ x503;
  assign n12126 = n9792 & n9827;
  assign n12127 = n9788 & n9811;
  assign n12128 = ~n12126 & ~n12127;
  assign n12129 = ~n9802 & n11412;
  assign n12130 = ~n9664 & n9812;
  assign n12131 = n9476 & n11876;
  assign n12132 = n9827 & ~n12131;
  assign n12133 = ~n9795 & n11397;
  assign n12134 = ~n12132 & ~n12133;
  assign n12135 = n9470 ^ n8590;
  assign n12136 = n12135 ^ n9227;
  assign n12137 = n12136 ^ n9470;
  assign n12138 = ~n9048 & ~n12137;
  assign n12139 = n12138 ^ n12135;
  assign n12140 = n9795 & n12139;
  assign n12141 = ~n9788 & ~n9824;
  assign n12142 = ~n9472 & ~n11857;
  assign n12143 = ~n12141 & ~n12142;
  assign n12144 = ~n9800 & ~n12143;
  assign n12145 = n9819 & n12144;
  assign n12146 = ~n9802 & ~n12145;
  assign n12147 = ~n12140 & ~n12146;
  assign n12148 = n12134 & n12147;
  assign n12149 = ~n12130 & n12148;
  assign n12150 = ~n12129 & n12149;
  assign n12151 = n12128 & n12150;
  assign n12152 = n12151 ^ n9557;
  assign n12153 = n12152 ^ x504;
  assign n12154 = n12125 & ~n12153;
  assign n12155 = n12124 & n12154;
  assign n12156 = n12091 & n12155;
  assign n12157 = ~n12092 & n12123;
  assign n12158 = n12125 & n12153;
  assign n12159 = n12157 & n12158;
  assign n12160 = n12091 & n12159;
  assign n12161 = n12089 & n12090;
  assign n12162 = n12092 & ~n12123;
  assign n12163 = ~n12125 & ~n12153;
  assign n12164 = n12162 & n12163;
  assign n12165 = n12161 & n12164;
  assign n12166 = ~n12160 & ~n12165;
  assign n12167 = ~n12156 & n12166;
  assign n12168 = n12124 & n12163;
  assign n12169 = n12161 & n12168;
  assign n12170 = n12092 & n12123;
  assign n12171 = ~n12125 & n12153;
  assign n12172 = n12170 & n12171;
  assign n12173 = n12157 & n12163;
  assign n12174 = ~n12172 & ~n12173;
  assign n12175 = n12091 & ~n12174;
  assign n12176 = ~n12169 & ~n12175;
  assign n12177 = ~n12089 & n12090;
  assign n12178 = n12124 & n12158;
  assign n12179 = n12154 & n12162;
  assign n12180 = ~n12178 & ~n12179;
  assign n12181 = n12177 & ~n12180;
  assign n12182 = n12154 & n12170;
  assign n12183 = ~n12159 & ~n12182;
  assign n12184 = n12161 & ~n12183;
  assign n12185 = ~n12181 & ~n12184;
  assign n12186 = ~n12168 & n12174;
  assign n12187 = n12177 & ~n12186;
  assign n12188 = ~n12089 & ~n12090;
  assign n12189 = ~n12159 & ~n12179;
  assign n12190 = n12188 & ~n12189;
  assign n12191 = n12162 & n12171;
  assign n12192 = n12158 & n12162;
  assign n12193 = n12124 & n12171;
  assign n12194 = ~n12192 & ~n12193;
  assign n12195 = ~n12182 & n12194;
  assign n12196 = ~n12191 & n12195;
  assign n12197 = n12091 & ~n12196;
  assign n12198 = n12163 & n12170;
  assign n12199 = ~n12193 & ~n12198;
  assign n12200 = n12161 & ~n12199;
  assign n12201 = n12090 ^ n12089;
  assign n12202 = n12154 & n12157;
  assign n12203 = ~n12192 & ~n12202;
  assign n12204 = ~n12201 & ~n12203;
  assign n12205 = n12158 & n12170;
  assign n12206 = ~n12202 & ~n12205;
  assign n12207 = ~n12191 & n12206;
  assign n12208 = n12177 & ~n12207;
  assign n12209 = n12157 & n12171;
  assign n12210 = ~n12198 & ~n12209;
  assign n12211 = ~n12168 & n12210;
  assign n12212 = ~n12164 & n12211;
  assign n12213 = n12188 & ~n12212;
  assign n12214 = ~n12208 & ~n12213;
  assign n12215 = ~n12204 & n12214;
  assign n12216 = ~n12200 & n12215;
  assign n12217 = ~n12197 & n12216;
  assign n12218 = ~n12190 & n12217;
  assign n12219 = ~n12187 & n12218;
  assign n12220 = n12185 & n12219;
  assign n12221 = n12176 & n12220;
  assign n12222 = n12167 & n12221;
  assign n12223 = n12222 ^ n9663;
  assign n12224 = n12223 ^ x563;
  assign n12229 = ~n12087 & ~n12224;
  assign n12230 = n11634 & n12229;
  assign n12231 = ~n12228 & ~n12230;
  assign n12088 = n12087 ^ n11856;
  assign n12225 = n12224 ^ n12088;
  assign n12226 = ~n11634 & ~n12225;
  assign n12232 = n12231 ^ n12226;
  assign n12233 = n11392 & ~n12232;
  assign n12234 = ~n11046 & n11391;
  assign n12235 = ~n11634 & ~n11856;
  assign n12236 = ~n12224 & n12235;
  assign n12237 = n12224 ^ n12087;
  assign n12238 = n11856 & ~n12237;
  assign n12239 = ~n11856 & ~n12087;
  assign n12240 = n11634 & ~n12239;
  assign n12241 = n12224 & n12240;
  assign n12242 = ~n12238 & ~n12241;
  assign n12243 = ~n12236 & n12242;
  assign n12244 = n12234 & n12243;
  assign n12245 = ~n12233 & ~n12244;
  assign n12246 = n11046 & n11391;
  assign n12247 = n12224 & n12227;
  assign n12248 = ~n11856 & n12087;
  assign n12249 = ~n12224 & n12248;
  assign n12250 = n11634 & n12249;
  assign n12251 = ~n12247 & ~n12250;
  assign n12252 = n11856 & n12229;
  assign n12253 = n12088 & ~n12224;
  assign n12254 = n12253 ^ n11856;
  assign n12255 = ~n11634 & ~n12254;
  assign n12256 = ~n12252 & ~n12255;
  assign n12257 = n12251 & n12256;
  assign n12258 = n12246 & ~n12257;
  assign n12259 = ~n11046 & ~n11391;
  assign n12260 = ~n11634 & ~n12088;
  assign n12261 = ~n12224 & n12260;
  assign n12262 = ~n11634 & n11856;
  assign n12263 = ~n12237 & n12262;
  assign n12264 = n12224 & n12239;
  assign n12265 = ~n12087 & n12224;
  assign n12266 = ~n12249 & ~n12265;
  assign n12267 = n11634 & ~n12266;
  assign n12268 = ~n12264 & ~n12267;
  assign n12269 = ~n12263 & n12268;
  assign n12270 = ~n12261 & n12269;
  assign n12271 = n12259 & ~n12270;
  assign n12272 = ~n12258 & ~n12271;
  assign n12273 = n12245 & n12272;
  assign n12274 = n12273 ^ n10458;
  assign n12275 = n12274 ^ x630;
  assign n12276 = n11855 ^ x568;
  assign n12277 = n11395 & n11600;
  assign n12278 = ~n11583 & ~n11601;
  assign n12279 = n11563 & ~n12278;
  assign n12280 = ~n12277 & ~n12279;
  assign n12281 = n11590 & ~n11615;
  assign n12282 = n11578 & ~n12281;
  assign n12283 = n11428 & n11573;
  assign n12284 = ~n11610 & ~n12283;
  assign n12285 = n11563 & ~n12284;
  assign n12286 = ~n12282 & ~n12285;
  assign n12287 = n12280 & n12286;
  assign n12288 = n11563 & n11615;
  assign n12289 = ~n11561 & ~n11600;
  assign n12290 = ~n11617 & n12289;
  assign n12291 = n11578 & ~n12290;
  assign n12292 = ~n12288 & ~n12291;
  assign n12293 = n11563 & n11589;
  assign n12294 = n11395 & n11610;
  assign n12295 = ~n12293 & ~n12294;
  assign n12296 = n11574 & n11592;
  assign n12297 = n12295 & ~n12296;
  assign n12298 = n11563 & ~n12289;
  assign n12299 = ~n11579 & ~n11594;
  assign n12300 = ~n11599 & ~n12299;
  assign n12301 = ~n12298 & ~n12300;
  assign n12302 = n11395 & n11601;
  assign n12303 = ~n11395 & ~n11589;
  assign n12304 = n11612 & ~n12283;
  assign n12305 = ~n11592 & n12304;
  assign n12306 = ~n12303 & ~n12305;
  assign n12307 = ~n11570 & ~n12306;
  assign n12308 = ~n11617 & n12307;
  assign n12309 = n11394 & ~n12308;
  assign n12310 = ~n12302 & ~n12309;
  assign n12311 = n12301 & n12310;
  assign n12312 = n12297 & n12311;
  assign n12313 = n12292 & n12312;
  assign n12314 = n12287 & n12313;
  assign n12315 = ~n11598 & n12314;
  assign n12316 = n12315 ^ n10109;
  assign n12317 = n12316 ^ x573;
  assign n12318 = n12276 & n12317;
  assign n12319 = n11700 ^ x514;
  assign n12320 = n12018 ^ x519;
  assign n12321 = ~n12319 & n12320;
  assign n12322 = n11886 ^ x518;
  assign n12323 = n10502 & n10642;
  assign n12324 = n10503 & n10648;
  assign n12325 = ~n12323 & ~n12324;
  assign n12326 = ~n10637 & n10639;
  assign n12327 = ~n10647 & ~n10652;
  assign n12328 = n10619 & ~n12327;
  assign n12329 = ~n10645 & ~n10654;
  assign n12330 = ~n10624 & ~n12329;
  assign n12331 = ~n10622 & ~n10669;
  assign n12332 = n10503 & ~n12331;
  assign n12333 = ~n12330 & ~n12332;
  assign n12334 = n10619 & n11152;
  assign n12335 = ~n10627 & ~n11158;
  assign n12336 = n10630 & ~n12335;
  assign n12337 = n10659 & n12327;
  assign n12338 = n10639 & ~n12337;
  assign n12339 = ~n12336 & ~n12338;
  assign n12340 = ~n12334 & n12339;
  assign n12341 = n12333 & n12340;
  assign n12342 = ~n10618 & n12341;
  assign n12343 = ~n11144 & n12342;
  assign n12344 = ~n11893 & n12343;
  assign n12345 = ~n12328 & n12344;
  assign n12346 = ~n12326 & n12345;
  assign n12347 = n12325 & n12346;
  assign n12348 = n11156 & n12347;
  assign n12349 = ~n10653 & n12348;
  assign n12350 = n12349 ^ n8328;
  assign n12351 = n12350 ^ x517;
  assign n12352 = n12322 & ~n12351;
  assign n12353 = ~n10764 & n10796;
  assign n12354 = ~n10788 & n12353;
  assign n12355 = n10749 & ~n12354;
  assign n12356 = n10796 & n11738;
  assign n12357 = n10763 & ~n12356;
  assign n12358 = ~n12355 & ~n12357;
  assign n12359 = ~n10747 & n10779;
  assign n12360 = n10754 & ~n12359;
  assign n12361 = ~n10754 & n11216;
  assign n12362 = ~n10756 & n10785;
  assign n12363 = ~n10749 & n12362;
  assign n12364 = ~n12361 & ~n12363;
  assign n12365 = ~n10691 & n12364;
  assign n12366 = n10791 & n11208;
  assign n12367 = n10693 & ~n12366;
  assign n12368 = ~n12365 & ~n12367;
  assign n12369 = ~n12360 & n12368;
  assign n12370 = n12358 & n12369;
  assign n12371 = n10771 & n12370;
  assign n12372 = ~n10748 & n12371;
  assign n12373 = n12372 ^ n8544;
  assign n12374 = n12373 ^ x516;
  assign n12375 = n11789 ^ x515;
  assign n12376 = ~n12374 & n12375;
  assign n12377 = ~n12352 & n12376;
  assign n12378 = ~n12374 & ~n12375;
  assign n12379 = ~n12351 & n12378;
  assign n12380 = n12351 & n12375;
  assign n12381 = n12351 ^ n12322;
  assign n12382 = n12380 & n12381;
  assign n12383 = n12382 ^ n12381;
  assign n12384 = n12374 & n12383;
  assign n12385 = ~n12379 & ~n12384;
  assign n12386 = ~n12377 & n12385;
  assign n12387 = n12321 & ~n12386;
  assign n12388 = n12319 & n12320;
  assign n12389 = n12352 & n12376;
  assign n12390 = n12374 & ~n12375;
  assign n12391 = n12352 & n12390;
  assign n12392 = n12351 & n12378;
  assign n12393 = ~n12391 & ~n12392;
  assign n12394 = n12322 & n12351;
  assign n12395 = ~n12376 & n12394;
  assign n12396 = ~n12322 & ~n12351;
  assign n12397 = ~n12376 & ~n12390;
  assign n12398 = n12396 & n12397;
  assign n12399 = ~n12395 & ~n12398;
  assign n12400 = n12393 & n12399;
  assign n12401 = ~n12389 & n12400;
  assign n12402 = n12388 & ~n12401;
  assign n12403 = ~n12387 & ~n12402;
  assign n12404 = n12319 & ~n12320;
  assign n12406 = ~n12378 & ~n12380;
  assign n12405 = n12390 ^ n12351;
  assign n12407 = n12406 ^ n12405;
  assign n12408 = ~n12322 & n12407;
  assign n12409 = n12408 ^ n12406;
  assign n12410 = n12404 & n12409;
  assign n12411 = ~n12319 & ~n12320;
  assign n12412 = n12374 & n12380;
  assign n12413 = ~n12375 & n12396;
  assign n12414 = ~n12380 & ~n12397;
  assign n12415 = n12322 & ~n12414;
  assign n12416 = ~n12413 & ~n12415;
  assign n12417 = ~n12412 & n12416;
  assign n12418 = n12411 & ~n12417;
  assign n12419 = ~n12410 & ~n12418;
  assign n12420 = n12403 & n12419;
  assign n12421 = n12420 ^ n10181;
  assign n12422 = n12421 ^ x572;
  assign n12423 = n11923 ^ x526;
  assign n12424 = n10811 ^ x531;
  assign n12425 = n12423 & n12424;
  assign n12426 = n9838 ^ x530;
  assign n12427 = n11913 ^ x527;
  assign n12428 = n12426 & n12427;
  assign n12429 = ~n11110 & ~n11692;
  assign n12430 = n11128 & ~n12429;
  assign n12431 = n11102 & ~n11118;
  assign n12432 = ~n12110 & ~n12431;
  assign n12433 = n11102 & ~n11114;
  assign n12434 = n11049 & ~n12433;
  assign n12435 = ~n12432 & ~n12434;
  assign n12436 = ~n11105 & n12435;
  assign n12437 = n11047 & ~n12436;
  assign n12438 = ~n12430 & ~n12437;
  assign n12439 = n11049 & n11091;
  assign n12440 = n11126 & ~n11687;
  assign n12441 = ~n11090 & n12440;
  assign n12442 = n11118 & ~n12441;
  assign n12443 = ~n12439 & ~n12442;
  assign n12444 = ~n11082 & ~n11125;
  assign n12445 = n11088 & ~n12444;
  assign n12446 = n11086 & ~n12093;
  assign n12447 = n11128 & ~n12446;
  assign n12448 = ~n11105 & n12429;
  assign n12449 = n11088 & ~n12448;
  assign n12450 = ~n12447 & ~n12449;
  assign n12451 = ~n11687 & n12450;
  assign n12452 = ~n11047 & ~n12451;
  assign n12453 = ~n12445 & ~n12452;
  assign n12454 = n12443 & n12453;
  assign n12455 = n12438 & n12454;
  assign n12456 = n12097 & n12455;
  assign n12457 = n11094 & n12456;
  assign n12458 = n12457 ^ n9095;
  assign n12459 = n12458 ^ x528;
  assign n12460 = n11490 & n11535;
  assign n12461 = n11494 & ~n11527;
  assign n12462 = ~n12460 & ~n12461;
  assign n12463 = ~n11512 & ~n11518;
  assign n12464 = n11656 & n11659;
  assign n12465 = ~n11505 & n12464;
  assign n12466 = ~n11526 & n12465;
  assign n12467 = n11523 & ~n12466;
  assign n12468 = n11492 & ~n11997;
  assign n12469 = ~n11503 & n11659;
  assign n12470 = ~n11519 & n12002;
  assign n12471 = ~n11499 & n12470;
  assign n12472 = ~n12469 & ~n12471;
  assign n12473 = ~n11508 & ~n12472;
  assign n12474 = n11491 & ~n12473;
  assign n12475 = ~n12468 & ~n12474;
  assign n12476 = ~n12467 & n12475;
  assign n12477 = ~n12463 & n12476;
  assign n12478 = n12462 & n12477;
  assign n12479 = n11502 & n12478;
  assign n12480 = n11985 & n12479;
  assign n12481 = n11648 & n12480;
  assign n12482 = n12481 ^ n9127;
  assign n12483 = n12482 ^ x529;
  assign n12484 = n12459 & n12483;
  assign n12485 = n12428 & n12484;
  assign n12486 = n12425 & n12485;
  assign n12487 = ~n12423 & ~n12424;
  assign n12488 = ~n12459 & ~n12483;
  assign n12489 = n12428 & n12488;
  assign n12490 = n12487 & n12489;
  assign n12491 = ~n12486 & ~n12490;
  assign n12492 = ~n12426 & n12427;
  assign n12493 = n12459 & ~n12483;
  assign n12494 = n12492 & n12493;
  assign n12495 = n12425 & n12494;
  assign n12496 = ~n12423 & n12424;
  assign n12497 = n12426 & ~n12427;
  assign n12498 = n12493 & n12497;
  assign n12499 = ~n12426 & ~n12427;
  assign n12500 = n12488 & n12499;
  assign n12501 = ~n12498 & ~n12500;
  assign n12502 = n12496 & ~n12501;
  assign n12503 = ~n12495 & ~n12502;
  assign n12504 = n12428 & n12493;
  assign n12505 = n12496 & n12504;
  assign n12506 = n12423 & ~n12424;
  assign n12507 = n12493 & n12499;
  assign n12508 = n12506 & n12507;
  assign n12509 = ~n12505 & ~n12508;
  assign n12510 = ~n12459 & n12483;
  assign n12511 = n12499 & n12510;
  assign n12512 = n12496 & n12511;
  assign n12513 = n12428 & n12510;
  assign n12514 = n12484 & n12492;
  assign n12515 = ~n12513 & ~n12514;
  assign n12516 = n12487 & ~n12515;
  assign n12517 = ~n12512 & ~n12516;
  assign n12518 = n12492 & n12510;
  assign n12519 = n12487 & n12518;
  assign n12520 = n12425 & ~n12515;
  assign n12521 = ~n12519 & ~n12520;
  assign n12522 = n12496 & n12514;
  assign n12523 = n12424 ^ n12423;
  assign n12524 = n12497 & n12510;
  assign n12525 = ~n12489 & ~n12518;
  assign n12526 = ~n12524 & n12525;
  assign n12527 = n12523 & ~n12526;
  assign n12528 = ~n12522 & ~n12527;
  assign n12529 = n12488 & n12492;
  assign n12530 = n12484 & n12497;
  assign n12531 = n12484 & n12499;
  assign n12532 = ~n12530 & ~n12531;
  assign n12533 = ~n12494 & n12532;
  assign n12534 = ~n12529 & n12533;
  assign n12535 = n12506 & ~n12534;
  assign n12536 = ~n12425 & ~n12487;
  assign n12537 = n12488 & n12497;
  assign n12538 = ~n12511 & ~n12537;
  assign n12539 = ~n12487 & n12538;
  assign n12540 = ~n12504 & ~n12530;
  assign n12541 = ~n12425 & n12540;
  assign n12542 = ~n12539 & ~n12541;
  assign n12543 = n12501 & ~n12542;
  assign n12544 = ~n12536 & ~n12543;
  assign n12545 = ~n12535 & ~n12544;
  assign n12546 = n12528 & n12545;
  assign n12547 = n12521 & n12546;
  assign n12548 = n12517 & n12547;
  assign n12549 = n12509 & n12548;
  assign n12550 = n12503 & n12549;
  assign n12551 = n12491 & n12550;
  assign n12552 = n12551 ^ n10715;
  assign n12553 = n12552 ^ x571;
  assign n12554 = n12422 & n12553;
  assign n12555 = ~n12155 & n12203;
  assign n12556 = n12188 & ~n12555;
  assign n12557 = ~n12164 & ~n12191;
  assign n12558 = n12091 & ~n12557;
  assign n12559 = ~n12159 & ~n12192;
  assign n12560 = n12177 & ~n12559;
  assign n12561 = n12161 & n12209;
  assign n12562 = ~n12168 & ~n12191;
  assign n12563 = ~n12201 & ~n12562;
  assign n12564 = ~n12182 & n12199;
  assign n12565 = n12188 & ~n12564;
  assign n12566 = n12174 & n12210;
  assign n12567 = n12177 & ~n12566;
  assign n12568 = ~n12565 & ~n12567;
  assign n12569 = ~n12563 & n12568;
  assign n12570 = n12161 & ~n12180;
  assign n12571 = ~n12182 & ~n12205;
  assign n12572 = ~n12178 & n12571;
  assign n12573 = ~n12173 & n12572;
  assign n12574 = ~n12168 & n12573;
  assign n12575 = n12091 & ~n12574;
  assign n12576 = ~n12570 & ~n12575;
  assign n12577 = n12569 & n12576;
  assign n12578 = ~n12561 & n12577;
  assign n12579 = ~n12560 & n12578;
  assign n12580 = n12166 & n12579;
  assign n12581 = n12185 & n12580;
  assign n12582 = ~n12558 & n12581;
  assign n12583 = ~n12556 & n12582;
  assign n12584 = n12583 ^ n10744;
  assign n12585 = n12584 ^ x570;
  assign n12586 = n11390 ^ x569;
  assign n12587 = ~n12585 & n12586;
  assign n12588 = n12554 & n12587;
  assign n12589 = n12318 & n12588;
  assign n12590 = n12276 & ~n12317;
  assign n12591 = n12588 & n12590;
  assign n12592 = ~n12276 & ~n12317;
  assign n12593 = ~n12422 & n12553;
  assign n12594 = n12587 & n12593;
  assign n12595 = n12592 & n12594;
  assign n12596 = n12422 & ~n12553;
  assign n12597 = n12585 & ~n12586;
  assign n12598 = n12596 & n12597;
  assign n12599 = n12318 & n12598;
  assign n12600 = ~n12422 & ~n12553;
  assign n12601 = n12585 & n12586;
  assign n12602 = n12600 & n12601;
  assign n12603 = n12554 & n12601;
  assign n12604 = ~n12602 & ~n12603;
  assign n12605 = n12590 & ~n12604;
  assign n12606 = ~n12599 & ~n12605;
  assign n12607 = ~n12595 & n12606;
  assign n12608 = ~n12591 & n12607;
  assign n12609 = ~n12276 & n12317;
  assign n12610 = ~n12585 & ~n12586;
  assign n12611 = n12593 & n12610;
  assign n12612 = n12596 & n12610;
  assign n12613 = ~n12611 & ~n12612;
  assign n12614 = n12609 & ~n12613;
  assign n12615 = n12590 & n12594;
  assign n12616 = n12597 & n12600;
  assign n12617 = n12554 & n12597;
  assign n12618 = ~n12616 & ~n12617;
  assign n12619 = n12609 & ~n12618;
  assign n12620 = ~n12615 & ~n12619;
  assign n12621 = n12317 ^ n12276;
  assign n12622 = n12593 & n12601;
  assign n12623 = n12621 & n12622;
  assign n12624 = ~n12612 & ~n12616;
  assign n12625 = n12593 & n12597;
  assign n12626 = n12554 & n12610;
  assign n12627 = ~n12625 & ~n12626;
  assign n12628 = n12624 & n12627;
  assign n12629 = n12592 & ~n12628;
  assign n12630 = ~n12623 & ~n12629;
  assign n12631 = n12587 & n12596;
  assign n12632 = n12587 & n12600;
  assign n12633 = n12596 & n12601;
  assign n12634 = ~n12632 & ~n12633;
  assign n12635 = ~n12631 & n12634;
  assign n12636 = ~n12276 & ~n12635;
  assign n12637 = n12600 & n12610;
  assign n12638 = ~n12611 & ~n12637;
  assign n12639 = ~n12612 & n12638;
  assign n12640 = n12590 & ~n12639;
  assign n12641 = ~n12622 & ~n12633;
  assign n12642 = ~n12594 & n12641;
  assign n12643 = n12618 & n12642;
  assign n12644 = ~n12637 & n12643;
  assign n12645 = n12318 & ~n12644;
  assign n12646 = ~n12640 & ~n12645;
  assign n12647 = ~n12636 & n12646;
  assign n12648 = n12630 & n12647;
  assign n12649 = n12620 & n12648;
  assign n12650 = ~n12614 & n12649;
  assign n12651 = n12608 & n12650;
  assign n12652 = ~n12589 & n12651;
  assign n12653 = n12652 ^ n10811;
  assign n12654 = n12653 ^ x629;
  assign n12655 = ~n12275 & n12654;
  assign n12656 = n10287 ^ n9839;
  assign n12657 = n10993 & n11001;
  assign n12658 = ~n11030 & ~n12657;
  assign n12659 = ~n11021 & ~n11031;
  assign n12660 = n12658 & n12659;
  assign n12661 = n12656 & ~n12660;
  assign n12662 = n10985 & n11015;
  assign n12663 = ~n10995 & ~n12662;
  assign n12664 = n11017 & n12663;
  assign n12665 = n11007 & ~n12664;
  assign n12666 = ~n12661 & ~n12665;
  assign n12667 = ~n11005 & ~n11035;
  assign n12668 = ~n11000 & n12667;
  assign n12669 = ~n11031 & n12668;
  assign n12670 = n10288 & ~n12669;
  assign n12671 = ~n10994 & ~n11002;
  assign n12672 = ~n10986 & n12671;
  assign n12673 = ~n10989 & n12672;
  assign n12674 = ~n10288 & n12673;
  assign n12675 = ~n10989 & ~n12662;
  assign n12676 = ~n10994 & n12675;
  assign n12677 = ~n11008 & n12676;
  assign n12678 = ~n11020 & n12677;
  assign n12679 = ~n12674 & ~n12678;
  assign n12680 = n9839 & n12679;
  assign n12681 = ~n11016 & n12672;
  assign n12682 = n10992 & ~n12681;
  assign n12683 = ~n11008 & n12668;
  assign n12684 = n11007 & ~n12683;
  assign n12685 = ~n12682 & ~n12684;
  assign n12686 = ~n12680 & n12685;
  assign n12687 = ~n12670 & n12686;
  assign n12688 = n12666 & n12687;
  assign n12689 = n12688 ^ n10863;
  assign n12690 = n12689 ^ x553;
  assign n12691 = n11793 & ~n11818;
  assign n12692 = ~n11812 & n11823;
  assign n12693 = ~n12691 & ~n12692;
  assign n12694 = n11798 & n11834;
  assign n12695 = n11680 & n11807;
  assign n12696 = ~n11811 & ~n12695;
  assign n12697 = n11824 & ~n12696;
  assign n12698 = ~n12694 & ~n12697;
  assign n12699 = ~n11820 & ~n11842;
  assign n12700 = n12696 & n12699;
  assign n12701 = ~n11801 & n12700;
  assign n12702 = n11798 & ~n12701;
  assign n12703 = ~n11808 & ~n11833;
  assign n12704 = ~n11817 & n12703;
  assign n12705 = ~n11795 & n12704;
  assign n12706 = ~n11842 & n12705;
  assign n12707 = ~n11801 & n12706;
  assign n12708 = n11824 & ~n12707;
  assign n12709 = ~n12702 & ~n12708;
  assign n12710 = ~n11820 & n12696;
  assign n12711 = ~n11834 & n12710;
  assign n12712 = ~n11808 & n12711;
  assign n12713 = ~n11736 & n12712;
  assign n12714 = n11791 & ~n12713;
  assign n12715 = n11795 & ~n11812;
  assign n12716 = n11680 & n11800;
  assign n12717 = ~n11835 & n12703;
  assign n12718 = ~n12716 & n12717;
  assign n12719 = ~n11803 & n12718;
  assign n12720 = ~n11736 & n12719;
  assign n12721 = n11793 & ~n12720;
  assign n12722 = ~n12715 & ~n12721;
  assign n12723 = ~n12714 & n12722;
  assign n12724 = n12709 & n12723;
  assign n12725 = n12698 & n12724;
  assign n12726 = n12693 & n12725;
  assign n12727 = n12726 ^ n10917;
  assign n12728 = n12727 ^ x552;
  assign n12729 = ~n12690 & n12728;
  assign n12730 = n11563 & n11596;
  assign n12731 = n11395 & n11615;
  assign n12732 = n11579 & n11592;
  assign n12733 = ~n12731 & ~n12732;
  assign n12734 = ~n12730 & n12733;
  assign n12735 = n11583 & n11592;
  assign n12736 = ~n11393 & n12283;
  assign n12737 = ~n12735 & ~n12736;
  assign n12738 = n11395 & n11617;
  assign n12739 = n11592 & ~n12281;
  assign n12740 = ~n12738 & ~n12739;
  assign n12741 = n11561 & ~n11599;
  assign n12742 = n11563 & n11570;
  assign n12743 = ~n12741 & ~n12742;
  assign n12744 = ~n11583 & n11620;
  assign n12745 = n11578 & ~n12744;
  assign n12746 = ~n11594 & ~n11596;
  assign n12747 = n11394 & ~n12746;
  assign n12748 = ~n12745 & ~n12747;
  assign n12749 = n12743 & n12748;
  assign n12750 = n12740 & n12749;
  assign n12751 = n12737 & n12750;
  assign n12752 = n12734 & n12751;
  assign n12753 = n11577 & n12752;
  assign n12754 = n12287 & n12753;
  assign n12755 = n12754 ^ n10892;
  assign n12756 = n12755 ^ x551;
  assign n12757 = n12027 & n12033;
  assign n12758 = n12029 & n12062;
  assign n12759 = ~n12757 & ~n12758;
  assign n12760 = ~n11887 & n12039;
  assign n12761 = n12023 & n12033;
  assign n12762 = ~n12760 & ~n12761;
  assign n12763 = n12062 & n12064;
  assign n12764 = n12027 & n12063;
  assign n12765 = ~n12763 & ~n12764;
  assign n12766 = n12762 & n12765;
  assign n12767 = ~n11887 & n12051;
  assign n12768 = n12062 & ~n12077;
  assign n12769 = ~n12767 & ~n12768;
  assign n12770 = n12066 & n12071;
  assign n12771 = n11915 & ~n12770;
  assign n12772 = n12042 & ~n12047;
  assign n12773 = n12027 & ~n12772;
  assign n12774 = n12028 & n12038;
  assign n12775 = ~n12021 & ~n12040;
  assign n12776 = ~n12069 & n12775;
  assign n12777 = ~n12052 & n12776;
  assign n12778 = ~n12063 & n12777;
  assign n12779 = ~n12774 & n12778;
  assign n12780 = n12023 & ~n12779;
  assign n12781 = ~n12773 & ~n12780;
  assign n12782 = ~n12771 & n12781;
  assign n12783 = n12769 & n12782;
  assign n12784 = n12766 & n12783;
  assign n12785 = n12759 & n12784;
  assign n12786 = n12037 & n12785;
  assign n12787 = n12786 ^ n9786;
  assign n12788 = n12787 ^ x554;
  assign n12789 = n12756 & n12788;
  assign n12790 = n12729 & n12789;
  assign n12791 = n12690 & ~n12728;
  assign n12792 = n12756 & ~n12788;
  assign n12793 = n12791 & n12792;
  assign n12794 = ~n12790 & ~n12793;
  assign n12795 = n11178 & n11352;
  assign n12796 = n11324 & n11370;
  assign n12797 = n11314 & n11348;
  assign n12798 = ~n12796 & ~n12797;
  assign n12799 = n11312 & n11324;
  assign n12800 = n11178 & n11354;
  assign n12801 = ~n12799 & ~n12800;
  assign n12802 = ~n11177 & n11374;
  assign n12803 = ~n11324 & n11363;
  assign n12804 = n11339 & ~n12803;
  assign n12805 = ~n12802 & ~n12804;
  assign n12806 = ~n11316 & ~n11369;
  assign n12807 = ~n11321 & n12806;
  assign n12808 = n11337 & ~n12807;
  assign n12809 = n12805 & ~n12808;
  assign n12810 = n11358 & ~n11363;
  assign n12811 = n11324 & n11365;
  assign n12812 = ~n12810 & ~n12811;
  assign n12813 = n11143 & n11334;
  assign n12814 = n11314 & ~n11330;
  assign n12815 = ~n12813 & ~n12814;
  assign n12816 = n12812 & n12815;
  assign n12817 = n12809 & n12816;
  assign n12818 = n12801 & n12817;
  assign n12819 = n11356 & n12818;
  assign n12820 = n12798 & n12819;
  assign n12821 = n11332 & n12820;
  assign n12822 = ~n12795 & n12821;
  assign n12823 = n11318 & n12822;
  assign n12824 = ~n11344 & n12823;
  assign n12825 = n12824 ^ n9469;
  assign n12826 = n12825 ^ x555;
  assign n12827 = ~n12498 & ~n12531;
  assign n12828 = n12425 & ~n12827;
  assign n12829 = ~n12500 & ~n12524;
  assign n12830 = ~n12494 & n12829;
  assign n12831 = n12506 & ~n12830;
  assign n12832 = n12506 & n12530;
  assign n12833 = ~n12536 & n12537;
  assign n12834 = ~n12832 & ~n12833;
  assign n12835 = n12425 & n12507;
  assign n12836 = ~n12498 & ~n12511;
  assign n12837 = ~n12494 & n12836;
  assign n12838 = n12487 & ~n12837;
  assign n12839 = n12506 & ~n12515;
  assign n12840 = ~n12504 & ~n12529;
  assign n12841 = n12523 & ~n12840;
  assign n12842 = ~n12839 & ~n12841;
  assign n12843 = ~n12518 & n12533;
  assign n12844 = n12829 & n12843;
  assign n12845 = n12496 & ~n12844;
  assign n12846 = ~n12485 & ~n12518;
  assign n12847 = ~n12425 & n12846;
  assign n12848 = ~n12489 & ~n12529;
  assign n12849 = ~n12487 & n12848;
  assign n12850 = ~n12847 & ~n12849;
  assign n12851 = ~n12514 & ~n12850;
  assign n12852 = ~n12536 & ~n12851;
  assign n12853 = ~n12845 & ~n12852;
  assign n12854 = n12842 & n12853;
  assign n12855 = n12491 & n12854;
  assign n12856 = ~n12838 & n12855;
  assign n12857 = ~n12835 & n12856;
  assign n12858 = n12834 & n12857;
  assign n12859 = ~n12831 & n12858;
  assign n12860 = ~n12828 & n12859;
  assign n12861 = n12860 ^ n10841;
  assign n12862 = n12861 ^ x550;
  assign n12863 = ~n12826 & ~n12862;
  assign n12864 = ~n12794 & n12863;
  assign n12865 = n12690 & n12728;
  assign n12866 = ~n12756 & n12788;
  assign n12867 = n12865 & n12866;
  assign n12868 = ~n12756 & ~n12788;
  assign n12869 = n12791 & n12868;
  assign n12870 = ~n12867 & ~n12869;
  assign n12871 = n12826 & ~n12862;
  assign n12872 = ~n12870 & n12871;
  assign n12873 = ~n12864 & ~n12872;
  assign n12874 = ~n12690 & ~n12728;
  assign n12875 = n12868 & n12874;
  assign n12876 = n12826 & n12862;
  assign n12877 = n12875 & n12876;
  assign n12878 = n12866 & n12874;
  assign n12879 = n12792 & n12865;
  assign n12880 = ~n12878 & ~n12879;
  assign n12881 = n12871 & ~n12880;
  assign n12882 = ~n12877 & ~n12881;
  assign n12883 = n12789 & n12791;
  assign n12884 = n12862 & n12883;
  assign n12885 = ~n12826 & n12862;
  assign n12886 = n12789 & n12874;
  assign n12887 = ~n12879 & ~n12886;
  assign n12888 = ~n12793 & n12887;
  assign n12889 = n12885 & ~n12888;
  assign n12890 = ~n12794 & n12871;
  assign n12891 = n12865 & n12868;
  assign n12892 = n12876 & n12891;
  assign n12893 = n12729 & n12866;
  assign n12894 = n12863 & n12893;
  assign n12895 = ~n12892 & ~n12894;
  assign n12896 = ~n12890 & n12895;
  assign n12897 = ~n12867 & ~n12875;
  assign n12898 = n12885 & ~n12897;
  assign n12899 = n12862 ^ n12826;
  assign n12900 = n12789 & n12865;
  assign n12901 = n12792 & n12874;
  assign n12902 = ~n12900 & ~n12901;
  assign n12903 = ~n12899 & ~n12902;
  assign n12904 = ~n12869 & ~n12891;
  assign n12905 = ~n12878 & n12904;
  assign n12906 = n12863 & ~n12905;
  assign n12907 = ~n12903 & ~n12906;
  assign n12908 = n12729 & n12792;
  assign n12909 = ~n12886 & ~n12908;
  assign n12910 = n12871 & ~n12909;
  assign n12911 = n12791 & n12866;
  assign n12912 = n12729 & n12868;
  assign n12913 = ~n12911 & ~n12912;
  assign n12914 = n12876 & n12893;
  assign n12915 = n12913 & ~n12914;
  assign n12916 = n12862 & ~n12915;
  assign n12917 = ~n12910 & ~n12916;
  assign n12918 = n12907 & n12917;
  assign n12919 = ~n12898 & n12918;
  assign n12920 = n12896 & n12919;
  assign n12921 = ~n12889 & n12920;
  assign n12922 = ~n12884 & n12921;
  assign n12923 = n12882 & n12922;
  assign n12924 = n12873 & n12923;
  assign n12925 = n12924 ^ n10983;
  assign n12926 = n12925 ^ x632;
  assign n12927 = n11793 & n11823;
  assign n12928 = n11797 & ~n12927;
  assign n12929 = n12696 & n12703;
  assign n12930 = n11793 & ~n12929;
  assign n12931 = n12711 & n12717;
  assign n12932 = n11824 & ~n12931;
  assign n12933 = ~n12930 & ~n12932;
  assign n12934 = n11791 & ~n12707;
  assign n12935 = ~n11803 & n11818;
  assign n12936 = ~n11834 & n12935;
  assign n12937 = ~n11811 & n12936;
  assign n12938 = ~n11736 & n12937;
  assign n12939 = ~n11842 & n12938;
  assign n12940 = n11798 & ~n12939;
  assign n12941 = ~n12934 & ~n12940;
  assign n12942 = n12933 & n12941;
  assign n12943 = n12693 & n12942;
  assign n12944 = n12928 & n12943;
  assign n12945 = ~n11825 & n12944;
  assign n12946 = n12945 ^ n10613;
  assign n12947 = n12946 ^ x588;
  assign n12948 = n12506 & ~n12846;
  assign n12949 = ~n12507 & ~n12530;
  assign n12950 = n12496 & ~n12949;
  assign n12951 = n12487 & n12524;
  assign n12952 = n12494 & ~n12536;
  assign n12953 = ~n12951 & ~n12952;
  assign n12954 = n12829 & n12840;
  assign n12955 = ~n12537 & n12954;
  assign n12956 = n12506 & ~n12955;
  assign n12957 = ~n12459 & n12496;
  assign n12958 = n12427 & n12957;
  assign n12959 = ~n12956 & ~n12958;
  assign n12960 = ~n12514 & n12525;
  assign n12961 = n12425 & ~n12960;
  assign n12962 = ~n12487 & n12829;
  assign n12963 = n12501 & ~n12531;
  assign n12964 = ~n12537 & n12963;
  assign n12965 = ~n12425 & n12964;
  assign n12966 = ~n12962 & ~n12965;
  assign n12967 = ~n12536 & n12966;
  assign n12968 = ~n12961 & ~n12967;
  assign n12969 = n12959 & n12968;
  assign n12970 = n12953 & n12969;
  assign n12971 = ~n12950 & n12970;
  assign n12972 = n12517 & n12971;
  assign n12973 = ~n12948 & n12972;
  assign n12974 = n12509 & n12973;
  assign n12975 = ~n12828 & n12974;
  assign n12976 = n12975 ^ n10567;
  assign n12977 = n12976 ^ x587;
  assign n12978 = n12947 & ~n12977;
  assign n12979 = ~n10986 & ~n10995;
  assign n12980 = n11020 & ~n12979;
  assign n12981 = n11003 & n11017;
  assign n12982 = n12656 & ~n12981;
  assign n12983 = ~n12980 & ~n12982;
  assign n12984 = n10992 & ~n11036;
  assign n12985 = n10288 & n11025;
  assign n12986 = ~n12984 & ~n12985;
  assign n12987 = n12983 & n12986;
  assign n12988 = n9839 & ~n12658;
  assign n12989 = n11007 & n11028;
  assign n12990 = ~n12988 & ~n12989;
  assign n12991 = n12987 & n12990;
  assign n12992 = n10998 & n12991;
  assign n12993 = n12992 ^ n10589;
  assign n12994 = n12993 ^ x590;
  assign n12995 = n11178 & n11316;
  assign n12996 = ~n11355 & ~n12995;
  assign n12997 = n11312 & n11337;
  assign n12998 = ~n11358 & ~n11374;
  assign n12999 = n11314 & ~n12998;
  assign n13000 = ~n12997 & ~n12999;
  assign n13001 = ~n11177 & n11352;
  assign n13002 = ~n11329 & n12806;
  assign n13003 = ~n11370 & n13002;
  assign n13004 = n11337 & ~n13003;
  assign n13005 = ~n13001 & ~n13004;
  assign n13006 = n11314 & n11354;
  assign n13007 = ~n11327 & ~n11365;
  assign n13008 = ~n11321 & n13007;
  assign n13009 = n11178 & ~n13008;
  assign n13010 = n11314 & n11344;
  assign n13011 = ~n11334 & ~n11374;
  assign n13012 = n11324 & ~n13011;
  assign n13013 = ~n13010 & ~n13012;
  assign n13014 = n12798 & n13013;
  assign n13015 = ~n11322 & n13014;
  assign n13016 = ~n13009 & n13015;
  assign n13017 = ~n13006 & n13016;
  assign n13018 = n13005 & n13017;
  assign n13019 = n12801 & n13018;
  assign n13020 = ~n11350 & n13019;
  assign n13021 = n13000 & n13020;
  assign n13022 = n12996 & n13021;
  assign n13023 = n11342 & n13022;
  assign n13024 = ~n12795 & n13023;
  assign n13025 = n13024 ^ n10531;
  assign n13026 = n13025 ^ x589;
  assign n13027 = n12994 & ~n13026;
  assign n13028 = n12978 & n13027;
  assign n13029 = n12352 & n12375;
  assign n13030 = ~n12322 & ~n12406;
  assign n13031 = ~n13029 & ~n13030;
  assign n13032 = n12393 & n13031;
  assign n13033 = n12411 & ~n13032;
  assign n13034 = ~n12375 & n12394;
  assign n13035 = n12374 & n12396;
  assign n13036 = ~n12322 & ~n12397;
  assign n13037 = ~n13035 & ~n13036;
  assign n13038 = ~n13034 & n13037;
  assign n13039 = n12404 & ~n13038;
  assign n13040 = ~n13033 & ~n13039;
  assign n13041 = ~n12374 & ~n12381;
  assign n13042 = ~n12322 & n12412;
  assign n13043 = ~n13041 & ~n13042;
  assign n13044 = ~n12351 & ~n12397;
  assign n13045 = n13043 & ~n13044;
  assign n13046 = n12388 & ~n13045;
  assign n13047 = ~n12351 & n12374;
  assign n13048 = n12375 & n13047;
  assign n13049 = n12322 & n12397;
  assign n13050 = ~n13048 & ~n13049;
  assign n13051 = n12352 & ~n12374;
  assign n13052 = n12351 & n13036;
  assign n13053 = ~n13051 & ~n13052;
  assign n13054 = n13050 & n13053;
  assign n13055 = n12321 & ~n13054;
  assign n13056 = ~n13046 & ~n13055;
  assign n13057 = n13040 & n13056;
  assign n13058 = ~n12389 & n13057;
  assign n13059 = n13058 ^ n10472;
  assign n13060 = n13059 ^ x591;
  assign n13061 = n12155 & n12161;
  assign n13062 = n12188 & n12205;
  assign n13063 = ~n12182 & ~n12202;
  assign n13064 = n12189 & n13063;
  assign n13065 = n12177 & ~n13064;
  assign n13066 = n12091 & ~n12203;
  assign n13067 = ~n12561 & ~n13066;
  assign n13068 = ~n12159 & n12180;
  assign n13069 = ~n12164 & n13068;
  assign n13070 = n12091 & ~n13069;
  assign n13071 = n12123 ^ n12092;
  assign n13072 = ~n12125 & ~n13071;
  assign n13073 = n12177 & n13072;
  assign n13074 = ~n13070 & ~n13073;
  assign n13075 = n12161 & ~n12571;
  assign n13076 = ~n12188 & n12199;
  assign n13077 = ~n12173 & ~n12200;
  assign n13078 = ~n12209 & n13077;
  assign n13079 = ~n12164 & n13078;
  assign n13080 = ~n13076 & ~n13079;
  assign n13081 = ~n12191 & ~n13080;
  assign n13082 = ~n12201 & ~n13081;
  assign n13083 = ~n13075 & ~n13082;
  assign n13084 = n13074 & n13083;
  assign n13085 = n13067 & n13084;
  assign n13086 = ~n13065 & n13085;
  assign n13087 = ~n13062 & n13086;
  assign n13088 = n12176 & n13087;
  assign n13089 = ~n12556 & n13088;
  assign n13090 = ~n13061 & n13089;
  assign n13091 = n13090 ^ n10501;
  assign n13092 = n13091 ^ x586;
  assign n13093 = ~n13060 & n13092;
  assign n13094 = n13028 & n13093;
  assign n13095 = ~n12947 & ~n12977;
  assign n13096 = ~n12994 & n13026;
  assign n13097 = n13095 & n13096;
  assign n13098 = n13060 & n13092;
  assign n13099 = n13097 & n13098;
  assign n13100 = ~n13094 & ~n13099;
  assign n13101 = ~n12994 & ~n13026;
  assign n13102 = n13095 & n13101;
  assign n13103 = ~n12947 & n12977;
  assign n13104 = n13096 & n13103;
  assign n13105 = n12947 & n12977;
  assign n13106 = n12994 & n13026;
  assign n13107 = n13105 & n13106;
  assign n13108 = ~n13104 & ~n13107;
  assign n13109 = ~n13102 & n13108;
  assign n13110 = ~n13060 & ~n13092;
  assign n13111 = ~n13109 & n13110;
  assign n13112 = n12978 & n13096;
  assign n13113 = n13027 & n13095;
  assign n13114 = ~n13112 & ~n13113;
  assign n13115 = n13060 & ~n13092;
  assign n13116 = ~n13114 & n13115;
  assign n13117 = ~n13111 & ~n13116;
  assign n13118 = n13027 & n13103;
  assign n13119 = n13115 & n13118;
  assign n13120 = n13095 & n13106;
  assign n13121 = n12978 & n13101;
  assign n13122 = ~n13120 & ~n13121;
  assign n13123 = n13110 & ~n13122;
  assign n13124 = ~n13119 & ~n13123;
  assign n13125 = n13096 & n13105;
  assign n13126 = ~n13118 & ~n13125;
  assign n13127 = n13098 & ~n13126;
  assign n13128 = n13028 & n13110;
  assign n13129 = n13097 & n13115;
  assign n13130 = ~n13128 & ~n13129;
  assign n13131 = n12978 & n13106;
  assign n13132 = n13027 & n13105;
  assign n13133 = ~n13125 & ~n13132;
  assign n13134 = ~n13131 & n13133;
  assign n13135 = n13115 & ~n13134;
  assign n13136 = n13101 & n13105;
  assign n13137 = n13115 & n13136;
  assign n13138 = n13101 & n13103;
  assign n13139 = ~n13132 & ~n13138;
  assign n13140 = n13092 & ~n13139;
  assign n13141 = ~n13137 & ~n13140;
  assign n13142 = n13093 & ~n13108;
  assign n13143 = n13103 & n13106;
  assign n13144 = ~n13138 & ~n13143;
  assign n13145 = n13110 & ~n13144;
  assign n13146 = n13114 & ~n13120;
  assign n13147 = ~n13098 & n13146;
  assign n13148 = n13122 & ~n13131;
  assign n13149 = ~n13093 & n13148;
  assign n13150 = ~n13147 & ~n13149;
  assign n13151 = n13092 & n13150;
  assign n13152 = ~n13145 & ~n13151;
  assign n13153 = ~n13142 & n13152;
  assign n13154 = n13141 & n13153;
  assign n13155 = ~n13135 & n13154;
  assign n13156 = n13130 & n13155;
  assign n13157 = ~n13127 & n13156;
  assign n13158 = n13124 & n13157;
  assign n13159 = n13117 & n13158;
  assign n13160 = n13100 & n13159;
  assign n13161 = n13160 ^ n10688;
  assign n13162 = n13161 ^ x631;
  assign n13163 = ~n12926 & ~n13162;
  assign n13164 = n12655 & n13163;
  assign n13165 = n12223 ^ x561;
  assign n13166 = n12787 ^ x556;
  assign n13167 = ~n13165 & n13166;
  assign n13168 = n12411 & n13054;
  assign n13169 = n12321 & ~n13032;
  assign n13170 = ~n13168 & ~n13169;
  assign n13171 = n12404 & n13045;
  assign n13172 = ~n12389 & n13038;
  assign n13173 = n12388 & ~n13172;
  assign n13174 = ~n13171 & ~n13173;
  assign n13175 = n13170 & n13174;
  assign n13176 = n13175 ^ n8589;
  assign n13177 = n13176 ^ x558;
  assign n13178 = n12825 ^ x557;
  assign n13179 = ~n13177 & n13178;
  assign n13180 = n11045 ^ x560;
  assign n13181 = n12511 & ~n12536;
  assign n13182 = n12515 & n12532;
  assign n13183 = ~n12529 & n13182;
  assign n13184 = ~n12537 & n13183;
  assign n13185 = n12487 & ~n13184;
  assign n13186 = ~n13181 & ~n13185;
  assign n13187 = ~n12524 & n12840;
  assign n13188 = n12425 & ~n13187;
  assign n13189 = ~n12513 & n12827;
  assign n13190 = n12506 & ~n13189;
  assign n13191 = n12459 ^ n12426;
  assign n13192 = n13191 ^ n12483;
  assign n13193 = n12427 & n13192;
  assign n13194 = n12496 & n13193;
  assign n13195 = ~n13190 & ~n13194;
  assign n13196 = ~n13188 & n13195;
  assign n13197 = n13186 & n13196;
  assign n13198 = ~n12950 & n13197;
  assign n13199 = ~n12948 & n13198;
  assign n13200 = ~n12831 & n13199;
  assign n13201 = n12503 & n13200;
  assign n13202 = n12491 & n13201;
  assign n13203 = ~n12828 & n13202;
  assign n13204 = n13203 ^ n9226;
  assign n13205 = n13204 ^ x559;
  assign n13206 = ~n13180 & n13205;
  assign n13207 = n13179 & n13206;
  assign n13208 = n13167 & n13207;
  assign n13209 = n13165 & ~n13166;
  assign n13210 = ~n13177 & ~n13178;
  assign n13211 = n13206 & n13210;
  assign n13212 = n13180 & ~n13205;
  assign n13213 = n13210 & n13212;
  assign n13214 = ~n13211 & ~n13213;
  assign n13215 = n13209 & ~n13214;
  assign n13216 = ~n13208 & ~n13215;
  assign n13217 = n13166 ^ n13165;
  assign n13218 = n13179 & n13212;
  assign n13219 = n13217 & n13218;
  assign n13220 = n13177 & ~n13178;
  assign n13221 = n13206 & n13220;
  assign n13222 = n13212 & n13220;
  assign n13223 = ~n13221 & ~n13222;
  assign n13224 = ~n13207 & n13223;
  assign n13225 = n13209 & ~n13224;
  assign n13226 = n13177 & n13178;
  assign n13227 = n13180 & n13205;
  assign n13228 = n13226 & n13227;
  assign n13229 = n13209 & n13228;
  assign n13230 = n13165 & n13166;
  assign n13231 = n13210 & n13227;
  assign n13232 = ~n13221 & ~n13231;
  assign n13233 = n13230 & ~n13232;
  assign n13234 = ~n13229 & ~n13233;
  assign n13235 = ~n13165 & ~n13166;
  assign n13236 = n13179 & n13227;
  assign n13237 = n13206 & n13226;
  assign n13238 = ~n13236 & ~n13237;
  assign n13239 = n13235 & ~n13238;
  assign n13240 = ~n13180 & ~n13205;
  assign n13241 = n13179 & n13240;
  assign n13242 = n13212 & n13226;
  assign n13243 = ~n13241 & ~n13242;
  assign n13244 = n13230 & ~n13243;
  assign n13245 = ~n13239 & ~n13244;
  assign n13246 = n13167 & n13228;
  assign n13247 = n13220 & n13227;
  assign n13248 = n13210 & n13240;
  assign n13249 = ~n13247 & ~n13248;
  assign n13250 = n13230 & ~n13249;
  assign n13251 = ~n13246 & ~n13250;
  assign n13252 = n13207 & n13230;
  assign n13253 = ~n13231 & n13243;
  assign n13254 = ~n13222 & n13253;
  assign n13255 = ~n13248 & n13254;
  assign n13256 = n13235 & ~n13255;
  assign n13257 = ~n13252 & ~n13256;
  assign n13258 = ~n13230 & ~n13235;
  assign n13259 = n13220 & n13240;
  assign n13260 = ~n13258 & n13259;
  assign n13261 = n13226 & n13240;
  assign n13262 = n13258 & n13261;
  assign n13263 = n13223 & ~n13231;
  assign n13264 = ~n13247 & n13263;
  assign n13265 = n13167 & ~n13264;
  assign n13266 = ~n13262 & ~n13265;
  assign n13267 = ~n13260 & n13266;
  assign n13268 = n13257 & n13267;
  assign n13269 = n13251 & n13268;
  assign n13270 = n13245 & n13269;
  assign n13271 = n13234 & n13270;
  assign n13272 = ~n13225 & n13271;
  assign n13273 = ~n13219 & n13272;
  assign n13274 = n13216 & n13273;
  assign n13275 = n13274 ^ n9838;
  assign n13276 = n13275 ^ x628;
  assign n13277 = n12421 ^ x574;
  assign n13278 = n12021 & n12027;
  assign n13279 = n12023 & n12029;
  assign n13280 = ~n13278 & ~n13279;
  assign n13281 = n12027 & n12045;
  assign n13282 = ~n12041 & ~n12774;
  assign n13283 = ~n12064 & n13282;
  assign n13284 = ~n12070 & n13283;
  assign n13285 = n12053 & n13284;
  assign n13286 = ~n12039 & n13285;
  assign n13287 = n11915 & ~n13286;
  assign n13288 = ~n13281 & ~n13287;
  assign n13289 = n12062 & ~n12074;
  assign n13290 = ~n12057 & n12075;
  assign n13291 = n12023 & ~n13290;
  assign n13292 = ~n12040 & ~n12774;
  assign n13293 = ~n12069 & n13292;
  assign n13294 = ~n12062 & n13293;
  assign n13295 = ~n12039 & n12776;
  assign n13296 = ~n12027 & n13295;
  assign n13297 = ~n13294 & ~n13296;
  assign n13298 = ~n12047 & ~n13297;
  assign n13299 = ~n11887 & ~n13298;
  assign n13300 = ~n13291 & ~n13299;
  assign n13301 = ~n13289 & n13300;
  assign n13302 = n13288 & n13301;
  assign n13303 = n12036 & n13302;
  assign n13304 = n12759 & n13303;
  assign n13305 = n13280 & n13304;
  assign n13306 = n13305 ^ n10220;
  assign n13307 = n13306 ^ x579;
  assign n13308 = n13277 & ~n13307;
  assign n13309 = n11818 & ~n11835;
  assign n13310 = ~n11842 & n13309;
  assign n13311 = n11793 & ~n13310;
  assign n13312 = ~n11801 & n12936;
  assign n13313 = n11824 & ~n13312;
  assign n13314 = ~n13311 & ~n13313;
  assign n13315 = n11826 & ~n11835;
  assign n13316 = ~n11791 & n13315;
  assign n13317 = ~n11834 & n12717;
  assign n13318 = ~n11798 & n13317;
  assign n13319 = ~n13316 & ~n13318;
  assign n13320 = ~n12716 & ~n13319;
  assign n13321 = n12699 & n13320;
  assign n13322 = ~n11812 & ~n13321;
  assign n13323 = n13314 & ~n13322;
  assign n13324 = n11806 & n13323;
  assign n13325 = n12698 & n13324;
  assign n13326 = n12928 & n13325;
  assign n13327 = ~n11825 & n13326;
  assign n13328 = n13327 ^ n9946;
  assign n13329 = n13328 ^ x578;
  assign n13330 = ~n11177 & n11344;
  assign n13331 = n11337 & n11348;
  assign n13332 = ~n13330 & ~n13331;
  assign n13333 = ~n11339 & n13007;
  assign n13334 = n11314 & ~n13333;
  assign n13335 = n11340 & n12807;
  assign n13336 = ~n11327 & n13335;
  assign n13337 = ~n11312 & n13336;
  assign n13338 = n11324 & ~n13337;
  assign n13339 = ~n13334 & ~n13338;
  assign n13340 = ~n11337 & ~n11358;
  assign n13341 = ~n11339 & n11375;
  assign n13342 = ~n13340 & ~n13341;
  assign n13343 = ~n11370 & ~n13342;
  assign n13344 = ~n11374 & n13343;
  assign n13345 = ~n11363 & ~n13344;
  assign n13346 = n13339 & ~n13345;
  assign n13347 = n13332 & n13346;
  assign n13348 = ~n11336 & n13347;
  assign n13349 = n13000 & n13348;
  assign n13350 = n12996 & n13349;
  assign n13351 = ~n11322 & n13350;
  assign n13352 = ~n12795 & n13351;
  assign n13353 = n11318 & n13352;
  assign n13354 = n13353 ^ n9981;
  assign n13355 = n13354 ^ x577;
  assign n13356 = ~n13329 & n13355;
  assign n13357 = n9839 & n11005;
  assign n13358 = ~n11000 & n12675;
  assign n13359 = n11036 & n13358;
  assign n13360 = ~n11031 & n13359;
  assign n13361 = n11007 & ~n13360;
  assign n13362 = ~n13357 & ~n13361;
  assign n13363 = ~n11002 & n11032;
  assign n13364 = n11020 & ~n13363;
  assign n13365 = ~n12657 & n12663;
  assign n13366 = n10288 & ~n13365;
  assign n13367 = ~n13364 & ~n13366;
  assign n13368 = ~n11008 & n12659;
  assign n13369 = n10992 & ~n13368;
  assign n13370 = ~n10985 & ~n11020;
  assign n13371 = n10986 & n10992;
  assign n13372 = n11017 & ~n13371;
  assign n13373 = ~n10994 & n13372;
  assign n13374 = ~n11008 & n13373;
  assign n13375 = ~n13370 & ~n13374;
  assign n13376 = n12656 & n13375;
  assign n13377 = ~n13369 & ~n13376;
  assign n13378 = n13367 & n13377;
  assign n13379 = n13362 & n13378;
  assign n13380 = n11012 & n13379;
  assign n13381 = n10998 & n13380;
  assign n13382 = n13381 ^ n10145;
  assign n13383 = n13382 ^ x576;
  assign n13384 = n12316 ^ x575;
  assign n13385 = n13383 & n13384;
  assign n13386 = n13356 & n13385;
  assign n13387 = n13329 & n13355;
  assign n13388 = ~n13383 & n13384;
  assign n13389 = n13387 & n13388;
  assign n13390 = ~n13386 & ~n13389;
  assign n13391 = n13308 & ~n13390;
  assign n13392 = ~n13329 & ~n13355;
  assign n13393 = ~n13383 & ~n13384;
  assign n13394 = n13392 & n13393;
  assign n13395 = ~n13277 & n13307;
  assign n13396 = ~n13308 & ~n13395;
  assign n13397 = n13394 & ~n13396;
  assign n13398 = n13277 & n13307;
  assign n13399 = n13329 & ~n13355;
  assign n13400 = n13385 & n13399;
  assign n13401 = n13398 & n13400;
  assign n13402 = ~n13277 & ~n13307;
  assign n13403 = n13388 & n13392;
  assign n13404 = n13402 & n13403;
  assign n13405 = n13383 & ~n13384;
  assign n13406 = n13399 & n13405;
  assign n13407 = ~n13396 & n13406;
  assign n13408 = ~n13404 & ~n13407;
  assign n13409 = ~n13401 & n13408;
  assign n13410 = ~n13397 & n13409;
  assign n13411 = n13356 & n13405;
  assign n13412 = ~n13396 & n13411;
  assign n13413 = n13393 & n13399;
  assign n13414 = n13308 & n13413;
  assign n13415 = n13387 & n13393;
  assign n13416 = n13395 & n13415;
  assign n13417 = ~n13414 & ~n13416;
  assign n13418 = ~n13412 & n13417;
  assign n13419 = n13385 & n13392;
  assign n13420 = n13308 & n13419;
  assign n13421 = n13398 & n13403;
  assign n13422 = ~n13420 & ~n13421;
  assign n13423 = ~n13394 & ~n13415;
  assign n13424 = n13402 & ~n13423;
  assign n13425 = n13422 & ~n13424;
  assign n13426 = n13308 & n13415;
  assign n13427 = n13356 & n13393;
  assign n13428 = n13384 ^ n13383;
  assign n13429 = n13355 ^ n13329;
  assign n13430 = n13429 ^ n13384;
  assign n13431 = n13428 & ~n13430;
  assign n13432 = ~n13389 & ~n13431;
  assign n13433 = ~n13427 & n13432;
  assign n13434 = n13398 & ~n13433;
  assign n13435 = ~n13426 & ~n13434;
  assign n13436 = n13392 & n13405;
  assign n13437 = ~n13413 & ~n13436;
  assign n13438 = n13402 & ~n13437;
  assign n13439 = n13356 & n13388;
  assign n13440 = n13385 & n13387;
  assign n13441 = ~n13439 & ~n13440;
  assign n13442 = ~n13395 & n13441;
  assign n13443 = ~n13400 & n13442;
  assign n13444 = n13388 & n13399;
  assign n13445 = ~n13439 & ~n13444;
  assign n13446 = ~n13386 & n13445;
  assign n13447 = ~n13419 & n13446;
  assign n13448 = n13395 & ~n13447;
  assign n13449 = ~n13402 & ~n13448;
  assign n13450 = ~n13443 & ~n13449;
  assign n13451 = ~n13438 & ~n13450;
  assign n13452 = n13435 & n13451;
  assign n13453 = n13425 & n13452;
  assign n13454 = n13418 & n13453;
  assign n13455 = n13410 & n13454;
  assign n13456 = ~n13391 & n13455;
  assign n13457 = n13456 ^ n10286;
  assign n13458 = n13457 ^ x633;
  assign n13459 = ~n13276 & ~n13458;
  assign n13460 = n13164 & n13459;
  assign n13461 = ~n12926 & n13162;
  assign n13462 = n12275 & ~n12654;
  assign n13463 = n13461 & n13462;
  assign n13464 = n13276 & ~n13458;
  assign n13465 = n13463 & n13464;
  assign n13466 = ~n13460 & ~n13465;
  assign n13467 = ~n13276 & n13458;
  assign n13468 = n13463 & n13467;
  assign n13469 = n13276 & n13458;
  assign n13470 = n12926 & ~n13162;
  assign n13471 = n12655 & n13470;
  assign n13472 = n13469 & n13471;
  assign n13473 = ~n13468 & ~n13472;
  assign n13474 = n12655 & n13461;
  assign n13475 = n13467 & n13474;
  assign n13476 = n12275 & n12654;
  assign n13477 = n13461 & n13476;
  assign n13478 = n13464 & n13477;
  assign n13479 = ~n13475 & ~n13478;
  assign n13480 = n12926 & n13162;
  assign n13481 = n13462 & n13480;
  assign n13482 = n13163 & n13462;
  assign n13483 = ~n12275 & ~n12654;
  assign n13484 = n13470 & n13483;
  assign n13485 = ~n13482 & ~n13484;
  assign n13486 = ~n13481 & n13485;
  assign n13487 = n13459 & ~n13486;
  assign n13488 = n13470 & n13476;
  assign n13489 = ~n13471 & ~n13488;
  assign n13490 = ~n13464 & ~n13467;
  assign n13491 = ~n13489 & ~n13490;
  assign n13492 = n13480 & n13483;
  assign n13493 = n13461 & n13483;
  assign n13494 = n13462 & n13470;
  assign n13495 = n13163 & n13483;
  assign n13496 = ~n13494 & ~n13495;
  assign n13497 = ~n13493 & n13496;
  assign n13498 = ~n13492 & n13497;
  assign n13499 = ~n13490 & ~n13498;
  assign n13500 = n13476 & n13480;
  assign n13501 = ~n13474 & ~n13500;
  assign n13502 = n12655 & n13480;
  assign n13503 = n13163 & n13476;
  assign n13504 = ~n13502 & ~n13503;
  assign n13505 = n13501 & n13504;
  assign n13506 = n13459 & ~n13505;
  assign n13507 = ~n13164 & ~n13493;
  assign n13508 = ~n13477 & ~n13502;
  assign n13509 = n13486 & n13508;
  assign n13510 = n13507 & n13509;
  assign n13511 = n13469 & ~n13510;
  assign n13512 = ~n13506 & ~n13511;
  assign n13513 = ~n13499 & n13512;
  assign n13514 = ~n13491 & n13513;
  assign n13515 = ~n13487 & n13514;
  assign n13516 = n13479 & n13515;
  assign n13517 = n13473 & n13516;
  assign n13518 = n13466 & n13517;
  assign n13519 = n13518 ^ n12689;
  assign n13520 = n13519 ^ x649;
  assign n13521 = ~n13222 & ~n13259;
  assign n13522 = n13167 & ~n13521;
  assign n13523 = n13209 & n13248;
  assign n13524 = ~n13213 & ~n13221;
  assign n13525 = n13167 & ~n13524;
  assign n13526 = ~n13523 & ~n13525;
  assign n13527 = ~n13211 & ~n13231;
  assign n13528 = n13249 & n13527;
  assign n13529 = n13235 & ~n13528;
  assign n13530 = n13167 & n13236;
  assign n13531 = ~n13228 & ~n13241;
  assign n13532 = ~n13218 & n13531;
  assign n13533 = n13167 & ~n13532;
  assign n13534 = ~n13236 & n13243;
  assign n13535 = n13209 & ~n13534;
  assign n13536 = ~n13533 & ~n13535;
  assign n13537 = ~n13237 & ~n13261;
  assign n13538 = ~n13218 & n13537;
  assign n13539 = ~n13241 & n13538;
  assign n13540 = n13230 & ~n13539;
  assign n13541 = ~n13259 & n13527;
  assign n13542 = ~n13247 & n13541;
  assign n13543 = n13230 & ~n13542;
  assign n13544 = ~n13242 & n13538;
  assign n13545 = n13235 & ~n13544;
  assign n13546 = ~n13543 & ~n13545;
  assign n13547 = ~n13540 & n13546;
  assign n13548 = n13536 & n13547;
  assign n13549 = ~n13530 & n13548;
  assign n13550 = ~n13229 & n13549;
  assign n13551 = ~n13529 & n13550;
  assign n13552 = n13526 & n13551;
  assign n13553 = ~n13522 & n13552;
  assign n13554 = ~n13225 & n13553;
  assign n13555 = n13554 ^ n11886;
  assign n13556 = n13555 ^ x616;
  assign n13557 = n13028 & n13115;
  assign n13558 = n13110 & n13112;
  assign n13559 = n13115 & n13138;
  assign n13560 = ~n13558 & ~n13559;
  assign n13561 = ~n13557 & n13560;
  assign n13562 = n13098 & n13112;
  assign n13563 = n13110 & n13113;
  assign n13564 = ~n13562 & ~n13563;
  assign n13565 = ~n13120 & ~n13136;
  assign n13566 = n13110 & ~n13565;
  assign n13567 = ~n13098 & ~n13110;
  assign n13568 = n13118 & ~n13567;
  assign n13569 = ~n13566 & ~n13568;
  assign n13570 = ~n13121 & ~n13138;
  assign n13571 = n13093 & ~n13570;
  assign n13572 = ~n13102 & ~n13131;
  assign n13573 = n13092 & ~n13572;
  assign n13574 = ~n13571 & ~n13573;
  assign n13575 = n13108 & n13133;
  assign n13576 = n13115 & ~n13575;
  assign n13577 = ~n13104 & ~n13132;
  assign n13578 = ~n13143 & n13577;
  assign n13579 = ~n13098 & n13578;
  assign n13580 = ~n13121 & ~n13143;
  assign n13581 = ~n13136 & n13580;
  assign n13582 = ~n13093 & n13581;
  assign n13583 = ~n13579 & ~n13582;
  assign n13584 = n13092 & n13583;
  assign n13585 = ~n13576 & ~n13584;
  assign n13586 = n13574 & n13585;
  assign n13587 = n13569 & n13586;
  assign n13588 = n13564 & n13587;
  assign n13589 = n13561 & n13588;
  assign n13590 = n13117 & n13589;
  assign n13591 = n13100 & n13590;
  assign n13592 = n13591 ^ n11913;
  assign n13593 = n13592 ^ x621;
  assign n13594 = n13556 & ~n13593;
  assign n13595 = n12875 & ~n12899;
  assign n13596 = ~n12878 & ~n12893;
  assign n13597 = n12876 & ~n13596;
  assign n13598 = ~n13595 & ~n13597;
  assign n13599 = n12863 & ~n12913;
  assign n13600 = n12904 & ~n12911;
  assign n13601 = ~n12867 & n13600;
  assign n13602 = n12885 & ~n13601;
  assign n13603 = ~n12879 & ~n12900;
  assign n13604 = ~n12883 & n13603;
  assign n13605 = ~n12908 & n13604;
  assign n13606 = n12871 & ~n13605;
  assign n13607 = n12887 & ~n12908;
  assign n13608 = ~n12883 & n13607;
  assign n13609 = n12876 & ~n13608;
  assign n13610 = ~n13606 & ~n13609;
  assign n13611 = n12794 & ~n12883;
  assign n13612 = ~n12901 & n13611;
  assign n13613 = n12863 & ~n13612;
  assign n13614 = ~n12869 & n13596;
  assign n13615 = ~n12875 & n13614;
  assign n13616 = n12871 & ~n13615;
  assign n13617 = ~n12790 & n13607;
  assign n13618 = n12885 & ~n13617;
  assign n13619 = ~n13616 & ~n13618;
  assign n13620 = ~n13613 & n13619;
  assign n13621 = n13610 & n13620;
  assign n13622 = ~n13602 & n13621;
  assign n13623 = ~n13599 & n13622;
  assign n13624 = n13598 & n13623;
  assign n13625 = n12895 & n13624;
  assign n13626 = n13625 ^ n11950;
  assign n13627 = n13626 ^ x618;
  assign n13628 = n13387 & n13405;
  assign n13629 = n13308 & n13628;
  assign n13630 = n13398 & ~n13445;
  assign n13631 = ~n13629 & ~n13630;
  assign n13632 = ~n13411 & ~n13419;
  assign n13633 = n13402 & ~n13632;
  assign n13634 = ~n13419 & ~n13440;
  assign n13635 = n13390 & n13634;
  assign n13636 = ~n13413 & n13635;
  assign n13637 = n13395 & ~n13636;
  assign n13638 = ~n13415 & ~n13431;
  assign n13639 = n13402 & ~n13638;
  assign n13640 = ~n13637 & ~n13639;
  assign n13641 = n13307 & n13427;
  assign n13642 = ~n13400 & n13445;
  assign n13643 = n13308 & ~n13642;
  assign n13644 = ~n13406 & n13423;
  assign n13645 = ~n13386 & n13644;
  assign n13646 = n13398 & ~n13645;
  assign n13647 = ~n13643 & ~n13646;
  assign n13648 = ~n13641 & n13647;
  assign n13649 = n13640 & n13648;
  assign n13650 = ~n13633 & n13649;
  assign n13651 = n13631 & n13650;
  assign n13652 = n13410 & n13651;
  assign n13653 = ~n13391 & n13652;
  assign n13654 = n13653 ^ n11982;
  assign n13655 = n13654 ^ x619;
  assign n13656 = ~n12243 & n12259;
  assign n13657 = n11392 & n12257;
  assign n13658 = ~n13656 & ~n13657;
  assign n13659 = ~n12232 & n12246;
  assign n13660 = n12234 & ~n12270;
  assign n13661 = ~n13659 & ~n13660;
  assign n13662 = n13658 & n13661;
  assign n13663 = n13662 ^ n11923;
  assign n13664 = n13663 ^ x620;
  assign n13665 = n12993 ^ x544;
  assign n13666 = n12755 ^ x549;
  assign n13667 = n13665 & n13666;
  assign n13668 = n12065 & n13283;
  assign n13669 = ~n12069 & n13668;
  assign n13670 = n12023 & ~n13669;
  assign n13671 = n12053 & n12065;
  assign n13672 = ~n12774 & n13671;
  assign n13673 = n12062 & ~n13672;
  assign n13674 = ~n13670 & ~n13673;
  assign n13675 = ~n11887 & n12040;
  assign n13676 = ~n12029 & n12076;
  assign n13677 = n12027 & ~n13676;
  assign n13678 = ~n12025 & n12077;
  assign n13679 = n11915 & ~n13678;
  assign n13680 = ~n13677 & ~n13679;
  assign n13681 = ~n13675 & n13680;
  assign n13682 = n13674 & n13681;
  assign n13683 = ~n12044 & n13682;
  assign n13684 = n12766 & n13683;
  assign n13685 = n13280 & n13684;
  assign n13686 = n13685 ^ n11459;
  assign n13687 = n13686 ^ x547;
  assign n13688 = ~n12172 & ~n12193;
  assign n13689 = n12161 & ~n13688;
  assign n13690 = ~n12205 & ~n12209;
  assign n13691 = ~n12090 & ~n13690;
  assign n13692 = ~n13689 & ~n13691;
  assign n13693 = n12188 & ~n12562;
  assign n13694 = ~n12164 & n12571;
  assign n13695 = n12177 & ~n13694;
  assign n13696 = n12180 & ~n13061;
  assign n13697 = ~n12155 & ~n12178;
  assign n13698 = ~n12188 & n13697;
  assign n13699 = ~n13696 & ~n13698;
  assign n13700 = n13063 & ~n13699;
  assign n13701 = ~n12201 & ~n13700;
  assign n13702 = ~n13695 & ~n13701;
  assign n13703 = ~n13693 & n13702;
  assign n13704 = n13692 & n13703;
  assign n13705 = ~n12560 & n13704;
  assign n13706 = ~n12187 & n13705;
  assign n13707 = ~n12558 & n13706;
  assign n13708 = n12167 & n13707;
  assign n13709 = n13067 & n13708;
  assign n13710 = n13709 ^ n11486;
  assign n13711 = n13710 ^ x546;
  assign n13712 = ~n13687 & n13711;
  assign n13713 = n13059 ^ x545;
  assign n13714 = n12861 ^ x548;
  assign n13715 = ~n13713 & ~n13714;
  assign n13716 = n13712 & n13715;
  assign n13717 = n13667 & n13716;
  assign n13718 = ~n13665 & n13666;
  assign n13719 = ~n13713 & n13714;
  assign n13720 = n13712 & n13719;
  assign n13721 = n13718 & n13720;
  assign n13722 = n13665 & ~n13666;
  assign n13723 = n13687 & ~n13711;
  assign n13724 = n13719 & n13723;
  assign n13725 = ~n13716 & ~n13724;
  assign n13726 = n13722 & ~n13725;
  assign n13727 = ~n13721 & ~n13726;
  assign n13728 = ~n13665 & ~n13666;
  assign n13729 = ~n13687 & ~n13711;
  assign n13730 = n13719 & n13729;
  assign n13731 = ~n13716 & ~n13730;
  assign n13732 = n13728 & ~n13731;
  assign n13733 = n13687 & n13711;
  assign n13734 = n13719 & n13733;
  assign n13735 = n13715 & n13729;
  assign n13736 = ~n13734 & ~n13735;
  assign n13737 = n13667 & ~n13736;
  assign n13738 = n13715 & n13733;
  assign n13739 = ~n13720 & ~n13738;
  assign n13740 = n13728 & ~n13739;
  assign n13741 = ~n13737 & ~n13740;
  assign n13742 = n13665 & n13730;
  assign n13743 = n13713 & ~n13714;
  assign n13744 = n13712 & n13743;
  assign n13745 = n13723 & n13743;
  assign n13746 = ~n13744 & ~n13745;
  assign n13747 = n13713 & n13714;
  assign n13748 = n13712 & n13747;
  assign n13749 = n13733 & n13743;
  assign n13750 = ~n13748 & ~n13749;
  assign n13751 = n13729 & n13747;
  assign n13752 = n13715 & n13723;
  assign n13753 = ~n13734 & ~n13752;
  assign n13754 = ~n13751 & n13753;
  assign n13755 = n13750 & n13754;
  assign n13756 = n13746 & n13755;
  assign n13757 = n13718 & ~n13756;
  assign n13758 = ~n13742 & ~n13757;
  assign n13759 = n13733 & n13747;
  assign n13760 = n13729 & n13743;
  assign n13761 = ~n13759 & ~n13760;
  assign n13762 = n13750 & n13761;
  assign n13763 = ~n13720 & n13762;
  assign n13764 = n13722 & ~n13763;
  assign n13765 = n13723 & n13747;
  assign n13766 = ~n13667 & n13746;
  assign n13767 = ~n13759 & n13766;
  assign n13768 = ~n13765 & n13767;
  assign n13769 = ~n13749 & n13761;
  assign n13770 = ~n13765 & n13769;
  assign n13771 = n13667 & ~n13770;
  assign n13772 = ~n13728 & ~n13771;
  assign n13773 = ~n13768 & ~n13772;
  assign n13774 = ~n13764 & ~n13773;
  assign n13775 = n13758 & n13774;
  assign n13776 = n13741 & n13775;
  assign n13777 = ~n13732 & n13776;
  assign n13778 = n13727 & n13777;
  assign n13779 = ~n13717 & n13778;
  assign n13780 = n13779 ^ n12018;
  assign n13781 = n13780 ^ x617;
  assign n13782 = n13664 & ~n13781;
  assign n13783 = ~n13655 & n13782;
  assign n13784 = n13627 & n13783;
  assign n13785 = n13594 & n13784;
  assign n13786 = n13556 & n13593;
  assign n13787 = ~n13627 & n13655;
  assign n13788 = n13664 & n13781;
  assign n13789 = n13787 & n13788;
  assign n13790 = n13786 & n13789;
  assign n13791 = ~n13556 & n13593;
  assign n13792 = n13627 & n13655;
  assign n13793 = ~n13664 & ~n13781;
  assign n13794 = n13792 & n13793;
  assign n13795 = n13791 & n13794;
  assign n13796 = ~n13556 & ~n13593;
  assign n13797 = n13627 & ~n13655;
  assign n13798 = ~n13664 & n13781;
  assign n13799 = n13797 & n13798;
  assign n13800 = ~n13789 & ~n13799;
  assign n13801 = n13796 & ~n13800;
  assign n13802 = ~n13795 & ~n13801;
  assign n13803 = ~n13790 & n13802;
  assign n13804 = n13782 & n13787;
  assign n13805 = ~n13627 & ~n13655;
  assign n13806 = n13793 & n13805;
  assign n13807 = ~n13804 & ~n13806;
  assign n13808 = n13791 & ~n13807;
  assign n13809 = n13798 & n13805;
  assign n13810 = n13594 & n13809;
  assign n13811 = n13782 & n13792;
  assign n13812 = n13786 & n13811;
  assign n13813 = ~n13810 & ~n13812;
  assign n13814 = n13788 & n13805;
  assign n13815 = n13556 & n13814;
  assign n13816 = n13788 & n13792;
  assign n13817 = n13792 & n13798;
  assign n13818 = ~n13794 & ~n13809;
  assign n13819 = n13796 & ~n13818;
  assign n13820 = n13787 & n13793;
  assign n13821 = ~n13806 & ~n13820;
  assign n13822 = n13786 & ~n13821;
  assign n13823 = ~n13819 & ~n13822;
  assign n13824 = ~n13783 & n13823;
  assign n13825 = ~n13817 & n13824;
  assign n13826 = ~n13816 & n13825;
  assign n13827 = n13796 & ~n13826;
  assign n13828 = ~n13815 & ~n13827;
  assign n13829 = n13788 & n13797;
  assign n13830 = n13787 & n13798;
  assign n13831 = ~n13789 & ~n13830;
  assign n13832 = ~n13627 & n13783;
  assign n13833 = n13831 & ~n13832;
  assign n13834 = ~n13817 & n13833;
  assign n13835 = ~n13829 & n13834;
  assign n13836 = n13791 & ~n13835;
  assign n13837 = ~n13816 & ~n13830;
  assign n13838 = n13793 & n13797;
  assign n13839 = ~n13811 & ~n13838;
  assign n13840 = ~n13804 & n13839;
  assign n13841 = n13837 & n13840;
  assign n13842 = n13594 & ~n13841;
  assign n13843 = ~n13799 & n13824;
  assign n13844 = n13786 & ~n13843;
  assign n13845 = ~n13842 & ~n13844;
  assign n13846 = ~n13836 & n13845;
  assign n13847 = n13828 & n13846;
  assign n13848 = n13813 & n13847;
  assign n13849 = ~n13808 & n13848;
  assign n13850 = n13803 & n13849;
  assign n13851 = ~n13785 & n13850;
  assign n13852 = n13851 ^ n12787;
  assign n13853 = n13852 ^ x650;
  assign n13854 = n13520 & n13853;
  assign n13855 = n12262 & n12265;
  assign n13856 = ~n11856 & n12237;
  assign n13857 = ~n12224 & n12227;
  assign n13858 = ~n11634 & n12248;
  assign n13859 = ~n13857 & ~n13858;
  assign n13860 = ~n13856 & n13859;
  assign n13861 = n11392 & ~n13860;
  assign n13862 = n12087 & n12224;
  assign n13863 = ~n11634 & n13862;
  assign n13864 = n11634 & n13856;
  assign n13865 = ~n12087 & n12262;
  assign n13866 = ~n13864 & ~n13865;
  assign n13867 = ~n13863 & n13866;
  assign n13868 = ~n12238 & n13867;
  assign n13869 = n12234 & ~n13868;
  assign n13870 = ~n13861 & ~n13869;
  assign n13871 = ~n12087 & n12227;
  assign n13872 = n11634 & n12248;
  assign n13873 = n12224 & n13872;
  assign n13874 = ~n13871 & ~n13873;
  assign n13875 = ~n11634 & ~n12266;
  assign n13876 = n13874 & ~n13875;
  assign n13877 = ~n12261 & n13876;
  assign n13878 = n12246 & ~n13877;
  assign n13879 = n12224 & n12262;
  assign n13880 = n11634 & ~n12254;
  assign n13881 = ~n13879 & ~n13880;
  assign n13882 = ~n12261 & n13881;
  assign n13883 = n12259 & ~n13882;
  assign n13884 = ~n13878 & ~n13883;
  assign n13885 = n13870 & n13884;
  assign n13886 = ~n13855 & n13885;
  assign n13887 = n13886 ^ n11205;
  assign n13888 = n13887 ^ x639;
  assign n13889 = n12925 ^ x634;
  assign n13890 = ~n13888 & n13889;
  assign n13891 = n13718 & n13759;
  assign n13892 = ~n13745 & n13750;
  assign n13893 = n13728 & ~n13892;
  assign n13894 = ~n13891 & ~n13893;
  assign n13895 = ~n13717 & n13894;
  assign n13896 = ~n13745 & ~n13748;
  assign n13897 = n13667 & ~n13896;
  assign n13898 = n13728 & n13759;
  assign n13899 = ~n13716 & ~n13720;
  assign n13900 = n13718 & ~n13899;
  assign n13901 = ~n13898 & ~n13900;
  assign n13902 = n13728 & ~n13736;
  assign n13903 = ~n13724 & ~n13738;
  assign n13904 = ~n13749 & ~n13751;
  assign n13905 = ~n13744 & n13904;
  assign n13906 = n13903 & n13905;
  assign n13907 = ~n13745 & n13906;
  assign n13908 = n13722 & ~n13907;
  assign n13909 = ~n13902 & ~n13908;
  assign n13910 = ~n13735 & n13905;
  assign n13911 = ~n13724 & n13910;
  assign n13912 = n13718 & ~n13911;
  assign n13913 = ~n13720 & ~n13760;
  assign n13914 = n13665 & ~n13913;
  assign n13915 = n13753 & ~n13765;
  assign n13916 = n13667 & ~n13915;
  assign n13917 = ~n13914 & ~n13916;
  assign n13918 = ~n13912 & n13917;
  assign n13919 = n13909 & n13918;
  assign n13920 = n13901 & n13919;
  assign n13921 = ~n13897 & n13920;
  assign n13922 = ~n13732 & n13921;
  assign n13923 = n13895 & n13922;
  assign n13924 = n13923 ^ n11559;
  assign n13925 = n13924 ^ x637;
  assign n13926 = n13328 ^ x580;
  assign n13927 = n12976 ^ x585;
  assign n13928 = n13926 & ~n13927;
  assign n13929 = ~n12386 & n12411;
  assign n13930 = n12388 & ~n12409;
  assign n13931 = ~n13929 & ~n13930;
  assign n13932 = ~n12401 & n12404;
  assign n13933 = n12321 & n12417;
  assign n13934 = ~n13932 & ~n13933;
  assign n13935 = n13931 & n13934;
  assign n13936 = n13935 ^ n11057;
  assign n13937 = n13936 ^ x582;
  assign n13938 = n13306 ^ x581;
  assign n13939 = ~n13937 & ~n13938;
  assign n13940 = n11395 & n11589;
  assign n13941 = ~n11599 & n11610;
  assign n13942 = ~n13940 & ~n13941;
  assign n13943 = n11563 & ~n12299;
  assign n13944 = ~n11588 & ~n11601;
  assign n13945 = n11394 & ~n13944;
  assign n13946 = ~n11574 & ~n11588;
  assign n13947 = ~n11570 & n13946;
  assign n13948 = n11578 & ~n13947;
  assign n13949 = ~n13945 & ~n13948;
  assign n13950 = ~n13943 & n13949;
  assign n13951 = n13942 & n13950;
  assign n13952 = n12737 & n13951;
  assign n13953 = n11568 & n13952;
  assign n13954 = n12734 & n13953;
  assign n13955 = n12297 & n13954;
  assign n13956 = n12280 & n13955;
  assign n13957 = n12292 & n13956;
  assign n13958 = ~n11598 & n13957;
  assign n13959 = n13958 ^ n11078;
  assign n13960 = n13959 ^ x583;
  assign n13961 = n13091 ^ x584;
  assign n13962 = ~n13960 & n13961;
  assign n13963 = n13939 & n13962;
  assign n13964 = n13928 & n13963;
  assign n13965 = ~n13937 & n13938;
  assign n13966 = n13961 & n13965;
  assign n13967 = n13960 & n13966;
  assign n13968 = n13937 & n13938;
  assign n13969 = n13960 & ~n13961;
  assign n13970 = n13968 & n13969;
  assign n13971 = ~n13967 & ~n13970;
  assign n13972 = n13928 & ~n13971;
  assign n13973 = ~n13926 & n13927;
  assign n13974 = n13962 & n13968;
  assign n13975 = ~n13960 & ~n13961;
  assign n13976 = n13965 & n13975;
  assign n13977 = ~n13974 & ~n13976;
  assign n13978 = n13973 & ~n13977;
  assign n13979 = ~n13972 & ~n13978;
  assign n13980 = ~n13960 & n13966;
  assign n13981 = n13928 & n13980;
  assign n13982 = ~n13928 & ~n13973;
  assign n13983 = n13939 & n13969;
  assign n13984 = ~n13982 & n13983;
  assign n13985 = ~n13981 & ~n13984;
  assign n13986 = n13926 & n13927;
  assign n13987 = n13965 & n13969;
  assign n13988 = ~n13970 & ~n13987;
  assign n13989 = ~n13980 & n13988;
  assign n13990 = n13986 & ~n13989;
  assign n13991 = n13937 & ~n13938;
  assign n13992 = n13975 & n13991;
  assign n13993 = n13926 & n13992;
  assign n13994 = n13960 & n13961;
  assign n13995 = n13939 & n13994;
  assign n13996 = n13939 & n13975;
  assign n13997 = ~n13995 & ~n13996;
  assign n13998 = ~n13963 & n13997;
  assign n13999 = ~n13974 & n13998;
  assign n14000 = n13986 & ~n13999;
  assign n14001 = ~n13993 & ~n14000;
  assign n14002 = ~n13926 & ~n13927;
  assign n14003 = ~n13970 & ~n13974;
  assign n14004 = ~n13980 & n14003;
  assign n14005 = n13962 & n13991;
  assign n14006 = n13991 & n13994;
  assign n14007 = ~n13996 & ~n14006;
  assign n14008 = ~n14005 & n14007;
  assign n14009 = ~n13983 & n14008;
  assign n14010 = n14004 & n14009;
  assign n14011 = ~n13995 & n14010;
  assign n14012 = n14002 & n14011;
  assign n14013 = ~n13976 & ~n14005;
  assign n14014 = n13928 & ~n14013;
  assign n14015 = n13971 & n14008;
  assign n14016 = n13973 & ~n14015;
  assign n14017 = ~n14014 & ~n14016;
  assign n14018 = ~n14012 & n14017;
  assign n14019 = n14001 & n14018;
  assign n14020 = ~n13990 & n14019;
  assign n14021 = n13985 & n14020;
  assign n14022 = n13979 & n14021;
  assign n14023 = ~n13964 & n14022;
  assign n14024 = n14023 ^ n11142;
  assign n14025 = n14024 ^ x638;
  assign n14026 = ~n13925 & n14025;
  assign n14027 = ~n13214 & ~n13258;
  assign n14028 = n13245 & ~n14027;
  assign n14029 = ~n13242 & ~n13259;
  assign n14030 = ~n13207 & n14029;
  assign n14031 = n13249 & n14030;
  assign n14032 = n13209 & ~n14031;
  assign n14033 = ~n13218 & n13223;
  assign n14034 = ~n13248 & n14033;
  assign n14035 = n13235 & ~n14034;
  assign n14036 = ~n14032 & ~n14035;
  assign n14037 = n13230 & ~n13238;
  assign n14038 = n13167 & ~n13255;
  assign n14039 = ~n14037 & ~n14038;
  assign n14040 = n14036 & n14039;
  assign n14041 = n13251 & n14040;
  assign n14042 = n13216 & n14041;
  assign n14043 = n14028 & n14042;
  assign n14044 = ~n13530 & n14043;
  assign n14045 = ~n13229 & n14044;
  assign n14046 = n14045 ^ n11425;
  assign n14047 = n14046 ^ x636;
  assign n14048 = n13457 ^ x635;
  assign n14049 = ~n14047 & n14048;
  assign n14050 = n14026 & n14049;
  assign n14051 = n13890 & n14050;
  assign n14052 = ~n13888 & ~n13889;
  assign n14053 = n13925 & ~n14025;
  assign n14054 = n14049 & n14053;
  assign n14055 = n13925 & n14025;
  assign n14056 = n14047 & n14048;
  assign n14057 = n14055 & n14056;
  assign n14058 = ~n14054 & ~n14057;
  assign n14059 = n14052 & ~n14058;
  assign n14060 = ~n14051 & ~n14059;
  assign n14061 = n13888 & ~n13889;
  assign n14062 = ~n14058 & n14061;
  assign n14063 = n13888 & n13889;
  assign n14064 = n14053 & n14056;
  assign n14065 = n14049 & n14055;
  assign n14066 = ~n14064 & ~n14065;
  assign n14067 = n14063 & ~n14066;
  assign n14068 = ~n13925 & ~n14025;
  assign n14069 = n14047 & ~n14048;
  assign n14070 = n14068 & n14069;
  assign n14071 = ~n14047 & ~n14048;
  assign n14072 = n14026 & n14071;
  assign n14073 = ~n14070 & ~n14072;
  assign n14074 = n14055 & n14069;
  assign n14075 = n14055 & n14071;
  assign n14076 = ~n14074 & ~n14075;
  assign n14077 = n14073 & n14076;
  assign n14078 = n14052 & ~n14077;
  assign n14079 = ~n14052 & ~n14063;
  assign n14080 = n14026 & n14056;
  assign n14081 = n14056 & n14068;
  assign n14082 = ~n14080 & ~n14081;
  assign n14083 = ~n14079 & ~n14082;
  assign n14084 = n14073 & ~n14075;
  assign n14085 = n14063 & ~n14084;
  assign n14086 = n14049 & n14068;
  assign n14087 = ~n14080 & ~n14086;
  assign n14088 = n14053 & n14071;
  assign n14089 = ~n14064 & ~n14088;
  assign n14090 = n14076 & n14089;
  assign n14091 = n14087 & n14090;
  assign n14092 = n13890 & ~n14091;
  assign n14093 = ~n14085 & ~n14092;
  assign n14094 = ~n14083 & n14093;
  assign n14095 = ~n13890 & ~n14063;
  assign n14096 = n14068 & n14071;
  assign n14097 = ~n14095 & n14096;
  assign n14098 = n14026 & n14069;
  assign n14099 = n14053 & n14069;
  assign n14100 = ~n14074 & ~n14096;
  assign n14101 = ~n14099 & n14100;
  assign n14102 = ~n14098 & n14101;
  assign n14103 = ~n14081 & n14102;
  assign n14104 = ~n14050 & n14103;
  assign n14105 = n14061 & ~n14104;
  assign n14106 = ~n14097 & ~n14105;
  assign n14107 = n14094 & n14106;
  assign n14108 = ~n14078 & n14107;
  assign n14109 = ~n14067 & n14108;
  assign n14110 = ~n14062 & n14109;
  assign n14111 = n14060 & n14110;
  assign n14112 = n14111 ^ n12755;
  assign n14113 = n14112 ^ x647;
  assign n14114 = n12871 & n12879;
  assign n14115 = n12863 & n12891;
  assign n14116 = ~n14114 & ~n14115;
  assign n14117 = n12869 & n12885;
  assign n14118 = n12871 & n12893;
  assign n14119 = ~n14117 & ~n14118;
  assign n14120 = ~n12898 & n14119;
  assign n14121 = n12876 & n12912;
  assign n14122 = n12871 & n12901;
  assign n14123 = ~n14121 & ~n14122;
  assign n14124 = n12863 & ~n12887;
  assign n14125 = ~n12790 & ~n12912;
  assign n14126 = ~n12883 & n14125;
  assign n14127 = n12871 & ~n14126;
  assign n14128 = ~n14124 & ~n14127;
  assign n14129 = n12885 & n12893;
  assign n14130 = ~n12875 & ~n12911;
  assign n14131 = ~n12878 & n14130;
  assign n14132 = ~n12899 & ~n14131;
  assign n14133 = ~n12879 & n13611;
  assign n14134 = ~n12885 & n14133;
  assign n14135 = n12728 ^ n12690;
  assign n14136 = n14135 ^ n12788;
  assign n14137 = n12756 & n14136;
  assign n14138 = ~n12876 & ~n14137;
  assign n14139 = ~n14134 & ~n14138;
  assign n14140 = n12862 & n14139;
  assign n14141 = ~n14132 & ~n14140;
  assign n14142 = ~n14129 & n14141;
  assign n14143 = n14128 & n14142;
  assign n14144 = n14123 & n14143;
  assign n14145 = n14120 & n14144;
  assign n14146 = n14116 & n14145;
  assign n14147 = n12873 & n14146;
  assign n14148 = n14147 ^ n11789;
  assign n14149 = n14148 ^ x609;
  assign n14150 = ~n12625 & ~n12637;
  assign n14151 = n12592 & ~n14150;
  assign n14152 = n12318 & n12622;
  assign n14153 = n12590 & n12598;
  assign n14154 = n12609 & n12626;
  assign n14155 = ~n14153 & ~n14154;
  assign n14156 = ~n14152 & n14155;
  assign n14157 = n12621 & n12625;
  assign n14158 = n12592 & ~n12618;
  assign n14159 = ~n14157 & ~n14158;
  assign n14160 = n12318 & ~n12635;
  assign n14161 = n12588 & n12592;
  assign n14162 = n12590 & n12611;
  assign n14163 = ~n14161 & ~n14162;
  assign n14164 = ~n12602 & ~n12631;
  assign n14165 = n12592 & ~n14164;
  assign n14166 = ~n12626 & n12638;
  assign n14167 = n12318 & ~n14166;
  assign n14168 = ~n14165 & ~n14167;
  assign n14169 = n12590 & ~n12634;
  assign n14170 = ~n12603 & ~n12616;
  assign n14171 = ~n12632 & n14170;
  assign n14172 = ~n12594 & n14171;
  assign n14173 = n12609 & ~n14172;
  assign n14174 = ~n14169 & ~n14173;
  assign n14175 = n14168 & n14174;
  assign n14176 = n14163 & n14175;
  assign n14177 = n12608 & n14176;
  assign n14178 = ~n14160 & n14177;
  assign n14179 = n14159 & n14178;
  assign n14180 = n14156 & n14179;
  assign n14181 = ~n14151 & n14180;
  assign n14182 = ~n12614 & n14181;
  assign n14183 = n14182 ^ n11764;
  assign n14184 = n14183 ^ x604;
  assign n14185 = n14149 & n14184;
  assign n14186 = n12259 & n13868;
  assign n14187 = n11392 & n13877;
  assign n14188 = ~n14186 & ~n14187;
  assign n14189 = ~n13855 & n13860;
  assign n14190 = n12246 & ~n14189;
  assign n14191 = n12234 & ~n13882;
  assign n14192 = ~n14190 & ~n14191;
  assign n14193 = n14188 & n14192;
  assign n14194 = n14193 ^ n11644;
  assign n14195 = n14194 ^ x606;
  assign n14196 = n13968 & n13975;
  assign n14197 = n13982 & n14196;
  assign n14198 = ~n13974 & ~n13987;
  assign n14199 = ~n13976 & n14198;
  assign n14200 = ~n13995 & n14199;
  assign n14201 = n13973 & ~n14200;
  assign n14202 = n13928 & n14011;
  assign n14203 = ~n14201 & ~n14202;
  assign n14204 = n13971 & ~n13980;
  assign n14205 = n14002 & ~n14204;
  assign n14206 = n13961 ^ n13960;
  assign n14207 = n13938 & n14206;
  assign n14208 = n14207 ^ n14206;
  assign n14209 = ~n13926 & n14208;
  assign n14210 = n13986 & ~n14009;
  assign n14211 = ~n14209 & ~n14210;
  assign n14212 = ~n14205 & n14211;
  assign n14213 = n14203 & n14212;
  assign n14214 = ~n13990 & n14213;
  assign n14215 = ~n14197 & n14214;
  assign n14216 = n14215 ^ n11700;
  assign n14217 = n14216 ^ x608;
  assign n14218 = n14195 & n14217;
  assign n14219 = n13728 & n13730;
  assign n14220 = ~n13730 & ~n13752;
  assign n14221 = n13718 & ~n14220;
  assign n14222 = ~n14219 & ~n14221;
  assign n14223 = ~n13760 & n13903;
  assign n14224 = n13728 & ~n14223;
  assign n14225 = n13736 & ~n13765;
  assign n14226 = n13718 & ~n14225;
  assign n14227 = ~n14224 & ~n14226;
  assign n14228 = n13722 & ~n13755;
  assign n14229 = n13739 & n13761;
  assign n14230 = ~n13730 & n14229;
  assign n14231 = ~n13745 & n14230;
  assign n14232 = n13667 & ~n14231;
  assign n14233 = ~n14228 & ~n14232;
  assign n14234 = n14227 & n14233;
  assign n14235 = n13727 & n14234;
  assign n14236 = n14222 & n14235;
  assign n14237 = n13895 & n14236;
  assign n14238 = ~n13744 & n14237;
  assign n14239 = n14238 ^ n11678;
  assign n14240 = n14239 ^ x605;
  assign n14241 = n13308 & n13444;
  assign n14242 = n13398 & n13628;
  assign n14243 = ~n14241 & ~n14242;
  assign n14244 = n13307 & n13406;
  assign n14245 = n13402 & ~n13644;
  assign n14246 = ~n14244 & ~n14245;
  assign n14247 = n13308 & n13403;
  assign n14248 = ~n13396 & n13427;
  assign n14249 = ~n14247 & ~n14248;
  assign n14250 = ~n13394 & n13634;
  assign n14251 = ~n13436 & n14250;
  assign n14252 = n13398 & ~n14251;
  assign n14253 = ~n13389 & n13442;
  assign n14254 = ~n13403 & n13634;
  assign n14255 = ~n13400 & n14254;
  assign n14256 = n13395 & ~n14255;
  assign n14257 = ~n13402 & ~n14256;
  assign n14258 = ~n14253 & ~n14257;
  assign n14259 = ~n14252 & ~n14258;
  assign n14260 = n14249 & n14259;
  assign n14261 = n14246 & n14260;
  assign n14262 = n14243 & n14261;
  assign n14263 = ~n13633 & n14262;
  assign n14264 = n13418 & n14263;
  assign n14265 = n13631 & n14264;
  assign n14266 = ~n13391 & n14265;
  assign n14267 = n14266 ^ n11733;
  assign n14268 = n14267 ^ x607;
  assign n14269 = n14240 & ~n14268;
  assign n14270 = n14218 & n14269;
  assign n14271 = n14185 & n14270;
  assign n14272 = ~n14149 & n14184;
  assign n14273 = n14240 & n14268;
  assign n14274 = n14218 & n14273;
  assign n14275 = n14195 & ~n14217;
  assign n14276 = n14269 & n14275;
  assign n14277 = ~n14274 & ~n14276;
  assign n14278 = n14272 & ~n14277;
  assign n14279 = n14149 & ~n14184;
  assign n14280 = n14217 ^ n14195;
  assign n14281 = n14280 ^ n14268;
  assign n14282 = n14268 ^ n14240;
  assign n14283 = n14281 & ~n14282;
  assign n14284 = n14279 & n14283;
  assign n14285 = ~n14278 & ~n14284;
  assign n14286 = ~n14240 & ~n14268;
  assign n14287 = ~n14195 & ~n14217;
  assign n14288 = n14286 & n14287;
  assign n14289 = n14272 & n14288;
  assign n14290 = ~n14149 & ~n14184;
  assign n14291 = ~n14240 & n14268;
  assign n14292 = n14218 & n14291;
  assign n14293 = n14275 & n14291;
  assign n14294 = ~n14292 & ~n14293;
  assign n14295 = n14290 & ~n14294;
  assign n14296 = ~n14289 & ~n14295;
  assign n14297 = ~n14195 & n14217;
  assign n14298 = n14269 & n14297;
  assign n14299 = n14272 & n14298;
  assign n14300 = n14269 & n14287;
  assign n14301 = n14290 & n14300;
  assign n14302 = ~n14299 & ~n14301;
  assign n14303 = n14149 & n14288;
  assign n14304 = n14185 & n14292;
  assign n14305 = n14218 & n14286;
  assign n14306 = ~n14293 & ~n14305;
  assign n14307 = ~n14300 & n14306;
  assign n14308 = n14272 & ~n14307;
  assign n14309 = ~n14304 & ~n14308;
  assign n14310 = n14184 ^ n14149;
  assign n14311 = n14291 & n14297;
  assign n14312 = n14310 & n14311;
  assign n14313 = n14273 & n14275;
  assign n14314 = ~n14270 & ~n14313;
  assign n14315 = n14279 & ~n14314;
  assign n14316 = n14287 & n14291;
  assign n14317 = ~n14305 & ~n14316;
  assign n14318 = n14273 & n14297;
  assign n14319 = ~n14276 & ~n14318;
  assign n14320 = ~n14298 & n14319;
  assign n14321 = n14317 & n14320;
  assign n14322 = ~n14310 & ~n14321;
  assign n14323 = ~n14315 & ~n14322;
  assign n14324 = ~n14312 & n14323;
  assign n14325 = n14309 & n14324;
  assign n14326 = ~n14303 & n14325;
  assign n14327 = n14302 & n14326;
  assign n14328 = n14296 & n14327;
  assign n14329 = n14285 & n14328;
  assign n14330 = ~n14271 & n14329;
  assign n14331 = n14330 ^ n12727;
  assign n14332 = n14331 ^ x648;
  assign n14333 = ~n14113 & ~n14332;
  assign n14334 = n13854 & n14333;
  assign n14335 = n13093 & n13097;
  assign n14336 = n13100 & ~n14335;
  assign n14337 = ~n13113 & ~n13136;
  assign n14338 = n13092 & ~n14337;
  assign n14339 = ~n13125 & n13139;
  assign n14340 = n13110 & ~n14339;
  assign n14341 = ~n14338 & ~n14340;
  assign n14342 = n13115 & ~n13580;
  assign n14343 = n13109 & ~n13143;
  assign n14344 = n13093 & ~n14343;
  assign n14345 = ~n13107 & ~n13120;
  assign n14346 = ~n13567 & ~n14345;
  assign n14347 = ~n14344 & ~n14346;
  assign n14348 = ~n14342 & n14347;
  assign n14349 = n14341 & n14348;
  assign n14350 = ~n13135 & n14349;
  assign n14351 = n13130 & n14350;
  assign n14352 = ~n13127 & n14351;
  assign n14353 = n13564 & n14352;
  assign n14354 = n14336 & n14353;
  assign n14355 = n13561 & n14354;
  assign n14356 = n14355 ^ n11176;
  assign n14357 = n14356 ^ x597;
  assign n14358 = n14024 ^ x592;
  assign n14359 = ~n14357 & ~n14358;
  assign n14360 = n12862 & n12878;
  assign n14361 = ~n12891 & ~n12900;
  assign n14362 = ~n12878 & n14361;
  assign n14363 = n12871 & ~n14362;
  assign n14364 = ~n14360 & ~n14363;
  assign n14365 = n12883 & ~n12899;
  assign n14366 = n12866 ^ n12792;
  assign n14367 = n12728 & n14366;
  assign n14368 = n12690 & n14367;
  assign n14369 = n14368 ^ n12792;
  assign n14370 = n12876 & n14369;
  assign n14371 = ~n12790 & n13604;
  assign n14372 = n12885 & ~n14371;
  assign n14373 = ~n12875 & ~n14137;
  assign n14374 = n12863 & ~n14373;
  assign n14375 = ~n14372 & ~n14374;
  assign n14376 = ~n14370 & n14375;
  assign n14377 = ~n14365 & n14376;
  assign n14378 = n14364 & n14377;
  assign n14379 = n14123 & n14378;
  assign n14380 = n14120 & n14379;
  assign n14381 = n14116 & n14380;
  assign n14382 = n12896 & n14381;
  assign n14383 = n14382 ^ n11309;
  assign n14384 = n14383 ^ x594;
  assign n14385 = n13308 & n13427;
  assign n14386 = ~n13396 & n13413;
  assign n14387 = ~n14385 & ~n14386;
  assign n14388 = n13395 & n13436;
  assign n14389 = n13390 & ~n13628;
  assign n14390 = ~n13400 & n14389;
  assign n14391 = ~n13419 & n14390;
  assign n14392 = n13402 & ~n14391;
  assign n14393 = n13307 & n13411;
  assign n14394 = n13386 & ~n13396;
  assign n14395 = ~n14393 & ~n14394;
  assign n14396 = ~n13396 & ~n13442;
  assign n14397 = ~n13440 & ~n13444;
  assign n14398 = ~n13403 & n14397;
  assign n14399 = ~n13308 & n14398;
  assign n14400 = n14396 & ~n14399;
  assign n14401 = n13423 & ~n13439;
  assign n14402 = ~n13419 & n14401;
  assign n14403 = n13398 & ~n14402;
  assign n14404 = ~n14400 & ~n14403;
  assign n14405 = n14395 & n14404;
  assign n14406 = ~n14392 & n14405;
  assign n14407 = ~n14388 & n14406;
  assign n14408 = n14387 & n14407;
  assign n14409 = n14243 & n14408;
  assign n14410 = n13425 & n14409;
  assign n14411 = n13409 & n14410;
  assign n14412 = n14411 ^ n11269;
  assign n14413 = n14412 ^ x596;
  assign n14414 = ~n14384 & n14413;
  assign n14415 = n13887 ^ x593;
  assign n14416 = n12590 & n12617;
  assign n14417 = n12318 & n12631;
  assign n14418 = n12592 & n12598;
  assign n14419 = ~n14417 & ~n14418;
  assign n14420 = ~n14416 & n14419;
  assign n14421 = n12621 & n12637;
  assign n14422 = ~n12622 & ~n12632;
  assign n14423 = ~n12612 & n14422;
  assign n14424 = n12592 & ~n14423;
  assign n14425 = ~n12631 & ~n12632;
  assign n14426 = n12590 & ~n14425;
  assign n14427 = ~n12594 & n12634;
  assign n14428 = ~n12602 & n14427;
  assign n14429 = n12609 & ~n14428;
  assign n14430 = ~n12611 & n14170;
  assign n14431 = ~n12625 & n14430;
  assign n14432 = n12318 & ~n14431;
  assign n14433 = ~n14429 & ~n14432;
  assign n14434 = ~n14426 & n14433;
  assign n14435 = ~n14424 & n14434;
  assign n14436 = ~n14421 & n14435;
  assign n14437 = ~n14161 & n14436;
  assign n14438 = n14420 & n14437;
  assign n14439 = n14156 & n14438;
  assign n14440 = ~n14151 & n14439;
  assign n14441 = n12620 & n14440;
  assign n14442 = n12607 & n14441;
  assign n14443 = ~n12589 & n14442;
  assign n14444 = n14443 ^ n11237;
  assign n14445 = n14444 ^ x595;
  assign n14446 = ~n14415 & n14445;
  assign n14447 = n14414 & n14446;
  assign n14448 = n14359 & n14447;
  assign n14449 = ~n14357 & n14358;
  assign n14450 = ~n14415 & ~n14445;
  assign n14451 = n14414 & n14450;
  assign n14452 = n14449 & n14451;
  assign n14453 = ~n14448 & ~n14452;
  assign n14454 = n14357 & ~n14358;
  assign n14455 = n14384 & n14413;
  assign n14456 = n14415 & ~n14445;
  assign n14457 = n14455 & n14456;
  assign n14458 = n14454 & n14457;
  assign n14459 = n14357 & n14358;
  assign n14460 = ~n14413 & n14456;
  assign n14461 = ~n14384 & n14460;
  assign n14462 = n14459 & n14461;
  assign n14463 = ~n14458 & ~n14462;
  assign n14464 = n14453 & n14463;
  assign n14465 = n14457 & n14459;
  assign n14466 = ~n14413 & n14450;
  assign n14467 = ~n14384 & n14466;
  assign n14468 = n14454 & n14467;
  assign n14469 = ~n14465 & ~n14468;
  assign n14470 = n14415 & n14445;
  assign n14471 = ~n14413 & n14470;
  assign n14472 = n14384 & n14471;
  assign n14473 = n14450 & n14455;
  assign n14474 = n14454 & n14473;
  assign n14475 = ~n14384 & n14471;
  assign n14476 = n14459 & n14475;
  assign n14477 = n14359 & n14461;
  assign n14478 = ~n14476 & ~n14477;
  assign n14479 = ~n14474 & n14478;
  assign n14480 = ~n14359 & ~n14459;
  assign n14481 = n14384 & n14466;
  assign n14482 = ~n14480 & n14481;
  assign n14483 = n14446 & n14455;
  assign n14484 = ~n14413 & n14446;
  assign n14485 = n14384 & n14484;
  assign n14486 = ~n14483 & ~n14485;
  assign n14487 = ~n14447 & n14486;
  assign n14488 = n14459 & ~n14487;
  assign n14489 = ~n14482 & ~n14488;
  assign n14490 = n14414 & n14470;
  assign n14491 = n14449 & n14490;
  assign n14492 = n14414 & n14456;
  assign n14493 = ~n14384 & n14484;
  assign n14494 = ~n14447 & ~n14493;
  assign n14495 = ~n14492 & n14494;
  assign n14496 = ~n14483 & n14495;
  assign n14497 = n14454 & ~n14496;
  assign n14498 = ~n14473 & ~n14485;
  assign n14499 = n14455 & n14470;
  assign n14500 = n14384 & n14460;
  assign n14501 = ~n14499 & ~n14500;
  assign n14502 = n14498 & n14501;
  assign n14503 = ~n14467 & n14502;
  assign n14504 = n14449 & ~n14503;
  assign n14505 = ~n14475 & n14501;
  assign n14506 = ~n14451 & n14505;
  assign n14507 = n14359 & ~n14506;
  assign n14508 = ~n14504 & ~n14507;
  assign n14509 = ~n14497 & n14508;
  assign n14510 = ~n14491 & n14509;
  assign n14511 = n14489 & n14510;
  assign n14512 = n14479 & n14511;
  assign n14513 = ~n14472 & n14512;
  assign n14514 = n14469 & n14513;
  assign n14515 = n14464 & n14514;
  assign n14516 = n14515 ^ n12825;
  assign n14517 = n14516 ^ x651;
  assign n14518 = n13663 ^ x622;
  assign n14519 = n12653 ^ x627;
  assign n14520 = n14518 & n14519;
  assign n14521 = n13275 ^ x626;
  assign n14522 = n13667 & n13759;
  assign n14523 = n13718 & ~n13762;
  assign n14524 = ~n14522 & ~n14523;
  assign n14525 = ~n13748 & ~n13760;
  assign n14526 = ~n13744 & n14525;
  assign n14527 = ~n13765 & n14526;
  assign n14528 = n13722 & ~n14527;
  assign n14529 = ~n13720 & n13911;
  assign n14530 = n13728 & ~n14529;
  assign n14531 = n13722 & ~n14220;
  assign n14532 = ~n13737 & ~n14531;
  assign n14533 = n13903 & n14532;
  assign n14534 = n13665 & ~n14533;
  assign n14535 = ~n14530 & ~n14534;
  assign n14536 = ~n14528 & n14535;
  assign n14537 = n14524 & n14536;
  assign n14538 = n13901 & n14537;
  assign n14539 = ~n13897 & n14538;
  assign n14540 = n14222 & n14539;
  assign n14541 = ~n13717 & n14540;
  assign n14542 = n14541 ^ n12482;
  assign n14543 = n14542 ^ x625;
  assign n14544 = n14521 & ~n14543;
  assign n14545 = n13592 ^ x623;
  assign n14546 = ~n13974 & ~n14196;
  assign n14547 = n13928 & ~n14546;
  assign n14548 = n13969 & n13991;
  assign n14549 = n14008 & ~n14548;
  assign n14550 = n14002 & ~n14549;
  assign n14551 = ~n14547 & ~n14550;
  assign n14552 = n13966 & n13973;
  assign n14553 = n13968 & n13994;
  assign n14554 = ~n13987 & ~n14553;
  assign n14555 = ~n13980 & n14554;
  assign n14556 = ~n13976 & n14555;
  assign n14557 = n13986 & ~n14556;
  assign n14558 = ~n13926 & n14196;
  assign n14559 = ~n13928 & ~n14005;
  assign n14560 = ~n13992 & n14559;
  assign n14561 = ~n13986 & ~n14548;
  assign n14562 = ~n14560 & ~n14561;
  assign n14563 = ~n13983 & ~n14562;
  assign n14564 = ~n13995 & n14563;
  assign n14565 = n13926 & ~n14564;
  assign n14566 = ~n13973 & n14555;
  assign n14567 = ~n14006 & ~n14548;
  assign n14568 = ~n14002 & n14567;
  assign n14569 = ~n13926 & ~n14568;
  assign n14570 = ~n13995 & ~n14569;
  assign n14571 = ~n14566 & ~n14570;
  assign n14572 = ~n14565 & ~n14571;
  assign n14573 = ~n14558 & n14572;
  assign n14574 = ~n14557 & n14573;
  assign n14575 = ~n14552 & n14574;
  assign n14576 = n14551 & n14575;
  assign n14577 = n13979 & n14576;
  assign n14578 = ~n13964 & n14577;
  assign n14579 = n14578 ^ n12458;
  assign n14580 = n14579 ^ x624;
  assign n14581 = n14545 & n14580;
  assign n14582 = n14544 & n14581;
  assign n14583 = n14520 & n14582;
  assign n14584 = n14518 & ~n14519;
  assign n14585 = ~n14521 & ~n14543;
  assign n14586 = n14581 & n14585;
  assign n14587 = n14545 & ~n14580;
  assign n14588 = n14544 & n14587;
  assign n14589 = ~n14586 & ~n14588;
  assign n14590 = n14584 & ~n14589;
  assign n14591 = ~n14583 & ~n14590;
  assign n14592 = ~n14518 & ~n14519;
  assign n14593 = ~n14521 & n14543;
  assign n14594 = n14581 & n14593;
  assign n14595 = ~n14582 & ~n14594;
  assign n14596 = n14592 & ~n14595;
  assign n14597 = n14521 & n14543;
  assign n14598 = n14581 & n14597;
  assign n14599 = n14587 & n14593;
  assign n14600 = ~n14598 & ~n14599;
  assign n14601 = n14584 & ~n14600;
  assign n14602 = ~n14596 & ~n14601;
  assign n14603 = n14520 & n14586;
  assign n14604 = ~n14518 & n14519;
  assign n14605 = ~n14545 & ~n14580;
  assign n14606 = n14597 & n14605;
  assign n14607 = n14593 & n14605;
  assign n14608 = ~n14545 & n14580;
  assign n14609 = n14597 & n14608;
  assign n14610 = n14585 & n14608;
  assign n14611 = ~n14609 & ~n14610;
  assign n14612 = ~n14607 & n14611;
  assign n14613 = ~n14606 & n14612;
  assign n14614 = n14604 & ~n14613;
  assign n14615 = ~n14603 & ~n14614;
  assign n14616 = ~n14520 & ~n14592;
  assign n14617 = n14587 & n14597;
  assign n14618 = ~n14599 & ~n14617;
  assign n14619 = ~n14616 & ~n14618;
  assign n14620 = n14584 & ~n14611;
  assign n14622 = n14585 & n14587;
  assign n14636 = n14584 & n14606;
  assign n14637 = n14589 & ~n14594;
  assign n14638 = n14604 & ~n14637;
  assign n14639 = ~n14636 & ~n14638;
  assign n14640 = ~n14622 & n14639;
  assign n14621 = n14544 & n14605;
  assign n14623 = n14593 & n14608;
  assign n14624 = n14544 & n14608;
  assign n14625 = ~n14623 & ~n14624;
  assign n14626 = ~n14622 & n14625;
  assign n14627 = ~n14520 & n14626;
  assign n14628 = n14585 & n14605;
  assign n14629 = ~n14622 & ~n14623;
  assign n14630 = n14592 & ~n14629;
  assign n14631 = ~n14628 & ~n14630;
  assign n14632 = ~n14624 & n14631;
  assign n14633 = ~n14607 & n14632;
  assign n14634 = ~n14627 & ~n14633;
  assign n14635 = ~n14621 & ~n14634;
  assign n14641 = n14640 ^ n14635;
  assign n14642 = ~n14616 & n14641;
  assign n14643 = n14642 ^ n14640;
  assign n14644 = ~n14620 & n14643;
  assign n14645 = ~n14619 & n14644;
  assign n14646 = n14615 & n14645;
  assign n14647 = n14602 & n14646;
  assign n14648 = n14591 & n14647;
  assign n14649 = n14648 ^ n12861;
  assign n14650 = n14649 ^ x646;
  assign n14651 = n14517 & n14650;
  assign n14652 = n14334 & n14651;
  assign n14653 = ~n14113 & n14332;
  assign n14654 = ~n13520 & n13853;
  assign n14655 = n14653 & n14654;
  assign n14656 = ~n14517 & n14650;
  assign n14657 = n14655 & n14656;
  assign n14658 = ~n14652 & ~n14657;
  assign n14659 = n14113 & n14332;
  assign n14660 = n13854 & n14659;
  assign n14661 = n14517 & ~n14650;
  assign n14662 = n14660 & n14661;
  assign n14663 = n14333 & n14654;
  assign n14664 = ~n14517 & ~n14650;
  assign n14665 = n14663 & n14664;
  assign n14666 = ~n14662 & ~n14665;
  assign n14667 = n14658 & n14666;
  assign n14668 = ~n13520 & ~n13853;
  assign n14669 = n14333 & n14668;
  assign n14670 = n14661 & n14669;
  assign n14671 = n14659 & n14668;
  assign n14672 = n14651 & n14671;
  assign n14673 = n14655 & n14661;
  assign n14674 = ~n14672 & ~n14673;
  assign n14675 = ~n14670 & n14674;
  assign n14676 = n13854 & n14653;
  assign n14677 = ~n14669 & ~n14676;
  assign n14678 = n14656 & ~n14677;
  assign n14679 = n14113 & ~n14332;
  assign n14680 = n14654 & n14679;
  assign n14681 = n14651 & n14680;
  assign n14682 = n13520 & ~n13853;
  assign n14683 = n14679 & n14682;
  assign n14684 = ~n14671 & ~n14680;
  assign n14685 = ~n14683 & n14684;
  assign n14686 = n14661 & ~n14685;
  assign n14687 = ~n14681 & ~n14686;
  assign n14688 = n14659 & n14682;
  assign n14689 = ~n14680 & ~n14688;
  assign n14690 = n14664 & ~n14689;
  assign n14691 = n14333 & n14682;
  assign n14692 = n14668 & n14679;
  assign n14693 = ~n14691 & ~n14692;
  assign n14694 = n14654 & n14659;
  assign n14695 = n13854 & n14679;
  assign n14696 = ~n14688 & ~n14695;
  assign n14697 = ~n14694 & n14696;
  assign n14698 = n14693 & n14697;
  assign n14699 = n14656 & ~n14698;
  assign n14700 = ~n14683 & ~n14694;
  assign n14701 = n14653 & n14682;
  assign n14702 = n14653 & n14668;
  assign n14703 = ~n14676 & ~n14702;
  assign n14704 = ~n14701 & n14703;
  assign n14705 = n14700 & n14704;
  assign n14706 = n14650 ^ n14517;
  assign n14707 = ~n14705 & ~n14706;
  assign n14708 = ~n14334 & ~n14691;
  assign n14709 = n14661 & ~n14708;
  assign n14710 = ~n14707 & ~n14709;
  assign n14711 = ~n14699 & n14710;
  assign n14712 = ~n14690 & n14711;
  assign n14713 = n14687 & n14712;
  assign n14714 = ~n14678 & n14713;
  assign n14715 = n14675 & n14714;
  assign n14716 = n14667 & n14715;
  assign n14717 = n14716 ^ n14148;
  assign n14718 = n14717 ^ x705;
  assign n14719 = n14239 ^ x603;
  assign n14720 = n14412 ^ x598;
  assign n14721 = n14719 & ~n14720;
  assign n14722 = n14356 ^ x599;
  assign n14723 = n13926 & ~n14198;
  assign n14724 = n13973 & ~n14004;
  assign n14725 = ~n14723 & ~n14724;
  assign n14726 = n13986 & n14553;
  assign n14727 = n13997 & ~n14005;
  assign n14728 = n14002 & ~n14727;
  assign n14729 = n13997 & n14559;
  assign n14730 = ~n14548 & n14729;
  assign n14731 = ~n13992 & n14567;
  assign n14732 = ~n13986 & n14731;
  assign n14733 = ~n14730 & ~n14732;
  assign n14734 = n13926 & n14733;
  assign n14735 = n13971 & ~n14553;
  assign n14736 = ~n13976 & n14735;
  assign n14737 = n14002 & ~n14736;
  assign n14738 = ~n13963 & n14731;
  assign n14739 = n13973 & ~n14738;
  assign n14740 = ~n14737 & ~n14739;
  assign n14741 = ~n14734 & n14740;
  assign n14742 = ~n13964 & n14741;
  assign n14743 = ~n14728 & n14742;
  assign n14744 = ~n14726 & n14743;
  assign n14745 = n14725 & n14744;
  assign n14746 = ~n14197 & n14745;
  assign n14747 = n13985 & n14746;
  assign n14748 = n14747 ^ n12122;
  assign n14749 = n14748 ^ x601;
  assign n14750 = ~n14722 & n14749;
  assign n14751 = ~n13207 & ~n13237;
  assign n14752 = n13167 & ~n14751;
  assign n14753 = ~n13211 & n13238;
  assign n14754 = ~n13222 & n14753;
  assign n14755 = n13209 & ~n14754;
  assign n14756 = ~n14752 & ~n14755;
  assign n14757 = ~n13249 & n13258;
  assign n14758 = ~n13228 & ~n13261;
  assign n14759 = n13230 & ~n14758;
  assign n14760 = ~n13247 & n14030;
  assign n14761 = n13235 & ~n14760;
  assign n14762 = ~n14759 & ~n14761;
  assign n14763 = ~n14757 & n14762;
  assign n14764 = n14756 & n14763;
  assign n14765 = ~n13522 & n14764;
  assign n14766 = n13234 & n14765;
  assign n14767 = ~n13219 & n14766;
  assign n14768 = n14028 & n14767;
  assign n14769 = ~n13530 & n14768;
  assign n14770 = n14769 ^ n12152;
  assign n14771 = n14770 ^ x600;
  assign n14772 = n14183 ^ x602;
  assign n14773 = n14771 & ~n14772;
  assign n14774 = n14750 & n14773;
  assign n14775 = n14721 & n14774;
  assign n14776 = n14719 & n14720;
  assign n14777 = n14722 & ~n14749;
  assign n14778 = n14773 & n14777;
  assign n14779 = n14776 & n14778;
  assign n14780 = ~n14719 & n14720;
  assign n14781 = ~n14771 & n14772;
  assign n14782 = n14777 & n14781;
  assign n14783 = n14780 & n14782;
  assign n14784 = ~n14779 & ~n14783;
  assign n14785 = ~n14775 & n14784;
  assign n14786 = n14776 & n14782;
  assign n14787 = n14722 & n14749;
  assign n14788 = n14781 & n14787;
  assign n14789 = n14773 & n14787;
  assign n14790 = ~n14788 & ~n14789;
  assign n14791 = n14720 & ~n14790;
  assign n14792 = ~n14786 & ~n14791;
  assign n14793 = ~n14771 & ~n14772;
  assign n14794 = n14787 & n14793;
  assign n14795 = n14780 & n14794;
  assign n14796 = ~n14719 & ~n14720;
  assign n14797 = n14771 & n14772;
  assign n14798 = n14787 & n14797;
  assign n14799 = n14777 & n14797;
  assign n14800 = ~n14794 & ~n14799;
  assign n14801 = ~n14778 & n14800;
  assign n14802 = ~n14798 & n14801;
  assign n14803 = n14796 & ~n14802;
  assign n14804 = ~n14795 & ~n14803;
  assign n14805 = ~n14722 & ~n14749;
  assign n14806 = n14797 & n14805;
  assign n14807 = n14750 & n14797;
  assign n14808 = n14750 & n14793;
  assign n14809 = ~n14807 & ~n14808;
  assign n14810 = ~n14806 & n14809;
  assign n14811 = n14721 & ~n14810;
  assign n14812 = n14721 & n14782;
  assign n14813 = n14750 & n14781;
  assign n14814 = n14773 & n14805;
  assign n14815 = ~n14813 & ~n14814;
  assign n14816 = n14796 & ~n14815;
  assign n14817 = n14781 & n14805;
  assign n14818 = ~n14774 & ~n14817;
  assign n14819 = n14776 & ~n14818;
  assign n14820 = ~n14816 & ~n14819;
  assign n14821 = n14720 ^ n14719;
  assign n14822 = ~n14809 & ~n14821;
  assign n14823 = n14780 & n14805;
  assign n14824 = n14777 & n14793;
  assign n14825 = ~n14778 & ~n14824;
  assign n14826 = ~n14788 & n14825;
  assign n14827 = n14721 & ~n14826;
  assign n14828 = ~n14823 & ~n14827;
  assign n14829 = ~n14822 & n14828;
  assign n14830 = n14820 & n14829;
  assign n14831 = ~n14812 & n14830;
  assign n14832 = ~n14811 & n14831;
  assign n14833 = n14804 & n14832;
  assign n14834 = n14792 & n14833;
  assign n14835 = n14785 & n14834;
  assign n14836 = n14835 ^ n12584;
  assign n14837 = n14836 ^ x666;
  assign n14838 = n14588 & n14604;
  assign n14839 = n14584 & n14628;
  assign n14840 = ~n14838 & ~n14839;
  assign n14841 = ~n14610 & ~n14621;
  assign n14842 = ~n14616 & ~n14841;
  assign n14843 = n14840 & ~n14842;
  assign n14844 = n14595 & ~n14623;
  assign n14845 = n14604 & ~n14844;
  assign n14846 = n14604 & ~n14841;
  assign n14847 = n14584 & n14607;
  assign n14848 = n14600 & ~n14606;
  assign n14849 = n14592 & ~n14848;
  assign n14850 = ~n14847 & ~n14849;
  assign n14851 = ~n14846 & n14850;
  assign n14852 = n14599 & n14604;
  assign n14853 = ~n14636 & ~n14852;
  assign n14854 = n14609 & n14616;
  assign n14855 = ~n14617 & ~n14622;
  assign n14856 = n14600 & n14855;
  assign n14857 = n14520 & ~n14856;
  assign n14858 = ~n14854 & ~n14857;
  assign n14859 = ~n14588 & n14595;
  assign n14860 = n14592 & ~n14859;
  assign n14861 = n14520 & ~n14625;
  assign n14862 = ~n14586 & n14595;
  assign n14863 = ~n14622 & n14862;
  assign n14864 = n14584 & ~n14863;
  assign n14865 = ~n14861 & ~n14864;
  assign n14866 = ~n14860 & n14865;
  assign n14867 = n14858 & n14866;
  assign n14868 = n14853 & n14867;
  assign n14869 = n14851 & n14868;
  assign n14870 = ~n14845 & n14869;
  assign n14871 = n14843 & n14870;
  assign n14872 = n14871 ^ n12552;
  assign n14873 = n14872 ^ x667;
  assign n14874 = ~n14837 & ~n14873;
  assign n14875 = n14216 ^ x610;
  assign n14876 = n13780 ^ x615;
  assign n14877 = ~n14875 & ~n14876;
  assign n14878 = n13555 ^ x614;
  assign n14907 = n14148 ^ x611;
  assign n14879 = n12592 & n12626;
  assign n14880 = n12621 & ~n12624;
  assign n14881 = ~n14879 & ~n14880;
  assign n14882 = ~n12276 & n12625;
  assign n14883 = n12609 & n12637;
  assign n14884 = ~n14882 & ~n14883;
  assign n14885 = ~n12598 & ~n12602;
  assign n14886 = n12318 & ~n14885;
  assign n14887 = ~n12617 & n12627;
  assign n14888 = ~n12637 & n14887;
  assign n14889 = n12318 & ~n14888;
  assign n14890 = n12604 & n14425;
  assign n14891 = n12592 & ~n14890;
  assign n14892 = ~n12603 & n14427;
  assign n14893 = n12590 & ~n14892;
  assign n14894 = ~n12588 & n12642;
  assign n14895 = n12609 & ~n14894;
  assign n14896 = ~n14893 & ~n14895;
  assign n14897 = ~n14891 & n14896;
  assign n14898 = ~n14889 & n14897;
  assign n14899 = ~n14886 & n14898;
  assign n14900 = n14884 & n14899;
  assign n14901 = n14881 & n14900;
  assign n14902 = n14420 & n14901;
  assign n14903 = n14163 & n14902;
  assign n14904 = ~n12589 & n14903;
  assign n14905 = n14904 ^ n12373;
  assign n14906 = n14905 ^ x612;
  assign n14908 = n14907 ^ n14906;
  assign n14909 = ~n14878 & n14908;
  assign n14910 = n13093 & ~n13122;
  assign n14911 = n13133 & n14337;
  assign n14912 = ~n13102 & n14911;
  assign n14913 = ~n13104 & n14912;
  assign n14914 = n13098 & ~n14913;
  assign n14915 = ~n14910 & ~n14914;
  assign n14916 = n13131 & ~n13567;
  assign n14917 = ~n13112 & n13148;
  assign n14918 = ~n13107 & n14917;
  assign n14919 = ~n13132 & n14918;
  assign n14920 = n13115 & ~n14919;
  assign n14921 = ~n13104 & n13139;
  assign n14922 = ~n13118 & n14921;
  assign n14923 = ~n13093 & n14922;
  assign n14924 = ~n13107 & n13144;
  assign n14925 = ~n13125 & n14924;
  assign n14926 = n13093 & ~n14925;
  assign n14927 = ~n13110 & ~n14926;
  assign n14928 = ~n14923 & ~n14927;
  assign n14929 = ~n14920 & ~n14928;
  assign n14930 = ~n14916 & n14929;
  assign n14931 = n14915 & n14930;
  assign n14932 = n13560 & n14931;
  assign n14933 = n14336 & n14932;
  assign n14934 = n13124 & n14933;
  assign n14935 = n14934 ^ n12350;
  assign n14936 = n14935 ^ x613;
  assign n14937 = n14878 & n14936;
  assign n14938 = ~n14907 & n14937;
  assign n14939 = n14906 ^ n14878;
  assign n14940 = n14907 & ~n14936;
  assign n14941 = n14939 & n14940;
  assign n14942 = ~n14938 & ~n14941;
  assign n14943 = ~n14909 & n14942;
  assign n14944 = n14877 & ~n14943;
  assign n14945 = n14875 & n14876;
  assign n14946 = n14906 & ~n14907;
  assign n14947 = ~n14936 & n14946;
  assign n14948 = n14936 & n14939;
  assign n14949 = n14907 & n14948;
  assign n14950 = ~n14907 & ~n14939;
  assign n14951 = ~n14878 & ~n14906;
  assign n14952 = ~n14936 & n14951;
  assign n14953 = ~n14950 & ~n14952;
  assign n14954 = ~n14949 & n14953;
  assign n14955 = ~n14947 & n14954;
  assign n14956 = n14945 & ~n14955;
  assign n14957 = ~n14944 & ~n14956;
  assign n14958 = n14875 & ~n14876;
  assign n14959 = n14936 ^ n14906;
  assign n14960 = n14951 & ~n14959;
  assign n14961 = n14960 ^ n14959;
  assign n14962 = ~n14907 & ~n14961;
  assign n14963 = n14907 & n14937;
  assign n14964 = ~n14940 & ~n14946;
  assign n14965 = ~n14878 & ~n14964;
  assign n14966 = ~n14963 & ~n14965;
  assign n14967 = ~n14962 & n14966;
  assign n14968 = n14958 & n14967;
  assign n14969 = ~n14875 & n14876;
  assign n14970 = n14936 & ~n14939;
  assign n14971 = n14906 & n14940;
  assign n14972 = ~n14970 & ~n14971;
  assign n14973 = ~n14962 & n14972;
  assign n14974 = n14969 & ~n14973;
  assign n14975 = ~n14968 & ~n14974;
  assign n14976 = n14957 & n14975;
  assign n14977 = n14976 ^ n12421;
  assign n14978 = n14977 ^ x668;
  assign n14979 = n14359 & n14457;
  assign n14980 = n14359 & n14472;
  assign n14981 = n14459 & n14500;
  assign n14982 = ~n14980 & ~n14981;
  assign n14983 = n14494 & n14498;
  assign n14984 = ~n14359 & n14983;
  assign n14985 = ~n14481 & n14486;
  assign n14986 = ~n14459 & n14985;
  assign n14987 = ~n14984 & ~n14986;
  assign n14988 = ~n14480 & n14987;
  assign n14989 = n14487 & n14505;
  assign n14990 = ~n14457 & n14989;
  assign n14991 = n14449 & ~n14990;
  assign n14992 = ~n14988 & ~n14991;
  assign n14993 = ~n14480 & n14492;
  assign n14994 = ~n14461 & ~n14483;
  assign n14995 = ~n14490 & ~n14500;
  assign n14996 = ~n14472 & n14995;
  assign n14997 = n14994 & n14996;
  assign n14998 = ~n14499 & n14997;
  assign n14999 = n14454 & ~n14998;
  assign n15000 = ~n14993 & ~n14999;
  assign n15001 = n14992 & n15000;
  assign n15002 = n14982 & n15001;
  assign n15003 = ~n14979 & n15002;
  assign n15004 = n14479 & n15003;
  assign n15005 = n14453 & n15004;
  assign n15006 = n14469 & n15005;
  assign n15007 = n15006 ^ n11390;
  assign n15008 = n15007 ^ x665;
  assign n15009 = ~n14978 & ~n15008;
  assign n15010 = n14874 & n15009;
  assign n15011 = ~n14096 & ~n14098;
  assign n15012 = n14063 & ~n15011;
  assign n15013 = ~n14062 & ~n15012;
  assign n15014 = ~n14070 & ~n14088;
  assign n15015 = ~n14079 & ~n15014;
  assign n15016 = ~n14072 & ~n14075;
  assign n15017 = n14052 & ~n15016;
  assign n15018 = ~n15015 & ~n15017;
  assign n15019 = n14061 & ~n14082;
  assign n15020 = ~n14098 & ~n14099;
  assign n15021 = ~n14074 & ~n14088;
  assign n15022 = n15020 & n15021;
  assign n15023 = n13890 & ~n15022;
  assign n15024 = n13890 & n14054;
  assign n15025 = n13890 & n14057;
  assign n15026 = n14061 & n14070;
  assign n15027 = ~n15025 & ~n15026;
  assign n15028 = n14050 & ~n14095;
  assign n15029 = n14063 & n14099;
  assign n15030 = ~n15028 & ~n15029;
  assign n15031 = n13889 ^ n13888;
  assign n15032 = n14086 & n15031;
  assign n15033 = n14052 & ~n14087;
  assign n15034 = ~n15032 & ~n15033;
  assign n15035 = n15030 & n15034;
  assign n15036 = ~n14066 & ~n14079;
  assign n15037 = n14061 & ~n14076;
  assign n15038 = ~n15036 & ~n15037;
  assign n15039 = n15035 & n15038;
  assign n15040 = n15027 & n15039;
  assign n15041 = ~n15024 & n15040;
  assign n15042 = ~n15023 & n15041;
  assign n15043 = ~n15019 & n15042;
  assign n15044 = n15018 & n15043;
  assign n15045 = n15013 & n15044;
  assign n15046 = n15045 ^ n12316;
  assign n15047 = n15046 ^ x669;
  assign n15048 = n14272 & n14316;
  assign n15049 = n14273 & n14287;
  assign n15050 = ~n14298 & ~n15049;
  assign n15051 = ~n14270 & n15050;
  assign n15052 = n14290 & ~n15051;
  assign n15053 = n14290 & n14318;
  assign n15054 = n14275 & n14286;
  assign n15055 = ~n14310 & n15054;
  assign n15056 = ~n15053 & ~n15055;
  assign n15057 = n14286 & n14297;
  assign n15058 = ~n14305 & ~n15057;
  assign n15059 = ~n14293 & n15058;
  assign n15060 = n14279 & ~n15059;
  assign n15061 = n14290 & n14311;
  assign n15062 = n14272 & ~n15058;
  assign n15063 = ~n15061 & ~n15062;
  assign n15064 = ~n14313 & ~n14318;
  assign n15065 = n14310 & ~n15064;
  assign n15066 = ~n14276 & ~n15049;
  assign n15067 = ~n14288 & n15066;
  assign n15068 = n14279 & ~n15067;
  assign n15069 = ~n14274 & ~n15049;
  assign n15070 = ~n14292 & ~n14316;
  assign n15071 = ~n14300 & n15070;
  assign n15072 = n15069 & n15071;
  assign n15073 = ~n14298 & n15072;
  assign n15074 = n14185 & ~n15073;
  assign n15075 = ~n15068 & ~n15074;
  assign n15076 = ~n15065 & n15075;
  assign n15077 = n15063 & n15076;
  assign n15078 = ~n15060 & n15077;
  assign n15079 = n15056 & n15078;
  assign n15080 = ~n14278 & n15079;
  assign n15081 = ~n15052 & n15080;
  assign n15082 = n14296 & n15081;
  assign n15083 = ~n14271 & n15082;
  assign n15084 = ~n15048 & n15083;
  assign n15085 = n15084 ^ n11855;
  assign n15086 = n15085 ^ x664;
  assign n15087 = ~n15047 & ~n15086;
  assign n15088 = n15010 & n15087;
  assign n15089 = n15047 & ~n15086;
  assign n15090 = n14978 & ~n15008;
  assign n15091 = n14837 & n15090;
  assign n15092 = n14873 & n15091;
  assign n15093 = n15089 & n15092;
  assign n15094 = ~n15088 & ~n15093;
  assign n15095 = ~n14978 & n15008;
  assign n15096 = n14874 & n15095;
  assign n15097 = ~n15047 & n15086;
  assign n15098 = n15096 & n15097;
  assign n15099 = n14837 & n14873;
  assign n15100 = n15095 & n15099;
  assign n15101 = n14837 & ~n14873;
  assign n15102 = n14978 & n15008;
  assign n15103 = n15101 & n15102;
  assign n15104 = ~n15100 & ~n15103;
  assign n15105 = n15087 & ~n15104;
  assign n15106 = ~n15098 & ~n15105;
  assign n15107 = n15047 & n15086;
  assign n15108 = n15010 & n15107;
  assign n15109 = n14874 & n15102;
  assign n15110 = n15087 & n15109;
  assign n15111 = n15099 & n15102;
  assign n15112 = n15095 & n15101;
  assign n15113 = ~n15111 & ~n15112;
  assign n15114 = n15089 & ~n15113;
  assign n15115 = ~n15110 & ~n15114;
  assign n15116 = ~n15108 & n15115;
  assign n15117 = n15096 & n15107;
  assign n15118 = n15097 & n15109;
  assign n15119 = ~n15117 & ~n15118;
  assign n15120 = ~n14837 & n14873;
  assign n15121 = n15009 & n15120;
  assign n15122 = n15008 ^ n14873;
  assign n15123 = ~n14837 & ~n15122;
  assign n15124 = ~n15121 & ~n15123;
  assign n15125 = n15089 & ~n15124;
  assign n15126 = n15095 & n15120;
  assign n15127 = ~n15111 & ~n15126;
  assign n15128 = n15009 & n15101;
  assign n15129 = ~n15092 & ~n15128;
  assign n15130 = n15127 & n15129;
  assign n15131 = n15087 & ~n15130;
  assign n15132 = n15009 & n15099;
  assign n15133 = ~n14873 & n15091;
  assign n15134 = ~n15132 & ~n15133;
  assign n15135 = n15102 & n15120;
  assign n15136 = ~n15100 & ~n15135;
  assign n15137 = ~n15121 & ~n15128;
  assign n15138 = n15136 & n15137;
  assign n15139 = n15134 & n15138;
  assign n15140 = n15097 & ~n15139;
  assign n15141 = n14978 ^ n14837;
  assign n15142 = ~n15008 & n15141;
  assign n15143 = ~n15126 & ~n15142;
  assign n15144 = ~n15103 & n15143;
  assign n15145 = n15107 & ~n15144;
  assign n15146 = ~n15140 & ~n15145;
  assign n15147 = ~n15131 & n15146;
  assign n15148 = ~n15125 & n15147;
  assign n15149 = n15119 & n15148;
  assign n15150 = n15116 & n15149;
  assign n15151 = n15106 & n15150;
  assign n15152 = n15094 & n15151;
  assign n15153 = n15152 ^ n14183;
  assign n15154 = n15153 ^ x700;
  assign n15155 = ~n14718 & n15154;
  assign n15156 = n15007 ^ x663;
  assign n15157 = n14793 & n14805;
  assign n15158 = ~n14806 & ~n15157;
  assign n15159 = n14721 & ~n15158;
  assign n15160 = n14780 & n14799;
  assign n15161 = n14796 & ~n14800;
  assign n15162 = ~n15160 & ~n15161;
  assign n15163 = ~n15159 & n15162;
  assign n15164 = n14782 & ~n14821;
  assign n15165 = n14776 & ~n14801;
  assign n15166 = ~n15164 & ~n15165;
  assign n15167 = n14789 & n14796;
  assign n15168 = n14790 & ~n14824;
  assign n15169 = n14780 & ~n15168;
  assign n15170 = ~n15167 & ~n15169;
  assign n15171 = ~n14808 & ~n14813;
  assign n15172 = n14721 & ~n15171;
  assign n15173 = n14721 & n14798;
  assign n15174 = n14780 & ~n15158;
  assign n15175 = ~n15173 & ~n15174;
  assign n15176 = ~n14812 & n15175;
  assign n15177 = n14780 & ~n14809;
  assign n15178 = ~n14774 & n14815;
  assign n15179 = n14776 & ~n15178;
  assign n15180 = ~n15177 & ~n15179;
  assign n15181 = n14807 & ~n14821;
  assign n15182 = ~n14778 & ~n14794;
  assign n15183 = n14721 & ~n15182;
  assign n15184 = ~n14814 & n14818;
  assign n15185 = n14796 & ~n15184;
  assign n15186 = ~n15183 & ~n15185;
  assign n15187 = ~n15181 & n15186;
  assign n15188 = n15180 & n15187;
  assign n15189 = n15176 & n15188;
  assign n15190 = ~n15172 & n15189;
  assign n15191 = n15170 & n15190;
  assign n15192 = n15166 & n15191;
  assign n15193 = n15163 & n15192;
  assign n15194 = n15193 ^ n12223;
  assign n15195 = n15194 ^ x659;
  assign n15196 = n13786 & n13820;
  assign n15197 = n13594 & ~n13831;
  assign n15198 = ~n15196 & ~n15197;
  assign n15199 = n13791 & n13809;
  assign n15200 = n13594 & n13794;
  assign n15201 = ~n15199 & ~n15200;
  assign n15202 = ~n13785 & n15201;
  assign n15203 = n13594 & n13806;
  assign n15204 = ~n13820 & ~n13832;
  assign n15205 = n13796 & ~n15204;
  assign n15206 = ~n15203 & ~n15205;
  assign n15207 = ~n13814 & ~n13817;
  assign n15208 = n13839 & n15207;
  assign n15209 = n13796 & ~n15208;
  assign n15210 = ~n13784 & n13837;
  assign n15211 = ~n13838 & n15210;
  assign n15212 = n13791 & ~n15211;
  assign n15213 = ~n15209 & ~n15212;
  assign n15214 = ~n13799 & ~n13816;
  assign n15215 = n13594 & ~n15214;
  assign n15216 = ~n13809 & n15207;
  assign n15217 = ~n13784 & n15216;
  assign n15218 = ~n13829 & n15217;
  assign n15219 = ~n13804 & n15218;
  assign n15220 = n13786 & ~n15219;
  assign n15221 = ~n15215 & ~n15220;
  assign n15222 = n15213 & n15221;
  assign n15223 = n13813 & n15222;
  assign n15224 = ~n13808 & n15223;
  assign n15225 = n15206 & n15224;
  assign n15226 = n15202 & n15225;
  assign n15227 = n15198 & n15226;
  assign n15228 = n13802 & n15227;
  assign n15229 = n15228 ^ n12086;
  assign n15230 = n15229 ^ x660;
  assign n15231 = n15195 & n15230;
  assign n15232 = n14061 & n14080;
  assign n15233 = n14073 & n15020;
  assign n15234 = ~n14065 & n15233;
  assign n15235 = ~n13889 & ~n15234;
  assign n15236 = ~n15232 & ~n15235;
  assign n15237 = ~n14079 & n14086;
  assign n15238 = ~n14057 & ~n14081;
  assign n15239 = ~n14075 & n15238;
  assign n15240 = n14089 & n15239;
  assign n15241 = n14063 & ~n15240;
  assign n15242 = n14082 & n14101;
  assign n15243 = ~n14072 & n15242;
  assign n15244 = n13890 & ~n15243;
  assign n15245 = ~n15241 & ~n15244;
  assign n15246 = ~n15237 & n15245;
  assign n15247 = n15236 & n15246;
  assign n15248 = n15013 & n15247;
  assign n15249 = n14060 & n15248;
  assign n15250 = ~n15024 & n15249;
  assign n15251 = n15250 ^ n11633;
  assign n15252 = n15251 ^ x661;
  assign n15253 = n15085 ^ x662;
  assign n15254 = n15252 & ~n15253;
  assign n15255 = n15231 & n15254;
  assign n15256 = ~n15195 & n15230;
  assign n15257 = ~n15252 & ~n15253;
  assign n15258 = n15256 & n15257;
  assign n15259 = ~n15255 & ~n15258;
  assign n15260 = n15156 & ~n15259;
  assign n15261 = ~n13488 & ~n13493;
  assign n15262 = n13459 & ~n15261;
  assign n15263 = ~n13463 & ~n13484;
  assign n15264 = n13469 & ~n15263;
  assign n15265 = ~n15262 & ~n15264;
  assign n15266 = n13469 & n13482;
  assign n15267 = ~n13477 & ~n13488;
  assign n15268 = n13469 & ~n15267;
  assign n15269 = ~n13471 & ~n13503;
  assign n15270 = n13467 & ~n15269;
  assign n15271 = ~n15268 & ~n15270;
  assign n15272 = ~n15266 & n15271;
  assign n15273 = ~n13474 & ~n13492;
  assign n15274 = n13489 & n15273;
  assign n15275 = n13486 & n15274;
  assign n15276 = ~n13463 & n15275;
  assign n15277 = n13464 & n15276;
  assign n15278 = ~n13164 & ~n13494;
  assign n15279 = n15263 & n15278;
  assign n15280 = n13501 & n15279;
  assign n15281 = n13459 & ~n15280;
  assign n15282 = ~n15277 & ~n15281;
  assign n15283 = ~n13164 & n15273;
  assign n15284 = n13469 & ~n15283;
  assign n15285 = ~n13481 & ~n13494;
  assign n15286 = ~n13493 & n15285;
  assign n15287 = ~n13477 & n15286;
  assign n15288 = n15263 & n15287;
  assign n15289 = n13467 & ~n15288;
  assign n15290 = ~n15284 & ~n15289;
  assign n15291 = n15282 & n15290;
  assign n15292 = n15272 & n15291;
  assign n15293 = n15265 & n15292;
  assign n15294 = n15293 ^ n11045;
  assign n15295 = n15294 ^ x658;
  assign n15296 = n15156 & ~n15295;
  assign n15297 = ~n15195 & ~n15230;
  assign n15298 = n15254 & n15297;
  assign n15299 = n15195 & ~n15230;
  assign n15300 = ~n15252 & n15299;
  assign n15301 = ~n15256 & ~n15300;
  assign n15302 = n15253 & ~n15301;
  assign n15303 = n15252 ^ n15230;
  assign n15304 = n15253 ^ n15230;
  assign n15305 = n15303 & ~n15304;
  assign n15306 = n15195 & n15305;
  assign n15307 = ~n15302 & ~n15306;
  assign n15308 = ~n15298 & n15307;
  assign n15309 = n15296 & ~n15308;
  assign n15310 = ~n15260 & ~n15309;
  assign n15311 = ~n15156 & ~n15295;
  assign n15312 = n15252 & n15253;
  assign n15313 = ~n15195 & n15312;
  assign n15314 = n15231 & n15257;
  assign n15315 = ~n15298 & ~n15314;
  assign n15316 = ~n15313 & n15315;
  assign n15317 = n15230 ^ n15195;
  assign n15318 = n15253 ^ n15252;
  assign n15319 = ~n15303 & ~n15318;
  assign n15320 = ~n15317 & n15319;
  assign n15321 = n15316 & ~n15320;
  assign n15322 = ~n15302 & n15321;
  assign n15323 = n15311 & ~n15322;
  assign n15324 = ~n15156 & n15295;
  assign n15325 = n15231 & n15252;
  assign n15326 = n15253 & n15300;
  assign n15327 = ~n15325 & ~n15326;
  assign n15328 = n15316 & n15327;
  assign n15329 = ~n15258 & n15328;
  assign n15330 = n15324 & n15329;
  assign n15331 = n15156 & n15295;
  assign n15332 = n15231 & n15253;
  assign n15333 = n15299 & n15312;
  assign n15334 = ~n15254 & n15297;
  assign n15335 = ~n15333 & ~n15334;
  assign n15336 = ~n15332 & n15335;
  assign n15337 = n15331 & ~n15336;
  assign n15338 = ~n15330 & ~n15337;
  assign n15339 = ~n15323 & n15338;
  assign n15340 = n15310 & n15339;
  assign n15341 = n15340 ^ n14194;
  assign n15342 = n15341 ^ x702;
  assign n15343 = n14592 & n14624;
  assign n15344 = ~n14620 & ~n15343;
  assign n15345 = n14607 & ~n14616;
  assign n15346 = n14520 & n14609;
  assign n15347 = ~n14606 & ~n14628;
  assign n15348 = n14604 & ~n15347;
  assign n15349 = ~n15346 & ~n15348;
  assign n15350 = ~n15345 & n15349;
  assign n15351 = n14518 & n14594;
  assign n15352 = n14520 & n14599;
  assign n15353 = ~n15351 & ~n15352;
  assign n15354 = ~n14616 & n14622;
  assign n15355 = ~n14586 & ~n14598;
  assign n15356 = n14604 & ~n15355;
  assign n15357 = ~n15354 & ~n15356;
  assign n15358 = ~n14617 & ~n14624;
  assign n15359 = n14584 & ~n15358;
  assign n15360 = n14600 & ~n14609;
  assign n15361 = n14592 & ~n15360;
  assign n15362 = ~n15359 & ~n15361;
  assign n15363 = n15357 & n15362;
  assign n15364 = n15353 & n15363;
  assign n15365 = n15350 & n15364;
  assign n15366 = n14591 & n15365;
  assign n15367 = ~n14845 & n15366;
  assign n15368 = n14843 & n15367;
  assign n15369 = n15344 & n15368;
  assign n15370 = n15369 ^ n12976;
  assign n15371 = n15370 ^ x681;
  assign n15372 = n14185 & n14300;
  assign n15373 = ~n14271 & ~n15372;
  assign n15374 = ~n14310 & ~n15064;
  assign n15375 = ~n15049 & ~n15057;
  assign n15376 = ~n14292 & n15375;
  assign n15377 = n14272 & ~n15376;
  assign n15378 = ~n15374 & ~n15377;
  assign n15379 = n14293 & n14310;
  assign n15380 = ~n14300 & n14317;
  assign n15381 = n14279 & ~n15380;
  assign n15382 = ~n14288 & ~n14311;
  assign n15383 = ~n14292 & ~n15054;
  assign n15384 = n15382 & n15383;
  assign n15385 = n14185 & ~n15384;
  assign n15386 = n15058 & n15383;
  assign n15387 = ~n14270 & n15386;
  assign n15388 = n14290 & ~n15387;
  assign n15389 = ~n15385 & ~n15388;
  assign n15390 = ~n15381 & n15389;
  assign n15391 = ~n15379 & n15390;
  assign n15392 = n15378 & n15391;
  assign n15393 = n14302 & n15392;
  assign n15394 = n14285 & n15393;
  assign n15395 = n15373 & n15394;
  assign n15396 = ~n15048 & n15395;
  assign n15397 = n15396 ^ n13328;
  assign n15398 = n15397 ^ x676;
  assign n15399 = n15371 & ~n15398;
  assign n15400 = n14943 & n14969;
  assign n15401 = ~n14955 & n14958;
  assign n15402 = ~n15400 & ~n15401;
  assign n15403 = n14877 & ~n14973;
  assign n15404 = n14945 & ~n14967;
  assign n15405 = ~n15403 & ~n15404;
  assign n15406 = n15402 & n15405;
  assign n15407 = n15406 ^ n13936;
  assign n15408 = n15407 ^ x678;
  assign n15409 = n14052 & ~n15021;
  assign n15410 = n13890 & ~n14077;
  assign n15411 = ~n15409 & ~n15410;
  assign n15412 = ~n14072 & ~n14099;
  assign n15413 = ~n14079 & ~n15412;
  assign n15414 = n13890 & ~n14087;
  assign n15415 = n15011 & n15239;
  assign n15416 = n14066 & n15415;
  assign n15417 = n14061 & ~n15416;
  assign n15418 = ~n14065 & n15238;
  assign n15419 = ~n14052 & n15418;
  assign n15420 = ~n14050 & n14087;
  assign n15421 = ~n14063 & n15420;
  assign n15422 = ~n15419 & ~n15421;
  assign n15423 = ~n14054 & ~n15422;
  assign n15424 = ~n14079 & ~n15423;
  assign n15425 = ~n15417 & ~n15424;
  assign n15426 = ~n15414 & n15425;
  assign n15427 = n15027 & n15426;
  assign n15428 = ~n15024 & n15427;
  assign n15429 = ~n15413 & n15428;
  assign n15430 = n15411 & n15429;
  assign n15431 = ~n15012 & n15430;
  assign n15432 = n15431 ^ n13959;
  assign n15433 = n15432 ^ x679;
  assign n15434 = n15408 & n15433;
  assign n15435 = n13791 & n13829;
  assign n15436 = n13796 & n13804;
  assign n15437 = n13594 & n13820;
  assign n15438 = ~n15436 & ~n15437;
  assign n15439 = ~n15435 & n15438;
  assign n15440 = n13796 & n13809;
  assign n15441 = ~n13811 & n15207;
  assign n15442 = n13594 & ~n15441;
  assign n15443 = ~n15440 & ~n15442;
  assign n15444 = n13840 & n15216;
  assign n15445 = n13791 & ~n15444;
  assign n15446 = ~n13814 & ~n13829;
  assign n15447 = n15214 & n15446;
  assign n15448 = n13796 & ~n15447;
  assign n15449 = n13835 & n13839;
  assign n15450 = n13786 & ~n15449;
  assign n15451 = ~n15448 & ~n15450;
  assign n15452 = ~n15445 & n15451;
  assign n15453 = n15443 & n15452;
  assign n15454 = ~n13795 & n15453;
  assign n15455 = n15206 & n15454;
  assign n15456 = n15439 & n15455;
  assign n15457 = n15198 & n15456;
  assign n15458 = ~n13785 & n15457;
  assign n15459 = n15458 ^ n13306;
  assign n15460 = n15459 ^ x677;
  assign n15461 = ~n14798 & ~n14824;
  assign n15462 = ~n14821 & ~n15461;
  assign n15463 = ~n14789 & ~n15157;
  assign n15464 = ~n14778 & n15463;
  assign n15465 = n14780 & ~n15464;
  assign n15466 = ~n15462 & ~n15465;
  assign n15467 = n14720 & n14807;
  assign n15468 = n14790 & n14800;
  assign n15469 = n14721 & ~n15468;
  assign n15470 = ~n14808 & n14818;
  assign n15471 = ~n14806 & n15470;
  assign n15472 = ~n14720 & n15471;
  assign n15473 = ~n14808 & ~n14817;
  assign n15474 = ~n14796 & n15473;
  assign n15475 = ~n14821 & ~n15474;
  assign n15476 = n14815 & ~n15475;
  assign n15477 = ~n15472 & ~n15476;
  assign n15478 = ~n15469 & ~n15477;
  assign n15479 = ~n15467 & n15478;
  assign n15480 = n15466 & n15479;
  assign n15481 = n15163 & n15480;
  assign n15482 = n14785 & n15481;
  assign n15483 = ~n14812 & n15482;
  assign n15484 = n15483 ^ n13091;
  assign n15485 = n15484 ^ x680;
  assign n15486 = ~n15460 & ~n15485;
  assign n15487 = n15434 & n15486;
  assign n15488 = n15399 & n15487;
  assign n15489 = ~n15408 & n15433;
  assign n15490 = n15486 & n15489;
  assign n15491 = ~n15460 & n15485;
  assign n15492 = n15408 & ~n15433;
  assign n15493 = n15491 & n15492;
  assign n15494 = ~n15490 & ~n15493;
  assign n15495 = n15399 & ~n15494;
  assign n15496 = ~n15488 & ~n15495;
  assign n15497 = ~n15408 & ~n15433;
  assign n15498 = n15491 & n15497;
  assign n15499 = n15399 & n15498;
  assign n15500 = n15371 & n15398;
  assign n15501 = n15460 & ~n15485;
  assign n15502 = n15434 & n15501;
  assign n15503 = n15489 & n15501;
  assign n15504 = n15460 & n15485;
  assign n15505 = n15492 & n15504;
  assign n15506 = ~n15503 & ~n15505;
  assign n15507 = ~n15502 & n15506;
  assign n15508 = n15500 & ~n15507;
  assign n15509 = ~n15499 & ~n15508;
  assign n15510 = n15398 ^ n15371;
  assign n15511 = n15497 & n15501;
  assign n15512 = ~n15510 & n15511;
  assign n15513 = ~n15371 & n15398;
  assign n15514 = n15489 & n15491;
  assign n15515 = n15486 & n15492;
  assign n15516 = ~n15514 & ~n15515;
  assign n15517 = n15434 & n15491;
  assign n15518 = n15497 & n15504;
  assign n15519 = ~n15517 & ~n15518;
  assign n15520 = ~n15487 & ~n15498;
  assign n15521 = n15506 & n15520;
  assign n15522 = n15519 & n15521;
  assign n15523 = n15516 & n15522;
  assign n15524 = n15513 & n15523;
  assign n15525 = n15492 & n15501;
  assign n15526 = n15519 & ~n15525;
  assign n15527 = ~n15502 & n15526;
  assign n15528 = n15399 & ~n15527;
  assign n15529 = ~n15524 & ~n15528;
  assign n15530 = n15516 & n15520;
  assign n15531 = n15500 & ~n15530;
  assign n15532 = ~n15371 & ~n15398;
  assign n15533 = n15434 & n15504;
  assign n15534 = n15494 & ~n15533;
  assign n15535 = n15521 & n15534;
  assign n15536 = n15532 & ~n15535;
  assign n15537 = ~n15531 & ~n15536;
  assign n15538 = n15529 & n15537;
  assign n15539 = ~n15512 & n15538;
  assign n15540 = n15509 & n15539;
  assign n15541 = n15496 & n15540;
  assign n15542 = n15541 ^ n14216;
  assign n15543 = n15542 ^ x704;
  assign n15544 = ~n15342 & n15543;
  assign n15545 = n14977 ^ x670;
  assign n15546 = n15459 ^ x675;
  assign n15547 = ~n15545 & ~n15546;
  assign n15548 = n13467 & n13492;
  assign n15549 = n13469 & n13495;
  assign n15550 = ~n15548 & ~n15549;
  assign n15551 = ~n13481 & n13504;
  assign n15552 = n13469 & ~n15551;
  assign n15553 = n13507 & n15285;
  assign n15554 = ~n13471 & n15553;
  assign n15555 = n13501 & n15554;
  assign n15556 = n13464 & ~n15555;
  assign n15557 = ~n15552 & ~n15556;
  assign n15558 = n13485 & n13508;
  assign n15559 = ~n13492 & n15558;
  assign n15560 = n13459 & ~n15559;
  assign n15561 = ~n13500 & n13507;
  assign n15562 = ~n13481 & n15561;
  assign n15563 = ~n13488 & n15562;
  assign n15564 = n13467 & ~n15563;
  assign n15565 = ~n15560 & ~n15564;
  assign n15566 = n15557 & n15565;
  assign n15567 = n13466 & n15566;
  assign n15568 = n15271 & n15567;
  assign n15569 = n15550 & n15568;
  assign n15570 = n15265 & n15569;
  assign n15571 = n15570 ^ n13382;
  assign n15572 = n15571 ^ x672;
  assign n15573 = n15397 ^ x674;
  assign n15574 = n15572 & ~n15573;
  assign n15575 = n15046 ^ x671;
  assign n15576 = n14449 & n14471;
  assign n15577 = ~n14979 & ~n15576;
  assign n15578 = ~n14492 & ~n14499;
  assign n15579 = ~n14466 & n15578;
  assign n15580 = ~n14447 & n15579;
  assign n15581 = n14449 & ~n15580;
  assign n15582 = n14454 & ~n14989;
  assign n15583 = ~n15581 & ~n15582;
  assign n15584 = n14359 & ~n14996;
  assign n15585 = ~n14485 & ~n14499;
  assign n15586 = n14459 & ~n15585;
  assign n15587 = ~n14451 & ~n14493;
  assign n15588 = ~n14459 & ~n14483;
  assign n15589 = ~n14359 & ~n14473;
  assign n15590 = ~n14481 & n15589;
  assign n15591 = ~n15588 & ~n15590;
  assign n15592 = n15587 & ~n15591;
  assign n15593 = ~n14480 & ~n15592;
  assign n15594 = ~n15586 & ~n15593;
  assign n15595 = ~n15584 & n15594;
  assign n15596 = n15583 & n15595;
  assign n15597 = n15577 & n15596;
  assign n15598 = n14469 & n15597;
  assign n15599 = n14464 & n15598;
  assign n15600 = n15599 ^ n13354;
  assign n15601 = n15600 ^ x673;
  assign n15602 = ~n15575 & ~n15601;
  assign n15603 = n15574 & n15602;
  assign n15604 = n15547 & n15603;
  assign n15605 = ~n15545 & n15546;
  assign n15606 = ~n15575 & n15601;
  assign n15607 = ~n15572 & ~n15573;
  assign n15608 = n15606 & n15607;
  assign n15609 = ~n15572 & n15573;
  assign n15610 = n15602 & n15609;
  assign n15611 = ~n15608 & ~n15610;
  assign n15612 = n15605 & ~n15611;
  assign n15613 = ~n15604 & ~n15612;
  assign n15614 = n15545 & ~n15546;
  assign n15615 = n15573 ^ n15572;
  assign n15616 = n15575 & n15601;
  assign n15617 = ~n15615 & n15616;
  assign n15618 = n15614 & n15617;
  assign n15619 = n15606 & n15609;
  assign n15620 = n15614 & n15619;
  assign n15621 = n15572 & n15573;
  assign n15622 = n15606 & n15621;
  assign n15623 = ~n15608 & ~n15622;
  assign n15624 = n15547 & ~n15623;
  assign n15625 = ~n15620 & ~n15624;
  assign n15626 = n15602 & n15621;
  assign n15627 = ~n15608 & ~n15626;
  assign n15628 = n15614 & ~n15627;
  assign n15629 = n15546 ^ n15545;
  assign n15630 = n15574 & n15606;
  assign n15631 = n15629 & n15630;
  assign n15632 = n15572 & n15616;
  assign n15633 = n15609 & n15616;
  assign n15634 = n15575 & ~n15601;
  assign n15635 = n15607 & n15634;
  assign n15636 = ~n15633 & ~n15635;
  assign n15637 = ~n15632 & n15636;
  assign n15638 = ~n15610 & n15637;
  assign n15639 = n15547 & ~n15638;
  assign n15640 = ~n15631 & ~n15639;
  assign n15641 = n15546 & ~n15636;
  assign n15642 = n15574 & n15634;
  assign n15643 = n15621 & n15634;
  assign n15644 = ~n15642 & ~n15643;
  assign n15645 = n15614 & ~n15644;
  assign n15646 = n15609 & n15634;
  assign n15647 = ~n15642 & ~n15646;
  assign n15648 = ~n15622 & n15647;
  assign n15649 = n15605 & ~n15648;
  assign n15650 = n15545 & n15546;
  assign n15651 = n15574 & n15616;
  assign n15652 = ~n15643 & ~n15651;
  assign n15653 = n15602 & n15607;
  assign n15654 = ~n15619 & ~n15653;
  assign n15655 = ~n15603 & ~n15610;
  assign n15656 = n15654 & n15655;
  assign n15657 = n15652 & n15656;
  assign n15658 = n15650 & ~n15657;
  assign n15659 = ~n15649 & ~n15658;
  assign n15660 = ~n15645 & n15659;
  assign n15661 = ~n15641 & n15660;
  assign n15662 = n15640 & n15661;
  assign n15663 = ~n15628 & n15662;
  assign n15664 = n15625 & n15663;
  assign n15665 = ~n15618 & n15664;
  assign n15666 = n15613 & n15665;
  assign n15667 = n15666 ^ n14267;
  assign n15668 = n15667 ^ x703;
  assign n15669 = n15544 & ~n15668;
  assign n15670 = ~n13799 & ~n13830;
  assign n15671 = n13791 & ~n15670;
  assign n15672 = ~n13794 & ~n13838;
  assign n15673 = ~n13814 & n15672;
  assign n15674 = n13796 & ~n15673;
  assign n15675 = ~n15671 & ~n15674;
  assign n15676 = n13594 & n13804;
  assign n15677 = ~n13806 & n13840;
  assign n15678 = n13786 & ~n15677;
  assign n15679 = ~n13816 & n15207;
  assign n15680 = n13786 & ~n15679;
  assign n15681 = ~n13783 & ~n13811;
  assign n15682 = n13791 & ~n15681;
  assign n15683 = ~n15680 & ~n15682;
  assign n15684 = n13796 & ~n13837;
  assign n15685 = ~n13789 & n15446;
  assign n15686 = ~n13809 & n15685;
  assign n15687 = n13594 & ~n15686;
  assign n15688 = ~n15684 & ~n15687;
  assign n15689 = n15683 & n15688;
  assign n15690 = n13803 & n15689;
  assign n15691 = ~n15678 & n15690;
  assign n15692 = ~n15676 & n15691;
  assign n15693 = n15675 & n15692;
  assign n15694 = n15439 & n15693;
  assign n15695 = n15202 & n15694;
  assign n15696 = n15695 ^ n13686;
  assign n15697 = n15696 ^ x643;
  assign n15698 = n14780 & n14807;
  assign n15699 = n14720 & n14774;
  assign n15700 = ~n15698 & ~n15699;
  assign n15701 = ~n14813 & ~n15157;
  assign n15702 = n14776 & ~n15701;
  assign n15703 = n14721 & ~n14800;
  assign n15704 = ~n15702 & ~n15703;
  assign n15705 = n15700 & n15704;
  assign n15706 = n14817 & ~n14821;
  assign n15707 = n14809 & ~n14824;
  assign n15708 = n14796 & ~n15707;
  assign n15709 = ~n14788 & ~n14798;
  assign n15710 = n14776 & ~n15709;
  assign n15711 = ~n14778 & n14790;
  assign n15712 = n14796 & ~n15711;
  assign n15713 = ~n15710 & ~n15712;
  assign n15714 = n14799 & ~n14821;
  assign n15715 = ~n14794 & n14825;
  assign n15716 = n14780 & ~n15715;
  assign n15717 = ~n14824 & n15470;
  assign n15718 = n14721 & ~n15717;
  assign n15719 = ~n15716 & ~n15718;
  assign n15720 = ~n15714 & n15719;
  assign n15721 = n15713 & n15720;
  assign n15722 = n14784 & n15721;
  assign n15723 = ~n15708 & n15722;
  assign n15724 = ~n15706 & n15723;
  assign n15725 = n15705 & n15724;
  assign n15726 = n15176 & n15725;
  assign n15727 = n15726 ^ n13710;
  assign n15728 = n15727 ^ x642;
  assign n15729 = n15697 & n15728;
  assign n15730 = n14936 ^ n14907;
  assign n15731 = n14906 & ~n15730;
  assign n15732 = ~n14878 & n15731;
  assign n15733 = n14906 & n14936;
  assign n15734 = n14878 & n15733;
  assign n15735 = ~n14950 & ~n15734;
  assign n15736 = n14942 & n15735;
  assign n15737 = n14969 & n15736;
  assign n15738 = n14936 & n14951;
  assign n15739 = n15738 ^ n15733;
  assign n15740 = ~n14907 & n15739;
  assign n15741 = n15740 ^ n15733;
  assign n15742 = n14942 & ~n15741;
  assign n15743 = ~n15732 & n15742;
  assign n15744 = n14945 & ~n15743;
  assign n15745 = ~n15737 & ~n15744;
  assign n15746 = n14878 & ~n14964;
  assign n15747 = ~n15738 & ~n15746;
  assign n15748 = n14877 & ~n15747;
  assign n15749 = n14878 & n14906;
  assign n15750 = n14907 & n15749;
  assign n15751 = n14907 ^ n14878;
  assign n15752 = n14936 & ~n15751;
  assign n15753 = n15752 ^ n14907;
  assign n15754 = ~n14906 & ~n15753;
  assign n15755 = ~n15750 & ~n15754;
  assign n15756 = n14958 & ~n15755;
  assign n15757 = ~n15748 & ~n15756;
  assign n15758 = n15745 & n15757;
  assign n15759 = ~n15732 & n15758;
  assign n15760 = n15759 ^ n13059;
  assign n15761 = n15760 ^ x641;
  assign n15762 = n14649 ^ x644;
  assign n15763 = n15761 & ~n15762;
  assign n15764 = n15729 & n15763;
  assign n15765 = n13469 & ~n15285;
  assign n15766 = n13467 & ~n13485;
  assign n15767 = ~n15765 & ~n15766;
  assign n15768 = n13459 & n15276;
  assign n15769 = n13469 & n13474;
  assign n15770 = n13490 & ~n15769;
  assign n15771 = ~n13501 & ~n15770;
  assign n15772 = n13496 & ~n13503;
  assign n15773 = n15263 & n15772;
  assign n15774 = ~n13488 & n15773;
  assign n15775 = n13464 & ~n15774;
  assign n15776 = ~n15771 & ~n15775;
  assign n15777 = ~n15768 & n15776;
  assign n15778 = n15767 & n15777;
  assign n15779 = n13473 & n15778;
  assign n15780 = n15550 & n15779;
  assign n15781 = n15272 & n15780;
  assign n15782 = n15781 ^ n12993;
  assign n15783 = n15782 ^ x640;
  assign n15784 = n14112 ^ x645;
  assign n15785 = n15783 & n15784;
  assign n15786 = n15697 & ~n15728;
  assign n15787 = n15763 & n15786;
  assign n15788 = n15785 & n15787;
  assign n15789 = ~n15783 & n15784;
  assign n15790 = ~n15697 & n15728;
  assign n15791 = ~n15761 & n15762;
  assign n15792 = n15790 & n15791;
  assign n15793 = ~n15697 & ~n15728;
  assign n15794 = ~n15761 & ~n15762;
  assign n15795 = n15793 & n15794;
  assign n15796 = ~n15792 & ~n15795;
  assign n15797 = n15789 & ~n15796;
  assign n15798 = ~n15788 & ~n15797;
  assign n15799 = n15761 & n15762;
  assign n15800 = n15790 & n15799;
  assign n15801 = n15789 & n15800;
  assign n15802 = n15783 & ~n15784;
  assign n15803 = n15791 & n15793;
  assign n15804 = n15802 & n15803;
  assign n15805 = ~n15801 & ~n15804;
  assign n15806 = n15729 & n15791;
  assign n15807 = n15729 & n15794;
  assign n15808 = ~n15806 & ~n15807;
  assign n15809 = n15785 & ~n15808;
  assign n15810 = n15805 & ~n15809;
  assign n15811 = n15789 & n15806;
  assign n15812 = ~n15783 & ~n15784;
  assign n15813 = n15763 & n15793;
  assign n15814 = n15812 & n15813;
  assign n15815 = ~n15811 & ~n15814;
  assign n15816 = ~n15785 & ~n15812;
  assign n15817 = n15786 & n15791;
  assign n15818 = n15790 & n15794;
  assign n15819 = ~n15817 & ~n15818;
  assign n15820 = ~n15816 & ~n15819;
  assign n15821 = n15729 & n15799;
  assign n15822 = n15763 & n15790;
  assign n15823 = ~n15821 & ~n15822;
  assign n15824 = n15786 & n15799;
  assign n15825 = n15796 & ~n15824;
  assign n15826 = n15823 & n15825;
  assign n15827 = ~n15807 & n15826;
  assign n15828 = n15802 & ~n15827;
  assign n15829 = ~n15820 & ~n15828;
  assign n15830 = ~n15800 & ~n15813;
  assign n15831 = n15785 & ~n15830;
  assign n15832 = n15793 & n15799;
  assign n15833 = n15786 & n15794;
  assign n15834 = ~n15817 & ~n15833;
  assign n15835 = ~n15832 & n15834;
  assign n15836 = n15789 & ~n15835;
  assign n15837 = ~n15787 & n15823;
  assign n15838 = ~n15803 & n15837;
  assign n15839 = n15812 & ~n15838;
  assign n15840 = ~n15836 & ~n15839;
  assign n15841 = ~n15831 & n15840;
  assign n15842 = n15829 & n15841;
  assign n15843 = n15815 & n15842;
  assign n15844 = n15810 & n15843;
  assign n15845 = n15798 & n15844;
  assign n15846 = ~n15764 & n15845;
  assign n15847 = n15846 ^ n14239;
  assign n15848 = n15847 ^ x701;
  assign n15849 = n15669 & ~n15848;
  assign n15850 = n15155 & n15849;
  assign n15851 = ~n14718 & ~n15154;
  assign n15852 = ~n15543 & ~n15848;
  assign n15853 = n15342 & n15852;
  assign n15854 = n15668 & n15853;
  assign n15855 = n15851 & n15854;
  assign n15856 = ~n15850 & ~n15855;
  assign n15857 = n14718 & ~n15154;
  assign n15858 = n15849 & n15857;
  assign n15859 = n15543 & n15668;
  assign n15860 = n15342 & n15859;
  assign n15861 = ~n15848 & n15860;
  assign n15862 = n15851 & n15861;
  assign n15863 = ~n15858 & ~n15862;
  assign n15864 = n14718 & n15154;
  assign n15865 = ~n15342 & n15848;
  assign n15866 = ~n15543 & n15865;
  assign n15867 = n15668 & n15866;
  assign n15868 = n15342 & ~n15668;
  assign n15869 = ~n15543 & n15868;
  assign n15870 = n15848 & n15869;
  assign n15871 = n15543 & n15868;
  assign n15872 = n15848 & n15871;
  assign n15873 = ~n15668 & n15866;
  assign n15874 = ~n15872 & ~n15873;
  assign n15875 = ~n15870 & n15874;
  assign n15876 = ~n15867 & n15875;
  assign n15877 = n15864 & ~n15876;
  assign n15878 = n15342 & ~n15543;
  assign n15879 = n15668 & n15878;
  assign n15880 = n15848 & n15879;
  assign n15881 = n15852 & n15868;
  assign n15882 = ~n15342 & n15852;
  assign n15883 = n15668 & n15882;
  assign n15884 = ~n15881 & ~n15883;
  assign n15885 = ~n15880 & n15884;
  assign n15886 = n15857 & ~n15885;
  assign n15887 = ~n15877 & ~n15886;
  assign n15888 = ~n15342 & n15859;
  assign n15889 = ~n15848 & n15888;
  assign n15890 = ~n15881 & ~n15889;
  assign n15891 = n15851 & ~n15890;
  assign n15892 = ~n15668 & n15882;
  assign n15893 = ~n15848 & n15871;
  assign n15894 = ~n15883 & ~n15893;
  assign n15895 = ~n15892 & n15894;
  assign n15896 = n15155 & ~n15895;
  assign n15897 = n15859 & n15865;
  assign n15898 = n15857 & n15897;
  assign n15899 = n15854 & n15864;
  assign n15900 = ~n15898 & ~n15899;
  assign n15901 = n15543 & n15865;
  assign n15902 = ~n15668 & n15901;
  assign n15903 = ~n15867 & ~n15902;
  assign n15904 = n15851 & ~n15903;
  assign n15905 = n15155 & n15897;
  assign n15906 = n15155 & n15872;
  assign n15907 = n15861 & n15864;
  assign n15908 = ~n15906 & ~n15907;
  assign n15909 = n15848 & n15860;
  assign n15910 = ~n15870 & ~n15909;
  assign n15911 = ~n15902 & n15910;
  assign n15912 = n15857 & ~n15911;
  assign n15913 = n15851 & ~n15874;
  assign n15914 = ~n15912 & ~n15913;
  assign n15915 = n15155 & ~n15910;
  assign n15916 = ~n15889 & ~n15892;
  assign n15917 = n15864 & ~n15916;
  assign n15918 = ~n15915 & ~n15917;
  assign n15919 = n15914 & n15918;
  assign n15920 = n15908 & n15919;
  assign n15921 = ~n15905 & n15920;
  assign n15922 = ~n15904 & n15921;
  assign n15923 = n15900 & n15922;
  assign n15924 = ~n15896 & n15923;
  assign n15925 = ~n15891 & n15924;
  assign n15926 = n15887 & n15925;
  assign n15927 = n15863 & n15926;
  assign n15928 = n15856 & n15927;
  assign n15929 = n15928 ^ n15085;
  assign n15930 = n15929 ^ x760;
  assign n15931 = n15296 & n15322;
  assign n15932 = ~n15308 & n15311;
  assign n15933 = ~n15931 & ~n15932;
  assign n15934 = n15324 & ~n15336;
  assign n15935 = ~n15329 & n15331;
  assign n15936 = ~n15934 & ~n15935;
  assign n15937 = n15933 & n15936;
  assign n15938 = n15259 & n15937;
  assign n15939 = n15938 ^ n13887;
  assign n15940 = n15939 ^ x735;
  assign n15941 = n14664 & ~n14700;
  assign n15942 = n14656 & ~n14689;
  assign n15943 = n14661 & n14701;
  assign n15944 = ~n15942 & ~n15943;
  assign n15945 = ~n15941 & n15944;
  assign n15946 = n14661 & n14680;
  assign n15947 = ~n14678 & ~n15946;
  assign n15948 = ~n14334 & ~n14702;
  assign n15949 = ~n14671 & ~n14694;
  assign n15950 = n15948 & n15949;
  assign n15951 = n14656 & ~n15950;
  assign n15952 = n13853 ^ n13520;
  assign n15953 = ~n14113 & n15952;
  assign n15954 = n14664 & n15953;
  assign n15955 = ~n15951 & ~n15954;
  assign n15956 = ~n14676 & ~n14691;
  assign n15957 = n15948 & n15956;
  assign n15958 = ~n14663 & n15957;
  assign n15959 = n14651 & ~n15958;
  assign n15960 = ~n14660 & ~n14692;
  assign n15961 = ~n14706 & ~n15960;
  assign n15962 = n14696 & n14700;
  assign n15963 = n14661 & ~n15962;
  assign n15964 = ~n15961 & ~n15963;
  assign n15965 = ~n15959 & n15964;
  assign n15966 = n15955 & n15965;
  assign n15967 = n15947 & n15966;
  assign n15968 = n14675 & n15967;
  assign n15969 = n15945 & n15968;
  assign n15970 = n15969 ^ n12925;
  assign n15971 = n15970 ^ x730;
  assign n15972 = ~n15940 & n15971;
  assign n15973 = ~n15525 & ~n15533;
  assign n15974 = ~n15518 & n15973;
  assign n15975 = n15399 & ~n15974;
  assign n15976 = n15486 & n15497;
  assign n15977 = ~n15493 & ~n15976;
  assign n15978 = n15513 & ~n15977;
  assign n15979 = ~n15515 & ~n15517;
  assign n15980 = n15500 & ~n15979;
  assign n15981 = ~n15978 & ~n15980;
  assign n15982 = ~n15518 & n15977;
  assign n15983 = n15500 & ~n15982;
  assign n15984 = ~n15503 & n15516;
  assign n15985 = n15399 & ~n15984;
  assign n15986 = ~n15983 & ~n15985;
  assign n15987 = n15523 & n15532;
  assign n15988 = n15521 & n15973;
  assign n15989 = n15513 & ~n15988;
  assign n15990 = ~n15987 & ~n15989;
  assign n15991 = n15986 & n15990;
  assign n15992 = ~n15488 & n15991;
  assign n15993 = n15981 & n15992;
  assign n15994 = n15509 & n15993;
  assign n15995 = ~n15975 & n15994;
  assign n15996 = n15995 ^ n14024;
  assign n15997 = n15996 ^ x734;
  assign n15998 = n15294 ^ x656;
  assign n15999 = ~n14592 & ~n14855;
  assign n16000 = ~n14594 & ~n14598;
  assign n16001 = n14584 & ~n16000;
  assign n16002 = ~n14582 & ~n14586;
  assign n16003 = n14592 & ~n16002;
  assign n16004 = ~n16001 & ~n16003;
  assign n16005 = ~n15999 & n16004;
  assign n16006 = n14518 & n14621;
  assign n16007 = ~n14595 & n14604;
  assign n16008 = ~n16006 & ~n16007;
  assign n16009 = ~n14616 & n14623;
  assign n16010 = n14520 & ~n14589;
  assign n16011 = ~n16009 & ~n16010;
  assign n16012 = n16008 & n16011;
  assign n16013 = n16005 & n16012;
  assign n16014 = n15350 & n16013;
  assign n16015 = n14851 & n16014;
  assign n16016 = n15344 & n16015;
  assign n16017 = n16016 ^ n13204;
  assign n16018 = n16017 ^ x655;
  assign n16019 = ~n15998 & n16018;
  assign n16020 = n14958 & n15743;
  assign n16021 = n14876 & n15732;
  assign n16022 = n14877 & ~n15736;
  assign n16023 = ~n16021 & ~n16022;
  assign n16024 = ~n16020 & n16023;
  assign n16025 = n14969 & ~n15747;
  assign n16026 = n14945 & ~n15755;
  assign n16027 = ~n16025 & ~n16026;
  assign n16028 = n16024 & n16027;
  assign n16029 = n16028 ^ n13176;
  assign n16030 = n16029 ^ x654;
  assign n16031 = n14516 ^ x653;
  assign n16032 = n16030 & ~n16031;
  assign n16033 = n16019 & n16032;
  assign n16034 = n15194 ^ x657;
  assign n16035 = n13852 ^ x652;
  assign n16036 = ~n16034 & ~n16035;
  assign n16037 = n15998 & ~n16018;
  assign n16038 = ~n16030 & n16031;
  assign n16039 = n16037 & n16038;
  assign n16040 = n16036 & n16039;
  assign n16041 = n16030 & n16031;
  assign n16042 = n16037 & n16041;
  assign n16043 = n16036 & n16042;
  assign n16044 = ~n16040 & ~n16043;
  assign n16045 = n16034 & n16035;
  assign n16046 = n16039 & n16045;
  assign n16047 = n15998 & n16018;
  assign n16048 = ~n16030 & ~n16031;
  assign n16049 = n16047 & n16048;
  assign n16050 = n16036 & n16049;
  assign n16051 = ~n16046 & ~n16050;
  assign n16052 = n16034 & ~n16035;
  assign n16053 = n16037 & n16048;
  assign n16054 = ~n16033 & ~n16053;
  assign n16055 = n16052 & ~n16054;
  assign n16056 = n16051 & ~n16055;
  assign n16057 = ~n16034 & n16035;
  assign n16058 = n16033 & n16057;
  assign n16059 = n16019 & n16041;
  assign n16060 = n16038 & n16047;
  assign n16061 = ~n16059 & ~n16060;
  assign n16062 = n16052 & ~n16061;
  assign n16063 = ~n16058 & ~n16062;
  assign n16064 = ~n15998 & ~n16018;
  assign n16065 = n16041 & n16064;
  assign n16066 = n16036 & n16065;
  assign n16067 = ~n16052 & ~n16057;
  assign n16068 = n16032 & n16064;
  assign n16069 = n16032 & n16047;
  assign n16070 = ~n16068 & ~n16069;
  assign n16071 = ~n16067 & ~n16070;
  assign n16072 = ~n16066 & ~n16071;
  assign n16073 = n16038 & n16064;
  assign n16074 = ~n16042 & ~n16073;
  assign n16075 = ~n16067 & ~n16074;
  assign n16076 = n16041 & n16047;
  assign n16077 = n16048 & n16064;
  assign n16078 = ~n16049 & ~n16077;
  assign n16079 = ~n16076 & n16078;
  assign n16080 = n16057 & ~n16079;
  assign n16081 = ~n16075 & ~n16080;
  assign n16082 = n16032 & n16037;
  assign n16083 = n16061 & ~n16082;
  assign n16084 = n16036 & ~n16083;
  assign n16085 = n16019 & n16048;
  assign n16086 = ~n16065 & ~n16085;
  assign n16087 = ~n16060 & n16086;
  assign n16088 = ~n16053 & n16087;
  assign n16089 = n16070 & n16088;
  assign n16090 = n16045 & ~n16089;
  assign n16091 = ~n16084 & ~n16090;
  assign n16092 = n16081 & n16091;
  assign n16093 = n16072 & n16092;
  assign n16094 = n16063 & n16093;
  assign n16095 = n16056 & n16094;
  assign n16096 = n16044 & n16095;
  assign n16097 = ~n16033 & n16096;
  assign n16098 = n16097 ^ n14046;
  assign n16099 = n16098 ^ x732;
  assign n16100 = ~n15997 & ~n16099;
  assign n16101 = n15614 & n15622;
  assign n16102 = n15629 & n15635;
  assign n16103 = ~n16101 & ~n16102;
  assign n16104 = n15607 & n15616;
  assign n16105 = n15652 & ~n16104;
  assign n16106 = n15605 & ~n16105;
  assign n16107 = ~n15646 & n15654;
  assign n16108 = ~n15630 & n16107;
  assign n16109 = n15650 & ~n16108;
  assign n16110 = n15614 & ~n15655;
  assign n16111 = n15574 & n15575;
  assign n16112 = ~n15646 & ~n16111;
  assign n16113 = ~n15633 & n16112;
  assign n16114 = n15547 & ~n16113;
  assign n16115 = n15575 & n15650;
  assign n16116 = n15572 & n16115;
  assign n16117 = ~n16114 & ~n16116;
  assign n16118 = ~n15547 & ~n15603;
  assign n16119 = ~n15626 & ~n15653;
  assign n16120 = ~n15605 & n16119;
  assign n16121 = ~n16118 & ~n16120;
  assign n16122 = ~n15622 & ~n16121;
  assign n16123 = ~n15545 & ~n16122;
  assign n16124 = n16117 & ~n16123;
  assign n16125 = ~n15628 & n16124;
  assign n16126 = ~n16110 & n16125;
  assign n16127 = n15613 & n16126;
  assign n16128 = ~n16109 & n16127;
  assign n16129 = ~n16106 & n16128;
  assign n16130 = n16103 & n16129;
  assign n16131 = ~n15618 & n16130;
  assign n16132 = n16131 ^ n13457;
  assign n16133 = n16132 ^ x731;
  assign n16134 = n15785 & n15792;
  assign n16135 = n15812 & ~n15834;
  assign n16136 = ~n16134 & ~n16135;
  assign n16137 = ~n15787 & ~n15822;
  assign n16138 = n15802 & ~n16137;
  assign n16139 = n15823 & n15830;
  assign n16140 = n15812 & ~n16139;
  assign n16141 = ~n15764 & ~n15824;
  assign n16142 = ~n15818 & n16141;
  assign n16143 = ~n15806 & n16142;
  assign n16144 = ~n15813 & n16143;
  assign n16145 = n15802 & ~n16144;
  assign n16146 = ~n16140 & ~n16145;
  assign n16147 = ~n15795 & ~n15832;
  assign n16148 = ~n15821 & n16147;
  assign n16149 = ~n15787 & n16148;
  assign n16150 = ~n15813 & n16149;
  assign n16151 = n15785 & ~n16150;
  assign n16152 = ~n15792 & ~n15807;
  assign n16153 = n15812 & ~n16152;
  assign n16154 = ~n15822 & n16141;
  assign n16155 = ~n15833 & n16154;
  assign n16156 = ~n15803 & n16155;
  assign n16157 = ~n15807 & n16156;
  assign n16158 = n15789 & ~n16157;
  assign n16159 = ~n16153 & ~n16158;
  assign n16160 = ~n16151 & n16159;
  assign n16161 = n16146 & n16160;
  assign n16162 = ~n16138 & n16161;
  assign n16163 = n16136 & n16162;
  assign n16164 = n15810 & n16163;
  assign n16165 = ~n15811 & n16164;
  assign n16166 = n16165 ^ n13924;
  assign n16167 = n16166 ^ x733;
  assign n16168 = n16133 & ~n16167;
  assign n16169 = n16100 & n16168;
  assign n16170 = n15972 & n16169;
  assign n16171 = n15940 & n15971;
  assign n16172 = n15997 & n16099;
  assign n16173 = ~n16133 & n16167;
  assign n16174 = n16172 & n16173;
  assign n16175 = n16100 & n16173;
  assign n16176 = ~n16174 & ~n16175;
  assign n16177 = n16171 & ~n16176;
  assign n16178 = ~n16170 & ~n16177;
  assign n16179 = n16099 ^ n15997;
  assign n16180 = n16168 & n16179;
  assign n16181 = n16171 & n16180;
  assign n16182 = n15940 & ~n15971;
  assign n16183 = ~n15997 & n16099;
  assign n16184 = n16133 & n16167;
  assign n16185 = n16183 & n16184;
  assign n16186 = n16168 & n16172;
  assign n16187 = ~n16185 & ~n16186;
  assign n16188 = ~n16169 & n16187;
  assign n16189 = n16182 & ~n16188;
  assign n16190 = ~n16181 & ~n16189;
  assign n16191 = ~n15940 & ~n15971;
  assign n16192 = n16173 & n16183;
  assign n16193 = n15997 & ~n16099;
  assign n16194 = n16173 & n16193;
  assign n16195 = ~n16192 & ~n16194;
  assign n16196 = n16191 & ~n16195;
  assign n16197 = ~n16133 & ~n16167;
  assign n16198 = n16183 & n16197;
  assign n16199 = n16172 & n16197;
  assign n16200 = ~n16198 & ~n16199;
  assign n16201 = n15972 & ~n16200;
  assign n16202 = ~n16196 & ~n16201;
  assign n16203 = n16172 & n16184;
  assign n16204 = n16191 & n16203;
  assign n16205 = n16182 & n16192;
  assign n16206 = ~n16204 & ~n16205;
  assign n16207 = n16182 & n16203;
  assign n16208 = n16100 & n16197;
  assign n16209 = n16171 & n16208;
  assign n16210 = ~n16207 & ~n16209;
  assign n16211 = n15972 & n16174;
  assign n16212 = n16193 & n16197;
  assign n16213 = n16191 & n16212;
  assign n16214 = ~n16211 & ~n16213;
  assign n16215 = n16100 & n16184;
  assign n16216 = ~n16199 & ~n16212;
  assign n16217 = ~n16215 & n16216;
  assign n16218 = n16182 & ~n16217;
  assign n16219 = n16184 & n16193;
  assign n16220 = ~n16192 & ~n16219;
  assign n16221 = ~n16198 & n16220;
  assign n16222 = n16171 & ~n16221;
  assign n16223 = ~n16215 & ~n16219;
  assign n16224 = ~n16186 & n16223;
  assign n16225 = ~n16191 & n16224;
  assign n16226 = ~n16180 & ~n16215;
  assign n16227 = ~n15972 & n16226;
  assign n16228 = ~n16225 & ~n16227;
  assign n16229 = ~n16208 & ~n16228;
  assign n16230 = ~n15940 & ~n16229;
  assign n16231 = ~n16222 & ~n16230;
  assign n16232 = ~n16218 & n16231;
  assign n16233 = n16214 & n16232;
  assign n16234 = n16210 & n16233;
  assign n16235 = n16206 & n16234;
  assign n16236 = n16202 & n16235;
  assign n16237 = n16190 & n16236;
  assign n16238 = n16178 & n16237;
  assign n16239 = n16238 ^ n15046;
  assign n16240 = n16239 ^ x765;
  assign n16241 = n15930 & n16240;
  assign n16242 = n15760 ^ x687;
  assign n16243 = n15484 ^ x682;
  assign n16244 = ~n16242 & n16243;
  assign n16245 = n15782 ^ x686;
  assign n16246 = n14274 & ~n14310;
  assign n16247 = n14185 & n14293;
  assign n16248 = ~n16246 & ~n16247;
  assign n16249 = ~n15057 & n15071;
  assign n16250 = n14290 & ~n16249;
  assign n16251 = n14317 & n15382;
  assign n16252 = n14149 & ~n16251;
  assign n16253 = ~n16250 & ~n16252;
  assign n16254 = n14240 & n14281;
  assign n16255 = n14279 & n16254;
  assign n16256 = n14320 & n15384;
  assign n16257 = n14272 & ~n16256;
  assign n16258 = ~n16255 & ~n16257;
  assign n16259 = n16253 & n16258;
  assign n16260 = n16248 & n16259;
  assign n16261 = ~n15052 & n16260;
  assign n16262 = n15373 & n16261;
  assign n16263 = ~n15048 & n16262;
  assign n16264 = n16263 ^ n12946;
  assign n16265 = n16264 ^ x684;
  assign n16266 = n16245 & n16265;
  assign n16267 = n15370 ^ x683;
  assign n16268 = n14359 & n14493;
  assign n16269 = n14454 & ~n14996;
  assign n16270 = ~n16268 & ~n16269;
  assign n16271 = ~n14480 & ~n14498;
  assign n16272 = n14994 & n14995;
  assign n16273 = ~n14481 & n16272;
  assign n16274 = n14449 & ~n16273;
  assign n16275 = ~n16271 & ~n16274;
  assign n16276 = ~n14467 & ~n14483;
  assign n16277 = n14459 & ~n16276;
  assign n16278 = n14486 & n15587;
  assign n16279 = n14454 & ~n16278;
  assign n16280 = ~n14359 & n15578;
  assign n16281 = ~n14459 & n14501;
  assign n16282 = ~n16280 & ~n16281;
  assign n16283 = ~n14480 & n16282;
  assign n16284 = ~n16279 & ~n16283;
  assign n16285 = ~n16277 & n16284;
  assign n16286 = n16275 & n16285;
  assign n16287 = n16270 & n16286;
  assign n16288 = n15577 & n16287;
  assign n16289 = n14478 & n16288;
  assign n16290 = n14464 & n16289;
  assign n16291 = n16290 ^ n13025;
  assign n16292 = n16291 ^ x685;
  assign n16293 = ~n16267 & n16292;
  assign n16294 = n16266 & n16293;
  assign n16295 = ~n16245 & n16265;
  assign n16296 = n16293 & n16295;
  assign n16297 = ~n16294 & ~n16296;
  assign n16298 = n16244 & ~n16297;
  assign n16299 = n16242 & ~n16243;
  assign n16300 = n16267 & ~n16292;
  assign n16301 = n16266 & n16300;
  assign n16302 = ~n16245 & ~n16265;
  assign n16303 = n16267 & n16292;
  assign n16304 = n16302 & n16303;
  assign n16305 = n16266 & n16303;
  assign n16306 = ~n16304 & ~n16305;
  assign n16307 = ~n16301 & n16306;
  assign n16308 = n16299 & ~n16307;
  assign n16309 = ~n16298 & ~n16308;
  assign n16310 = ~n16242 & ~n16243;
  assign n16311 = ~n16267 & ~n16292;
  assign n16312 = n16295 & n16311;
  assign n16313 = n16245 & ~n16265;
  assign n16314 = n16311 & n16313;
  assign n16315 = ~n16312 & ~n16314;
  assign n16316 = n16310 & ~n16315;
  assign n16317 = n16244 & n16314;
  assign n16318 = n16302 & n16311;
  assign n16319 = n16243 & n16318;
  assign n16320 = ~n16317 & ~n16319;
  assign n16321 = n16303 & n16313;
  assign n16322 = n16299 & n16321;
  assign n16323 = n16266 & n16311;
  assign n16324 = n16242 & n16243;
  assign n16325 = ~n16310 & ~n16324;
  assign n16326 = n16323 & ~n16325;
  assign n16327 = ~n16322 & ~n16326;
  assign n16328 = n16320 & n16327;
  assign n16329 = n16296 & n16310;
  assign n16330 = n16293 & n16313;
  assign n16331 = n16293 & n16302;
  assign n16332 = ~n16330 & ~n16331;
  assign n16333 = n16324 & ~n16332;
  assign n16334 = n16304 & n16310;
  assign n16335 = n16295 & n16300;
  assign n16336 = n16324 & n16335;
  assign n16337 = ~n16334 & ~n16336;
  assign n16338 = n16315 & ~n16323;
  assign n16339 = ~n16296 & n16338;
  assign n16340 = n16299 & ~n16339;
  assign n16341 = n16300 & n16313;
  assign n16342 = ~n16335 & ~n16341;
  assign n16343 = ~n16304 & n16342;
  assign n16344 = ~n16301 & n16343;
  assign n16345 = n16244 & ~n16344;
  assign n16346 = n16300 & n16302;
  assign n16347 = ~n16321 & ~n16346;
  assign n16348 = ~n16324 & n16347;
  assign n16349 = n16295 & n16303;
  assign n16350 = ~n16346 & ~n16349;
  assign n16351 = ~n16310 & n16350;
  assign n16352 = ~n16348 & ~n16351;
  assign n16353 = ~n16305 & ~n16352;
  assign n16354 = ~n16325 & ~n16353;
  assign n16355 = ~n16345 & ~n16354;
  assign n16356 = ~n16340 & n16355;
  assign n16357 = n16337 & n16356;
  assign n16358 = ~n16333 & n16357;
  assign n16359 = ~n16329 & n16358;
  assign n16360 = n16328 & n16359;
  assign n16361 = ~n16316 & n16360;
  assign n16362 = n16309 & n16361;
  assign n16363 = n16362 ^ n14935;
  assign n16364 = n16363 ^ x709;
  assign n16365 = n16036 & n16085;
  assign n16366 = n16067 & ~n16078;
  assign n16367 = n16054 & ~n16068;
  assign n16368 = ~n16082 & n16367;
  assign n16369 = n16057 & ~n16368;
  assign n16370 = ~n16366 & ~n16369;
  assign n16371 = ~n15998 & n16038;
  assign n16372 = ~n16076 & ~n16371;
  assign n16373 = ~n16059 & n16372;
  assign n16374 = n16052 & ~n16373;
  assign n16375 = ~n16033 & ~n16065;
  assign n16376 = n16045 & ~n16375;
  assign n16377 = ~n16374 & ~n16376;
  assign n16378 = n16036 & n16069;
  assign n16379 = ~n16059 & ~n16076;
  assign n16380 = n16036 & ~n16379;
  assign n16381 = ~n16039 & n16061;
  assign n16382 = ~n16042 & n16381;
  assign n16383 = n16045 & ~n16382;
  assign n16384 = ~n16380 & ~n16383;
  assign n16385 = ~n16060 & n16372;
  assign n16386 = n16057 & ~n16385;
  assign n16387 = ~n16082 & ~n16085;
  assign n16388 = ~n16068 & n16387;
  assign n16389 = ~n16053 & n16388;
  assign n16390 = n16052 & ~n16389;
  assign n16391 = ~n16386 & ~n16390;
  assign n16392 = n16384 & n16391;
  assign n16393 = n16044 & n16392;
  assign n16394 = ~n16378 & n16393;
  assign n16395 = n16377 & n16394;
  assign n16396 = n16370 & n16395;
  assign n16397 = ~n16365 & n16396;
  assign n16398 = n16397 ^ n13555;
  assign n16399 = n16398 ^ x710;
  assign n16400 = n15089 & n15109;
  assign n16401 = ~n14837 & n15090;
  assign n16402 = ~n15087 & ~n15107;
  assign n16403 = n16401 & ~n16402;
  assign n16404 = n14873 & n16403;
  assign n16405 = ~n16400 & ~n16404;
  assign n16406 = n15089 & ~n15136;
  assign n16407 = ~n14873 & n16401;
  assign n16408 = n15129 & ~n16407;
  assign n16409 = ~n15109 & n16408;
  assign n16410 = n15097 & ~n16409;
  assign n16411 = ~n15089 & ~n15107;
  assign n16412 = ~n15137 & ~n16411;
  assign n16413 = n15089 & n15090;
  assign n16414 = ~n14873 & n16413;
  assign n16415 = ~n16412 & ~n16414;
  assign n16416 = n15107 & n15132;
  assign n16417 = n15087 & ~n15134;
  assign n16418 = ~n16416 & ~n16417;
  assign n16419 = ~n15126 & ~n15135;
  assign n16420 = n15104 & n16419;
  assign n16421 = n15097 & ~n16420;
  assign n16422 = ~n15109 & n15113;
  assign n16423 = ~n15087 & n16422;
  assign n16424 = ~n15103 & n15127;
  assign n16425 = ~n15107 & n16424;
  assign n16426 = ~n16423 & ~n16425;
  assign n16427 = ~n15096 & ~n16426;
  assign n16428 = ~n16402 & ~n16427;
  assign n16429 = ~n16421 & ~n16428;
  assign n16430 = n16418 & n16429;
  assign n16431 = n16415 & n16430;
  assign n16432 = ~n16410 & n16431;
  assign n16433 = ~n16406 & n16432;
  assign n16434 = n16405 & n16433;
  assign n16435 = n15094 & n16434;
  assign n16436 = n16435 ^ n14905;
  assign n16437 = n16436 ^ x708;
  assign n16438 = ~n16399 & ~n16437;
  assign n16439 = ~n16364 & n16438;
  assign n16440 = n14717 ^ x707;
  assign n16445 = n16399 ^ n16364;
  assign n16441 = ~n16364 & n16437;
  assign n16442 = n16437 ^ n16399;
  assign n16443 = n16441 & n16442;
  assign n16444 = n16443 ^ n16442;
  assign n16446 = n16445 ^ n16444;
  assign n16447 = ~n16440 & ~n16446;
  assign n16448 = n16447 ^ n16445;
  assign n16449 = ~n16439 & n16448;
  assign n16450 = n15542 ^ x706;
  assign n16451 = n15802 & n15821;
  assign n16452 = n15785 & n15822;
  assign n16453 = ~n16451 & ~n16452;
  assign n16454 = n15764 & n15812;
  assign n16455 = n15789 & n15813;
  assign n16456 = ~n15789 & n15800;
  assign n16457 = n15808 & ~n15817;
  assign n16458 = ~n15803 & n16457;
  assign n16459 = n15802 & ~n16458;
  assign n16460 = ~n16456 & ~n16459;
  assign n16461 = n15823 & n16141;
  assign n16462 = n15789 & ~n16461;
  assign n16463 = ~n15807 & n15834;
  assign n16464 = ~n15812 & n16463;
  assign n16465 = n15808 & n15819;
  assign n16466 = ~n15785 & n16465;
  assign n16467 = ~n16464 & ~n16466;
  assign n16468 = ~n15832 & ~n16467;
  assign n16469 = ~n15816 & ~n16468;
  assign n16470 = ~n16462 & ~n16469;
  assign n16471 = n16460 & n16470;
  assign n16472 = ~n16134 & n16471;
  assign n16473 = ~n16455 & n16472;
  assign n16474 = ~n16454 & n16473;
  assign n16475 = n16453 & n16474;
  assign n16476 = ~n16138 & n16475;
  assign n16477 = n15798 & n16476;
  assign n16478 = n15815 & n16477;
  assign n16479 = n16478 ^ n13780;
  assign n16480 = n16479 ^ x711;
  assign n16481 = n16450 & ~n16480;
  assign n16482 = n16449 & n16481;
  assign n16483 = ~n16450 & n16480;
  assign n16484 = n16399 & n16441;
  assign n16485 = n16364 & ~n16437;
  assign n16486 = n16440 & n16485;
  assign n16487 = n16364 & n16399;
  assign n16488 = n16364 ^ x708;
  assign n16489 = n16488 ^ n16436;
  assign n16490 = n16487 & ~n16489;
  assign n16491 = n16490 ^ n16489;
  assign n16492 = ~n16440 & ~n16491;
  assign n16493 = ~n16439 & ~n16492;
  assign n16494 = ~n16486 & n16493;
  assign n16495 = ~n16484 & n16494;
  assign n16496 = n16483 & ~n16495;
  assign n16497 = ~n16482 & ~n16496;
  assign n16498 = ~n16364 & ~n16399;
  assign n16499 = ~n16440 & n16498;
  assign n16500 = n16440 ^ n16437;
  assign n16501 = n16399 & ~n16500;
  assign n16502 = ~n16438 & n16440;
  assign n16503 = n16364 & n16502;
  assign n16504 = ~n16501 & ~n16503;
  assign n16505 = ~n16499 & n16504;
  assign n16506 = ~n16450 & ~n16480;
  assign n16507 = ~n16505 & n16506;
  assign n16508 = n16450 & n16480;
  assign n16509 = n16399 & ~n16437;
  assign n16510 = ~n16364 & n16440;
  assign n16511 = n16509 & n16510;
  assign n16512 = ~n16399 & n16441;
  assign n16513 = n16512 ^ n16487;
  assign n16514 = n16440 & n16513;
  assign n16515 = n16514 ^ n16487;
  assign n16516 = ~n16511 & ~n16515;
  assign n16517 = n16437 & n16487;
  assign n16518 = ~n16364 & n16399;
  assign n16519 = n16518 ^ n16437;
  assign n16520 = ~n16440 & ~n16519;
  assign n16521 = ~n16517 & ~n16520;
  assign n16522 = n16516 & n16521;
  assign n16523 = n16508 & ~n16522;
  assign n16524 = ~n16507 & ~n16523;
  assign n16525 = n16497 & n16524;
  assign n16526 = n16525 ^ n14977;
  assign n16527 = n16526 ^ x764;
  assign n16528 = n15939 ^ x689;
  assign n16529 = ~n14663 & ~n14701;
  assign n16530 = ~n14669 & n16529;
  assign n16531 = n14651 & ~n16530;
  assign n16532 = n14656 & n14701;
  assign n16533 = ~n16531 & ~n16532;
  assign n16534 = n14661 & ~n14700;
  assign n16535 = ~n14692 & n15956;
  assign n16536 = n14664 & ~n16535;
  assign n16537 = n14651 & n14695;
  assign n16538 = n14664 & n14671;
  assign n16539 = ~n16537 & ~n16538;
  assign n16540 = n14685 & ~n14692;
  assign n16541 = n14656 & ~n16540;
  assign n16542 = n14664 & ~n14697;
  assign n16543 = ~n16541 & ~n16542;
  assign n16544 = ~n14660 & n15949;
  assign n16545 = n14651 & ~n16544;
  assign n16546 = n14693 & n16529;
  assign n16547 = n14661 & ~n16546;
  assign n16548 = ~n16545 & ~n16547;
  assign n16549 = n16543 & n16548;
  assign n16550 = n16539 & n16549;
  assign n16551 = ~n16536 & n16550;
  assign n16552 = ~n16534 & n16551;
  assign n16553 = n16533 & n16552;
  assign n16554 = n15947 & n16553;
  assign n16555 = n14667 & n16554;
  assign n16556 = n16555 ^ n14383;
  assign n16557 = n16556 ^ x690;
  assign n16558 = n16528 & n16557;
  assign n16559 = n15605 & n15653;
  assign n16560 = n15650 & ~n16112;
  assign n16561 = ~n16559 & ~n16560;
  assign n16562 = n15626 & n15629;
  assign n16563 = n15545 & n15635;
  assign n16564 = ~n16562 & ~n16563;
  assign n16565 = ~n15610 & ~n15630;
  assign n16566 = n15614 & ~n16565;
  assign n16567 = ~n15619 & n15648;
  assign n16568 = ~n15617 & n16567;
  assign n16569 = ~n15635 & n16568;
  assign n16570 = n15547 & ~n16569;
  assign n16571 = n15606 ^ n15602;
  assign n16572 = ~n15573 & n16571;
  assign n16573 = n15572 & n16572;
  assign n16574 = n16573 ^ n15606;
  assign n16575 = n15650 & n16574;
  assign n16576 = ~n15633 & n16105;
  assign n16577 = n15614 & ~n16576;
  assign n16578 = n15601 ^ n15572;
  assign n16579 = n15575 & n16578;
  assign n16580 = n15605 & n16579;
  assign n16581 = ~n16577 & ~n16580;
  assign n16582 = ~n16575 & n16581;
  assign n16583 = ~n16570 & n16582;
  assign n16584 = ~n16566 & n16583;
  assign n16585 = n16564 & n16584;
  assign n16586 = n16561 & n16585;
  assign n16587 = n15613 & n16586;
  assign n16588 = n16587 ^ n14412;
  assign n16589 = n16588 ^ x692;
  assign n16590 = n15107 & ~n15127;
  assign n16591 = n15106 & ~n16590;
  assign n16592 = n15100 & n15107;
  assign n16593 = ~n15010 & n15129;
  assign n16594 = ~n15132 & n16593;
  assign n16595 = n15089 & ~n16594;
  assign n16596 = ~n15097 & ~n15107;
  assign n16597 = n15121 & ~n16596;
  assign n16598 = n15134 & ~n16407;
  assign n16599 = n15107 & ~n16598;
  assign n16600 = ~n15112 & ~n15135;
  assign n16601 = ~n15103 & n16600;
  assign n16602 = ~n15109 & n16601;
  assign n16603 = n15089 & ~n16602;
  assign n16604 = ~n15096 & ~n15121;
  assign n16605 = ~n15091 & n16604;
  assign n16606 = n15087 & ~n16605;
  assign n16607 = ~n16603 & ~n16606;
  assign n16608 = ~n16599 & n16607;
  assign n16609 = ~n16597 & n16608;
  assign n16610 = n15087 & ~n16419;
  assign n16611 = n14873 & n16401;
  assign n16612 = n15129 & ~n16611;
  assign n16613 = ~n15126 & n16612;
  assign n16614 = ~n15112 & n16613;
  assign n16615 = n15097 & ~n16614;
  assign n16616 = ~n16610 & ~n16615;
  assign n16617 = n16609 & n16616;
  assign n16618 = ~n16595 & n16617;
  assign n16619 = ~n16592 & n16618;
  assign n16620 = n15119 & n16619;
  assign n16621 = n16591 & n16620;
  assign n16622 = n16621 ^ n14444;
  assign n16623 = n16622 ^ x691;
  assign n16624 = ~n16589 & n16623;
  assign n16625 = n16558 & n16624;
  assign n16626 = n15996 ^ x688;
  assign n16627 = n16321 & n16324;
  assign n16628 = ~n16318 & ~n16323;
  assign n16629 = n16299 & ~n16628;
  assign n16630 = ~n16627 & ~n16629;
  assign n16631 = n16243 & n16349;
  assign n16632 = n16301 & ~n16325;
  assign n16633 = ~n16631 & ~n16632;
  assign n16634 = ~n16301 & ~n16346;
  assign n16635 = ~n16341 & n16634;
  assign n16636 = n16244 & ~n16635;
  assign n16637 = ~n16297 & n16299;
  assign n16638 = n16244 & n16331;
  assign n16639 = ~n16316 & ~n16638;
  assign n16640 = ~n16305 & ~n16335;
  assign n16641 = n16310 & ~n16640;
  assign n16642 = n16306 & n16342;
  assign n16643 = n16299 & ~n16642;
  assign n16644 = ~n16641 & ~n16643;
  assign n16645 = ~n16294 & ~n16330;
  assign n16646 = ~n16318 & n16645;
  assign n16647 = n16244 & ~n16646;
  assign n16648 = ~n16324 & n16645;
  assign n16649 = n16315 & ~n16318;
  assign n16650 = ~n16330 & n16649;
  assign n16651 = ~n16310 & n16650;
  assign n16652 = ~n16648 & ~n16651;
  assign n16653 = ~n16325 & n16652;
  assign n16654 = ~n16647 & ~n16653;
  assign n16655 = n16644 & n16654;
  assign n16656 = n16639 & n16655;
  assign n16657 = ~n16637 & n16656;
  assign n16658 = ~n16636 & n16657;
  assign n16659 = n16633 & n16658;
  assign n16660 = n16630 & n16659;
  assign n16661 = n16337 & n16660;
  assign n16662 = n16661 ^ n14356;
  assign n16663 = n16662 ^ x693;
  assign n16664 = n16626 & ~n16663;
  assign n16665 = n16625 & n16664;
  assign n16666 = ~n16626 & n16663;
  assign n16667 = n16625 & n16666;
  assign n16668 = n16626 & n16663;
  assign n16669 = ~n16528 & n16557;
  assign n16670 = ~n16589 & ~n16623;
  assign n16671 = n16669 & n16670;
  assign n16672 = n16668 & n16671;
  assign n16673 = ~n16667 & ~n16672;
  assign n16674 = n16589 & n16623;
  assign n16675 = n16669 & n16674;
  assign n16676 = ~n16528 & ~n16557;
  assign n16677 = n16670 & n16676;
  assign n16678 = ~n16675 & ~n16677;
  assign n16679 = n16668 & ~n16678;
  assign n16680 = n16673 & ~n16679;
  assign n16681 = n16558 & n16670;
  assign n16682 = n16528 & ~n16557;
  assign n16683 = n16589 & ~n16623;
  assign n16684 = n16682 & n16683;
  assign n16685 = ~n16681 & ~n16684;
  assign n16686 = n16666 & ~n16685;
  assign n16687 = n16558 & n16683;
  assign n16688 = n16664 & n16687;
  assign n16689 = ~n16626 & ~n16663;
  assign n16690 = n16676 & n16683;
  assign n16691 = n16689 & n16690;
  assign n16692 = ~n16688 & ~n16691;
  assign n16693 = n16624 & n16669;
  assign n16694 = n16689 & n16693;
  assign n16695 = n16668 & n16690;
  assign n16696 = ~n16694 & ~n16695;
  assign n16697 = n16624 & n16682;
  assign n16698 = n16689 & n16697;
  assign n16699 = n16624 & n16676;
  assign n16700 = ~n16675 & ~n16699;
  assign n16701 = n16669 & n16683;
  assign n16702 = ~n16697 & ~n16701;
  assign n16703 = n16700 & n16702;
  assign n16704 = ~n16687 & n16703;
  assign n16705 = n16666 & ~n16704;
  assign n16706 = n16674 & n16676;
  assign n16707 = n16558 & n16674;
  assign n16708 = n16670 & n16682;
  assign n16709 = ~n16707 & ~n16708;
  assign n16710 = ~n16706 & n16709;
  assign n16711 = ~n16690 & n16710;
  assign n16712 = n16664 & ~n16711;
  assign n16713 = n16674 & n16682;
  assign n16714 = ~n16681 & ~n16713;
  assign n16715 = ~n16707 & n16714;
  assign n16716 = n16689 & ~n16715;
  assign n16717 = ~n16671 & ~n16701;
  assign n16718 = ~n16663 & ~n16717;
  assign n16719 = n16709 & ~n16713;
  assign n16720 = ~n16625 & n16719;
  assign n16721 = n16668 & ~n16720;
  assign n16722 = ~n16718 & ~n16721;
  assign n16723 = ~n16716 & n16722;
  assign n16724 = ~n16712 & n16723;
  assign n16725 = ~n16705 & n16724;
  assign n16726 = ~n16698 & n16725;
  assign n16727 = n16696 & n16726;
  assign n16728 = n16692 & n16727;
  assign n16729 = ~n16686 & n16728;
  assign n16730 = n16680 & n16729;
  assign n16731 = ~n16665 & n16730;
  assign n16732 = n16731 ^ n15007;
  assign n16733 = n16732 ^ x761;
  assign n16734 = n16527 & ~n16733;
  assign n16735 = n15153 ^ x698;
  assign n16736 = n16662 ^ x695;
  assign n16737 = n16735 & ~n16736;
  assign n16738 = n15513 & n15518;
  assign n16739 = n15489 & n15504;
  assign n16740 = ~n15502 & ~n16739;
  assign n16741 = n15500 & ~n16740;
  assign n16742 = ~n16738 & ~n16741;
  assign n16743 = n15487 & n15513;
  assign n16744 = ~n15498 & ~n15515;
  assign n16745 = n15532 & ~n16744;
  assign n16746 = ~n16743 & ~n16745;
  assign n16747 = n15506 & ~n15514;
  assign n16748 = ~n15976 & n16747;
  assign n16749 = n15399 & ~n16748;
  assign n16750 = ~n15460 & n15489;
  assign n16751 = n15513 & n16750;
  assign n16752 = ~n15490 & ~n15498;
  assign n16753 = n15500 & ~n16752;
  assign n16754 = ~n15502 & ~n15505;
  assign n16755 = n15513 & ~n16754;
  assign n16756 = ~n16753 & ~n16755;
  assign n16757 = n15371 & n15518;
  assign n16758 = ~n15503 & ~n15517;
  assign n16759 = ~n16739 & n16758;
  assign n16760 = n15973 & n16759;
  assign n16761 = n15532 & ~n16760;
  assign n16762 = ~n16757 & ~n16761;
  assign n16763 = n16756 & n16762;
  assign n16764 = ~n16751 & n16763;
  assign n16765 = ~n16749 & n16764;
  assign n16766 = n16746 & n16765;
  assign n16767 = ~n15512 & n16766;
  assign n16768 = n15981 & n16767;
  assign n16769 = n16742 & n16768;
  assign n16770 = n15496 & n16769;
  assign n16771 = n16770 ^ n14748;
  assign n16772 = n16771 ^ x697;
  assign n16773 = ~n16077 & ~n16082;
  assign n16774 = n16052 & ~n16773;
  assign n16775 = n16067 & n16076;
  assign n16776 = n16057 & ~n16074;
  assign n16777 = ~n16775 & ~n16776;
  assign n16778 = ~n16774 & n16777;
  assign n16779 = n16057 & ~n16088;
  assign n16780 = n16019 & n16038;
  assign n16781 = n16381 & ~n16780;
  assign n16782 = n16052 & ~n16781;
  assign n16783 = n16054 & ~n16085;
  assign n16784 = ~n16045 & n16783;
  assign n16785 = ~n16365 & n16367;
  assign n16786 = ~n16049 & n16785;
  assign n16787 = ~n16784 & ~n16786;
  assign n16788 = n16074 & ~n16787;
  assign n16789 = n16067 & ~n16788;
  assign n16790 = ~n16782 & ~n16789;
  assign n16791 = ~n16779 & n16790;
  assign n16792 = n16072 & n16791;
  assign n16793 = n16051 & n16792;
  assign n16794 = n16778 & n16793;
  assign n16795 = n16794 ^ n14770;
  assign n16796 = n16795 ^ x696;
  assign n16797 = ~n16772 & n16796;
  assign n16798 = n16737 & n16797;
  assign n16799 = n16588 ^ x694;
  assign n16800 = n15847 ^ x699;
  assign n16801 = ~n16799 & n16800;
  assign n16802 = n16798 & n16801;
  assign n16803 = n16799 & ~n16800;
  assign n16804 = n16772 & n16796;
  assign n16805 = n16737 & n16804;
  assign n16806 = ~n16735 & ~n16736;
  assign n16807 = n16772 & ~n16796;
  assign n16808 = n16806 & n16807;
  assign n16809 = ~n16805 & ~n16808;
  assign n16810 = n16803 & ~n16809;
  assign n16811 = ~n16802 & ~n16810;
  assign n16812 = ~n16799 & ~n16800;
  assign n16813 = n16798 & n16812;
  assign n16814 = n16735 & n16736;
  assign n16815 = n16807 & n16814;
  assign n16816 = n16799 & n16800;
  assign n16817 = n16815 & n16816;
  assign n16818 = ~n16735 & n16736;
  assign n16819 = n16804 & n16818;
  assign n16820 = n16801 & n16819;
  assign n16821 = ~n16817 & ~n16820;
  assign n16822 = ~n16813 & n16821;
  assign n16823 = ~n16772 & ~n16796;
  assign n16824 = n16737 & n16823;
  assign n16825 = n16816 & n16824;
  assign n16826 = n16801 & n16815;
  assign n16827 = n16797 & n16814;
  assign n16828 = n16807 & n16818;
  assign n16829 = ~n16827 & ~n16828;
  assign n16830 = n16812 & ~n16829;
  assign n16831 = ~n16826 & ~n16830;
  assign n16832 = ~n16825 & n16831;
  assign n16833 = n16812 & n16815;
  assign n16834 = n16804 & n16814;
  assign n16835 = n16801 & n16834;
  assign n16836 = n16803 & n16827;
  assign n16837 = ~n16835 & ~n16836;
  assign n16838 = ~n16833 & n16837;
  assign n16839 = n16737 & n16807;
  assign n16840 = n16797 & n16818;
  assign n16841 = n16814 & n16823;
  assign n16842 = ~n16840 & ~n16841;
  assign n16843 = ~n16839 & n16842;
  assign n16844 = n16803 & ~n16843;
  assign n16845 = n16806 & n16823;
  assign n16846 = ~n16824 & ~n16845;
  assign n16847 = ~n16840 & n16846;
  assign n16848 = ~n16808 & n16847;
  assign n16849 = n16801 & ~n16848;
  assign n16850 = ~n16844 & ~n16849;
  assign n16851 = n16736 ^ n16735;
  assign n16852 = n16851 ^ n16796;
  assign n16853 = ~n16772 & ~n16852;
  assign n16854 = n16816 & n16853;
  assign n16855 = n16804 & n16806;
  assign n16856 = ~n16819 & ~n16855;
  assign n16857 = n16799 & ~n16856;
  assign n16858 = n16818 & n16823;
  assign n16859 = n16797 & n16806;
  assign n16860 = ~n16839 & ~n16859;
  assign n16861 = ~n16845 & n16860;
  assign n16862 = ~n16858 & n16861;
  assign n16863 = n16812 & ~n16862;
  assign n16864 = ~n16857 & ~n16863;
  assign n16865 = ~n16854 & n16864;
  assign n16866 = n16850 & n16865;
  assign n16867 = n16838 & n16866;
  assign n16868 = n16832 & n16867;
  assign n16869 = n16822 & n16868;
  assign n16870 = n16811 & n16869;
  assign n16871 = n16870 ^ n14836;
  assign n16872 = n16871 ^ x762;
  assign n16873 = n15299 & ~n15318;
  assign n16874 = ~n15258 & ~n16873;
  assign n16875 = n15297 ^ n15231;
  assign n16876 = ~n15252 & n16875;
  assign n16877 = n16876 ^ n15231;
  assign n16878 = n15253 & n16877;
  assign n16879 = n15252 & n15256;
  assign n16880 = ~n15314 & ~n16879;
  assign n16881 = ~n16878 & n16880;
  assign n16882 = n16874 & n16881;
  assign n16883 = n15324 & n16882;
  assign n16884 = n16877 ^ n15256;
  assign n16885 = ~n15253 & n16884;
  assign n16886 = n16885 ^ n15256;
  assign n16887 = n16874 & ~n16886;
  assign n16888 = ~n15298 & n16887;
  assign n16889 = n15331 & ~n16888;
  assign n16890 = ~n16883 & ~n16889;
  assign n16891 = ~n16878 & ~n16879;
  assign n16892 = ~n15306 & n16891;
  assign n16893 = n15315 & n16892;
  assign n16894 = n15296 & ~n16893;
  assign n16895 = n15299 ^ n15195;
  assign n16896 = ~n15312 & ~n16895;
  assign n16897 = n16896 ^ n15195;
  assign n16898 = n16880 & n16897;
  assign n16899 = ~n15258 & n16898;
  assign n16900 = n15311 & ~n16899;
  assign n16901 = ~n16894 & ~n16900;
  assign n16902 = n16890 & n16901;
  assign n16903 = n16902 ^ n13663;
  assign n16904 = n16903 ^ x718;
  assign n16905 = n15135 & ~n16596;
  assign n16906 = ~n15134 & ~n16411;
  assign n16907 = ~n16905 & ~n16906;
  assign n16908 = n15112 & ~n16402;
  assign n16909 = n15127 & ~n15142;
  assign n16910 = n15097 & ~n16909;
  assign n16911 = ~n15086 & ~n16604;
  assign n16912 = ~n16910 & ~n16911;
  assign n16913 = ~n16908 & n16912;
  assign n16914 = n16907 & n16913;
  assign n16915 = n15116 & n16914;
  assign n16916 = n16405 & n16915;
  assign n16917 = n16591 & n16916;
  assign n16918 = n15094 & n16917;
  assign n16919 = n16918 ^ n12653;
  assign n16920 = n16919 ^ x723;
  assign n16921 = ~n16904 & ~n16920;
  assign n16922 = ~n16312 & ~n16335;
  assign n16923 = n16299 & ~n16922;
  assign n16924 = n16324 & ~n16628;
  assign n16925 = ~n16923 & ~n16924;
  assign n16926 = ~n16325 & n16331;
  assign n16927 = n16306 & ~n16323;
  assign n16928 = ~n16341 & n16927;
  assign n16929 = ~n16346 & n16928;
  assign n16930 = n16244 & ~n16929;
  assign n16931 = ~n16926 & ~n16930;
  assign n16932 = n16310 & n16330;
  assign n16933 = ~n16312 & ~n16321;
  assign n16934 = n16324 & ~n16933;
  assign n16935 = ~n16346 & n16645;
  assign n16936 = n16299 & ~n16935;
  assign n16937 = ~n16296 & ~n16341;
  assign n16938 = ~n16310 & n16937;
  assign n16939 = ~n16301 & n16348;
  assign n16940 = ~n16938 & ~n16939;
  assign n16941 = ~n16349 & ~n16940;
  assign n16942 = ~n16325 & ~n16941;
  assign n16943 = ~n16936 & ~n16942;
  assign n16944 = ~n16934 & n16943;
  assign n16945 = ~n16932 & n16944;
  assign n16946 = n16931 & n16945;
  assign n16947 = n16925 & n16946;
  assign n16948 = n16309 & n16947;
  assign n16949 = n16639 & n16948;
  assign n16950 = n16949 ^ n13592;
  assign n16951 = n16950 ^ x719;
  assign n16952 = n16057 & ~n16061;
  assign n16953 = ~n16065 & ~n16780;
  assign n16954 = n16067 & ~n16953;
  assign n16955 = n16052 & ~n16086;
  assign n16956 = ~n16049 & n16387;
  assign n16957 = n16057 & ~n16956;
  assign n16958 = ~n16955 & ~n16957;
  assign n16959 = n16070 & n16078;
  assign n16960 = n16045 & ~n16959;
  assign n16961 = ~n16053 & n16773;
  assign n16962 = n16036 & ~n16961;
  assign n16963 = ~n16960 & ~n16962;
  assign n16964 = n16958 & n16963;
  assign n16965 = ~n16954 & n16964;
  assign n16966 = ~n16952 & n16965;
  assign n16967 = ~n16040 & n16966;
  assign n16968 = n16063 & n16967;
  assign n16969 = n16056 & n16968;
  assign n16970 = n16778 & n16969;
  assign n16971 = n16970 ^ n13275;
  assign n16972 = n16971 ^ x722;
  assign n16973 = n15500 & n15525;
  assign n16974 = n15534 & n16758;
  assign n16975 = ~n15511 & n16974;
  assign n16976 = n15513 & ~n16975;
  assign n16977 = ~n16973 & ~n16976;
  assign n16978 = ~n15511 & ~n16750;
  assign n16979 = n16740 & n16978;
  assign n16980 = ~n15505 & n16979;
  assign n16981 = n15532 & ~n16980;
  assign n16982 = ~n15500 & n16978;
  assign n16983 = n15520 & ~n15976;
  assign n16984 = ~n15399 & n16983;
  assign n16985 = ~n16982 & ~n16984;
  assign n16986 = ~n15505 & ~n16985;
  assign n16987 = ~n15517 & n16986;
  assign n16988 = n15371 & ~n16987;
  assign n16989 = ~n16981 & ~n16988;
  assign n16990 = n16977 & n16989;
  assign n16991 = n16746 & n16990;
  assign n16992 = ~n15975 & n16991;
  assign n16993 = n16742 & n16992;
  assign n16994 = n16993 ^ n14579;
  assign n16995 = n16994 ^ x720;
  assign n16996 = ~n16972 & n16995;
  assign n16997 = n16951 & n16996;
  assign n16998 = n15803 & ~n15816;
  assign n16999 = n15789 & ~n15837;
  assign n17000 = n15806 & n15812;
  assign n17001 = n15819 & n16149;
  assign n17002 = ~n15764 & n17001;
  assign n17003 = n15802 & ~n17002;
  assign n17004 = ~n17000 & ~n17003;
  assign n17005 = ~n15818 & ~n15833;
  assign n17006 = n15785 & ~n17005;
  assign n17007 = ~n15795 & ~n15817;
  assign n17008 = ~n15807 & n17007;
  assign n17009 = n15789 & ~n17008;
  assign n17010 = ~n17006 & ~n17009;
  assign n17011 = ~n15800 & n16154;
  assign n17012 = ~n15785 & n17011;
  assign n17013 = ~n15821 & n15830;
  assign n17014 = ~n15807 & n17013;
  assign n17015 = ~n15812 & n17014;
  assign n17016 = ~n17012 & ~n17015;
  assign n17017 = ~n15816 & n17016;
  assign n17018 = n17010 & ~n17017;
  assign n17019 = n17004 & n17018;
  assign n17020 = ~n15811 & n17019;
  assign n17021 = ~n16999 & n17020;
  assign n17022 = ~n16998 & n17021;
  assign n17023 = n16136 & n17022;
  assign n17024 = n15805 & n17023;
  assign n17025 = n17024 ^ n14542;
  assign n17026 = n17025 ^ x721;
  assign n17027 = n16997 & n17026;
  assign n17028 = ~n16995 & n17026;
  assign n17029 = n16972 & n17028;
  assign n17030 = n16951 & n17029;
  assign n17031 = ~n17027 & ~n17030;
  assign n17032 = n16921 & ~n17031;
  assign n17033 = n16972 & n16995;
  assign n17034 = ~n16951 & n17033;
  assign n17035 = ~n17026 & n17034;
  assign n17036 = n16921 & n17035;
  assign n17037 = n16904 & ~n16920;
  assign n17038 = ~n16951 & n17029;
  assign n17039 = n17037 & n17038;
  assign n17040 = ~n16904 & n16920;
  assign n17041 = ~n16972 & n17028;
  assign n17042 = n16951 & n17041;
  assign n17043 = n16972 & ~n16995;
  assign n17044 = n16951 & ~n17026;
  assign n17045 = n17043 & n17044;
  assign n17046 = ~n17042 & ~n17045;
  assign n17047 = n17040 & ~n17046;
  assign n17048 = ~n17039 & ~n17047;
  assign n17049 = ~n16951 & ~n16972;
  assign n17050 = ~n16995 & n17049;
  assign n17051 = ~n17026 & n17050;
  assign n17052 = ~n17035 & ~n17051;
  assign n17053 = n17040 & ~n17052;
  assign n17054 = n16904 & n16920;
  assign n17055 = n16951 & n17033;
  assign n17056 = n17026 & n17055;
  assign n17057 = n16996 & n17044;
  assign n17058 = ~n17056 & ~n17057;
  assign n17059 = n17054 & ~n17058;
  assign n17060 = ~n17053 & ~n17059;
  assign n17061 = n17048 & n17060;
  assign n17062 = n17027 & n17054;
  assign n17063 = n16921 & ~n17046;
  assign n17064 = ~n17062 & ~n17063;
  assign n17065 = n17028 & n17049;
  assign n17066 = n17033 & n17044;
  assign n17067 = ~n17065 & ~n17066;
  assign n17068 = n17040 & ~n17067;
  assign n17069 = n17051 & n17054;
  assign n17070 = n16995 & n17049;
  assign n17071 = ~n17026 & n17070;
  assign n17072 = n17037 & n17071;
  assign n17073 = ~n17069 & ~n17072;
  assign n17074 = n17026 & n17070;
  assign n17075 = n17037 & n17074;
  assign n17076 = ~n16951 & n17043;
  assign n17077 = ~n17026 & n17076;
  assign n17078 = ~n17065 & ~n17077;
  assign n17079 = ~n17035 & n17078;
  assign n17080 = ~n17030 & n17079;
  assign n17081 = n17054 & ~n17080;
  assign n17082 = ~n17075 & ~n17081;
  assign n17083 = n17026 & n17034;
  assign n17084 = ~n16920 & n17083;
  assign n17085 = ~n17027 & ~n17038;
  assign n17086 = n17040 & ~n17085;
  assign n17087 = ~n17051 & ~n17066;
  assign n17088 = n16921 & ~n17087;
  assign n17089 = ~n16995 & n17044;
  assign n17090 = ~n16972 & n17089;
  assign n17091 = n17046 & ~n17057;
  assign n17092 = ~n17090 & n17091;
  assign n17093 = n17037 & ~n17092;
  assign n17094 = ~n17088 & ~n17093;
  assign n17095 = ~n17086 & n17094;
  assign n17096 = ~n17084 & n17095;
  assign n17097 = n17082 & n17096;
  assign n17098 = n17073 & n17097;
  assign n17099 = ~n17068 & n17098;
  assign n17100 = n17064 & n17099;
  assign n17101 = n17061 & n17100;
  assign n17102 = ~n17036 & n17101;
  assign n17103 = ~n17032 & n17102;
  assign n17104 = n17103 ^ n14872;
  assign n17105 = n17104 ^ x763;
  assign n17106 = n16872 & ~n17105;
  assign n17107 = n16734 & n17106;
  assign n17108 = n16241 & n17107;
  assign n17109 = ~n15930 & ~n16240;
  assign n17110 = ~n16872 & ~n17105;
  assign n17111 = n16733 & n17110;
  assign n17112 = n16527 & n17111;
  assign n17113 = n17109 & n17112;
  assign n17114 = ~n17108 & ~n17113;
  assign n17115 = n16527 & n16733;
  assign n17116 = ~n16872 & n17105;
  assign n17117 = n17115 & n17116;
  assign n17118 = n17109 & n17117;
  assign n17119 = n16734 & n17116;
  assign n17120 = n16241 & n17119;
  assign n17121 = n17106 & n17115;
  assign n17122 = n15930 & ~n16240;
  assign n17123 = n17121 & n17122;
  assign n17124 = ~n17120 & ~n17123;
  assign n17125 = ~n17118 & n17124;
  assign n17126 = ~n16527 & n16733;
  assign n17127 = n17106 & n17126;
  assign n17128 = ~n16240 & n17127;
  assign n17129 = n16872 & n17105;
  assign n17130 = n17115 & n17129;
  assign n17131 = ~n15930 & n16240;
  assign n17132 = ~n17122 & ~n17131;
  assign n17133 = n17130 & ~n17132;
  assign n17134 = ~n17128 & ~n17133;
  assign n17135 = n17116 & n17126;
  assign n17136 = ~n15930 & n17135;
  assign n17137 = ~n16527 & ~n16733;
  assign n17138 = n17106 & n17137;
  assign n17139 = n17131 & n17138;
  assign n17140 = ~n17136 & ~n17139;
  assign n17141 = n17116 & n17137;
  assign n17142 = n17110 & n17137;
  assign n17143 = ~n17141 & ~n17142;
  assign n17144 = n16241 & ~n17143;
  assign n17145 = n17129 & n17137;
  assign n17146 = n16734 & n17110;
  assign n17147 = ~n17119 & ~n17141;
  assign n17148 = ~n17146 & n17147;
  assign n17149 = ~n17145 & n17148;
  assign n17150 = ~n17122 & n17149;
  assign n17151 = ~n17107 & ~n17141;
  assign n17152 = ~n17145 & n17151;
  assign n17153 = ~n17117 & n17152;
  assign n17154 = ~n17131 & n17153;
  assign n17155 = ~n17150 & ~n17154;
  assign n17156 = ~n17132 & n17155;
  assign n17157 = n17126 & n17129;
  assign n17158 = ~n17121 & ~n17157;
  assign n17159 = ~n17111 & n17158;
  assign n17160 = n16241 & ~n17159;
  assign n17161 = n16734 & n17129;
  assign n17162 = ~n17142 & ~n17161;
  assign n17163 = ~n17138 & n17162;
  assign n17164 = ~n17145 & n17163;
  assign n17165 = n17109 & ~n17164;
  assign n17166 = ~n17160 & ~n17165;
  assign n17167 = ~n17156 & n17166;
  assign n17168 = ~n17144 & n17167;
  assign n17169 = n17140 & n17168;
  assign n17170 = n17134 & n17169;
  assign n17171 = ~n16527 & n17111;
  assign n17172 = n16240 ^ n15930;
  assign n17173 = n17171 & n17172;
  assign n17174 = n17170 & ~n17173;
  assign n17175 = n17125 & n17174;
  assign n17176 = n17114 & n17175;
  assign n17177 = n17176 ^ n15153;
  assign n17178 = ~n16399 & n16500;
  assign n17179 = n16516 & ~n17178;
  assign n17180 = n16508 & ~n17179;
  assign n17181 = ~n16438 & n16510;
  assign n17182 = n16364 & n17178;
  assign n17183 = ~n17181 & ~n17182;
  assign n17184 = ~n16501 & n17183;
  assign n17185 = n16506 & n17184;
  assign n17186 = ~n17180 & ~n17185;
  assign n17187 = ~n16437 & ~n16445;
  assign n17188 = ~n16440 & n16441;
  assign n17189 = ~n17187 & ~n17188;
  assign n17190 = n16440 & ~n16491;
  assign n17191 = n17189 & ~n17190;
  assign n17192 = n16481 & n17191;
  assign n17193 = n16519 ^ n16445;
  assign n17194 = ~n16440 & ~n17193;
  assign n17195 = n17194 ^ n16445;
  assign n17196 = n16483 & n17195;
  assign n17197 = ~n17192 & ~n17196;
  assign n17198 = n17186 & n17197;
  assign n17199 = n17198 ^ n16029;
  assign n17200 = n17199 ^ x750;
  assign n17201 = n16664 & n16684;
  assign n17202 = n16666 & n16701;
  assign n17203 = ~n17201 & ~n17202;
  assign n17204 = ~n16698 & n17203;
  assign n17205 = ~n16690 & ~n16699;
  assign n17206 = n16666 & ~n17205;
  assign n17207 = n16692 & ~n17206;
  assign n17208 = n16666 & n16707;
  assign n17209 = n16687 & n16689;
  assign n17210 = ~n17208 & ~n17209;
  assign n17211 = ~n16663 & n16706;
  assign n17212 = ~n16671 & n16700;
  assign n17213 = n16664 & ~n17212;
  assign n17214 = ~n16625 & ~n16708;
  assign n17215 = n16689 & ~n17214;
  assign n17216 = ~n17213 & ~n17215;
  assign n17217 = ~n17211 & n17216;
  assign n17218 = n16678 & ~n16713;
  assign n17219 = n16666 & ~n17218;
  assign n17220 = ~n16693 & n16709;
  assign n17221 = n16702 & n17220;
  assign n17222 = ~n16671 & n17221;
  assign n17223 = n16668 & ~n17222;
  assign n17224 = ~n17219 & ~n17223;
  assign n17225 = n17217 & n17224;
  assign n17226 = n16696 & n17225;
  assign n17227 = n17210 & n17226;
  assign n17228 = n17207 & n17227;
  assign n17229 = n17204 & n17228;
  assign n17230 = ~n16665 & n17229;
  assign n17231 = ~n16681 & n17230;
  assign n17232 = n17231 ^ n14516;
  assign n17233 = n17232 ^ x749;
  assign n17234 = n17200 & ~n17233;
  assign n17235 = n16971 ^ x724;
  assign n17236 = n16132 ^ x729;
  assign n17237 = ~n17235 & n17236;
  assign n17238 = n15970 ^ x728;
  assign n17239 = n16919 ^ x725;
  assign n17240 = ~n17238 & n17239;
  assign n17241 = n15324 & ~n16888;
  assign n17242 = n15331 & ~n16882;
  assign n17243 = ~n17241 & ~n17242;
  assign n17244 = n15296 & n16899;
  assign n17245 = n15311 & ~n16893;
  assign n17246 = ~n17244 & ~n17245;
  assign n17247 = n17243 & n17246;
  assign n17248 = n17247 ^ n12274;
  assign n17249 = n17248 ^ x726;
  assign n17250 = ~n16305 & ~n16349;
  assign n17251 = ~n16330 & n17250;
  assign n17252 = ~n16321 & n17251;
  assign n17253 = n16299 & ~n17252;
  assign n17254 = ~n16294 & ~n16331;
  assign n17255 = n16310 & ~n17254;
  assign n17256 = ~n16296 & ~n16314;
  assign n17257 = ~n16325 & ~n17256;
  assign n17258 = n16315 & n16645;
  assign n17259 = n16244 & ~n17258;
  assign n17260 = ~n17257 & ~n17259;
  assign n17261 = n16310 & ~n16635;
  assign n17262 = n16244 & ~n16634;
  assign n17263 = n16306 & ~n17262;
  assign n17264 = n16243 & ~n17263;
  assign n17265 = ~n17261 & ~n17264;
  assign n17266 = n17260 & n17265;
  assign n17267 = ~n17255 & n17266;
  assign n17268 = ~n17253 & n17267;
  assign n17269 = n16630 & n17268;
  assign n17270 = n16925 & n17269;
  assign n17271 = n16337 & n17270;
  assign n17272 = n17271 ^ n13161;
  assign n17273 = n17272 ^ x727;
  assign n17274 = ~n17249 & ~n17273;
  assign n17275 = n17240 & n17274;
  assign n17276 = n17238 & n17239;
  assign n17277 = n17249 & ~n17273;
  assign n17278 = n17276 & n17277;
  assign n17279 = ~n17275 & ~n17278;
  assign n17280 = n17237 & ~n17279;
  assign n17281 = ~n17238 & ~n17239;
  assign n17282 = ~n17249 & n17273;
  assign n17283 = n17281 & n17282;
  assign n17284 = n17237 & n17283;
  assign n17285 = n17240 & n17277;
  assign n17286 = n17235 & n17236;
  assign n17287 = n17285 & n17286;
  assign n17288 = ~n17284 & ~n17287;
  assign n17289 = n17235 & ~n17236;
  assign n17290 = n17238 & ~n17239;
  assign n17291 = n17282 & n17290;
  assign n17292 = n17249 & n17273;
  assign n17293 = n17240 & n17292;
  assign n17294 = n17274 & n17276;
  assign n17295 = ~n17293 & ~n17294;
  assign n17296 = ~n17278 & n17295;
  assign n17297 = n17277 & n17290;
  assign n17298 = ~n17283 & ~n17297;
  assign n17299 = n17290 & n17292;
  assign n17300 = n17274 & n17281;
  assign n17301 = ~n17299 & ~n17300;
  assign n17302 = n17298 & n17301;
  assign n17303 = n17296 & n17302;
  assign n17304 = ~n17291 & n17303;
  assign n17305 = n17289 & n17304;
  assign n17306 = n17240 & n17282;
  assign n17307 = ~n17291 & ~n17306;
  assign n17308 = n17281 & n17292;
  assign n17309 = n17274 & n17290;
  assign n17310 = ~n17308 & ~n17309;
  assign n17311 = n17307 & n17310;
  assign n17312 = ~n17297 & n17311;
  assign n17313 = n17237 & ~n17312;
  assign n17314 = ~n17305 & ~n17313;
  assign n17315 = n17295 & n17302;
  assign n17316 = ~n17306 & n17315;
  assign n17317 = n17286 & ~n17316;
  assign n17318 = ~n17235 & ~n17236;
  assign n17319 = n17249 ^ n17238;
  assign n17320 = n17319 ^ n17238;
  assign n17321 = n17320 ^ n17273;
  assign n17322 = ~n17239 & n17321;
  assign n17323 = n17322 ^ n17319;
  assign n17324 = n17318 & n17323;
  assign n17325 = ~n17317 & ~n17324;
  assign n17326 = n17314 & n17325;
  assign n17327 = n17288 & n17326;
  assign n17328 = ~n17280 & n17327;
  assign n17329 = n17328 ^ n15294;
  assign n17330 = n17329 ^ x752;
  assign n17331 = ~n17035 & ~n17074;
  assign n17332 = n17054 & ~n17331;
  assign n17333 = ~n17071 & ~n17083;
  assign n17334 = n17040 & ~n17333;
  assign n17335 = ~n17332 & ~n17334;
  assign n17336 = ~n16920 & n17074;
  assign n17337 = ~n17066 & ~n17090;
  assign n17338 = ~n17065 & n17337;
  assign n17339 = ~n17038 & n17338;
  assign n17340 = n17054 & ~n17339;
  assign n17341 = ~n17336 & ~n17340;
  assign n17342 = ~n16921 & ~n17054;
  assign n17343 = ~n17058 & n17342;
  assign n17344 = ~n17042 & n17052;
  assign n17345 = ~n17030 & n17344;
  assign n17346 = n17037 & ~n17345;
  assign n17347 = ~n17045 & ~n17090;
  assign n17348 = n17078 & n17347;
  assign n17349 = ~n17083 & n17348;
  assign n17350 = n16921 & ~n17349;
  assign n17351 = ~n17346 & ~n17350;
  assign n17352 = ~n17343 & n17351;
  assign n17353 = n17341 & n17352;
  assign n17354 = n17061 & n17353;
  assign n17355 = n17335 & n17354;
  assign n17356 = ~n17032 & n17355;
  assign n17357 = n17356 ^ n16017;
  assign n17358 = n17357 ^ x751;
  assign n17359 = n17330 & ~n17358;
  assign n17360 = n17234 & n17359;
  assign n17361 = n16801 & ~n16809;
  assign n17362 = n16803 & n16828;
  assign n17363 = ~n16824 & ~n16855;
  assign n17364 = n16812 & ~n17363;
  assign n17365 = ~n17362 & ~n17364;
  assign n17366 = ~n17361 & n17365;
  assign n17367 = n16812 & n16841;
  assign n17368 = n16803 & n16834;
  assign n17369 = ~n17367 & ~n17368;
  assign n17370 = n16801 & n16858;
  assign n17371 = n16812 & n16845;
  assign n17372 = ~n17370 & ~n17371;
  assign n17373 = n16812 & n16839;
  assign n17374 = n16800 ^ n16799;
  assign n17375 = n16819 & ~n17374;
  assign n17376 = ~n17373 & ~n17375;
  assign n17377 = n16803 & n16853;
  assign n17378 = ~n16827 & ~n16859;
  assign n17379 = n16801 & ~n17378;
  assign n17380 = n16829 & n16861;
  assign n17381 = n16816 & ~n17380;
  assign n17382 = ~n17379 & ~n17381;
  assign n17383 = ~n17377 & n17382;
  assign n17384 = n17376 & n17383;
  assign n17385 = n16821 & n17384;
  assign n17386 = n17372 & n17385;
  assign n17387 = n17369 & n17386;
  assign n17388 = n16832 & n17387;
  assign n17389 = n17366 & n17388;
  assign n17390 = n16811 & n17389;
  assign n17391 = n17390 ^ n15194;
  assign n17392 = n17391 ^ x753;
  assign n17393 = n16398 ^ x712;
  assign n17394 = n16950 ^ x717;
  assign n17395 = n17393 & ~n17394;
  assign n17396 = n14660 & n14664;
  assign n17397 = n14661 & ~n15956;
  assign n17398 = ~n17396 & ~n17397;
  assign n17399 = n14651 & ~n14689;
  assign n17400 = ~n14683 & ~n14695;
  assign n17401 = n14656 & ~n17400;
  assign n17402 = n14664 & ~n15957;
  assign n17403 = ~n14113 & n14656;
  assign n17404 = ~n13520 & n17403;
  assign n17405 = ~n17402 & ~n17404;
  assign n17406 = n15956 & n16529;
  assign n17407 = n14651 & ~n17406;
  assign n17408 = n14684 & ~n14695;
  assign n17409 = ~n14692 & n17408;
  assign n17410 = n14661 & ~n17409;
  assign n17411 = ~n17407 & ~n17410;
  assign n17412 = n17405 & n17411;
  assign n17413 = ~n17401 & n17412;
  assign n17414 = ~n17399 & n17413;
  assign n17415 = n17398 & n17414;
  assign n17416 = n14674 & n17415;
  assign n17417 = n16539 & n17416;
  assign n17418 = n15945 & n17417;
  assign n17419 = n17418 ^ n13626;
  assign n17420 = n17419 ^ x714;
  assign n17421 = n15545 & n15646;
  assign n17422 = n15614 & ~n15652;
  assign n17423 = ~n17421 & ~n17422;
  assign n17424 = ~n15642 & n15652;
  assign n17425 = ~n15635 & n17424;
  assign n17426 = n15547 & ~n17425;
  assign n17427 = ~n15630 & n15655;
  assign n17428 = n15546 & ~n17427;
  assign n17429 = ~n15622 & n16105;
  assign n17430 = n15650 & ~n17429;
  assign n17431 = ~n17428 & ~n17430;
  assign n17432 = n15547 & ~n15654;
  assign n17433 = ~n15617 & n15636;
  assign n17434 = ~n15626 & n17433;
  assign n17435 = n15605 & ~n17434;
  assign n17436 = ~n17432 & ~n17435;
  assign n17437 = n17431 & n17436;
  assign n17438 = ~n17426 & n17437;
  assign n17439 = n17423 & n17438;
  assign n17440 = n15625 & n17439;
  assign n17441 = ~n16110 & n17440;
  assign n17442 = ~n15618 & n17441;
  assign n17443 = n17442 ^ n13654;
  assign n17444 = n17443 ^ x715;
  assign n17445 = n17420 & ~n17444;
  assign n17446 = n16903 ^ x716;
  assign n17447 = n16479 ^ x713;
  assign n17448 = n17446 & n17447;
  assign n17449 = n17445 & n17448;
  assign n17450 = n17395 & n17449;
  assign n17451 = ~n17420 & n17444;
  assign n17452 = n17446 & ~n17447;
  assign n17453 = n17451 & n17452;
  assign n17454 = n17395 & n17453;
  assign n17455 = n17393 & n17394;
  assign n17456 = ~n17446 & ~n17447;
  assign n17457 = n17445 & n17456;
  assign n17458 = n17455 & n17457;
  assign n17459 = ~n17454 & ~n17458;
  assign n17460 = ~n17450 & n17459;
  assign n17461 = ~n17446 & n17447;
  assign n17462 = n17445 & n17461;
  assign n17463 = n17395 & n17462;
  assign n17464 = ~n17393 & ~n17394;
  assign n17465 = ~n17420 & ~n17444;
  assign n17466 = n17447 & n17465;
  assign n17467 = ~n17446 & n17466;
  assign n17468 = ~n17449 & ~n17467;
  assign n17469 = n17464 & ~n17468;
  assign n17470 = ~n17463 & ~n17469;
  assign n17471 = ~n17393 & n17394;
  assign n17472 = n17453 & n17471;
  assign n17473 = n17445 & n17452;
  assign n17474 = n17420 & n17444;
  assign n17475 = n17452 & n17474;
  assign n17476 = ~n17473 & ~n17475;
  assign n17477 = n17464 & ~n17476;
  assign n17478 = ~n17472 & ~n17477;
  assign n17479 = n17451 & n17456;
  assign n17480 = n17471 & n17479;
  assign n17481 = n17395 & n17457;
  assign n17482 = n17453 & n17455;
  assign n17483 = ~n17481 & ~n17482;
  assign n17484 = ~n17480 & n17483;
  assign n17485 = n17471 & n17473;
  assign n17486 = n17455 & n17479;
  assign n17487 = ~n17485 & ~n17486;
  assign n17488 = n17448 & n17451;
  assign n17489 = ~n17393 & n17488;
  assign n17490 = ~n17395 & ~n17471;
  assign n17491 = n17452 & n17465;
  assign n17492 = n17490 & n17491;
  assign n17493 = ~n17489 & ~n17492;
  assign n17494 = n17446 & n17466;
  assign n17495 = n17461 & n17474;
  assign n17496 = ~n17494 & ~n17495;
  assign n17497 = ~n17475 & n17496;
  assign n17498 = ~n17490 & ~n17497;
  assign n17499 = n17493 & ~n17498;
  assign n17500 = n17451 & n17461;
  assign n17501 = ~n17394 & n17500;
  assign n17502 = n17456 & n17474;
  assign n17503 = n17464 & n17502;
  assign n17504 = ~n17501 & ~n17503;
  assign n17505 = n17456 & n17465;
  assign n17506 = n17471 & n17505;
  assign n17507 = n17448 & n17474;
  assign n17508 = ~n17462 & ~n17507;
  assign n17509 = ~n17466 & n17508;
  assign n17510 = n17455 & ~n17509;
  assign n17511 = ~n17506 & ~n17510;
  assign n17512 = n17504 & n17511;
  assign n17513 = n17499 & n17512;
  assign n17514 = n17487 & n17513;
  assign n17515 = n17484 & n17514;
  assign n17516 = n17478 & n17515;
  assign n17517 = n17470 & n17516;
  assign n17518 = n17460 & n17517;
  assign n17519 = n17518 ^ n13852;
  assign n17520 = n17519 ^ x748;
  assign n17521 = ~n17392 & n17520;
  assign n17522 = n17360 & n17521;
  assign n17523 = ~n17200 & ~n17233;
  assign n17524 = ~n17330 & n17358;
  assign n17525 = n17523 & n17524;
  assign n17526 = n17392 & n17520;
  assign n17527 = n17525 & n17526;
  assign n17528 = ~n17522 & ~n17527;
  assign n17529 = n17200 & n17233;
  assign n17530 = n17524 & n17529;
  assign n17531 = n17359 & n17529;
  assign n17532 = ~n17530 & ~n17531;
  assign n17533 = ~n17392 & ~n17520;
  assign n17534 = ~n17532 & n17533;
  assign n17535 = ~n17330 & ~n17358;
  assign n17536 = n17529 & n17535;
  assign n17537 = n17526 & n17536;
  assign n17538 = n17523 & n17535;
  assign n17539 = ~n17360 & ~n17538;
  assign n17540 = n17392 & ~n17520;
  assign n17541 = ~n17539 & n17540;
  assign n17542 = ~n17537 & ~n17541;
  assign n17543 = ~n17525 & ~n17538;
  assign n17544 = n17533 & ~n17543;
  assign n17545 = n17330 & n17358;
  assign n17546 = n17234 & n17545;
  assign n17547 = n17526 & n17546;
  assign n17548 = ~n17200 & n17233;
  assign n17549 = n17524 & n17548;
  assign n17550 = ~n17531 & ~n17549;
  assign n17551 = n17540 & ~n17550;
  assign n17552 = ~n17547 & ~n17551;
  assign n17553 = n17523 & n17545;
  assign n17554 = n17526 & n17553;
  assign n17555 = n17545 & n17548;
  assign n17556 = n17520 ^ n17392;
  assign n17557 = n17555 & n17556;
  assign n17558 = ~n17554 & ~n17557;
  assign n17559 = n17234 & n17535;
  assign n17560 = ~n17521 & ~n17526;
  assign n17561 = n17559 & ~n17560;
  assign n17562 = ~n17546 & ~n17553;
  assign n17563 = ~n17536 & n17562;
  assign n17564 = n17533 & ~n17563;
  assign n17565 = n17529 & n17545;
  assign n17566 = n17535 & n17548;
  assign n17567 = ~n17565 & ~n17566;
  assign n17568 = n17556 & ~n17567;
  assign n17569 = ~n17564 & ~n17568;
  assign n17570 = ~n17561 & n17569;
  assign n17571 = n17359 & n17548;
  assign n17572 = ~n17392 & n17571;
  assign n17573 = n17234 & n17524;
  assign n17574 = n17540 & n17573;
  assign n17575 = ~n17572 & ~n17574;
  assign n17576 = n17359 & n17523;
  assign n17577 = ~n17573 & ~n17576;
  assign n17578 = n17521 & ~n17577;
  assign n17579 = ~n17530 & ~n17571;
  assign n17580 = ~n17566 & n17579;
  assign n17581 = n17526 & ~n17580;
  assign n17582 = ~n17578 & ~n17581;
  assign n17583 = n17575 & n17582;
  assign n17584 = n17570 & n17583;
  assign n17585 = n17558 & n17584;
  assign n17586 = n17552 & n17585;
  assign n17587 = ~n17544 & n17586;
  assign n17588 = n17542 & n17587;
  assign n17589 = ~n17534 & n17588;
  assign n17590 = n17528 & n17589;
  assign n17591 = n17590 ^ n16398;
  assign n17592 = n17591 ^ x808;
  assign n17593 = n16483 & ~n17184;
  assign n17594 = ~n16515 & ~n17178;
  assign n17595 = n16481 & ~n17594;
  assign n17596 = ~n17593 & ~n17595;
  assign n17597 = n16508 & ~n17191;
  assign n17598 = n16506 & n17195;
  assign n17599 = ~n17597 & ~n17598;
  assign n17600 = n17596 & n17599;
  assign n17601 = ~n16511 & n17600;
  assign n17602 = n17601 ^ n15760;
  assign n17603 = n17602 ^ x783;
  assign n17604 = ~n16815 & ~n16819;
  assign n17605 = n16803 & ~n17604;
  assign n17606 = ~n16824 & n16829;
  assign n17607 = n16801 & ~n17606;
  assign n17608 = ~n17605 & ~n17607;
  assign n17609 = n16803 & n16841;
  assign n17610 = n16801 & ~n16842;
  assign n17611 = ~n17609 & ~n17610;
  assign n17612 = n16816 & n16845;
  assign n17613 = ~n16834 & ~n16858;
  assign n17614 = ~n17374 & ~n17613;
  assign n17615 = ~n17612 & ~n17614;
  assign n17616 = ~n16808 & n16829;
  assign n17617 = n16812 & ~n17616;
  assign n17618 = ~n16805 & n16861;
  assign n17619 = ~n16816 & n17618;
  assign n17620 = ~n16798 & n16860;
  assign n17621 = ~n16855 & n17620;
  assign n17622 = ~n16803 & n17621;
  assign n17623 = ~n17619 & ~n17622;
  assign n17624 = n16799 & n17623;
  assign n17625 = ~n17617 & ~n17624;
  assign n17626 = n17615 & n17625;
  assign n17627 = n17611 & n17626;
  assign n17628 = n17608 & n17627;
  assign n17629 = n17366 & n17628;
  assign n17630 = n16822 & n17629;
  assign n17631 = n17630 ^ n15484;
  assign n17632 = n17631 ^ x778;
  assign n17633 = ~n17603 & ~n17632;
  assign n17634 = n17304 & n17318;
  assign n17635 = ~n17300 & n17307;
  assign n17636 = n17296 & n17635;
  assign n17637 = n17286 & ~n17636;
  assign n17638 = ~n17634 & ~n17637;
  assign n17639 = n17277 & n17281;
  assign n17640 = ~n17309 & ~n17639;
  assign n17641 = n17235 & ~n17640;
  assign n17642 = n17276 & n17282;
  assign n17643 = ~n17293 & ~n17642;
  assign n17644 = n17302 & n17643;
  assign n17645 = n17237 & ~n17644;
  assign n17646 = n17298 & n17643;
  assign n17647 = ~n17294 & n17646;
  assign n17648 = ~n17275 & n17647;
  assign n17649 = n17289 & ~n17648;
  assign n17650 = ~n17645 & ~n17649;
  assign n17651 = ~n17641 & n17650;
  assign n17652 = n17638 & n17651;
  assign n17653 = ~n17280 & n17652;
  assign n17654 = n17653 ^ n15782;
  assign n17655 = n17654 ^ x782;
  assign n17656 = n16664 & n16708;
  assign n17657 = ~n16625 & ~n16707;
  assign n17658 = n16689 & ~n17657;
  assign n17659 = ~n17656 & ~n17658;
  assign n17660 = n16668 & n16697;
  assign n17661 = n16666 & n16671;
  assign n17662 = ~n17660 & ~n17661;
  assign n17663 = ~n16677 & ~n16706;
  assign n17664 = n16666 & ~n17663;
  assign n17665 = ~n16693 & ~n16706;
  assign n17666 = n16702 & n17665;
  assign n17667 = ~n16681 & n17666;
  assign n17668 = n16664 & ~n17667;
  assign n17669 = ~n17664 & ~n17668;
  assign n17670 = n16678 & ~n16690;
  assign n17671 = ~n16671 & n17670;
  assign n17672 = n16689 & ~n17671;
  assign n17673 = ~n16701 & ~n16708;
  assign n17674 = ~n16687 & n17673;
  assign n17675 = n16700 & n17674;
  assign n17676 = ~n16713 & n17675;
  assign n17677 = n16668 & ~n17676;
  assign n17678 = ~n17672 & ~n17677;
  assign n17679 = n17669 & n17678;
  assign n17680 = n16673 & n17679;
  assign n17681 = ~n16686 & n17680;
  assign n17682 = n17662 & n17681;
  assign n17683 = n17659 & n17682;
  assign n17684 = n17210 & n17683;
  assign n17685 = n17204 & n17684;
  assign n17686 = ~n16665 & n17685;
  assign n17687 = n17686 ^ n16291;
  assign n17688 = n17687 ^ x781;
  assign n17689 = ~n17655 & n17688;
  assign n17690 = n15857 & n15880;
  assign n17691 = n15864 & ~n15890;
  assign n17692 = ~n17690 & ~n17691;
  assign n17693 = n15864 & n15893;
  assign n17694 = ~n15872 & ~n15909;
  assign n17695 = ~n15849 & n17694;
  assign n17696 = ~n15867 & n17695;
  assign n17697 = n15851 & ~n17696;
  assign n17698 = ~n17693 & ~n17697;
  assign n17699 = n15155 & ~n15911;
  assign n17700 = ~n15861 & ~n15880;
  assign n17701 = ~n15851 & n17700;
  assign n17702 = ~n15155 & n15894;
  assign n17703 = ~n17701 & ~n17702;
  assign n17704 = ~n17699 & ~n17703;
  assign n17705 = ~n15892 & ~n15902;
  assign n17706 = n15857 & ~n17705;
  assign n17707 = ~n15867 & n15911;
  assign n17708 = n15864 & ~n17707;
  assign n17709 = ~n15854 & n15890;
  assign n17710 = ~n15893 & n17709;
  assign n17711 = n15857 & ~n17710;
  assign n17712 = ~n17708 & ~n17711;
  assign n17713 = ~n17706 & n17712;
  assign n17714 = n17704 & n17713;
  assign n17715 = n17698 & n17714;
  assign n17716 = n17692 & n17715;
  assign n17717 = ~n15905 & n17716;
  assign n17718 = n15856 & n17717;
  assign n17719 = n15900 & n17718;
  assign n17720 = ~n15881 & n17719;
  assign n17721 = n17720 ^ n16264;
  assign n17722 = n17721 ^ x780;
  assign n17723 = n16921 & n17074;
  assign n17724 = ~n17051 & ~n17077;
  assign n17725 = ~n16920 & ~n17724;
  assign n17726 = ~n17723 & ~n17725;
  assign n17727 = ~n17038 & ~n17057;
  assign n17728 = ~n17342 & ~n17727;
  assign n17729 = ~n17030 & ~n17090;
  assign n17730 = n17040 & ~n17729;
  assign n17731 = ~n17027 & n17046;
  assign n17732 = n17054 & ~n17731;
  assign n17733 = ~n17042 & n17337;
  assign n17734 = ~n17056 & n17733;
  assign n17735 = n17037 & ~n17734;
  assign n17736 = ~n17732 & ~n17735;
  assign n17737 = ~n17730 & n17736;
  assign n17738 = ~n17728 & n17737;
  assign n17739 = n17726 & n17738;
  assign n17740 = n17073 & n17739;
  assign n17741 = ~n17068 & n17740;
  assign n17742 = n17048 & n17741;
  assign n17743 = n17335 & n17742;
  assign n17744 = ~n17036 & n17743;
  assign n17745 = ~n17032 & n17744;
  assign n17746 = n17745 ^ n15370;
  assign n17747 = n17746 ^ x779;
  assign n17748 = n17722 & ~n17747;
  assign n17749 = n17689 & n17748;
  assign n17750 = n17655 & n17688;
  assign n17751 = ~n17722 & ~n17747;
  assign n17752 = n17750 & n17751;
  assign n17753 = ~n17749 & ~n17752;
  assign n17754 = n17633 & ~n17753;
  assign n17755 = n17603 & ~n17632;
  assign n17756 = ~n17655 & ~n17688;
  assign n17757 = ~n17722 & n17747;
  assign n17758 = n17756 & n17757;
  assign n17759 = n17655 & ~n17688;
  assign n17760 = n17747 & n17759;
  assign n17761 = n17722 & n17760;
  assign n17762 = n17722 & n17747;
  assign n17763 = n17689 & n17762;
  assign n17764 = ~n17761 & ~n17763;
  assign n17765 = ~n17758 & n17764;
  assign n17766 = n17755 & ~n17765;
  assign n17767 = n17689 & n17757;
  assign n17768 = n17750 & n17762;
  assign n17769 = ~n17767 & ~n17768;
  assign n17770 = n17633 & ~n17769;
  assign n17771 = n17751 & n17759;
  assign n17772 = ~n17749 & ~n17771;
  assign n17773 = n17755 & ~n17772;
  assign n17774 = ~n17770 & ~n17773;
  assign n17775 = ~n17603 & n17632;
  assign n17776 = n17767 & n17775;
  assign n17777 = n17603 & n17632;
  assign n17778 = ~n17722 & n17760;
  assign n17779 = n17756 & n17762;
  assign n17780 = ~n17778 & ~n17779;
  assign n17781 = n17777 & ~n17780;
  assign n17782 = ~n17776 & ~n17781;
  assign n17783 = n17748 & n17756;
  assign n17784 = n17777 & n17783;
  assign n17785 = ~n17758 & ~n17761;
  assign n17786 = n17775 & ~n17785;
  assign n17787 = ~n17784 & ~n17786;
  assign n17788 = n17750 & n17757;
  assign n17789 = n17632 & n17788;
  assign n17790 = n17748 & n17759;
  assign n17791 = n17769 & ~n17790;
  assign n17792 = n17755 & ~n17791;
  assign n17793 = n17751 & n17756;
  assign n17794 = ~n17771 & ~n17793;
  assign n17795 = n17780 & n17794;
  assign n17796 = n17633 & ~n17795;
  assign n17797 = n17748 & n17750;
  assign n17798 = n17689 & n17751;
  assign n17799 = ~n17797 & ~n17798;
  assign n17800 = ~n17775 & n17799;
  assign n17801 = ~n17749 & n17800;
  assign n17802 = ~n17783 & ~n17790;
  assign n17803 = ~n17797 & n17802;
  assign n17804 = ~n17777 & n17803;
  assign n17805 = ~n17801 & ~n17804;
  assign n17806 = ~n17793 & ~n17805;
  assign n17807 = n17632 & ~n17806;
  assign n17808 = ~n17796 & ~n17807;
  assign n17809 = ~n17792 & n17808;
  assign n17810 = ~n17789 & n17809;
  assign n17811 = n17787 & n17810;
  assign n17812 = n17782 & n17811;
  assign n17813 = n17774 & n17812;
  assign n17814 = ~n17766 & n17813;
  assign n17815 = ~n17754 & n17814;
  assign n17816 = n17815 ^ n16950;
  assign n17817 = n17816 ^ x813;
  assign n17818 = ~n17592 & n17817;
  assign n17819 = n17329 ^ x754;
  assign n17820 = n16732 ^ x759;
  assign n17821 = ~n17819 & ~n17820;
  assign n17822 = n17391 ^ x755;
  assign n17823 = ~n16099 & n16168;
  assign n17824 = ~n16186 & ~n17823;
  assign n17825 = n16195 & n17824;
  assign n17826 = n16182 & ~n17825;
  assign n17827 = n16171 & n16212;
  assign n17828 = n16133 ^ n16099;
  assign n17829 = n16167 & ~n17828;
  assign n17830 = ~n16219 & ~n17829;
  assign n17831 = n15972 & ~n17830;
  assign n17832 = ~n17827 & ~n17831;
  assign n17833 = ~n17826 & n17832;
  assign n17834 = ~n16171 & ~n16191;
  assign n17835 = ~n16191 & n17823;
  assign n17836 = n17835 ^ n16168;
  assign n17837 = n16187 & ~n17836;
  assign n17838 = ~n16171 & n17824;
  assign n17839 = ~n17837 & ~n17838;
  assign n17840 = ~n16215 & ~n17839;
  assign n17841 = ~n17834 & ~n17840;
  assign n17842 = ~n16174 & ~n16198;
  assign n17843 = ~n15971 & ~n17842;
  assign n17844 = ~n17841 & ~n17843;
  assign n17845 = n17833 & n17844;
  assign n17846 = n16210 & n17845;
  assign n17847 = n16202 & n17846;
  assign n17848 = n16178 & n17847;
  assign n17849 = n17848 ^ n15251;
  assign n17850 = n17849 ^ x757;
  assign n17851 = n17822 & n17850;
  assign n17852 = n17395 & n17502;
  assign n17853 = n17457 & n17464;
  assign n17854 = ~n17852 & ~n17853;
  assign n17855 = n17475 & n17490;
  assign n17856 = ~n17462 & ~n17488;
  assign n17857 = n17471 & ~n17856;
  assign n17858 = ~n17855 & ~n17857;
  assign n17859 = n17854 & n17858;
  assign n17860 = ~n17490 & n17505;
  assign n17861 = n17464 & n17479;
  assign n17862 = ~n17860 & ~n17861;
  assign n17863 = n17395 & n17488;
  assign n17864 = ~n17491 & ~n17502;
  assign n17865 = n17455 & ~n17864;
  assign n17866 = ~n17863 & ~n17865;
  assign n17867 = n17395 & n17473;
  assign n17868 = ~n17394 & ~n17496;
  assign n17869 = ~n17867 & ~n17868;
  assign n17870 = n17455 & ~n17468;
  assign n17871 = n17490 & n17500;
  assign n17872 = ~n17500 & ~n17507;
  assign n17873 = ~n17491 & n17872;
  assign n17874 = ~n17475 & n17873;
  assign n17875 = n17471 & ~n17874;
  assign n17876 = ~n17871 & ~n17875;
  assign n17877 = ~n17870 & n17876;
  assign n17878 = n17869 & n17877;
  assign n17879 = n17866 & n17878;
  assign n17880 = n17862 & n17879;
  assign n17881 = n17459 & n17880;
  assign n17882 = n17487 & n17881;
  assign n17883 = n17470 & n17882;
  assign n17884 = n17859 & n17883;
  assign n17885 = n17884 ^ n15229;
  assign n17886 = n17885 ^ x756;
  assign n17887 = n17851 & n17886;
  assign n17888 = ~n17822 & ~n17850;
  assign n17889 = n15929 ^ x758;
  assign n17890 = n17886 & n17889;
  assign n17891 = n17888 & ~n17890;
  assign n17892 = ~n17887 & ~n17891;
  assign n17893 = n17822 & n17890;
  assign n17894 = ~n17886 & n17889;
  assign n17895 = n17850 & n17894;
  assign n17896 = ~n17893 & ~n17895;
  assign n17897 = n17892 & n17896;
  assign n17898 = n17821 & ~n17897;
  assign n17899 = n17819 & ~n17820;
  assign n17900 = n17889 ^ n17850;
  assign n17901 = n17822 & ~n17900;
  assign n17902 = ~n17886 & n17888;
  assign n17903 = n17886 & ~n17889;
  assign n17904 = n17850 & n17903;
  assign n17905 = ~n17894 & ~n17904;
  assign n17906 = ~n17822 & ~n17905;
  assign n17907 = ~n17902 & ~n17906;
  assign n17908 = ~n17901 & n17907;
  assign n17909 = n17899 & n17908;
  assign n17910 = ~n17898 & ~n17909;
  assign n17911 = n17819 & n17820;
  assign n17912 = n17888 & n17890;
  assign n17913 = ~n17886 & ~n17889;
  assign n17914 = ~n17822 & n17913;
  assign n17915 = ~n17912 & ~n17914;
  assign n17916 = ~n17822 & n17850;
  assign n17917 = ~n17886 & n17916;
  assign n17918 = n17850 & n17890;
  assign n17919 = n17822 & ~n17850;
  assign n17920 = ~n17890 & ~n17913;
  assign n17921 = n17919 & n17920;
  assign n17922 = ~n17918 & ~n17921;
  assign n17923 = ~n17917 & n17922;
  assign n17924 = n17915 & n17923;
  assign n17925 = n17911 & ~n17924;
  assign n17926 = ~n17819 & n17820;
  assign n17927 = n17903 & n17916;
  assign n17928 = n17851 & ~n17886;
  assign n17929 = ~n17927 & ~n17928;
  assign n17930 = n17888 & n17889;
  assign n17931 = ~n17850 & ~n17920;
  assign n17932 = ~n17930 & ~n17931;
  assign n17933 = n17929 & n17932;
  assign n17934 = n17926 & ~n17933;
  assign n17935 = ~n17925 & ~n17934;
  assign n17936 = n17910 & n17935;
  assign n17937 = n17936 ^ n16903;
  assign n17938 = n17937 ^ x812;
  assign n17939 = ~n15870 & ~n15902;
  assign n17940 = n15864 & ~n17939;
  assign n17941 = n15908 & ~n17940;
  assign n17942 = n17696 & n17709;
  assign n17943 = n15857 & ~n17942;
  assign n17944 = n15894 & ~n15897;
  assign n17945 = ~n15873 & n17944;
  assign n17946 = n15864 & ~n17945;
  assign n17947 = ~n17943 & ~n17946;
  assign n17948 = n15155 & n15867;
  assign n17949 = ~n15880 & ~n15892;
  assign n17950 = ~n15889 & ~n15893;
  assign n17951 = ~n15155 & n17950;
  assign n17952 = ~n15851 & n15890;
  assign n17953 = ~n17951 & ~n17952;
  assign n17954 = n17949 & ~n17953;
  assign n17955 = ~n15909 & n17954;
  assign n17956 = ~n14718 & ~n17955;
  assign n17957 = ~n17948 & ~n17956;
  assign n17958 = n17947 & n17957;
  assign n17959 = n17941 & n17958;
  assign n17960 = n15856 & n17959;
  assign n17961 = ~n15904 & n17960;
  assign n17962 = n15900 & n17961;
  assign n17963 = n17962 ^ n14331;
  assign n17964 = n17963 ^ x744;
  assign n17965 = n17283 & n17289;
  assign n17966 = n17285 & n17318;
  assign n17967 = ~n17965 & ~n17966;
  assign n17968 = n17289 & n17294;
  assign n17969 = n17276 & n17292;
  assign n17970 = ~n17300 & ~n17969;
  assign n17971 = ~n17297 & n17970;
  assign n17972 = ~n17291 & n17971;
  assign n17973 = ~n17275 & n17972;
  assign n17974 = n17643 & n17973;
  assign n17975 = n17318 & ~n17974;
  assign n17976 = n17236 ^ n17235;
  assign n17977 = ~n17299 & ~n17308;
  assign n17978 = n17640 & n17977;
  assign n17979 = n17976 & ~n17978;
  assign n17980 = n17237 & ~n17296;
  assign n17981 = ~n17979 & ~n17980;
  assign n17982 = ~n17278 & ~n17306;
  assign n17983 = n17235 & ~n17982;
  assign n17984 = ~n17308 & n17972;
  assign n17985 = n17286 & ~n17984;
  assign n17986 = ~n17983 & ~n17985;
  assign n17987 = n17981 & n17986;
  assign n17988 = ~n17975 & n17987;
  assign n17989 = ~n17968 & n17988;
  assign n17990 = n17288 & n17989;
  assign n17991 = n17967 & n17990;
  assign n17992 = n17991 ^ n13519;
  assign n17993 = n17992 ^ x745;
  assign n17994 = n16169 & n16191;
  assign n17995 = n15972 & n16203;
  assign n17996 = ~n16176 & n16182;
  assign n17997 = ~n17995 & ~n17996;
  assign n17998 = ~n17994 & n17997;
  assign n17999 = ~n16203 & n16216;
  assign n18000 = n16187 & n17999;
  assign n18001 = n16195 & n18000;
  assign n18002 = n16191 & ~n18001;
  assign n18003 = n16099 & n16184;
  assign n18004 = n16171 & n18003;
  assign n18005 = n16200 & ~n16219;
  assign n18006 = n16182 & ~n18005;
  assign n18007 = ~n18004 & ~n18006;
  assign n18008 = ~n18002 & n18007;
  assign n18009 = n16168 & n16183;
  assign n18010 = n16223 & ~n18009;
  assign n18011 = n15972 & ~n18010;
  assign n18012 = n16195 & ~n16212;
  assign n18013 = ~n15972 & n18012;
  assign n18014 = ~n16208 & n16216;
  assign n18015 = ~n16171 & n18014;
  assign n18016 = ~n18013 & ~n18015;
  assign n18017 = ~n16175 & ~n18016;
  assign n18018 = n15971 & ~n18017;
  assign n18019 = ~n18011 & ~n18018;
  assign n18020 = n18008 & n18019;
  assign n18021 = n17998 & n18020;
  assign n18022 = n16190 & n18021;
  assign n18023 = n18022 ^ n14112;
  assign n18024 = n18023 ^ x743;
  assign n18025 = n17993 & n18024;
  assign n18026 = n17519 ^ x746;
  assign n18027 = n18025 & n18026;
  assign n18028 = ~n17964 & n18027;
  assign n18029 = n17232 ^ x747;
  assign n18030 = n17056 & ~n17342;
  assign n18031 = n17054 & ~n17347;
  assign n18032 = ~n18030 & ~n18031;
  assign n18033 = n17040 & n17074;
  assign n18034 = ~n16920 & n17027;
  assign n18035 = ~n18033 & ~n18034;
  assign n18036 = ~n17030 & n17337;
  assign n18037 = n17037 & ~n18036;
  assign n18038 = ~n17071 & ~n17077;
  assign n18039 = n17054 & ~n18038;
  assign n18040 = ~n17057 & n17078;
  assign n18041 = n16921 & ~n18040;
  assign n18042 = ~n18039 & ~n18041;
  assign n18043 = n17040 & ~n17733;
  assign n18044 = n17727 & ~n18043;
  assign n18045 = ~n17083 & n18044;
  assign n18046 = ~n17051 & n18045;
  assign n18047 = n17342 & ~n18046;
  assign n18048 = n18042 & ~n18047;
  assign n18049 = ~n17332 & n18048;
  assign n18050 = ~n17036 & n18049;
  assign n18051 = ~n18037 & n18050;
  assign n18052 = n18035 & n18051;
  assign n18053 = n18032 & n18052;
  assign n18054 = n17064 & n18053;
  assign n18055 = n18054 ^ n14649;
  assign n18056 = n18055 ^ x742;
  assign n18057 = n18029 & n18056;
  assign n18058 = n18028 & n18057;
  assign n18059 = n17964 & ~n18026;
  assign n18060 = n18025 & n18059;
  assign n18061 = n18029 & ~n18056;
  assign n18062 = n18060 & n18061;
  assign n18063 = ~n18058 & ~n18062;
  assign n18064 = ~n18029 & n18056;
  assign n18065 = n18060 & n18064;
  assign n18066 = n17964 & n18027;
  assign n18067 = n18061 & n18066;
  assign n18068 = ~n18065 & ~n18067;
  assign n18069 = ~n17993 & n18026;
  assign n18070 = n17964 & n18069;
  assign n18071 = n18024 & n18070;
  assign n18072 = ~n17964 & ~n18026;
  assign n18073 = n18025 & n18072;
  assign n18074 = ~n18071 & ~n18073;
  assign n18075 = ~n18029 & ~n18056;
  assign n18076 = ~n18074 & n18075;
  assign n18077 = ~n17964 & n18069;
  assign n18078 = ~n18024 & n18077;
  assign n18079 = n17993 & ~n18024;
  assign n18080 = n18072 & n18079;
  assign n18081 = ~n18078 & ~n18080;
  assign n18082 = n18061 & ~n18081;
  assign n18083 = ~n18076 & ~n18082;
  assign n18084 = ~n18071 & ~n18079;
  assign n18085 = n18064 & ~n18084;
  assign n18086 = ~n17993 & n18059;
  assign n18087 = n18024 & n18086;
  assign n18088 = ~n18028 & ~n18087;
  assign n18089 = n18061 & ~n18088;
  assign n18090 = ~n18024 & n18070;
  assign n18091 = ~n17993 & n18072;
  assign n18092 = ~n18024 & n18091;
  assign n18093 = ~n18090 & ~n18092;
  assign n18094 = ~n18064 & ~n18093;
  assign n18095 = n18024 & n18077;
  assign n18096 = ~n18087 & ~n18095;
  assign n18097 = n18056 & ~n18096;
  assign n18098 = ~n18094 & ~n18097;
  assign n18099 = n18059 & n18079;
  assign n18100 = ~n18060 & ~n18099;
  assign n18101 = ~n18078 & n18100;
  assign n18102 = n18057 & ~n18101;
  assign n18103 = n18024 & n18091;
  assign n18104 = n18026 & n18079;
  assign n18105 = ~n17964 & n18104;
  assign n18106 = ~n18024 & n18086;
  assign n18107 = ~n18105 & ~n18106;
  assign n18108 = ~n18103 & n18107;
  assign n18109 = ~n18028 & n18108;
  assign n18110 = n18075 & ~n18109;
  assign n18111 = ~n18102 & ~n18110;
  assign n18112 = n18098 & n18111;
  assign n18113 = ~n18089 & n18112;
  assign n18114 = ~n18085 & n18113;
  assign n18115 = n18083 & n18114;
  assign n18116 = n18068 & n18115;
  assign n18117 = n18063 & n18116;
  assign n18118 = n18117 ^ n17419;
  assign n18119 = n18118 ^ x810;
  assign n18120 = ~n17938 & ~n18119;
  assign n18121 = n16526 ^ x766;
  assign n18122 = n17471 & n17502;
  assign n18123 = n17394 & n17473;
  assign n18124 = n17464 & n17505;
  assign n18125 = ~n18123 & ~n18124;
  assign n18126 = ~n18122 & n18125;
  assign n18127 = n17490 & ~n17856;
  assign n18128 = n17471 & ~n17509;
  assign n18129 = ~n18127 & ~n18128;
  assign n18130 = n17464 & n17466;
  assign n18131 = n17455 & ~n17872;
  assign n18132 = ~n17495 & n17872;
  assign n18133 = ~n17491 & n18132;
  assign n18134 = n17395 & ~n18133;
  assign n18135 = ~n18131 & ~n18134;
  assign n18136 = ~n18130 & n18135;
  assign n18137 = n18129 & n18136;
  assign n18138 = n17866 & n18137;
  assign n18139 = n17862 & n18138;
  assign n18140 = n18126 & n18139;
  assign n18141 = n17478 & n18140;
  assign n18142 = n17460 & n18141;
  assign n18143 = n18142 ^ n15459;
  assign n18144 = n18143 ^ x771;
  assign n18145 = ~n18121 & ~n18144;
  assign n18146 = ~n17306 & ~n17969;
  assign n18147 = ~n17294 & n18146;
  assign n18148 = n17318 & ~n18147;
  assign n18149 = n17289 & ~n17310;
  assign n18150 = ~n18148 & ~n18149;
  assign n18151 = n17235 & n17291;
  assign n18152 = ~n17285 & n17977;
  assign n18153 = ~n17291 & n18152;
  assign n18154 = n17237 & ~n18153;
  assign n18155 = ~n18151 & ~n18154;
  assign n18156 = n17298 & ~n17639;
  assign n18157 = n17286 & ~n18156;
  assign n18158 = n17237 & n17294;
  assign n18159 = ~n17278 & n17643;
  assign n18160 = ~n17285 & n18159;
  assign n18161 = n17237 & n17282;
  assign n18162 = ~n17289 & ~n18161;
  assign n18163 = ~n18160 & ~n18162;
  assign n18164 = ~n17275 & n18147;
  assign n18165 = n17286 & ~n18164;
  assign n18166 = ~n17297 & n17301;
  assign n18167 = ~n17308 & n18166;
  assign n18168 = n17318 & ~n18167;
  assign n18169 = ~n18165 & ~n18168;
  assign n18170 = ~n18163 & n18169;
  assign n18171 = ~n18158 & n18170;
  assign n18172 = ~n17280 & n18171;
  assign n18173 = ~n18157 & n18172;
  assign n18174 = n18155 & n18173;
  assign n18175 = n18150 & n18174;
  assign n18176 = n17967 & n18175;
  assign n18177 = n18176 ^ n15571;
  assign n18178 = n18177 ^ x768;
  assign n18179 = n16684 & n16689;
  assign n18180 = ~n16687 & n17665;
  assign n18181 = ~n16707 & n18180;
  assign n18182 = n16668 & ~n18181;
  assign n18183 = ~n18179 & ~n18182;
  assign n18184 = n16664 & n16713;
  assign n18185 = ~n16707 & n17674;
  assign n18186 = n16666 & ~n18185;
  assign n18187 = ~n16701 & n17663;
  assign n18188 = ~n16664 & n18187;
  assign n18189 = n17205 & n17665;
  assign n18190 = ~n16689 & n18189;
  assign n18191 = ~n18188 & ~n18190;
  assign n18192 = ~n16681 & ~n18191;
  assign n18193 = ~n16663 & ~n18192;
  assign n18194 = ~n18186 & ~n18193;
  assign n18195 = ~n18184 & n18194;
  assign n18196 = n18183 & n18195;
  assign n18197 = n17662 & n18196;
  assign n18198 = n17659 & n18197;
  assign n18199 = n16680 & n18198;
  assign n18200 = n17207 & n18199;
  assign n18201 = n18200 ^ n15600;
  assign n18202 = n18201 ^ x769;
  assign n18203 = n18178 & ~n18202;
  assign n18204 = ~n14718 & n15849;
  assign n18205 = ~n15883 & n17949;
  assign n18206 = n15864 & ~n18205;
  assign n18207 = ~n15873 & ~n15880;
  assign n18208 = n15155 & ~n18207;
  assign n18209 = ~n15881 & n15910;
  assign n18210 = ~n15892 & n18209;
  assign n18211 = n15851 & ~n18210;
  assign n18212 = ~n18208 & ~n18211;
  assign n18213 = ~n18206 & n18212;
  assign n18214 = ~n18204 & n18213;
  assign n18215 = ~n15861 & ~n15883;
  assign n18216 = ~n15889 & n18215;
  assign n18217 = n15155 & ~n18216;
  assign n18218 = n15874 & n17702;
  assign n18219 = ~n15854 & n18218;
  assign n18220 = n15857 & ~n18219;
  assign n18221 = ~n18217 & ~n18220;
  assign n18222 = n18214 & n18221;
  assign n18223 = ~n15898 & n18222;
  assign n18224 = n15863 & n18223;
  assign n18225 = n17692 & n18224;
  assign n18226 = n17941 & n18225;
  assign n18227 = ~n15905 & n18226;
  assign n18228 = ~n15904 & n18227;
  assign n18229 = n18228 ^ n15397;
  assign n18230 = n18229 ^ x770;
  assign n18231 = n16239 ^ x767;
  assign n18232 = ~n18230 & ~n18231;
  assign n18233 = n18203 & n18232;
  assign n18234 = n18145 & n18233;
  assign n18235 = n18121 & ~n18144;
  assign n18236 = ~n18178 & ~n18202;
  assign n18237 = n18232 & n18236;
  assign n18238 = n18230 & ~n18231;
  assign n18239 = n18203 & n18238;
  assign n18240 = ~n18237 & ~n18239;
  assign n18241 = n18235 & ~n18240;
  assign n18242 = ~n18234 & ~n18241;
  assign n18243 = n18121 & n18144;
  assign n18244 = n18178 & n18202;
  assign n18245 = ~n18230 & n18231;
  assign n18246 = n18244 & n18245;
  assign n18247 = n18230 & n18231;
  assign n18248 = n18236 & n18247;
  assign n18249 = ~n18178 & n18202;
  assign n18250 = n18245 & n18249;
  assign n18251 = ~n18248 & ~n18250;
  assign n18252 = ~n18246 & n18251;
  assign n18253 = n18243 & ~n18252;
  assign n18254 = n18238 & n18244;
  assign n18255 = n18235 & n18254;
  assign n18256 = ~n18121 & n18144;
  assign n18257 = ~n18235 & ~n18256;
  assign n18258 = n18247 & n18249;
  assign n18259 = n18252 & ~n18258;
  assign n18260 = ~n18256 & n18259;
  assign n18261 = n18244 & n18247;
  assign n18262 = n18203 & n18245;
  assign n18263 = ~n18246 & ~n18258;
  assign n18264 = ~n18262 & n18263;
  assign n18265 = ~n18261 & n18264;
  assign n18266 = ~n18235 & n18265;
  assign n18267 = ~n18260 & ~n18266;
  assign n18268 = ~n18257 & n18267;
  assign n18269 = n18238 & n18249;
  assign n18270 = ~n18237 & ~n18269;
  assign n18271 = n18232 & n18249;
  assign n18272 = ~n18239 & ~n18271;
  assign n18273 = n18270 & n18272;
  assign n18274 = n18243 & ~n18273;
  assign n18275 = n18236 & n18238;
  assign n18276 = ~n18271 & ~n18275;
  assign n18277 = n18240 & n18276;
  assign n18278 = n18256 & ~n18277;
  assign n18279 = ~n18274 & ~n18278;
  assign n18280 = ~n18268 & n18279;
  assign n18281 = n18203 & n18247;
  assign n18282 = n18121 & n18281;
  assign n18283 = n18236 & n18245;
  assign n18284 = n18232 & n18244;
  assign n18285 = ~n18254 & ~n18284;
  assign n18286 = ~n18262 & n18285;
  assign n18287 = n18251 & n18286;
  assign n18288 = ~n18269 & n18287;
  assign n18289 = ~n18283 & n18288;
  assign n18290 = n18145 & ~n18289;
  assign n18291 = ~n18282 & ~n18290;
  assign n18292 = n18280 & n18291;
  assign n18293 = ~n18255 & n18292;
  assign n18294 = ~n18253 & n18293;
  assign n18295 = n18242 & n18294;
  assign n18296 = n18295 ^ n17443;
  assign n18297 = n18296 ^ x811;
  assign n18298 = n17654 ^ x736;
  assign n18299 = n18023 ^ x741;
  assign n18300 = n18298 & n18299;
  assign n18301 = n16801 & n16855;
  assign n18302 = n16812 & n16834;
  assign n18303 = ~n18301 & ~n18302;
  assign n18304 = n16803 & ~n16846;
  assign n18305 = ~n16805 & ~n16859;
  assign n18306 = ~n16858 & n18305;
  assign n18307 = ~n16824 & n18306;
  assign n18308 = n16816 & ~n18307;
  assign n18309 = ~n16828 & ~n16840;
  assign n18310 = ~n16855 & n18309;
  assign n18311 = ~n17374 & ~n18310;
  assign n18312 = ~n18308 & ~n18311;
  assign n18313 = ~n18304 & n18312;
  assign n18314 = n18303 & n18313;
  assign n18315 = n17372 & n18314;
  assign n18316 = n17369 & n18315;
  assign n18317 = n16838 & n18316;
  assign n18318 = n17608 & n18317;
  assign n18319 = n16822 & n18318;
  assign n18320 = n16811 & n18319;
  assign n18321 = n18320 ^ n15727;
  assign n18322 = n18321 ^ x738;
  assign n18323 = ~n17444 & n17448;
  assign n18324 = n17471 & n18323;
  assign n18325 = ~n17490 & n17491;
  assign n18326 = ~n18324 & ~n18325;
  assign n18327 = n17468 & n17496;
  assign n18328 = n17395 & ~n18327;
  assign n18329 = ~n17494 & n17873;
  assign n18330 = n17464 & ~n18329;
  assign n18331 = ~n18328 & ~n18330;
  assign n18332 = ~n17394 & n17488;
  assign n18333 = ~n17467 & n18132;
  assign n18334 = ~n17457 & n18333;
  assign n18335 = n17455 & ~n18334;
  assign n18336 = ~n18332 & ~n18335;
  assign n18337 = n18331 & n18336;
  assign n18338 = n18326 & n18337;
  assign n18339 = n18126 & n18338;
  assign n18340 = n17484 & n18339;
  assign n18341 = n17859 & n18340;
  assign n18342 = n18341 ^ n15696;
  assign n18343 = n18342 ^ x739;
  assign n18344 = ~n18322 & n18343;
  assign n18345 = n17602 ^ x737;
  assign n18346 = n18055 ^ x740;
  assign n18347 = n18345 & n18346;
  assign n18348 = n18344 & n18347;
  assign n18349 = n18300 & n18348;
  assign n18350 = ~n18322 & ~n18343;
  assign n18351 = n18345 & ~n18346;
  assign n18352 = n18350 & n18351;
  assign n18353 = n18300 & n18352;
  assign n18354 = ~n18349 & ~n18353;
  assign n18355 = ~n18298 & n18299;
  assign n18356 = n18322 & ~n18343;
  assign n18357 = ~n18345 & n18346;
  assign n18358 = n18356 & n18357;
  assign n18359 = n18355 & n18358;
  assign n18360 = n18322 & n18343;
  assign n18361 = n18357 & n18360;
  assign n18362 = ~n18345 & ~n18346;
  assign n18363 = n18350 & n18362;
  assign n18364 = ~n18361 & ~n18363;
  assign n18365 = n18300 & ~n18364;
  assign n18366 = ~n18359 & ~n18365;
  assign n18367 = ~n18298 & ~n18299;
  assign n18368 = n18350 & n18357;
  assign n18369 = n18356 & n18362;
  assign n18370 = ~n18368 & ~n18369;
  assign n18371 = n18367 & ~n18370;
  assign n18372 = n18298 & ~n18299;
  assign n18373 = n18344 & n18357;
  assign n18374 = n18372 & n18373;
  assign n18375 = n18298 & n18369;
  assign n18376 = ~n18374 & ~n18375;
  assign n18377 = n18300 & n18360;
  assign n18378 = n18347 & n18377;
  assign n18379 = n18351 & n18377;
  assign n18380 = n18351 & n18356;
  assign n18381 = n18344 & n18351;
  assign n18382 = n18360 & n18362;
  assign n18383 = n18347 & n18360;
  assign n18384 = ~n18348 & ~n18383;
  assign n18385 = ~n18382 & n18384;
  assign n18386 = ~n18381 & n18385;
  assign n18387 = ~n18380 & n18386;
  assign n18388 = ~n18358 & n18387;
  assign n18389 = n18367 & ~n18388;
  assign n18390 = ~n18379 & ~n18389;
  assign n18391 = ~n18358 & ~n18368;
  assign n18392 = n18345 & n18360;
  assign n18393 = n18347 & n18356;
  assign n18394 = ~n18392 & ~n18393;
  assign n18395 = ~n18352 & n18394;
  assign n18396 = n18391 & n18395;
  assign n18397 = n18372 & ~n18396;
  assign n18398 = n18300 & n18368;
  assign n18399 = n18344 & n18362;
  assign n18400 = ~n18361 & ~n18399;
  assign n18401 = n18347 & n18350;
  assign n18402 = n18322 & n18351;
  assign n18403 = ~n18401 & ~n18402;
  assign n18404 = ~n18381 & n18403;
  assign n18405 = n18400 & n18404;
  assign n18406 = ~n18393 & n18405;
  assign n18407 = n18355 & ~n18406;
  assign n18408 = ~n18398 & ~n18407;
  assign n18409 = ~n18397 & n18408;
  assign n18410 = n18390 & n18409;
  assign n18411 = ~n18378 & n18410;
  assign n18412 = n18376 & n18411;
  assign n18413 = ~n18371 & n18412;
  assign n18414 = n18366 & n18413;
  assign n18415 = n18354 & n18414;
  assign n18416 = n18415 ^ n16479;
  assign n18417 = n18416 ^ x809;
  assign n18418 = n18297 & n18417;
  assign n18419 = n18120 & n18418;
  assign n18420 = n17818 & n18419;
  assign n18421 = n17592 & ~n17817;
  assign n18422 = ~n18297 & n18417;
  assign n18423 = n18120 & n18422;
  assign n18424 = n17938 & n18119;
  assign n18425 = ~n18297 & ~n18417;
  assign n18426 = n18424 & n18425;
  assign n18427 = ~n18423 & ~n18426;
  assign n18428 = n18421 & ~n18427;
  assign n18429 = ~n18420 & ~n18428;
  assign n18430 = ~n17938 & n18119;
  assign n18431 = n18297 & ~n18417;
  assign n18432 = n18430 & n18431;
  assign n18433 = n17818 & n18432;
  assign n18434 = ~n17592 & ~n17817;
  assign n18435 = n18423 & n18434;
  assign n18436 = n17817 ^ n17592;
  assign n18437 = n17938 & ~n18119;
  assign n18438 = n18425 & n18437;
  assign n18439 = ~n18436 & n18438;
  assign n18440 = ~n18435 & ~n18439;
  assign n18441 = n18418 & n18424;
  assign n18442 = n18422 & n18430;
  assign n18443 = ~n18441 & ~n18442;
  assign n18444 = n18434 & ~n18443;
  assign n18445 = n18440 & ~n18444;
  assign n18446 = n18431 & n18437;
  assign n18447 = n17818 & n18446;
  assign n18448 = n18418 & n18437;
  assign n18449 = n18418 & n18430;
  assign n18450 = ~n18448 & ~n18449;
  assign n18451 = n18434 & ~n18450;
  assign n18452 = ~n18447 & ~n18451;
  assign n18453 = n18421 & n18441;
  assign n18454 = n18120 & n18425;
  assign n18455 = n17818 & n18454;
  assign n18456 = ~n18453 & ~n18455;
  assign n18457 = n18422 & n18424;
  assign n18458 = n17818 & n18457;
  assign n18459 = n17592 & n17817;
  assign n18460 = n18454 & n18459;
  assign n18461 = ~n18458 & ~n18460;
  assign n18462 = n18422 & n18437;
  assign n18463 = n18459 & n18462;
  assign n18464 = n17818 & n18438;
  assign n18465 = ~n18463 & ~n18464;
  assign n18466 = n18426 & ~n18436;
  assign n18467 = n18432 & n18434;
  assign n18468 = ~n18466 & ~n18467;
  assign n18469 = n17818 & ~n18450;
  assign n18470 = n18424 & n18431;
  assign n18471 = n18120 & n18431;
  assign n18472 = ~n18470 & ~n18471;
  assign n18473 = ~n18442 & n18472;
  assign n18474 = ~n18448 & n18473;
  assign n18475 = n18459 & ~n18474;
  assign n18476 = n18425 & n18430;
  assign n18477 = ~n18446 & ~n18476;
  assign n18478 = ~n18470 & n18477;
  assign n18479 = ~n18462 & n18478;
  assign n18480 = ~n18419 & n18479;
  assign n18481 = n18421 & ~n18480;
  assign n18482 = ~n18475 & ~n18481;
  assign n18483 = ~n18469 & n18482;
  assign n18484 = n18468 & n18483;
  assign n18485 = n18465 & n18484;
  assign n18486 = n18461 & n18485;
  assign n18487 = n18456 & n18486;
  assign n18488 = n18452 & n18487;
  assign n18489 = n18445 & n18488;
  assign n18490 = ~n18433 & n18489;
  assign n18491 = n18429 & n18490;
  assign n18492 = n18491 ^ n17519;
  assign n18493 = n17964 & n18104;
  assign n18494 = ~n18080 & ~n18493;
  assign n18495 = n18064 & ~n18494;
  assign n18496 = n18057 & n18106;
  assign n18497 = n18061 & n18103;
  assign n18498 = ~n18496 & ~n18497;
  assign n18499 = ~n18495 & n18498;
  assign n18500 = n18075 & n18099;
  assign n18501 = ~n18092 & ~n18105;
  assign n18502 = ~n18078 & n18501;
  assign n18503 = ~n18057 & ~n18075;
  assign n18504 = ~n18502 & ~n18503;
  assign n18505 = ~n18060 & n18074;
  assign n18506 = ~n18095 & n18505;
  assign n18507 = n18075 & ~n18506;
  assign n18508 = ~n18028 & ~n18071;
  assign n18509 = n18494 & n18508;
  assign n18510 = ~n18106 & n18509;
  assign n18511 = ~n18090 & n18510;
  assign n18512 = n18061 & ~n18511;
  assign n18513 = ~n18507 & ~n18512;
  assign n18514 = n18064 & ~n18093;
  assign n18515 = ~n18064 & n18505;
  assign n18516 = ~n18057 & ~n18073;
  assign n18517 = n18096 & n18516;
  assign n18518 = ~n18066 & n18517;
  assign n18519 = ~n18515 & ~n18518;
  assign n18520 = n18056 & n18519;
  assign n18521 = ~n18514 & ~n18520;
  assign n18522 = n18513 & n18521;
  assign n18523 = n18063 & n18522;
  assign n18524 = ~n18504 & n18523;
  assign n18525 = ~n18500 & n18524;
  assign n18526 = n18499 & n18525;
  assign n18527 = n18526 ^ n14717;
  assign n18528 = n18527 ^ x801;
  assign n18529 = n17177 ^ x796;
  assign n18530 = ~n18528 & n18529;
  assign n18531 = n16483 & n16505;
  assign n18532 = ~n16449 & n16508;
  assign n18533 = ~n18531 & ~n18532;
  assign n18534 = ~n16495 & n16506;
  assign n18535 = n16481 & ~n16522;
  assign n18536 = ~n18534 & ~n18535;
  assign n18537 = n18533 & n18536;
  assign n18538 = n18537 ^ n15407;
  assign n18539 = n18538 ^ x774;
  assign n18540 = n17631 ^ x776;
  assign n18541 = n18539 & ~n18540;
  assign n18542 = ~n16186 & n16217;
  assign n18543 = n16195 & n18542;
  assign n18544 = n15972 & ~n18543;
  assign n18545 = ~n16180 & n16187;
  assign n18546 = ~n16212 & n18545;
  assign n18547 = n16182 & ~n18546;
  assign n18548 = n16194 & ~n17834;
  assign n18549 = n16168 & n16193;
  assign n18550 = ~n16198 & ~n18549;
  assign n18551 = n16188 & n18550;
  assign n18552 = n16171 & ~n18551;
  assign n18553 = n16200 & ~n16208;
  assign n18554 = n16223 & n18553;
  assign n18555 = n16191 & ~n18554;
  assign n18556 = ~n18552 & ~n18555;
  assign n18557 = ~n18548 & n18556;
  assign n18558 = ~n18547 & n18557;
  assign n18559 = ~n18544 & n18558;
  assign n18560 = n16206 & n18559;
  assign n18561 = n17998 & n18560;
  assign n18562 = n16178 & n18561;
  assign n18563 = n18562 ^ n15432;
  assign n18564 = n18563 ^ x775;
  assign n18565 = n18143 ^ x773;
  assign n18566 = n18564 & ~n18565;
  assign n18567 = n18541 & n18566;
  assign n18568 = n18229 ^ x772;
  assign n18569 = n17746 ^ x777;
  assign n18570 = ~n18568 & n18569;
  assign n18571 = ~n18568 & ~n18569;
  assign n18572 = ~n18570 & ~n18571;
  assign n18573 = n18567 & ~n18572;
  assign n18574 = n18568 & n18569;
  assign n18575 = ~n18539 & n18540;
  assign n18576 = ~n18564 & n18565;
  assign n18577 = n18575 & n18576;
  assign n18578 = ~n18539 & ~n18540;
  assign n18579 = n18564 & n18565;
  assign n18580 = n18578 & n18579;
  assign n18581 = ~n18577 & ~n18580;
  assign n18582 = n18574 & ~n18581;
  assign n18583 = ~n18573 & ~n18582;
  assign n18584 = n18566 & n18578;
  assign n18585 = n18570 & n18584;
  assign n18586 = ~n18571 & ~n18574;
  assign n18587 = n18541 & ~n18586;
  assign n18588 = n18576 & n18587;
  assign n18589 = ~n18585 & ~n18588;
  assign n18590 = n18541 & n18579;
  assign n18591 = n18574 & n18590;
  assign n18592 = n18576 & n18578;
  assign n18593 = n18570 & n18592;
  assign n18594 = ~n18591 & ~n18593;
  assign n18595 = n18566 & n18575;
  assign n18596 = n18570 & n18595;
  assign n18597 = n18574 & n18584;
  assign n18598 = ~n18596 & ~n18597;
  assign n18599 = n18539 & n18540;
  assign n18600 = n18566 & n18599;
  assign n18601 = ~n18564 & ~n18565;
  assign n18602 = n18599 & n18601;
  assign n18603 = n18578 & n18601;
  assign n18604 = ~n18602 & ~n18603;
  assign n18605 = ~n18600 & n18604;
  assign n18606 = n18574 & ~n18605;
  assign n18607 = n18575 & n18601;
  assign n18608 = ~n18568 & n18607;
  assign n18609 = n18576 & n18599;
  assign n18610 = ~n18580 & ~n18609;
  assign n18611 = ~n18602 & n18610;
  assign n18612 = n18570 & ~n18611;
  assign n18613 = ~n18608 & ~n18612;
  assign n18614 = ~n18606 & n18613;
  assign n18615 = n18568 & ~n18569;
  assign n18616 = ~n18595 & ~n18603;
  assign n18617 = ~n18609 & n18616;
  assign n18618 = n18564 ^ n18540;
  assign n18619 = n18564 ^ n18539;
  assign n18620 = n18619 ^ n18565;
  assign n18621 = n18618 & n18620;
  assign n18622 = n18617 & ~n18621;
  assign n18623 = ~n18600 & n18622;
  assign n18624 = n18615 & n18623;
  assign n18625 = n18575 & n18579;
  assign n18626 = ~n18621 & ~n18625;
  assign n18627 = n18571 & ~n18626;
  assign n18628 = ~n18624 & ~n18627;
  assign n18629 = n18614 & n18628;
  assign n18630 = n18598 & n18629;
  assign n18631 = n18594 & n18630;
  assign n18632 = n18589 & n18631;
  assign n18633 = n18583 & n18632;
  assign n18634 = n18633 ^ n15542;
  assign n18635 = n18634 ^ x800;
  assign n18636 = n18145 & n18258;
  assign n18637 = ~n18246 & ~n18248;
  assign n18638 = n18235 & ~n18637;
  assign n18639 = ~n18636 & ~n18638;
  assign n18640 = ~n18250 & ~n18261;
  assign n18641 = n18145 & ~n18640;
  assign n18642 = ~n18121 & n18262;
  assign n18643 = ~n18257 & n18283;
  assign n18644 = ~n18642 & ~n18643;
  assign n18645 = n18235 & n18258;
  assign n18646 = ~n18261 & ~n18281;
  assign n18647 = n18256 & ~n18646;
  assign n18648 = ~n18233 & n18251;
  assign n18649 = ~n18254 & ~n18262;
  assign n18650 = n18648 & n18649;
  assign n18651 = n18240 & n18650;
  assign n18652 = ~n18261 & n18651;
  assign n18653 = n18243 & ~n18652;
  assign n18654 = n18276 & n18285;
  assign n18655 = n18235 & ~n18654;
  assign n18656 = n18145 & ~n18270;
  assign n18657 = ~n18269 & ~n18271;
  assign n18658 = n18256 & ~n18657;
  assign n18659 = ~n18656 & ~n18658;
  assign n18660 = ~n18284 & n18659;
  assign n18661 = ~n18239 & n18660;
  assign n18662 = ~n18121 & ~n18661;
  assign n18663 = ~n18655 & ~n18662;
  assign n18664 = ~n18653 & n18663;
  assign n18665 = ~n18647 & n18664;
  assign n18666 = ~n18645 & n18665;
  assign n18667 = n18644 & n18666;
  assign n18668 = ~n18641 & n18667;
  assign n18669 = n18639 & n18668;
  assign n18670 = n18669 ^ n15667;
  assign n18671 = n18670 ^ x799;
  assign n18672 = n18635 & n18671;
  assign n18673 = n17822 & n17913;
  assign n18674 = n17886 & n17916;
  assign n18675 = ~n17850 & n17903;
  assign n18676 = ~n18674 & ~n18675;
  assign n18677 = ~n18673 & n18676;
  assign n18678 = n17911 & ~n18677;
  assign n18679 = ~n17886 & ~n17900;
  assign n18680 = n17886 & n17888;
  assign n18681 = n17822 & ~n17905;
  assign n18682 = ~n18680 & ~n18681;
  assign n18683 = ~n18679 & n18682;
  assign n18684 = n17899 & n18683;
  assign n18685 = ~n18678 & ~n18684;
  assign n18686 = n17850 ^ n17822;
  assign n18687 = n17894 & n18686;
  assign n18688 = n17820 & n18687;
  assign n18689 = n17822 & n17900;
  assign n18690 = n17915 & ~n18689;
  assign n18691 = n17926 & ~n18690;
  assign n18692 = ~n18688 & ~n18691;
  assign n18693 = n17888 & ~n17889;
  assign n18694 = n17890 & n17916;
  assign n18695 = ~n18693 & ~n18694;
  assign n18696 = ~n17850 & n17913;
  assign n18697 = n17851 & n17920;
  assign n18698 = ~n18696 & ~n18697;
  assign n18699 = n18695 & n18698;
  assign n18700 = n17915 & n18699;
  assign n18701 = n17821 & ~n18700;
  assign n18702 = n18692 & ~n18701;
  assign n18703 = n18685 & n18702;
  assign n18704 = n18703 ^ n15341;
  assign n18705 = n18704 ^ x798;
  assign n18706 = n18300 & n18381;
  assign n18707 = ~n18368 & ~n18399;
  assign n18708 = n18355 & ~n18707;
  assign n18709 = ~n18378 & ~n18708;
  assign n18710 = n18367 & n18381;
  assign n18711 = ~n18359 & ~n18710;
  assign n18712 = n18300 & ~n18391;
  assign n18713 = n18372 & ~n18400;
  assign n18714 = ~n18712 & ~n18713;
  assign n18715 = n18362 & n18377;
  assign n18716 = ~n18373 & ~n18382;
  assign n18717 = ~n18368 & n18716;
  assign n18718 = n18367 & ~n18717;
  assign n18719 = ~n18715 & ~n18718;
  assign n18720 = n18364 & n18384;
  assign n18721 = n18355 & ~n18720;
  assign n18722 = ~n18352 & ~n18372;
  assign n18723 = n18299 ^ n18298;
  assign n18724 = ~n18401 & n18723;
  assign n18725 = ~n18722 & ~n18724;
  assign n18726 = ~n18402 & ~n18725;
  assign n18727 = ~n18393 & n18726;
  assign n18728 = ~n18353 & ~n18380;
  assign n18729 = n18299 & n18728;
  assign n18730 = ~n18727 & ~n18729;
  assign n18731 = ~n18721 & ~n18730;
  assign n18732 = n18719 & n18731;
  assign n18733 = n18714 & n18732;
  assign n18734 = n18711 & n18733;
  assign n18735 = n18376 & n18734;
  assign n18736 = n18709 & n18735;
  assign n18737 = ~n18706 & n18736;
  assign n18738 = n18737 ^ n15847;
  assign n18739 = n18738 ^ x797;
  assign n18740 = n18705 & n18739;
  assign n18741 = n18672 & n18740;
  assign n18742 = n18530 & n18741;
  assign n18743 = n18528 & ~n18529;
  assign n18744 = n18635 & ~n18671;
  assign n18745 = ~n18705 & ~n18739;
  assign n18746 = n18744 & n18745;
  assign n18747 = n18743 & n18746;
  assign n18748 = ~n18742 & ~n18747;
  assign n18749 = ~n18530 & ~n18743;
  assign n18750 = n18740 & n18744;
  assign n18751 = n18749 & n18750;
  assign n18752 = ~n18528 & ~n18529;
  assign n18753 = n18705 & ~n18739;
  assign n18754 = n18672 & n18753;
  assign n18755 = ~n18635 & ~n18671;
  assign n18756 = n18753 & n18755;
  assign n18757 = ~n18754 & ~n18756;
  assign n18758 = n18752 & ~n18757;
  assign n18759 = ~n18751 & ~n18758;
  assign n18760 = n18748 & n18759;
  assign n18761 = n18528 & n18529;
  assign n18762 = ~n18635 & n18671;
  assign n18763 = ~n18705 & n18739;
  assign n18764 = n18762 & n18763;
  assign n18765 = ~n18741 & ~n18764;
  assign n18766 = n18761 & ~n18765;
  assign n18767 = n18744 & n18753;
  assign n18768 = n18745 & n18755;
  assign n18769 = ~n18767 & ~n18768;
  assign n18770 = n18743 & ~n18769;
  assign n18771 = ~n18766 & ~n18770;
  assign n18772 = n18753 & n18762;
  assign n18773 = ~n18764 & ~n18772;
  assign n18774 = ~n18529 & ~n18773;
  assign n18775 = n18672 & ~n18705;
  assign n18776 = n18752 & n18775;
  assign n18777 = ~n18774 & ~n18776;
  assign n18778 = n18771 & n18777;
  assign n18779 = n18740 & n18755;
  assign n18780 = n18672 & n18763;
  assign n18781 = n18740 & n18762;
  assign n18782 = ~n18780 & ~n18781;
  assign n18783 = ~n18779 & n18782;
  assign n18784 = ~n18749 & ~n18783;
  assign n18785 = n18744 & n18763;
  assign n18786 = n18749 & n18785;
  assign n18787 = n18755 & n18763;
  assign n18788 = n18745 & n18762;
  assign n18789 = ~n18754 & ~n18788;
  assign n18790 = ~n18787 & n18789;
  assign n18791 = ~n18756 & n18790;
  assign n18792 = n18761 & ~n18791;
  assign n18793 = ~n18746 & n18769;
  assign n18794 = ~n18788 & n18793;
  assign n18795 = n18530 & ~n18794;
  assign n18796 = ~n18792 & ~n18795;
  assign n18797 = ~n18786 & n18796;
  assign n18798 = ~n18784 & n18797;
  assign n18799 = n18778 & n18798;
  assign n18800 = n18760 & n18799;
  assign n18801 = n18800 ^ n15929;
  assign n18802 = n17360 & n17533;
  assign n18803 = n17540 & n17576;
  assign n18804 = ~n17531 & ~n17566;
  assign n18805 = n17526 & ~n18804;
  assign n18806 = ~n18803 & ~n18805;
  assign n18807 = ~n18802 & n18806;
  assign n18808 = ~n17392 & n17553;
  assign n18809 = n17525 & n17540;
  assign n18810 = ~n18808 & ~n18809;
  assign n18811 = n17521 & n17546;
  assign n18812 = ~n17538 & ~n17559;
  assign n18813 = n17533 & ~n18812;
  assign n18814 = ~n18811 & ~n18813;
  assign n18815 = n18810 & n18814;
  assign n18816 = ~n17549 & ~n17559;
  assign n18817 = n17526 & ~n18816;
  assign n18818 = ~n17360 & ~n17573;
  assign n18819 = n17556 & ~n18818;
  assign n18820 = n17533 & n17555;
  assign n18821 = n17533 & n17566;
  assign n18822 = n17562 & ~n17573;
  assign n18823 = ~n17538 & n18822;
  assign n18824 = n17526 & ~n18823;
  assign n18825 = n17330 ^ n17200;
  assign n18826 = n18825 ^ n17358;
  assign n18827 = n17233 & n18826;
  assign n18828 = n17556 & n18827;
  assign n18829 = ~n18824 & ~n18828;
  assign n18830 = ~n18821 & n18829;
  assign n18831 = ~n18820 & n18830;
  assign n18832 = ~n17534 & n18831;
  assign n18833 = ~n18819 & n18832;
  assign n18834 = ~n18817 & n18833;
  assign n18835 = n18815 & n18834;
  assign n18836 = n18807 & n18835;
  assign n18837 = n18836 ^ n16971;
  assign n18838 = n18743 & n18756;
  assign n18839 = ~n18779 & ~n18785;
  assign n18840 = n18530 & ~n18839;
  assign n18841 = ~n18838 & ~n18840;
  assign n18842 = ~n18529 & n18767;
  assign n18843 = n18743 & n18788;
  assign n18844 = ~n18842 & ~n18843;
  assign n18845 = n18746 & n18752;
  assign n18846 = n18782 & ~n18787;
  assign n18847 = n18749 & ~n18846;
  assign n18848 = ~n18845 & ~n18847;
  assign n18849 = n18844 & n18848;
  assign n18850 = n18530 & n18764;
  assign n18851 = n18671 ^ n18635;
  assign n18852 = n18745 & ~n18851;
  assign n18853 = ~n18756 & ~n18852;
  assign n18854 = ~n18754 & n18853;
  assign n18855 = n18761 & ~n18854;
  assign n18856 = ~n18772 & ~n18787;
  assign n18857 = n18765 & n18856;
  assign n18858 = ~n18530 & n18857;
  assign n18859 = ~n18772 & n18789;
  assign n18860 = ~n18746 & n18859;
  assign n18861 = ~n18743 & n18860;
  assign n18862 = ~n18858 & ~n18861;
  assign n18863 = ~n18749 & n18862;
  assign n18864 = ~n18855 & ~n18863;
  assign n18865 = ~n18850 & n18864;
  assign n18866 = n18849 & n18865;
  assign n18867 = n18841 & n18866;
  assign n18868 = n18760 & n18867;
  assign n18869 = n18868 ^ n18229;
  assign n18870 = ~n18609 & ~n18625;
  assign n18871 = n18570 & ~n18870;
  assign n18872 = n18541 & n18601;
  assign n18873 = n18574 & n18872;
  assign n18874 = n18571 & n18623;
  assign n18875 = ~n18607 & n18617;
  assign n18876 = n18581 & n18875;
  assign n18877 = n18574 & ~n18876;
  assign n18878 = ~n18874 & ~n18877;
  assign n18879 = ~n18584 & ~n18590;
  assign n18880 = n18605 & n18879;
  assign n18881 = n18570 & ~n18880;
  assign n18882 = ~n18607 & ~n18872;
  assign n18883 = n18626 & n18882;
  assign n18884 = ~n18592 & n18883;
  assign n18885 = n18615 & ~n18884;
  assign n18886 = ~n18881 & ~n18885;
  assign n18887 = n18878 & n18886;
  assign n18888 = ~n18873 & n18887;
  assign n18889 = n18594 & n18888;
  assign n18890 = ~n18871 & n18889;
  assign n18891 = n18890 ^ n15996;
  assign n18892 = n18837 ^ x820;
  assign n18893 = n18239 & n18256;
  assign n18894 = ~n18656 & ~n18893;
  assign n18895 = ~n18144 & n18275;
  assign n18896 = n18256 & ~n18270;
  assign n18897 = ~n18895 & ~n18896;
  assign n18898 = ~n18257 & n18284;
  assign n18899 = n18144 ^ n18121;
  assign n18900 = ~n18281 & ~n18283;
  assign n18901 = ~n18899 & ~n18900;
  assign n18902 = ~n18254 & n18648;
  assign n18903 = ~n18271 & n18902;
  assign n18904 = ~n18258 & n18903;
  assign n18905 = n18243 & ~n18904;
  assign n18906 = n18264 & ~n18269;
  assign n18907 = n18235 & ~n18906;
  assign n18908 = n18252 & ~n18262;
  assign n18909 = n18256 & ~n18908;
  assign n18910 = ~n18907 & ~n18909;
  assign n18911 = ~n18905 & n18910;
  assign n18912 = ~n18641 & n18911;
  assign n18913 = ~n18901 & n18912;
  assign n18914 = ~n18898 & n18913;
  assign n18915 = n18897 & n18914;
  assign n18916 = n18894 & n18915;
  assign n18917 = n18242 & n18916;
  assign n18918 = n18917 ^ n16132;
  assign n18919 = n18918 ^ x825;
  assign n18920 = n18892 & n18919;
  assign n18921 = n17897 & n17926;
  assign n18922 = ~n17908 & n17911;
  assign n18923 = ~n18921 & ~n18922;
  assign n18924 = n17899 & ~n17924;
  assign n18925 = n17821 & ~n17933;
  assign n18926 = ~n18924 & ~n18925;
  assign n18927 = n18923 & n18926;
  assign n18928 = n18927 ^ n17248;
  assign n18929 = n18928 ^ x822;
  assign n18930 = n17122 & n17135;
  assign n18931 = n17109 & n17145;
  assign n18932 = ~n18930 & ~n18931;
  assign n18933 = n16241 & n17138;
  assign n18934 = n17109 & n17171;
  assign n18935 = ~n18933 & ~n18934;
  assign n18936 = n17109 & n17119;
  assign n18937 = n16241 & ~n17162;
  assign n18938 = ~n18936 & ~n18937;
  assign n18939 = ~n17117 & ~n17157;
  assign n18940 = ~n17121 & ~n17135;
  assign n18941 = n18939 & n18940;
  assign n18942 = n16241 & ~n18941;
  assign n18943 = n17143 & ~n17146;
  assign n18944 = ~n17117 & n18943;
  assign n18945 = n17122 & ~n18944;
  assign n18946 = ~n18942 & ~n18945;
  assign n18947 = ~n17141 & ~n17161;
  assign n18948 = ~n17111 & n18947;
  assign n18949 = n17131 & ~n18948;
  assign n18950 = n17109 & n17135;
  assign n18951 = ~n17127 & ~n17130;
  assign n18952 = n17122 & ~n18951;
  assign n18953 = ~n18950 & ~n18952;
  assign n18954 = ~n17132 & n17157;
  assign n18955 = ~n17138 & ~n17146;
  assign n18956 = ~n17121 & n18955;
  assign n18957 = ~n15930 & ~n18956;
  assign n18958 = ~n18954 & ~n18957;
  assign n18959 = n18953 & n18958;
  assign n18960 = ~n18949 & n18959;
  assign n18961 = n18946 & n18960;
  assign n18962 = n18938 & n18961;
  assign n18963 = n18935 & n18962;
  assign n18964 = n18932 & n18963;
  assign n18965 = n17114 & n18964;
  assign n18966 = n18965 ^ n16919;
  assign n18967 = n18966 ^ x821;
  assign n18968 = ~n18929 & n18967;
  assign n18969 = n18057 & n18092;
  assign n18970 = n18061 & n18493;
  assign n18971 = ~n18969 & ~n18970;
  assign n18972 = ~n18028 & ~n18073;
  assign n18973 = ~n18095 & n18972;
  assign n18974 = n18064 & ~n18973;
  assign n18975 = ~n18066 & ~n18103;
  assign n18976 = ~n18503 & ~n18975;
  assign n18977 = ~n18090 & ~n18099;
  assign n18978 = n18081 & n18977;
  assign n18979 = n18075 & ~n18978;
  assign n18980 = n18074 & n18096;
  assign n18981 = n18061 & ~n18980;
  assign n18982 = ~n18979 & ~n18981;
  assign n18983 = ~n18976 & n18982;
  assign n18984 = ~n18064 & n18977;
  assign n18985 = ~n18092 & ~n18493;
  assign n18986 = ~n18057 & n18985;
  assign n18987 = ~n18984 & ~n18986;
  assign n18988 = n18107 & ~n18987;
  assign n18989 = n18056 & ~n18988;
  assign n18990 = n18983 & ~n18989;
  assign n18991 = ~n18974 & n18990;
  assign n18992 = n18971 & n18991;
  assign n18993 = ~n18065 & n18992;
  assign n18994 = n18083 & n18993;
  assign n18995 = n18063 & n18994;
  assign n18996 = n18995 ^ n15970;
  assign n18997 = n18996 ^ x824;
  assign n18998 = n18968 & n18997;
  assign n18999 = n17633 & n17758;
  assign n19000 = n17755 & n17797;
  assign n19001 = ~n18999 & ~n19000;
  assign n19002 = n17763 & n17777;
  assign n19003 = n17755 & n17798;
  assign n19004 = ~n19002 & ~n19003;
  assign n19005 = n17777 & n17778;
  assign n19006 = ~n17788 & n17802;
  assign n19007 = ~n17793 & n19006;
  assign n19008 = ~n17752 & n19007;
  assign n19009 = n17633 & ~n19008;
  assign n19010 = ~n19005 & ~n19009;
  assign n19011 = ~n17769 & n17775;
  assign n19012 = n17764 & n17780;
  assign n19013 = n17755 & ~n19012;
  assign n19014 = ~n17752 & n17800;
  assign n19015 = ~n17783 & n19014;
  assign n19016 = n17753 & ~n17771;
  assign n19017 = ~n17790 & n19016;
  assign n19018 = ~n17777 & n19017;
  assign n19019 = ~n19015 & ~n19018;
  assign n19020 = n17785 & ~n19019;
  assign n19021 = n17632 & ~n19020;
  assign n19022 = ~n19013 & ~n19021;
  assign n19023 = ~n19011 & n19022;
  assign n19024 = n19010 & n19023;
  assign n19025 = n19004 & n19024;
  assign n19026 = n17774 & n19025;
  assign n19027 = n19001 & n19026;
  assign n19028 = n19027 ^ n17272;
  assign n19029 = n19028 ^ x823;
  assign n19030 = n18998 & ~n19029;
  assign n19031 = n18920 & n19030;
  assign n19032 = ~n18892 & n18919;
  assign n19033 = ~n18929 & ~n18967;
  assign n19034 = n18997 & n19033;
  assign n19035 = n19029 & n19034;
  assign n19036 = n19032 & n19035;
  assign n19037 = n18892 & ~n18919;
  assign n19038 = n18929 & ~n18967;
  assign n19039 = n18997 & n19038;
  assign n19040 = ~n19029 & n19039;
  assign n19041 = n19037 & n19040;
  assign n19042 = ~n19036 & ~n19041;
  assign n19043 = ~n19031 & n19042;
  assign n19044 = ~n18997 & n19029;
  assign n19045 = n18968 & n19044;
  assign n19046 = n18920 & n19045;
  assign n19047 = n18929 & n18967;
  assign n19048 = n19044 & n19047;
  assign n19049 = n18997 & n19047;
  assign n19050 = ~n19029 & n19049;
  assign n19051 = ~n19048 & ~n19050;
  assign n19052 = n18920 & ~n19051;
  assign n19053 = ~n18997 & ~n19029;
  assign n19054 = n19047 & n19053;
  assign n19055 = ~n19030 & ~n19054;
  assign n19056 = n19032 & ~n19055;
  assign n19057 = ~n19052 & ~n19056;
  assign n19058 = ~n19046 & n19057;
  assign n19059 = n19038 & n19053;
  assign n19060 = n18920 & n19059;
  assign n19061 = n19038 & n19044;
  assign n19062 = ~n19029 & n19034;
  assign n19063 = ~n19061 & ~n19062;
  assign n19064 = n19032 & ~n19063;
  assign n19065 = ~n19060 & ~n19064;
  assign n19066 = n19032 & n19059;
  assign n19067 = ~n18892 & ~n18919;
  assign n19068 = n19029 & n19039;
  assign n19069 = ~n19062 & ~n19068;
  assign n19070 = ~n19030 & ~n19045;
  assign n19071 = ~n19061 & n19070;
  assign n19072 = ~n19050 & n19071;
  assign n19073 = n19069 & n19072;
  assign n19074 = ~n19035 & n19073;
  assign n19075 = ~n19059 & n19074;
  assign n19076 = n19067 & n19075;
  assign n19077 = ~n19066 & ~n19076;
  assign n19078 = n18919 ^ n18892;
  assign n19079 = n19029 & n19049;
  assign n19080 = ~n19045 & ~n19079;
  assign n19081 = n19078 & ~n19080;
  assign n19082 = n19033 & n19053;
  assign n19083 = ~n19054 & ~n19082;
  assign n19084 = n19063 & n19083;
  assign n19085 = ~n19050 & n19084;
  assign n19086 = n19037 & ~n19085;
  assign n19087 = ~n19039 & ~n19082;
  assign n19088 = n18920 & n19087;
  assign n19089 = n19088 ^ n18920;
  assign n19090 = ~n19086 & ~n19089;
  assign n19091 = ~n19081 & n19090;
  assign n19092 = n19077 & n19091;
  assign n19093 = n19065 & n19092;
  assign n19094 = n19058 & n19093;
  assign n19095 = n19043 & n19094;
  assign n19096 = n19095 ^ n17654;
  assign n19097 = n18570 & n18577;
  assign n19098 = n18571 & ~n18604;
  assign n19099 = ~n19097 & ~n19098;
  assign n19100 = n18579 & n18599;
  assign n19101 = n18574 & n19100;
  assign n19102 = n18609 & n18615;
  assign n19103 = ~n19101 & ~n19102;
  assign n19104 = n18571 & n18595;
  assign n19105 = n18581 & ~n18584;
  assign n19106 = n18615 & ~n19105;
  assign n19107 = ~n19104 & ~n19106;
  assign n19108 = n18574 & ~n18610;
  assign n19109 = ~n18590 & ~n18609;
  assign n19110 = n18570 & ~n19109;
  assign n19111 = ~n18590 & ~n18625;
  assign n19112 = ~n19100 & n19111;
  assign n19113 = ~n18592 & n19112;
  assign n19114 = n18571 & ~n19113;
  assign n19115 = ~n18567 & ~n18595;
  assign n19116 = n18604 & n19115;
  assign n19117 = n18574 & ~n19116;
  assign n19118 = ~n19114 & ~n19117;
  assign n19119 = n18567 & ~n18571;
  assign n19120 = ~n18600 & n18882;
  assign n19121 = n18586 & ~n19120;
  assign n19122 = ~n19119 & ~n19121;
  assign n19123 = n19118 & n19122;
  assign n19124 = ~n19110 & n19123;
  assign n19125 = ~n19108 & n19124;
  assign n19126 = n19107 & n19125;
  assign n19127 = n19103 & n19126;
  assign n19128 = n19099 & n19127;
  assign n19129 = n18589 & n19128;
  assign n19130 = n19129 ^ n16771;
  assign n19131 = n19033 & n19044;
  assign n19132 = ~n19040 & ~n19131;
  assign n19133 = n19032 & ~n19132;
  assign n19134 = ~n18920 & ~n19067;
  assign n19135 = n18968 & n19053;
  assign n19136 = ~n19134 & n19135;
  assign n19137 = n19067 & ~n19080;
  assign n19138 = ~n19136 & ~n19137;
  assign n19139 = ~n19133 & n19138;
  assign n19140 = n19059 & n19067;
  assign n19141 = n19029 ^ n18919;
  assign n19142 = n18998 & ~n19141;
  assign n19143 = n18892 & n19142;
  assign n19144 = ~n19140 & ~n19143;
  assign n19145 = n18998 & n19029;
  assign n19146 = n19067 & n19145;
  assign n19147 = n19037 & n19061;
  assign n19148 = ~n19146 & ~n19147;
  assign n19149 = n19054 & n19067;
  assign n19150 = ~n19069 & ~n19134;
  assign n19151 = ~n19149 & ~n19150;
  assign n19152 = n19037 & ~n19051;
  assign n19153 = n19032 & ~n19072;
  assign n19154 = ~n19152 & ~n19153;
  assign n19155 = ~n19048 & ~n19131;
  assign n19156 = ~n19059 & n19155;
  assign n19157 = n18920 & ~n19156;
  assign n19158 = ~n19035 & ~n19131;
  assign n19159 = n19037 & ~n19158;
  assign n19160 = ~n19082 & ~n19159;
  assign n19161 = n19134 & ~n19160;
  assign n19162 = ~n19157 & ~n19161;
  assign n19163 = n19154 & n19162;
  assign n19164 = n19151 & n19163;
  assign n19165 = n19148 & n19164;
  assign n19166 = n19144 & n19165;
  assign n19167 = n19043 & n19166;
  assign n19168 = n19139 & n19167;
  assign n19169 = n19168 ^ n17992;
  assign n19170 = n17632 & n17798;
  assign n19171 = n17633 & n17783;
  assign n19172 = ~n19170 & ~n19171;
  assign n19173 = n17777 & ~n17794;
  assign n19174 = ~n17778 & n17785;
  assign n19175 = ~n17768 & n19174;
  assign n19176 = n17755 & ~n19175;
  assign n19177 = ~n19173 & ~n19176;
  assign n19178 = n19172 & n19177;
  assign n19179 = n17632 ^ n17603;
  assign n19180 = n17797 & ~n19179;
  assign n19181 = ~n17752 & n17802;
  assign n19182 = n17775 & ~n19181;
  assign n19183 = n17767 & ~n19179;
  assign n19184 = ~n17758 & ~n17763;
  assign n19185 = ~n17788 & n19184;
  assign n19186 = ~n17768 & n19185;
  assign n19187 = n17775 & ~n19186;
  assign n19188 = ~n19183 & ~n19187;
  assign n19189 = n17633 & n17760;
  assign n19190 = n17764 & ~n17779;
  assign n19191 = n17777 & ~n19190;
  assign n19192 = n17753 & ~n17783;
  assign n19193 = n17755 & ~n19192;
  assign n19194 = ~n19191 & ~n19193;
  assign n19195 = ~n19189 & n19194;
  assign n19196 = n19188 & n19195;
  assign n19197 = n19001 & n19196;
  assign n19198 = ~n19182 & n19197;
  assign n19199 = ~n19180 & n19198;
  assign n19200 = n19178 & n19199;
  assign n19201 = ~n17754 & n19200;
  assign n19202 = n19201 ^ n16363;
  assign n19203 = n17899 & ~n18677;
  assign n19204 = n17926 & n18700;
  assign n19205 = ~n19203 & ~n19204;
  assign n19206 = n17821 & ~n18690;
  assign n19207 = n17911 & ~n18683;
  assign n19208 = ~n19206 & ~n19207;
  assign n19209 = n19205 & n19208;
  assign n19210 = ~n18687 & n19209;
  assign n19211 = n19210 ^ n15939;
  assign n19212 = n19211 ^ x831;
  assign n19213 = n18996 ^ x826;
  assign n19214 = n19212 & n19213;
  assign n19215 = ~n17546 & ~n17565;
  assign n19216 = ~n17525 & n19215;
  assign n19217 = n17540 & ~n19216;
  assign n19218 = n17555 & ~n17560;
  assign n19219 = ~n17530 & ~n17576;
  assign n19220 = n17526 & ~n19219;
  assign n19221 = n17577 & n17579;
  assign n19222 = n17533 & ~n19221;
  assign n19223 = ~n19220 & ~n19222;
  assign n19224 = ~n19218 & n19223;
  assign n19225 = n17540 & n17559;
  assign n19226 = ~n17565 & n18804;
  assign n19227 = ~n17553 & n19226;
  assign n19228 = ~n17549 & n19227;
  assign n19229 = n17521 & ~n19228;
  assign n19230 = ~n19225 & ~n19229;
  assign n19231 = n19224 & n19230;
  assign n19232 = n17552 & n19231;
  assign n19233 = ~n17544 & n19232;
  assign n19234 = ~n19217 & n19233;
  assign n19235 = n18807 & n19234;
  assign n19236 = ~n18820 & n19235;
  assign n19237 = n17528 & n19236;
  assign n19238 = ~n17538 & n19237;
  assign n19239 = n19238 ^ n16098;
  assign n19240 = n19239 ^ x828;
  assign n19241 = n18918 ^ x827;
  assign n19242 = ~n19240 & ~n19241;
  assign n19243 = n18891 ^ x830;
  assign n19244 = n18299 & n18369;
  assign n19245 = n18300 & n18393;
  assign n19246 = n18352 & n18372;
  assign n19247 = ~n19245 & ~n19246;
  assign n19248 = ~n19244 & n19247;
  assign n19249 = n18298 & n18358;
  assign n19250 = n18300 & ~n18400;
  assign n19251 = ~n19249 & ~n19250;
  assign n19252 = ~n18363 & n18403;
  assign n19253 = ~n18383 & n19252;
  assign n19254 = ~n18373 & n19253;
  assign n19255 = n18355 & ~n19254;
  assign n19256 = n18364 & n18394;
  assign n19257 = n18367 & ~n19256;
  assign n19258 = n18404 & n18716;
  assign n19259 = n18372 & ~n19258;
  assign n19260 = ~n19257 & ~n19259;
  assign n19261 = ~n19255 & n19260;
  assign n19262 = n19251 & n19261;
  assign n19263 = n18711 & n19262;
  assign n19264 = n19248 & n19263;
  assign n19265 = ~n18371 & n19264;
  assign n19266 = n18354 & n19265;
  assign n19267 = ~n18706 & n19266;
  assign n19268 = n19267 ^ n16166;
  assign n19269 = n19268 ^ x829;
  assign n19270 = ~n19243 & ~n19269;
  assign n19271 = n19242 & n19270;
  assign n19272 = n19214 & n19271;
  assign n19273 = ~n19212 & n19213;
  assign n19274 = ~n19240 & n19241;
  assign n19275 = n19243 & ~n19269;
  assign n19276 = n19274 & n19275;
  assign n19277 = n19273 & n19276;
  assign n19278 = ~n19212 & ~n19213;
  assign n19279 = n19242 & n19275;
  assign n19280 = n19240 & ~n19241;
  assign n19281 = n19270 & n19280;
  assign n19282 = ~n19279 & ~n19281;
  assign n19283 = n19278 & ~n19282;
  assign n19284 = ~n19277 & ~n19283;
  assign n19285 = ~n19272 & n19284;
  assign n19286 = ~n19243 & n19269;
  assign n19287 = n19274 & n19286;
  assign n19288 = n19273 & n19287;
  assign n19289 = n19212 & ~n19213;
  assign n19290 = n19281 & n19289;
  assign n19291 = ~n19288 & ~n19290;
  assign n19292 = n19240 & n19241;
  assign n19293 = n19269 ^ n19243;
  assign n19294 = n19292 & ~n19293;
  assign n19295 = n19214 & n19294;
  assign n19296 = n19291 & ~n19295;
  assign n19297 = n19287 & n19289;
  assign n19298 = n19271 & n19273;
  assign n19299 = ~n19297 & ~n19298;
  assign n19300 = n19243 & n19269;
  assign n19301 = n19292 & n19300;
  assign n19302 = ~n19287 & ~n19301;
  assign n19303 = n19278 & ~n19302;
  assign n19304 = n19280 & n19300;
  assign n19305 = n19273 & n19304;
  assign n19306 = n19286 & n19292;
  assign n19307 = n19214 & n19306;
  assign n19308 = ~n19305 & ~n19307;
  assign n19309 = n19275 & n19280;
  assign n19310 = n19289 & n19309;
  assign n19311 = ~n19214 & ~n19278;
  assign n19312 = n19270 & n19274;
  assign n19313 = ~n19311 & n19312;
  assign n19314 = ~n19269 & n19292;
  assign n19315 = n19280 & n19286;
  assign n19316 = ~n19279 & ~n19315;
  assign n19317 = ~n19314 & n19316;
  assign n19318 = n19273 & ~n19317;
  assign n19319 = ~n19313 & ~n19318;
  assign n19320 = n19274 & n19300;
  assign n19321 = ~n19213 & n19320;
  assign n19322 = n19243 & n19292;
  assign n19323 = n19316 & ~n19322;
  assign n19324 = n19289 & ~n19323;
  assign n19325 = ~n19309 & ~n19315;
  assign n19326 = ~n19214 & n19325;
  assign n19327 = n19242 & n19286;
  assign n19328 = n19242 & n19300;
  assign n19329 = ~n19309 & ~n19328;
  assign n19330 = ~n19327 & n19329;
  assign n19331 = ~n19278 & n19330;
  assign n19332 = ~n19326 & ~n19331;
  assign n19333 = ~n19311 & n19332;
  assign n19334 = ~n19324 & ~n19333;
  assign n19335 = ~n19321 & n19334;
  assign n19336 = n19319 & n19335;
  assign n19337 = ~n19310 & n19336;
  assign n19338 = n19308 & n19337;
  assign n19339 = ~n19303 & n19338;
  assign n19340 = n19299 & n19339;
  assign n19341 = n19296 & n19340;
  assign n19342 = n19285 & n19341;
  assign n19343 = n19342 ^ n17849;
  assign n19344 = n18355 & ~n18395;
  assign n19345 = n18298 & ~n18716;
  assign n19346 = ~n19344 & ~n19345;
  assign n19347 = ~n18348 & n18707;
  assign n19348 = ~n18380 & n19347;
  assign n19349 = ~n18393 & n19348;
  assign n19350 = n18372 & ~n19349;
  assign n19351 = n18391 & n19254;
  assign n19352 = n18367 & ~n19351;
  assign n19353 = ~n19350 & ~n19352;
  assign n19354 = n19346 & n19353;
  assign n19355 = n19248 & n19354;
  assign n19356 = n18366 & n19355;
  assign n19357 = n18709 & n19356;
  assign n19358 = ~n18706 & n19357;
  assign n19359 = n19358 ^ n17025;
  assign n19360 = n18891 ^ x784;
  assign n19361 = n17632 & n17768;
  assign n19362 = n17755 & ~n19006;
  assign n19363 = ~n19361 & ~n19362;
  assign n19364 = ~n17798 & n19016;
  assign n19365 = n17777 & ~n19364;
  assign n19366 = n17764 & ~n17771;
  assign n19367 = ~n17790 & n19366;
  assign n19368 = ~n17768 & n19367;
  assign n19369 = n17633 & ~n19368;
  assign n19370 = ~n17779 & n17794;
  assign n19371 = ~n17788 & n19370;
  assign n19372 = ~n17798 & n19371;
  assign n19373 = ~n17790 & n19372;
  assign n19374 = n17775 & ~n19373;
  assign n19375 = ~n19369 & ~n19374;
  assign n19376 = ~n19365 & n19375;
  assign n19377 = n19363 & n19376;
  assign n19378 = n17782 & n19377;
  assign n19379 = n19004 & n19378;
  assign n19380 = ~n17766 & n19379;
  assign n19381 = ~n17754 & n19380;
  assign n19382 = n19001 & n19381;
  assign n19383 = n19382 ^ n16662;
  assign n19384 = n19383 ^ x789;
  assign n19385 = ~n19360 & n19384;
  assign n19386 = n19211 ^ x785;
  assign n19387 = n17107 & n17109;
  assign n19388 = ~n17112 & ~n17117;
  assign n19389 = n16241 & ~n19388;
  assign n19390 = ~n19387 & ~n19389;
  assign n19391 = n17107 & n17122;
  assign n19392 = ~n17132 & ~n17162;
  assign n19393 = ~n19391 & ~n19392;
  assign n19394 = ~n17130 & ~n17157;
  assign n19395 = n16241 & ~n19394;
  assign n19396 = ~n17142 & ~n17146;
  assign n19397 = n17109 & ~n19396;
  assign n19398 = ~n19395 & ~n19397;
  assign n19399 = ~n17119 & ~n17138;
  assign n19400 = n17131 & ~n19399;
  assign n19401 = n17112 & n17122;
  assign n19402 = n17109 & ~n18939;
  assign n19403 = ~n19401 & ~n19402;
  assign n19404 = ~n17127 & n18940;
  assign n19405 = n17131 & ~n19404;
  assign n19406 = n16241 & ~n17152;
  assign n19407 = ~n19405 & ~n19406;
  assign n19408 = n19403 & n19407;
  assign n19409 = n18953 & n19408;
  assign n19410 = n18935 & n19409;
  assign n19411 = ~n17173 & n19410;
  assign n19412 = ~n19400 & n19411;
  assign n19413 = n19398 & n19412;
  assign n19414 = n19393 & n19413;
  assign n19415 = n19390 & n19414;
  assign n19416 = n18932 & n19415;
  assign n19417 = n19416 ^ n16622;
  assign n19418 = n19417 ^ x787;
  assign n19419 = n19386 & ~n19418;
  assign n19420 = ~n18121 & n18246;
  assign n19421 = ~n18257 & n18261;
  assign n19422 = ~n19420 & ~n19421;
  assign n19423 = n18235 & n18250;
  assign n19424 = ~n18250 & n18286;
  assign n19425 = n18270 & n19424;
  assign n19426 = n18243 & ~n19425;
  assign n19427 = n18145 & ~n18649;
  assign n19428 = ~n18239 & n18276;
  assign n19429 = ~n18262 & n19428;
  assign n19430 = n18235 & ~n19429;
  assign n19431 = ~n18248 & ~n18275;
  assign n19432 = ~n18233 & n19431;
  assign n19433 = ~n18283 & n19432;
  assign n19434 = ~n18284 & n19433;
  assign n19435 = n18256 & ~n19434;
  assign n19436 = ~n19430 & ~n19435;
  assign n19437 = ~n19427 & n19436;
  assign n19438 = n18894 & n19437;
  assign n19439 = ~n19426 & n19438;
  assign n19440 = ~n19423 & n19439;
  assign n19441 = n19422 & n19440;
  assign n19442 = n18639 & n19441;
  assign n19443 = ~n18901 & n19442;
  assign n19444 = n19443 ^ n16588;
  assign n19445 = n19444 ^ x788;
  assign n19446 = n18064 & n18092;
  assign n19447 = n18057 & n18493;
  assign n19448 = ~n19446 & ~n19447;
  assign n19449 = n18099 & ~n18503;
  assign n19450 = n18056 & n18078;
  assign n19451 = ~n18073 & ~n18087;
  assign n19452 = ~n18103 & n19451;
  assign n19453 = n18057 & ~n19452;
  assign n19454 = n18505 & n18977;
  assign n19455 = ~n18078 & n19454;
  assign n19456 = n18061 & ~n19455;
  assign n19457 = ~n19453 & ~n19456;
  assign n19458 = ~n18066 & n18093;
  assign n19459 = n18075 & ~n19458;
  assign n19460 = ~n18066 & n18508;
  assign n19461 = ~n18075 & n19460;
  assign n19462 = n18096 & n18972;
  assign n19463 = n18075 & ~n19462;
  assign n19464 = ~n18064 & ~n19463;
  assign n19465 = ~n19461 & ~n19464;
  assign n19466 = ~n19459 & ~n19465;
  assign n19467 = n19457 & n19466;
  assign n19468 = ~n18058 & n19467;
  assign n19469 = n18068 & n19468;
  assign n19470 = ~n19450 & n19469;
  assign n19471 = ~n19449 & n19470;
  assign n19472 = n19448 & n19471;
  assign n19473 = n18499 & n19472;
  assign n19474 = n19473 ^ n16556;
  assign n19475 = n19474 ^ x786;
  assign n19476 = ~n19445 & n19475;
  assign n19477 = n19419 & n19476;
  assign n19478 = n19385 & n19477;
  assign n19479 = n19360 & n19384;
  assign n19480 = ~n19386 & ~n19418;
  assign n19481 = n19445 & n19475;
  assign n19482 = n19480 & n19481;
  assign n19483 = ~n19386 & n19418;
  assign n19484 = ~n19445 & ~n19475;
  assign n19485 = n19483 & n19484;
  assign n19486 = ~n19482 & ~n19485;
  assign n19487 = n19479 & ~n19486;
  assign n19488 = ~n19478 & ~n19487;
  assign n19489 = n19476 & n19480;
  assign n19490 = n19479 & n19489;
  assign n19491 = n19445 & ~n19475;
  assign n19492 = n19480 & n19491;
  assign n19493 = ~n19384 & n19492;
  assign n19494 = ~n19490 & ~n19493;
  assign n19495 = n19479 & n19492;
  assign n19496 = n19483 & n19491;
  assign n19497 = ~n19384 & n19496;
  assign n19498 = ~n19495 & ~n19497;
  assign n19499 = ~n19360 & ~n19384;
  assign n19500 = n19481 & n19483;
  assign n19501 = n19419 & n19481;
  assign n19502 = n19386 & n19418;
  assign n19503 = n19475 ^ n19445;
  assign n19504 = n19502 & n19503;
  assign n19505 = ~n19477 & ~n19504;
  assign n19506 = ~n19501 & n19505;
  assign n19507 = ~n19485 & n19506;
  assign n19508 = ~n19500 & n19507;
  assign n19509 = n19499 & ~n19508;
  assign n19510 = n19360 & ~n19384;
  assign n19511 = n19476 & n19502;
  assign n19512 = n19480 & n19484;
  assign n19513 = n19419 & n19491;
  assign n19514 = n19481 & n19502;
  assign n19515 = n19484 & n19502;
  assign n19516 = ~n19514 & ~n19515;
  assign n19517 = ~n19513 & n19516;
  assign n19518 = ~n19512 & n19517;
  assign n19519 = ~n19489 & n19518;
  assign n19520 = ~n19511 & n19519;
  assign n19521 = n19510 & ~n19520;
  assign n19522 = ~n19509 & ~n19521;
  assign n19523 = ~n19501 & n19516;
  assign n19524 = n19385 & ~n19523;
  assign n19525 = n19419 & n19484;
  assign n19526 = n19476 & n19483;
  assign n19527 = ~n19501 & ~n19514;
  assign n19528 = ~n19526 & n19527;
  assign n19529 = ~n19525 & n19528;
  assign n19530 = ~n19385 & n19529;
  assign n19531 = ~n19496 & ~n19526;
  assign n19532 = ~n19500 & n19531;
  assign n19533 = ~n19512 & n19532;
  assign n19534 = n19385 & ~n19533;
  assign n19535 = ~n19479 & ~n19534;
  assign n19536 = ~n19530 & ~n19535;
  assign n19537 = ~n19524 & ~n19536;
  assign n19538 = n19522 & n19537;
  assign n19539 = n19498 & n19538;
  assign n19540 = n19494 & n19539;
  assign n19541 = n19488 & n19540;
  assign n19542 = n19541 ^ n18201;
  assign n19543 = n19479 & n19525;
  assign n19544 = n19385 & n19485;
  assign n19545 = ~n19543 & ~n19544;
  assign n19546 = n19385 & n19500;
  assign n19547 = n19499 & n19525;
  assign n19548 = ~n19546 & ~n19547;
  assign n19549 = ~n19384 & n19477;
  assign n19550 = n19483 ^ n19481;
  assign n19551 = n19499 & n19550;
  assign n19552 = ~n19549 & ~n19551;
  assign n19553 = ~n19504 & ~n19515;
  assign n19554 = n19510 & ~n19553;
  assign n19555 = n19506 & ~n19526;
  assign n19556 = ~n19492 & n19555;
  assign n19557 = n19385 & ~n19556;
  assign n19558 = ~n19554 & ~n19557;
  assign n19559 = n19552 & n19558;
  assign n19560 = n19479 & ~n19517;
  assign n19561 = ~n19482 & ~n19512;
  assign n19562 = ~n19526 & n19561;
  assign n19563 = ~n19510 & n19562;
  assign n19564 = ~n19489 & ~n19492;
  assign n19565 = ~n19525 & n19564;
  assign n19566 = ~n19479 & n19565;
  assign n19567 = ~n19563 & ~n19566;
  assign n19568 = ~n19500 & ~n19567;
  assign n19569 = n19360 & ~n19568;
  assign n19570 = ~n19560 & ~n19569;
  assign n19571 = n19559 & n19570;
  assign n19572 = n19548 & n19571;
  assign n19573 = n19545 & n19572;
  assign n19574 = n19573 ^ n17687;
  assign n19575 = n17521 & n17538;
  assign n19576 = n17577 & n19226;
  assign n19577 = n17526 & ~n19576;
  assign n19578 = ~n19575 & ~n19577;
  assign n19579 = n17556 & ~n17579;
  assign n19580 = ~n17525 & ~n17576;
  assign n19581 = n17533 & ~n19580;
  assign n19582 = ~n17546 & n18816;
  assign n19583 = ~n17392 & ~n19582;
  assign n19584 = ~n19581 & ~n19583;
  assign n19585 = ~n19579 & n19584;
  assign n19586 = n19578 & n19585;
  assign n19587 = n17542 & n19586;
  assign n19588 = n17558 & n19587;
  assign n19589 = ~n19217 & n19588;
  assign n19590 = ~n18820 & n19589;
  assign n19591 = ~n17534 & n19590;
  assign n19592 = n17528 & n19591;
  assign n19593 = n19592 ^ n16795;
  assign n19594 = n18769 & n18789;
  assign n19595 = ~n18750 & n19594;
  assign n19596 = n18761 & ~n19595;
  assign n19597 = ~n18780 & n18839;
  assign n19598 = n18749 & ~n19597;
  assign n19599 = n18745 ^ n18740;
  assign n19600 = ~n18851 & n19599;
  assign n19601 = n19600 ^ n18740;
  assign n19602 = n18765 & ~n19601;
  assign n19603 = n18743 & ~n19602;
  assign n19604 = ~n19598 & ~n19603;
  assign n19605 = ~n19596 & n19604;
  assign n19606 = ~n18752 & ~n18852;
  assign n19607 = ~n18530 & n18789;
  assign n19608 = ~n19606 & ~n19607;
  assign n19609 = n18856 & ~n19608;
  assign n19610 = ~n18767 & n19609;
  assign n19611 = ~n18528 & ~n19610;
  assign n19612 = n19605 & ~n19611;
  assign n19613 = n18841 & n19612;
  assign n19614 = n18748 & n19613;
  assign n19615 = n19614 ^ n17963;
  assign n19616 = ~n17132 & ~n18955;
  assign n19617 = ~n17130 & n18947;
  assign n19618 = n17122 & ~n19617;
  assign n19619 = ~n17127 & ~n17145;
  assign n19620 = n16241 & ~n19619;
  assign n19621 = ~n19618 & ~n19620;
  assign n19622 = ~n19616 & n19621;
  assign n19623 = n17109 & ~n18951;
  assign n19624 = ~n17142 & n18941;
  assign n19625 = ~n17145 & n19624;
  assign n19626 = n17131 & ~n19625;
  assign n19627 = ~n19623 & ~n19626;
  assign n19628 = n19622 & n19627;
  assign n19629 = n17171 & n19628;
  assign n19630 = ~n16240 & n19629;
  assign n19631 = n19630 ^ n19628;
  assign n19632 = n18938 & n19631;
  assign n19633 = n19390 & n19632;
  assign n19634 = n17125 & n19633;
  assign n19635 = n18932 & n19634;
  assign n19636 = n17114 & n19635;
  assign n19637 = n19636 ^ n16436;
  assign n19638 = n18421 & n18448;
  assign n19639 = n17818 & ~n18427;
  assign n19640 = ~n19638 & ~n19639;
  assign n19641 = ~n18419 & ~n18454;
  assign n19642 = n18421 & ~n19641;
  assign n19643 = n18421 & n18432;
  assign n19644 = ~n18423 & ~n18449;
  assign n19645 = ~n18457 & n19644;
  assign n19646 = n18459 & ~n19645;
  assign n19647 = ~n19643 & ~n19646;
  assign n19648 = ~n18436 & n18462;
  assign n19649 = ~n17817 & n18442;
  assign n19650 = ~n19648 & ~n19649;
  assign n19651 = ~n18441 & ~n18476;
  assign n19652 = n17818 & ~n19651;
  assign n19653 = ~n18446 & ~n18471;
  assign n19654 = ~n18470 & n19653;
  assign n19655 = ~n18426 & n19654;
  assign n19656 = n18459 & ~n19655;
  assign n19657 = n18472 & ~n18476;
  assign n19658 = ~n18438 & n19657;
  assign n19659 = n18434 & ~n19658;
  assign n19660 = ~n19656 & ~n19659;
  assign n19661 = ~n19652 & n19660;
  assign n19662 = n19650 & n19661;
  assign n19663 = n19647 & n19662;
  assign n19664 = ~n19642 & n19663;
  assign n19665 = n18456 & n19664;
  assign n19666 = n18452 & n19665;
  assign n19667 = n19640 & n19666;
  assign n19668 = ~n18433 & n19667;
  assign n19669 = n18429 & n19668;
  assign n19670 = n19669 ^ n17885;
  assign n19671 = ~n18572 & n18600;
  assign n19672 = ~n18592 & ~n18602;
  assign n19673 = ~n18595 & n19672;
  assign n19674 = n18574 & ~n19673;
  assign n19675 = ~n19671 & ~n19674;
  assign n19676 = n18581 & ~n19100;
  assign n19677 = n18571 & ~n19676;
  assign n19678 = n18541 & n18576;
  assign n19679 = ~n18574 & n19678;
  assign n19680 = n19111 & n19115;
  assign n19681 = ~n18607 & n19680;
  assign n19682 = ~n18584 & n19681;
  assign n19683 = n18615 & ~n19682;
  assign n19684 = ~n19679 & ~n19683;
  assign n19685 = ~n19677 & n19684;
  assign n19686 = n19675 & n19685;
  assign n19687 = ~n18593 & n19686;
  assign n19688 = n18598 & n19687;
  assign n19689 = ~n18873 & n19688;
  assign n19690 = n19103 & n19689;
  assign n19691 = n19099 & n19690;
  assign n19692 = ~n18871 & n19691;
  assign n19693 = n18583 & n19692;
  assign n19694 = n19693 ^ n16994;
  assign n19695 = n19032 & n19049;
  assign n19696 = ~n19131 & ~n19135;
  assign n19697 = n19051 & n19696;
  assign n19698 = ~n19034 & n19697;
  assign n19699 = n19067 & ~n19698;
  assign n19700 = n19037 & ~n19080;
  assign n19701 = ~n19068 & n19696;
  assign n19702 = n19078 & ~n19701;
  assign n19703 = n19069 & n19083;
  assign n19704 = ~n19061 & n19703;
  assign n19705 = n18920 & ~n19704;
  assign n19706 = ~n19702 & ~n19705;
  assign n19707 = ~n19700 & n19706;
  assign n19708 = ~n19699 & n19707;
  assign n19709 = ~n19695 & n19708;
  assign n19710 = n19042 & n19709;
  assign n19711 = n19148 & n19710;
  assign n19712 = n19144 & n19711;
  assign n19713 = n19057 & n19712;
  assign n19714 = n19713 ^ n18177;
  assign n19715 = n18765 & ~n18785;
  assign n19716 = n18752 & ~n19715;
  assign n19717 = ~n18754 & n19597;
  assign n19718 = n18530 & ~n19717;
  assign n19719 = ~n19716 & ~n19718;
  assign n19720 = ~n18767 & ~n18852;
  assign n19721 = ~n18788 & n19720;
  assign n19722 = n18743 & ~n19721;
  assign n19723 = ~n18741 & n18856;
  assign n19724 = n18761 & ~n19723;
  assign n19725 = ~n18788 & n18853;
  assign n19726 = n18530 & ~n19725;
  assign n19727 = n18761 & ~n19721;
  assign n19728 = ~n19726 & ~n19727;
  assign n19729 = n18765 & n18839;
  assign n19730 = n18743 & ~n19729;
  assign n19731 = ~n18746 & n18790;
  assign n19732 = n18752 & ~n19731;
  assign n19733 = ~n19730 & ~n19732;
  assign n19734 = n19728 & n19733;
  assign n19735 = ~n19724 & n19734;
  assign n19736 = ~n19722 & n19735;
  assign n19737 = n19719 & n19736;
  assign n19738 = ~n18751 & n19737;
  assign n19739 = n19738 ^ n17721;
  assign n19740 = n19289 & n19294;
  assign n19741 = ~n19304 & ~n19328;
  assign n19742 = n19273 & ~n19741;
  assign n19743 = ~n19310 & ~n19742;
  assign n19744 = n19214 & n19279;
  assign n19745 = n19271 & n19289;
  assign n19746 = n19275 & n19292;
  assign n19747 = ~n19312 & ~n19746;
  assign n19748 = n19273 & ~n19747;
  assign n19749 = ~n19745 & ~n19748;
  assign n19750 = ~n19744 & n19749;
  assign n19751 = n19278 & n19328;
  assign n19752 = n19273 & n19327;
  assign n19753 = n19214 & n19281;
  assign n19754 = ~n19752 & ~n19753;
  assign n19755 = ~n19751 & n19754;
  assign n19756 = ~n19213 & n19304;
  assign n19757 = n19273 & n19306;
  assign n19758 = ~n19756 & ~n19757;
  assign n19759 = ~n19306 & ~n19320;
  assign n19760 = ~n19328 & n19759;
  assign n19761 = n19214 & ~n19760;
  assign n19762 = ~n19311 & n19314;
  assign n19763 = ~n19276 & ~n19315;
  assign n19764 = n19289 & ~n19763;
  assign n19765 = ~n19762 & ~n19764;
  assign n19766 = ~n19761 & n19765;
  assign n19767 = n19758 & n19766;
  assign n19768 = ~n19303 & n19767;
  assign n19769 = n19299 & n19768;
  assign n19770 = n19755 & n19769;
  assign n19771 = n19750 & n19770;
  assign n19772 = n19743 & n19771;
  assign n19773 = ~n19740 & n19772;
  assign n19774 = n19285 & n19773;
  assign n19775 = n19774 ^ n18023;
  assign n19776 = n19593 ^ x792;
  assign n19777 = n19130 ^ x793;
  assign n19778 = n17177 ^ x794;
  assign n19779 = n19383 ^ x791;
  assign n19780 = n19778 & n19779;
  assign n19781 = ~n19777 & n19780;
  assign n19782 = ~n19776 & n19781;
  assign n19783 = n19444 ^ x790;
  assign n19784 = n18738 ^ x795;
  assign n19785 = ~n19783 & n19784;
  assign n19786 = n19782 & n19785;
  assign n19787 = n19776 & n19777;
  assign n19788 = ~n19779 & n19787;
  assign n19789 = n19778 & n19788;
  assign n19790 = n19783 & n19784;
  assign n19791 = n19789 & n19790;
  assign n19792 = ~n19786 & ~n19791;
  assign n19793 = n19780 & n19787;
  assign n19794 = n19785 & n19793;
  assign n19795 = ~n19783 & ~n19784;
  assign n19796 = n19789 & n19795;
  assign n19797 = n19783 & ~n19784;
  assign n19798 = ~n19777 & ~n19779;
  assign n19799 = ~n19776 & n19798;
  assign n19800 = ~n19778 & n19799;
  assign n19801 = n19776 & n19798;
  assign n19802 = n19778 & n19801;
  assign n19803 = ~n19800 & ~n19802;
  assign n19804 = n19797 & ~n19803;
  assign n19805 = ~n19796 & ~n19804;
  assign n19806 = ~n19794 & n19805;
  assign n19807 = n19778 & n19799;
  assign n19808 = n19795 & n19807;
  assign n19809 = ~n19776 & n19777;
  assign n19810 = ~n19779 & n19809;
  assign n19811 = ~n19778 & n19810;
  assign n19812 = ~n19789 & ~n19811;
  assign n19813 = n19797 & ~n19812;
  assign n19814 = ~n19808 & ~n19813;
  assign n19815 = n19778 & n19810;
  assign n19816 = n19790 & n19815;
  assign n19817 = ~n19778 & n19779;
  assign n19818 = n19809 & n19817;
  assign n19819 = ~n19777 & n19817;
  assign n19820 = n19776 & n19819;
  assign n19821 = ~n19818 & ~n19820;
  assign n19822 = n19785 & ~n19821;
  assign n19823 = n19776 & n19781;
  assign n19824 = n19797 & n19823;
  assign n19825 = n19785 & ~n19803;
  assign n19826 = ~n19824 & ~n19825;
  assign n19827 = n19787 & n19817;
  assign n19828 = ~n19818 & ~n19823;
  assign n19829 = ~n19782 & n19828;
  assign n19830 = ~n19827 & n19829;
  assign n19831 = n19795 & ~n19830;
  assign n19832 = ~n19820 & n19829;
  assign n19833 = n19790 & ~n19832;
  assign n19834 = ~n19831 & ~n19833;
  assign n19835 = n19785 & n19810;
  assign n19836 = ~n19776 & n19819;
  assign n19837 = n19780 & n19809;
  assign n19838 = ~n19827 & ~n19837;
  assign n19839 = ~n19836 & n19838;
  assign n19840 = n19797 & ~n19839;
  assign n19841 = ~n19778 & n19788;
  assign n19842 = ~n19778 & n19801;
  assign n19843 = ~n19841 & ~n19842;
  assign n19844 = ~n19785 & ~n19797;
  assign n19845 = ~n19843 & n19844;
  assign n19846 = ~n19840 & ~n19845;
  assign n19847 = ~n19835 & n19846;
  assign n19848 = n19834 & n19847;
  assign n19849 = n19826 & n19848;
  assign n19850 = ~n19822 & n19849;
  assign n19851 = ~n19816 & n19850;
  assign n19852 = n19814 & n19851;
  assign n19853 = n19806 & n19852;
  assign n19854 = n19792 & n19853;
  assign n19855 = n19854 ^ n17391;
  assign n19856 = n19273 & n19301;
  assign n19857 = ~n19320 & n19325;
  assign n19858 = n19214 & ~n19857;
  assign n19859 = ~n19856 & ~n19858;
  assign n19860 = n19278 & ~n19759;
  assign n19861 = ~n19213 & ~n19747;
  assign n19862 = ~n19860 & ~n19861;
  assign n19863 = n19214 & n19276;
  assign n19864 = ~n19311 & n19327;
  assign n19865 = ~n19863 & ~n19864;
  assign n19866 = ~n19287 & n19741;
  assign n19867 = n19289 & ~n19866;
  assign n19868 = ~n19312 & n19325;
  assign n19869 = n19273 & ~n19868;
  assign n19870 = ~n19867 & ~n19869;
  assign n19871 = n19865 & n19870;
  assign n19872 = n19862 & n19871;
  assign n19873 = n19308 & n19872;
  assign n19874 = n19291 & n19873;
  assign n19875 = n19755 & n19874;
  assign n19876 = n19859 & n19875;
  assign n19877 = ~n19740 & n19876;
  assign n19878 = n19285 & n19877;
  assign n19879 = n19878 ^ n16239;
  assign n19880 = n17937 ^ x814;
  assign n19881 = n18966 ^ x819;
  assign n19882 = n19880 & n19881;
  assign n19883 = ~n19880 & ~n19881;
  assign n19884 = ~n19882 & ~n19883;
  assign n19885 = n19694 ^ x816;
  assign n19886 = n18837 ^ x818;
  assign n19887 = n19359 ^ x817;
  assign n19888 = n17816 ^ x815;
  assign n19889 = ~n19887 & ~n19888;
  assign n19890 = n19886 & n19889;
  assign n19891 = ~n19885 & n19890;
  assign n19892 = ~n19884 & n19891;
  assign n19893 = n19880 & ~n19881;
  assign n19894 = ~n19885 & ~n19886;
  assign n19895 = n19889 & n19894;
  assign n19896 = n19893 & n19895;
  assign n19897 = ~n19880 & n19881;
  assign n19898 = n19885 & ~n19886;
  assign n19899 = n19887 & n19888;
  assign n19900 = n19898 & n19899;
  assign n19901 = ~n19887 & n19888;
  assign n19902 = n19886 & n19901;
  assign n19903 = n19885 & n19902;
  assign n19904 = ~n19900 & ~n19903;
  assign n19905 = n19897 & ~n19904;
  assign n19906 = ~n19896 & ~n19905;
  assign n19907 = ~n19892 & n19906;
  assign n19908 = n19887 & ~n19888;
  assign n19909 = n19894 & n19908;
  assign n19910 = ~n19884 & n19909;
  assign n19911 = n19886 & n19908;
  assign n19912 = ~n19885 & n19911;
  assign n19913 = ~n19895 & ~n19912;
  assign n19914 = n19897 & ~n19913;
  assign n19915 = ~n19910 & ~n19914;
  assign n19916 = n19886 ^ n19885;
  assign n19917 = n19901 & n19916;
  assign n19918 = n19897 & n19917;
  assign n19919 = n19889 & n19898;
  assign n19920 = n19885 & n19911;
  assign n19921 = ~n19919 & ~n19920;
  assign n19922 = n19893 & ~n19921;
  assign n19923 = ~n19918 & ~n19922;
  assign n19924 = n19885 & n19890;
  assign n19925 = ~n19881 & n19924;
  assign n19926 = n19886 & n19899;
  assign n19927 = n19885 & n19926;
  assign n19928 = n19898 & n19908;
  assign n19929 = ~n19927 & ~n19928;
  assign n19930 = n19897 & ~n19929;
  assign n19931 = ~n19925 & ~n19930;
  assign n19932 = ~n19884 & ~n19921;
  assign n19933 = n19894 & n19901;
  assign n19934 = n19894 & n19899;
  assign n19935 = ~n19927 & ~n19934;
  assign n19936 = ~n19933 & n19935;
  assign n19937 = n19883 & ~n19936;
  assign n19938 = n19888 & n19916;
  assign n19939 = ~n19882 & ~n19938;
  assign n19940 = n19904 & ~n19933;
  assign n19941 = ~n19934 & n19940;
  assign n19942 = ~n19893 & n19941;
  assign n19943 = ~n19939 & ~n19942;
  assign n19944 = n19880 & n19943;
  assign n19945 = ~n19937 & ~n19944;
  assign n19946 = ~n19932 & n19945;
  assign n19947 = n19931 & n19946;
  assign n19948 = n19923 & n19947;
  assign n19949 = n19915 & n19948;
  assign n19950 = n19907 & n19949;
  assign n19951 = n19950 ^ n17746;
  assign n19952 = n19897 & n19900;
  assign n19953 = ~n19884 & n19890;
  assign n19954 = ~n19952 & ~n19953;
  assign n19955 = n19883 & n19928;
  assign n19956 = n19893 & n19912;
  assign n19957 = ~n19955 & ~n19956;
  assign n19958 = n19954 & n19957;
  assign n19959 = ~n19882 & n19933;
  assign n19960 = ~n19895 & ~n19909;
  assign n19961 = n19882 & ~n19960;
  assign n19962 = n19883 & ~n19904;
  assign n19963 = ~n19885 & n19926;
  assign n19964 = ~n19934 & ~n19963;
  assign n19965 = ~n19884 & ~n19964;
  assign n19966 = n19898 & n19901;
  assign n19967 = ~n19903 & ~n19966;
  assign n19968 = n19882 & ~n19967;
  assign n19969 = ~n19965 & ~n19968;
  assign n19970 = ~n19962 & n19969;
  assign n19971 = ~n19917 & n19935;
  assign n19972 = n19893 & ~n19971;
  assign n19973 = ~n19909 & n19921;
  assign n19974 = ~n19912 & n19973;
  assign n19975 = n19897 & ~n19974;
  assign n19976 = ~n19972 & ~n19975;
  assign n19977 = n19970 & n19976;
  assign n19978 = ~n19961 & n19977;
  assign n19979 = ~n19959 & n19978;
  assign n19980 = n19958 & n19979;
  assign n19981 = n19923 & n19980;
  assign n19982 = n19981 ^ n18055;
  assign n19983 = n18920 & n19035;
  assign n19984 = ~n19063 & ~n19134;
  assign n19985 = ~n19983 & ~n19984;
  assign n19986 = ~n19048 & ~n19068;
  assign n19987 = n19032 & ~n19986;
  assign n19988 = ~n19050 & n19132;
  assign n19989 = n19067 & ~n19988;
  assign n19990 = ~n19987 & ~n19989;
  assign n19991 = n19037 & n19075;
  assign n19992 = n19990 & ~n19991;
  assign n19993 = n19985 & n19992;
  assign n19994 = n19065 & n19993;
  assign n19995 = n19058 & n19994;
  assign n19996 = n19139 & n19995;
  assign n19997 = n19996 ^ n17329;
  assign n19998 = n18634 ^ x802;
  assign n19999 = n18416 ^ x807;
  assign n20000 = ~n19998 & n19999;
  assign n20001 = n17591 ^ x806;
  assign n20002 = n19202 ^ x805;
  assign n20003 = n20001 & ~n20002;
  assign n20004 = n18527 ^ x803;
  assign n20005 = n19637 ^ x804;
  assign n20006 = ~n20004 & ~n20005;
  assign n20007 = n20003 & n20006;
  assign n20008 = ~n20001 & n20002;
  assign n20009 = n20008 ^ n20005;
  assign n20010 = n20009 ^ n20002;
  assign n20011 = n20009 ^ n20008;
  assign n20012 = n20010 & n20011;
  assign n20013 = ~n20004 & n20012;
  assign n20014 = n20013 ^ n20009;
  assign n20015 = ~n20007 & ~n20014;
  assign n20016 = n20000 & ~n20015;
  assign n20017 = ~n19998 & ~n19999;
  assign n20018 = n20005 ^ n20004;
  assign n20019 = n20005 ^ n20002;
  assign n20020 = n20018 & n20019;
  assign n20021 = n20001 & n20020;
  assign n20022 = n20021 ^ n20018;
  assign n20023 = n20002 ^ n20001;
  assign n20024 = n20004 ^ n20002;
  assign n20025 = ~n20018 & n20024;
  assign n20026 = ~n20023 & n20025;
  assign n20027 = ~n20022 & ~n20026;
  assign n20028 = n20017 & ~n20027;
  assign n20029 = ~n20016 & ~n20028;
  assign n20030 = n19998 & ~n19999;
  assign n20032 = ~n20001 & ~n20002;
  assign n20033 = n20001 & n20002;
  assign n20034 = ~n20032 & ~n20033;
  assign n20031 = n20005 ^ n20003;
  assign n20035 = n20034 ^ n20031;
  assign n20036 = ~n20004 & ~n20035;
  assign n20037 = n20036 ^ n20034;
  assign n20038 = n20030 & n20037;
  assign n20039 = n19998 & n19999;
  assign n20040 = ~n20004 & n20005;
  assign n20041 = n20001 & n20040;
  assign n20042 = n20004 & ~n20005;
  assign n20043 = n20033 & n20042;
  assign n20044 = ~n20041 & ~n20043;
  assign n20045 = n20004 & n20005;
  assign n20046 = n20045 ^ n20002;
  assign n20047 = ~n20006 & n20046;
  assign n20048 = ~n20001 & n20047;
  assign n20049 = n20048 ^ n20001;
  assign n20050 = n20044 & n20049;
  assign n20051 = n20039 & ~n20050;
  assign n20052 = ~n20038 & ~n20051;
  assign n20053 = n20029 & n20052;
  assign n20054 = n20053 ^ n16526;
  assign n20055 = n19795 & ~n19828;
  assign n20056 = n19790 & n19820;
  assign n20057 = n19785 & n19841;
  assign n20058 = n19782 & n19797;
  assign n20059 = ~n20057 & ~n20058;
  assign n20060 = ~n20056 & n20059;
  assign n20061 = ~n20055 & n20060;
  assign n20062 = ~n19793 & ~n19836;
  assign n20063 = n19844 & ~n20062;
  assign n20064 = ~n19815 & ~n19842;
  assign n20065 = ~n19807 & ~n19811;
  assign n20066 = n20064 & n20065;
  assign n20067 = n19790 & ~n20066;
  assign n20068 = ~n20063 & ~n20067;
  assign n20069 = ~n19820 & ~n19827;
  assign n20070 = n19797 & ~n20069;
  assign n20071 = n19828 & n19838;
  assign n20072 = n19785 & ~n20071;
  assign n20073 = n19778 ^ n19777;
  assign n20074 = ~n19779 & ~n20073;
  assign n20075 = n19797 & n20074;
  assign n20076 = ~n19841 & n20065;
  assign n20077 = ~n19802 & n20076;
  assign n20078 = n19795 & ~n20077;
  assign n20079 = ~n20075 & ~n20078;
  assign n20080 = ~n20072 & n20079;
  assign n20081 = ~n20070 & n20080;
  assign n20082 = n20068 & n20081;
  assign n20083 = n20061 & n20082;
  assign n20084 = n19826 & n20083;
  assign n20085 = n19792 & n20084;
  assign n20086 = n20085 ^ n17631;
  assign n20087 = ~n17817 & n18462;
  assign n20088 = ~n18450 & n18459;
  assign n20089 = ~n20087 & ~n20088;
  assign n20090 = ~n18433 & n20089;
  assign n20091 = ~n18457 & n19653;
  assign n20092 = n18421 & ~n20091;
  assign n20093 = ~n18448 & n18477;
  assign n20094 = ~n18419 & n20093;
  assign n20095 = n18434 & ~n20094;
  assign n20096 = ~n20092 & ~n20095;
  assign n20097 = ~n17817 & n18432;
  assign n20098 = ~n18442 & ~n18470;
  assign n20099 = n17818 & ~n20098;
  assign n20100 = ~n18441 & n18478;
  assign n20101 = n18459 & ~n20100;
  assign n20102 = ~n20099 & ~n20101;
  assign n20103 = ~n20097 & n20102;
  assign n20104 = n20096 & n20103;
  assign n20105 = ~n18444 & n20104;
  assign n20106 = n18465 & n20105;
  assign n20107 = n18461 & n20106;
  assign n20108 = n20090 & n20107;
  assign n20109 = n19640 & n20108;
  assign n20110 = n18429 & n20109;
  assign n20111 = n20110 ^ n18342;
  assign n20112 = ~n19891 & ~n19919;
  assign n20113 = n19897 & ~n20112;
  assign n20114 = n19880 & n19891;
  assign n20115 = ~n19933 & ~n19963;
  assign n20116 = ~n19920 & n20115;
  assign n20117 = ~n19917 & n20116;
  assign n20118 = n19882 & ~n20117;
  assign n20119 = ~n20114 & ~n20118;
  assign n20120 = ~n19884 & n19928;
  assign n20121 = n19893 & ~n19973;
  assign n20122 = ~n20120 & ~n20121;
  assign n20123 = n20119 & n20122;
  assign n20124 = n19904 & n20115;
  assign n20125 = n19897 & ~n20124;
  assign n20126 = ~n19912 & ~n19924;
  assign n20127 = n19883 & ~n20126;
  assign n20128 = ~n19883 & n20115;
  assign n20129 = ~n19927 & n20128;
  assign n20130 = ~n19900 & n20129;
  assign n20131 = ~n19893 & ~n19902;
  assign n20132 = ~n20124 & ~n20131;
  assign n20133 = n19935 & ~n20132;
  assign n20134 = ~n19966 & n20133;
  assign n20135 = ~n20130 & ~n20134;
  assign n20136 = ~n19881 & n20135;
  assign n20137 = ~n20127 & ~n20136;
  assign n20138 = ~n20125 & n20137;
  assign n20139 = n20123 & n20138;
  assign n20140 = n19915 & n20139;
  assign n20141 = ~n20113 & n20140;
  assign n20142 = n20141 ^ n17357;
  assign n20143 = n19897 & n19934;
  assign n20144 = ~n19884 & n19919;
  assign n20145 = ~n20143 & ~n20144;
  assign n20146 = ~n19881 & n19912;
  assign n20147 = ~n19909 & ~n19920;
  assign n20148 = n19893 & ~n20147;
  assign n20149 = ~n20146 & ~n20148;
  assign n20150 = n20145 & n20149;
  assign n20151 = ~n19880 & n19902;
  assign n20152 = ~n19924 & ~n19928;
  assign n20153 = n19882 & ~n20152;
  assign n20154 = ~n19920 & ~n19928;
  assign n20155 = n19897 & ~n20154;
  assign n20156 = n19940 & ~n19966;
  assign n20157 = n19893 & ~n20156;
  assign n20158 = ~n19882 & n19904;
  assign n20159 = ~n20128 & ~n20158;
  assign n20160 = n19935 & ~n20159;
  assign n20161 = ~n19884 & ~n20160;
  assign n20162 = ~n20157 & ~n20161;
  assign n20163 = ~n20155 & n20162;
  assign n20164 = ~n20113 & n20163;
  assign n20165 = ~n20153 & n20164;
  assign n20166 = ~n20151 & n20165;
  assign n20167 = n20150 & n20166;
  assign n20168 = n19907 & n20167;
  assign n20169 = n20168 ^ n17104;
  assign n20170 = n19289 & ~n19760;
  assign n20171 = n19273 & ~n19282;
  assign n20172 = ~n20170 & ~n20171;
  assign n20173 = n19287 & ~n19311;
  assign n20174 = n19316 & n19747;
  assign n20175 = ~n19304 & n20174;
  assign n20176 = ~n19327 & n20175;
  assign n20177 = ~n19276 & n20176;
  assign n20178 = n19278 & ~n20177;
  assign n20179 = ~n20173 & ~n20178;
  assign n20180 = n20172 & n20179;
  assign n20181 = ~n19272 & n20180;
  assign n20182 = n19296 & n20181;
  assign n20183 = n19750 & n20182;
  assign n20184 = n19859 & n20183;
  assign n20185 = n19743 & n20184;
  assign n20186 = ~n19740 & n20185;
  assign n20187 = n20186 ^ n18563;
  assign n20188 = n19785 & ~n20065;
  assign n20189 = n19836 & ~n19844;
  assign n20190 = ~n20188 & ~n20189;
  assign n20191 = n19790 & n19793;
  assign n20192 = n19797 & ~n19821;
  assign n20193 = ~n19823 & ~n19837;
  assign n20194 = n19844 & ~n20193;
  assign n20195 = n19785 & ~n19829;
  assign n20196 = ~n20194 & ~n20195;
  assign n20197 = n19795 & ~n20069;
  assign n20206 = n19788 & n19797;
  assign n20198 = ~n19811 & ~n19836;
  assign n20199 = ~n19790 & n20198;
  assign n20200 = ~n19800 & ~n19815;
  assign n20201 = ~n19841 & n20200;
  assign n20202 = ~n19795 & n20201;
  assign n20203 = ~n20199 & ~n20202;
  assign n20204 = ~n19807 & ~n20203;
  assign n20205 = n19844 & ~n20204;
  assign n20207 = n20206 ^ n20205;
  assign n20208 = ~n20197 & ~n20207;
  assign n20209 = n20196 & n20208;
  assign n20210 = n19806 & n20209;
  assign n20211 = ~n20192 & n20210;
  assign n20212 = ~n20191 & n20211;
  assign n20213 = n20190 & n20212;
  assign n20214 = n20060 & n20213;
  assign n20215 = n20214 ^ n18321;
  assign n20216 = ~n20005 & n20008;
  assign n20217 = n20003 & n20004;
  assign n20218 = ~n20216 & ~n20217;
  assign n20219 = ~n20041 & n20218;
  assign n20220 = n20005 & ~n20024;
  assign n20221 = ~n20001 & n20220;
  assign n20222 = n20219 & ~n20221;
  assign n20223 = n20000 & ~n20222;
  assign n20224 = ~n20032 & n20045;
  assign n20225 = ~n20004 & n20032;
  assign n20226 = ~n20005 & n20033;
  assign n20227 = ~n20225 & ~n20226;
  assign n20228 = ~n20007 & n20227;
  assign n20229 = ~n20224 & n20228;
  assign n20230 = n20039 & ~n20229;
  assign n20231 = ~n20223 & ~n20230;
  assign n20233 = n20008 & n20040;
  assign n20232 = n20004 & ~n20031;
  assign n20234 = n20233 ^ n20232;
  assign n20235 = ~n20221 & ~n20234;
  assign n20236 = ~n20007 & n20235;
  assign n20237 = n20017 & n20236;
  assign n20238 = n20003 & n20042;
  assign n20239 = n20002 & n20006;
  assign n20240 = n20005 & ~n20034;
  assign n20241 = ~n20239 & ~n20240;
  assign n20242 = ~n20238 & n20241;
  assign n20243 = ~n20221 & n20242;
  assign n20244 = n20030 & n20243;
  assign n20245 = ~n20237 & ~n20244;
  assign n20246 = n20231 & n20245;
  assign n20247 = n20246 ^ n17199;
  assign n20248 = ~n19793 & ~n19820;
  assign n20249 = n19795 & ~n20248;
  assign n20250 = ~n19782 & n19838;
  assign n20251 = n19790 & ~n20250;
  assign n20252 = ~n20249 & ~n20251;
  assign n20253 = ~n19818 & n19838;
  assign n20254 = n19797 & ~n20253;
  assign n20255 = n19797 & n19798;
  assign n20256 = n19790 & ~n20076;
  assign n20257 = ~n20255 & ~n20256;
  assign n20258 = n19812 & n20064;
  assign n20259 = n19795 & ~n20258;
  assign n20260 = ~n19802 & n19812;
  assign n20261 = ~n19837 & n20260;
  assign n20262 = ~n19819 & n20261;
  assign n20263 = n19785 & ~n20262;
  assign n20264 = ~n20259 & ~n20263;
  assign n20265 = n20257 & n20264;
  assign n20266 = n19792 & n20265;
  assign n20267 = ~n20254 & n20266;
  assign n20268 = n20252 & n20267;
  assign n20269 = n20061 & n20268;
  assign n20270 = n20269 ^ n16871;
  assign n20271 = n20000 & n20027;
  assign n20272 = ~n20015 & n20017;
  assign n20273 = ~n20271 & ~n20272;
  assign n20274 = n20030 & ~n20050;
  assign n20275 = ~n20037 & n20039;
  assign n20276 = ~n20274 & ~n20275;
  assign n20277 = n20273 & n20276;
  assign n20278 = n20277 ^ n18538;
  assign n20279 = n20001 & n20045;
  assign n20280 = n20228 & ~n20279;
  assign n20281 = n20030 & ~n20280;
  assign n20282 = n20000 & ~n20236;
  assign n20283 = ~n20281 & ~n20282;
  assign n20284 = n20017 & ~n20219;
  assign n20285 = n20039 & ~n20243;
  assign n20286 = ~n20284 & ~n20285;
  assign n20287 = n20283 & n20286;
  assign n20288 = ~n20221 & n20287;
  assign n20289 = n20288 ^ n17602;
  assign n20290 = n19385 & ~n19561;
  assign n20291 = n19548 & ~n20290;
  assign n20292 = n19489 & n19499;
  assign n20293 = n19479 & ~n19531;
  assign n20294 = ~n20292 & ~n20293;
  assign n20295 = ~n19477 & n19516;
  assign n20296 = n19499 & ~n20295;
  assign n20297 = n19510 & ~n19562;
  assign n20298 = ~n19360 & n19496;
  assign n20299 = ~n19501 & ~n19513;
  assign n20300 = n19385 & ~n20299;
  assign n20301 = ~n20298 & ~n20300;
  assign n20302 = ~n19500 & ~n19515;
  assign n20303 = ~n19501 & n20302;
  assign n20304 = n19479 & ~n20303;
  assign n20305 = ~n19510 & ~n19511;
  assign n20306 = ~n19504 & ~n19514;
  assign n20307 = ~n19477 & n20306;
  assign n20308 = ~n20305 & ~n20307;
  assign n20309 = ~n20304 & ~n20308;
  assign n20310 = n20301 & n20309;
  assign n20311 = ~n20297 & n20310;
  assign n20312 = ~n20296 & n20311;
  assign n20313 = n19494 & n20312;
  assign n20314 = n19545 & n20313;
  assign n20315 = n20294 & n20314;
  assign n20316 = n20291 & n20315;
  assign n20317 = n20316 ^ n17232;
  assign n20318 = n19492 & n19510;
  assign n20319 = ~n19525 & n20306;
  assign n20320 = n19385 & ~n20319;
  assign n20321 = ~n19384 & ~n19532;
  assign n20322 = n19501 & n19510;
  assign n20323 = ~n19479 & ~n20322;
  assign n20324 = ~n19515 & n20299;
  assign n20325 = ~n20323 & ~n20324;
  assign n20326 = ~n20321 & ~n20325;
  assign n20327 = ~n19511 & n20299;
  assign n20328 = n19499 & ~n20327;
  assign n20329 = n19477 & n19479;
  assign n20330 = ~n19510 & ~n20329;
  assign n20331 = ~n20295 & ~n20330;
  assign n20332 = ~n20328 & ~n20331;
  assign n20333 = n20326 & n20332;
  assign n20334 = ~n20320 & n20333;
  assign n20335 = ~n20318 & n20334;
  assign n20336 = n20294 & n20335;
  assign n20337 = n19488 & n20336;
  assign n20338 = n20291 & n20337;
  assign n20339 = n20338 ^ n16732;
  assign n20340 = ~n18436 & n18457;
  assign n20341 = ~n18426 & n18472;
  assign n20342 = n18450 & n20341;
  assign n20343 = n18421 & ~n20342;
  assign n20344 = ~n20340 & ~n20343;
  assign n20345 = n18434 & ~n19653;
  assign n20346 = ~n18419 & n19657;
  assign n20347 = n18459 & ~n20346;
  assign n20348 = n18479 & n19645;
  assign n20349 = n17818 & ~n20348;
  assign n20350 = ~n20347 & ~n20349;
  assign n20351 = ~n20345 & n20350;
  assign n20352 = n20344 & n20351;
  assign n20353 = ~n19642 & n20352;
  assign n20354 = n18445 & n20353;
  assign n20355 = n20090 & n20354;
  assign n20356 = n20355 ^ n18143;
  assign y0 = n17177;
  assign y1 = n18492;
  assign y2 = n17591;
  assign y3 = n18801;
  assign y4 = n18837;
  assign y5 = n18869;
  assign y6 = n18891;
  assign y7 = n19096;
  assign y8 = n19130;
  assign y9 = n19169;
  assign y10 = n19202;
  assign y11 = n19343;
  assign y12 = n19359;
  assign y13 = n19542;
  assign y14 = n19268;
  assign y15 = n19574;
  assign y16 = n19593;
  assign y17 = n19615;
  assign y18 = n19637;
  assign y19 = n19670;
  assign y20 = n19694;
  assign y21 = n19714;
  assign y22 = n19239;
  assign y23 = n19739;
  assign y24 = n19383;
  assign y25 = n19775;
  assign y26 = n18527;
  assign y27 = n19855;
  assign y28 = n17816;
  assign y29 = n19879;
  assign y30 = n18918;
  assign y31 = n19951;
  assign y32 = n19444;
  assign y33 = n19982;
  assign y34 = n18634;
  assign y35 = n19997;
  assign y36 = n17937;
  assign y37 = ~n20054;
  assign y38 = n18996;
  assign y39 = n20086;
  assign y40 = n19417;
  assign y41 = n20111;
  assign y42 = n18670;
  assign y43 = n20142;
  assign y44 = n18296;
  assign y45 = n20169;
  assign y46 = n19028;
  assign y47 = n20187;
  assign y48 = n19474;
  assign y49 = n20215;
  assign y50 = n18704;
  assign y51 = ~n20247;
  assign y52 = n18118;
  assign y53 = n20270;
  assign y54 = n18928;
  assign y55 = n20278;
  assign y56 = n19211;
  assign y57 = n20289;
  assign y58 = n18738;
  assign y59 = n20317;
  assign y60 = n18416;
  assign y61 = n20339;
  assign y62 = n18966;
  assign y63 = n20356;
endmodule
