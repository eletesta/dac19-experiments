module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, y0, y1, y2, y3, y4, y5, y6);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10;
  output y0, y1, y2, y3, y4, y5, y6;
  wire n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199;
  assign n12 = x8 & x9;
  assign n13 = x6 & x7;
  assign n14 = ~n12 & n13;
  assign n15 = ~x6 & ~x7;
  assign n16 = x10 & ~n15;
  assign n17 = ~n14 & n16;
  assign n19 = x3 ^ x2;
  assign n20 = x6 & ~n19;
  assign n21 = ~x7 & ~n20;
  assign n22 = x1 & x4;
  assign n23 = n22 ^ x0;
  assign n24 = n23 ^ x5;
  assign n25 = n24 ^ n23;
  assign n26 = x2 ^ x1;
  assign n27 = n26 ^ n23;
  assign n28 = n25 & n27;
  assign n29 = n28 ^ n23;
  assign n30 = ~x6 & ~n29;
  assign n31 = n21 & ~n30;
  assign n18 = x5 ^ x4;
  assign n32 = n31 ^ n18;
  assign n33 = n32 ^ n18;
  assign n34 = x4 ^ x3;
  assign n35 = x7 & n34;
  assign n36 = n35 ^ n18;
  assign n37 = n36 ^ n18;
  assign n38 = ~n33 & ~n37;
  assign n39 = n38 ^ n18;
  assign n40 = ~x8 & ~n39;
  assign n41 = n40 ^ n18;
  assign n42 = n41 ^ x9;
  assign n43 = n42 ^ n41;
  assign n44 = x6 ^ x5;
  assign n45 = n44 ^ n41;
  assign n46 = n43 & n45;
  assign n47 = n46 ^ n41;
  assign n48 = ~x10 & n47;
  assign n49 = ~n17 & ~n48;
  assign n50 = ~x7 & ~x8;
  assign n60 = x2 & x3;
  assign n61 = n60 ^ x4;
  assign n55 = x2 & x4;
  assign n53 = ~x0 & n22;
  assign n54 = n53 ^ x1;
  assign n56 = n55 ^ n54;
  assign n51 = x1 & x2;
  assign n52 = n51 ^ x3;
  assign n57 = n56 ^ n52;
  assign n58 = x5 & n57;
  assign n59 = n58 ^ n56;
  assign n62 = n61 ^ n59;
  assign n63 = n62 ^ n59;
  assign n64 = n59 ^ x9;
  assign n65 = n64 ^ n59;
  assign n66 = ~n63 & ~n65;
  assign n67 = n66 ^ n59;
  assign n68 = x6 & ~n67;
  assign n69 = n68 ^ n59;
  assign n70 = n50 & ~n69;
  assign n71 = x5 & x6;
  assign n72 = n71 ^ x7;
  assign n73 = x9 & n72;
  assign n74 = x4 & x5;
  assign n75 = n74 ^ x6;
  assign n76 = n75 ^ x8;
  assign n77 = n76 ^ n75;
  assign n78 = n77 ^ x9;
  assign n79 = x3 & x4;
  assign n80 = n79 ^ x5;
  assign n81 = n80 ^ x7;
  assign n82 = x7 & ~n81;
  assign n83 = n82 ^ n75;
  assign n84 = n83 ^ x7;
  assign n85 = n78 & ~n84;
  assign n86 = n85 ^ n82;
  assign n87 = n86 ^ x7;
  assign n88 = ~x9 & n87;
  assign n89 = n88 ^ x9;
  assign n90 = ~n73 & n89;
  assign n91 = ~x10 & ~n90;
  assign n92 = ~n70 & n91;
  assign n93 = x8 & n13;
  assign n94 = ~x9 & n93;
  assign n95 = ~x8 & ~n13;
  assign n96 = x10 & ~n95;
  assign n97 = ~n94 & n96;
  assign n98 = ~n92 & ~n97;
  assign n99 = x6 & n74;
  assign n100 = n60 & n99;
  assign n101 = ~x7 & ~n100;
  assign n102 = x5 ^ x2;
  assign n110 = n102 ^ x6;
  assign n103 = n102 ^ x2;
  assign n104 = n103 ^ n102;
  assign n105 = n104 ^ x6;
  assign n106 = n103 ^ x4;
  assign n107 = n106 ^ n103;
  assign n108 = n107 ^ n105;
  assign n109 = ~n105 & ~n108;
  assign n111 = n110 ^ n109;
  assign n112 = n111 ^ n105;
  assign n113 = x6 ^ x3;
  assign n114 = n109 ^ n105;
  assign n115 = ~n113 & ~n114;
  assign n116 = n115 ^ x6;
  assign n117 = ~n112 & ~n116;
  assign n118 = n117 ^ x6;
  assign n119 = n118 ^ x5;
  assign n120 = n119 ^ x6;
  assign n121 = n101 & n120;
  assign n122 = ~x0 & ~x5;
  assign n123 = x1 & ~n122;
  assign n124 = ~x3 & x5;
  assign n125 = n123 & ~n124;
  assign n133 = x3 & ~x6;
  assign n134 = n55 & n133;
  assign n126 = n44 ^ x6;
  assign n127 = n44 ^ x3;
  assign n128 = n127 ^ n44;
  assign n129 = ~n126 & ~n128;
  assign n130 = n129 ^ n44;
  assign n131 = x4 & n130;
  assign n132 = n131 ^ n44;
  assign n135 = n134 ^ n132;
  assign n136 = n125 & n135;
  assign n137 = n136 ^ n132;
  assign n138 = n121 & ~n137;
  assign n139 = ~x3 & n13;
  assign n140 = ~n138 & ~n139;
  assign n141 = ~x8 & ~n140;
  assign n142 = x7 & ~n99;
  assign n143 = ~n95 & n142;
  assign n144 = ~x7 & x8;
  assign n145 = ~n133 & ~n144;
  assign n146 = ~n15 & n74;
  assign n147 = ~n145 & n146;
  assign n148 = ~n143 & ~n147;
  assign n149 = ~n141 & n148;
  assign n150 = ~x9 & ~x10;
  assign n151 = ~n149 & n150;
  assign n152 = x10 ^ x9;
  assign n153 = n93 ^ x10;
  assign n154 = n153 ^ n93;
  assign n155 = x5 & n13;
  assign n156 = n155 ^ x8;
  assign n157 = n156 ^ n93;
  assign n158 = ~n154 & ~n157;
  assign n159 = n158 ^ n93;
  assign n160 = n152 & n159;
  assign n161 = n160 ^ x9;
  assign n162 = ~n151 & ~n161;
  assign n163 = ~x5 & ~x6;
  assign n164 = n50 & n163;
  assign n165 = ~x4 & n164;
  assign n166 = ~x2 & n74;
  assign n167 = n93 & n166;
  assign n168 = ~n165 & ~n167;
  assign n169 = ~x3 & n150;
  assign n170 = ~n168 & n169;
  assign n171 = n123 & n163;
  assign n172 = n60 & n171;
  assign n173 = n51 & n79;
  assign n174 = x4 & ~x5;
  assign n175 = ~x6 & ~n174;
  assign n176 = ~n173 & n175;
  assign n177 = ~n172 & ~n176;
  assign n178 = n101 & n177;
  assign n179 = ~x8 & ~n178;
  assign n180 = ~x2 & ~x3;
  assign n181 = n74 & ~n180;
  assign n182 = n13 & n181;
  assign n183 = ~x9 & ~n182;
  assign n184 = ~n179 & n183;
  assign n185 = x9 ^ x8;
  assign n186 = ~x9 & ~n79;
  assign n187 = ~n185 & n186;
  assign n188 = n187 ^ n185;
  assign n189 = n155 & ~n188;
  assign n190 = ~x10 & ~n189;
  assign n191 = ~n184 & n190;
  assign n192 = n125 & n134;
  assign n193 = n163 & ~n192;
  assign n194 = n50 & ~n100;
  assign n195 = ~n193 & n194;
  assign n196 = x8 & n182;
  assign n197 = n150 & ~n196;
  assign n198 = ~n195 & n197;
  assign n199 = n150 & n194;
  assign y0 = ~n49;
  assign y1 = ~n98;
  assign y2 = ~n162;
  assign y3 = ~n170;
  assign y4 = ~n191;
  assign y5 = ~n198;
  assign y6 = ~n199;
endmodule
