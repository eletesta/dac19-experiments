module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31;
  wire n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305, n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376;
  assign n5812 = x9 ^ x8;
  assign n5813 = x11 ^ x10;
  assign n5814 = n5812 & n5813;
  assign n46 = ~x27 & x28;
  assign n60 = ~x29 & x30;
  assign n150 = n46 & n60;
  assign n77 = x27 & ~x28;
  assign n78 = n60 & n77;
  assign n52 = x23 & x24;
  assign n75 = ~x25 & ~x26;
  assign n3332 = ~n52 & n75;
  assign n3333 = n78 & ~n3332;
  assign n3334 = ~n150 & ~n3333;
  assign n84 = ~x23 & x24;
  assign n137 = n75 & n84;
  assign n308 = n78 & n137;
  assign n102 = n52 & n75;
  assign n322 = n102 & n150;
  assign n3353 = ~n308 & ~n322;
  assign n151 = n137 & n150;
  assign n65 = x27 & x28;
  assign n73 = n60 & n65;
  assign n67 = x25 & ~x26;
  assign n119 = n52 & n67;
  assign n440 = n73 & n119;
  assign n3354 = ~n151 & ~n440;
  assign n3355 = n3353 & n3354;
  assign n3356 = n3334 & n3355;
  assign n97 = n67 & n84;
  assign n248 = n73 & n97;
  assign n49 = x23 & ~x24;
  assign n72 = n49 & n67;
  assign n74 = n72 & n73;
  assign n48 = ~x25 & x26;
  assign n1108 = ~x24 & n48;
  assign n1215 = n73 & n1108;
  assign n3345 = ~n74 & ~n1215;
  assign n3346 = ~n248 & n3345;
  assign n232 = n48 & n84;
  assign n504 = n73 & n232;
  assign n1135 = n73 & n102;
  assign n3089 = ~n504 & ~n1135;
  assign n323 = n73 & n137;
  assign n62 = ~x23 & ~x24;
  assign n68 = n62 & n67;
  assign n449 = n68 & n73;
  assign n3357 = ~n323 & ~n449;
  assign n3358 = n3089 & n3357;
  assign n3359 = n3346 & n3358;
  assign n3360 = n3356 & n3359;
  assign n182 = n49 & n75;
  assign n370 = n73 & n182;
  assign n1467 = ~x23 & ~x25;
  assign n1470 = x26 & ~n1467;
  assign n1471 = ~x24 & n1470;
  assign n1472 = n1471 ^ x26;
  assign n3300 = x25 & ~n62;
  assign n3301 = ~n1472 & ~n3300;
  assign n3302 = n150 & ~n3301;
  assign n3303 = ~n370 & ~n3302;
  assign n666 = n68 & n150;
  assign n50 = n48 & n49;
  assign n948 = n50 & n150;
  assign n353 = n78 & n182;
  assign n76 = n62 & n75;
  assign n640 = n73 & n76;
  assign n2526 = ~n353 & ~n640;
  assign n3361 = ~n948 & n2526;
  assign n3362 = ~n666 & n3361;
  assign n3363 = n3303 & n3362;
  assign n3364 = n3360 & n3363;
  assign n59 = ~x27 & ~x28;
  assign n91 = ~x29 & ~x30;
  assign n121 = n59 & n91;
  assign n122 = n119 & n121;
  assign n54 = x29 & x30;
  assign n81 = n54 & n65;
  assign n755 = n81 & n97;
  assign n3365 = ~n122 & ~n755;
  assign n53 = x25 & x26;
  assign n55 = n46 & n54;
  assign n56 = n53 & n55;
  assign n1475 = ~n75 & n84;
  assign n3366 = n81 & ~n1475;
  assign n3367 = ~n1470 & n3366;
  assign n3368 = ~n56 & ~n3367;
  assign n3369 = n3365 & n3368;
  assign n3370 = n3364 & n3369;
  assign n116 = n54 & n59;
  assign n524 = n116 & n119;
  assign n529 = n116 & n137;
  assign n2737 = ~n524 & ~n529;
  assign n655 = n75 & n121;
  assign n622 = x26 & n116;
  assign n108 = n54 & n77;
  assign n3371 = ~n53 & n108;
  assign n3372 = ~n622 & ~n3371;
  assign n3373 = ~n655 & n3372;
  assign n3374 = n2737 & n3373;
  assign n517 = n68 & n121;
  assign n197 = n102 & n116;
  assign n227 = n116 & n182;
  assign n3375 = ~n197 & ~n227;
  assign n3376 = ~n517 & n3375;
  assign n3377 = n3374 & n3376;
  assign n85 = n53 & n84;
  assign n361 = n73 & n85;
  assign n750 = n68 & n116;
  assign n1301 = ~n361 & ~n750;
  assign n82 = n52 & n53;
  assign n710 = n73 & n82;
  assign n117 = n72 & n116;
  assign n142 = n53 & n62;
  assign n841 = n73 & n142;
  assign n842 = ~n117 & ~n841;
  assign n3135 = ~n710 & n842;
  assign n3136 = n1301 & n3135;
  assign n152 = n76 & n116;
  assign n350 = n97 & n116;
  assign n2975 = ~n152 & ~n350;
  assign n147 = n48 & n52;
  assign n300 = n73 & n147;
  assign n114 = n49 & n53;
  assign n525 = n73 & n114;
  assign n3122 = ~n300 & ~n525;
  assign n3378 = n2975 & n3122;
  assign n3379 = n108 ^ n55;
  assign n3380 = n53 & n3379;
  assign n3381 = n3380 ^ n55;
  assign n3382 = n3378 & ~n3381;
  assign n3383 = n3136 & n3382;
  assign n3384 = n3377 & n3383;
  assign n3385 = n3370 & n3384;
  assign n63 = n48 & n62;
  assign n574 = ~x28 & n91;
  assign n575 = n63 & n574;
  assign n576 = ~x27 & n575;
  assign n134 = n50 & n81;
  assign n689 = n81 & n85;
  assign n1083 = ~n134 & ~n689;
  assign n409 = n81 & n114;
  assign n428 = n55 & n85;
  assign n850 = n55 & n142;
  assign n3081 = ~n428 & ~n850;
  assign n3082 = ~n409 & n3081;
  assign n3083 = n1083 & n3082;
  assign n3084 = ~n576 & n3083;
  assign n209 = n81 & n142;
  assign n330 = n81 & n232;
  assign n1058 = ~n209 & ~n330;
  assign n83 = n81 & n82;
  assign n758 = n81 & n147;
  assign n2654 = ~n83 & ~n758;
  assign n3318 = n1058 & n2654;
  assign n403 = n50 & n121;
  assign n61 = n59 & n60;
  assign n228 = n97 & n121;
  assign n11915 = ~n61 & ~n228;
  assign n11916 = ~n403 & n11915;
  assign n79 = n76 & n78;
  assign n610 = n72 & n121;
  assign n3450 = ~n79 & ~n610;
  assign n45 = x29 & ~x30;
  assign n66 = n45 & n65;
  assign n796 = x26 & n66;
  assign n5451 = ~x25 & n62;
  assign n11917 = n796 & ~n5451;
  assign n11918 = n3450 & ~n11917;
  assign n11919 = n11916 & n11918;
  assign n11920 = n3318 & n11919;
  assign n11921 = n3084 & n11920;
  assign n11922 = n3385 & n11921;
  assign n497 = n66 & n137;
  assign n262 = n66 & n182;
  assign n946 = n66 & n102;
  assign n1789 = ~n262 & ~n946;
  assign n3323 = ~n497 & n1789;
  assign n158 = n46 & n91;
  assign n761 = ~x26 & n52;
  assign n762 = n158 & n761;
  assign n763 = x25 & n762;
  assign n11743 = ~n763 & n3369;
  assign n11744 = n3323 & n11743;
  assign n11840 = n3384 & n11744;
  assign n47 = n45 & n46;
  assign n214 = x23 & n47;
  assign n439 = n47 & n137;
  assign n3412 = ~n214 & ~n439;
  assign n86 = n45 & n77;
  assign n499 = x23 & n67;
  assign n500 = n86 & n499;
  assign n646 = x26 & n62;
  assign n647 = n47 & n646;
  assign n3413 = ~n500 & ~n647;
  assign n470 = x24 & n75;
  assign n3414 = n86 & n470;
  assign n3415 = n3413 & ~n3414;
  assign n3416 = n3412 & n3415;
  assign n514 = n50 & n86;
  assign n920 = n66 & n76;
  assign n1164 = ~n514 & ~n920;
  assign n269 = n86 & n114;
  assign n751 = n86 & n142;
  assign n3417 = ~n269 & ~n751;
  assign n3418 = n1164 & n3417;
  assign n3419 = n3416 & n3418;
  assign n11841 = n3318 & n3419;
  assign n11842 = n11840 & n11841;
  assign n87 = n85 & n86;
  assign n558 = n66 & n97;
  assign n2721 = ~n87 & ~n558;
  assign n92 = n77 & n91;
  assign n416 = n85 & n92;
  assign n582 = n158 & n182;
  assign n3085 = ~n416 & ~n582;
  assign n3086 = n2721 & n3085;
  assign n186 = n86 & n182;
  assign n475 = n47 & n82;
  assign n3087 = ~n186 & ~n475;
  assign n3088 = n3086 & n3087;
  assign n69 = n66 & n68;
  assign n103 = n47 & n102;
  assign n2073 = ~n69 & ~n103;
  assign n111 = n47 & n85;
  assign n588 = n66 & n119;
  assign n2550 = ~n111 & ~n588;
  assign n2551 = n2073 & n2550;
  assign n278 = n86 & n232;
  assign n492 = n47 & n68;
  assign n3090 = ~n278 & ~n492;
  assign n3091 = n3089 & n3090;
  assign n3092 = n2551 & n3091;
  assign n3093 = n3088 & n3092;
  assign n3094 = n3084 & n3093;
  assign n509 = n114 & n158;
  assign n611 = ~n509 & ~n610;
  assign n1345 = n66 & n499;
  assign n1482 = ~x24 & n1345;
  assign n3095 = n611 & ~n1482;
  assign n3096 = n3094 & n3095;
  assign n975 = n102 & n158;
  assign n452 = n47 & n232;
  assign n4152 = ~n74 & ~n452;
  assign n4153 = ~n975 & n4152;
  assign n198 = n65 & n91;
  assign n199 = n182 & n198;
  assign n205 = x24 & n48;
  assign n206 = n158 & n205;
  assign n4154 = ~n199 & ~n206;
  assign n4155 = n4153 & n4154;
  assign n456 = n68 & n86;
  assign n457 = ~n228 & ~n456;
  assign n166 = n63 & n66;
  assign n549 = n47 & n97;
  assign n2292 = ~n166 & ~n549;
  assign n4156 = n457 & n2292;
  assign n812 = n63 & n86;
  assign n919 = n47 & n182;
  assign n2942 = ~n812 & ~n919;
  assign n201 = n47 & n76;
  assign n4157 = ~n201 & ~n403;
  assign n4158 = n2942 & n4157;
  assign n4159 = n4156 & n4158;
  assign n4160 = n4155 & n4159;
  assign n93 = n82 & n92;
  assign n3856 = ~n205 & ~n761;
  assign n3857 = n158 & n3856;
  assign n3858 = ~n93 & ~n3857;
  assign n402 = n85 & n158;
  assign n929 = n92 & n114;
  assign n999 = ~n402 & ~n929;
  assign n3859 = ~x23 & n75;
  assign n3860 = n198 & n3859;
  assign n3861 = n999 & ~n3860;
  assign n3862 = n3858 & n3861;
  assign n295 = n86 & n97;
  assign n296 = n86 & n147;
  assign n297 = ~n295 & ~n296;
  assign n787 = n82 & n86;
  assign n1197 = ~n449 & ~n787;
  assign n11843 = n297 & n1197;
  assign n215 = x24 & n67;
  assign n11844 = n73 & n215;
  assign n11845 = ~n1215 & ~n11844;
  assign n11846 = n11843 & n11845;
  assign n11847 = n3862 & n11846;
  assign n11848 = n4160 & n11847;
  assign n11849 = n3096 & n11848;
  assign n11850 = n11842 & n11849;
  assign n1055 = ~n666 & ~n751;
  assign n552 = n50 & n92;
  assign n1056 = ~n122 & ~n552;
  assign n1057 = n1055 & n1056;
  assign n1059 = n1057 & n1058;
  assign n293 = n119 & n150;
  assign n660 = n68 & n158;
  assign n937 = ~n293 & ~n660;
  assign n208 = n97 & n150;
  assign n1060 = n114 & n116;
  assign n1061 = ~n208 & ~n1060;
  assign n1062 = n937 & n1061;
  assign n469 = n63 & n121;
  assign n1063 = ~n201 & ~n469;
  assign n1064 = ~x23 & n53;
  assign n1065 = n61 & n1064;
  assign n1066 = n1063 & ~n1065;
  assign n1067 = n1062 & n1066;
  assign n1068 = n1059 & n1067;
  assign n417 = n92 & n137;
  assign n94 = n45 & n59;
  assign n115 = n94 & n114;
  assign n541 = n76 & n92;
  assign n602 = ~n115 & ~n541;
  assign n1069 = n602 & ~n919;
  assign n1070 = ~n417 & n1069;
  assign n1071 = n1068 & n1070;
  assign n550 = n50 & n116;
  assign n1072 = ~n524 & ~n550;
  assign n347 = n76 & n198;
  assign n1073 = ~n322 & ~n347;
  assign n1074 = n1072 & n1073;
  assign n277 = n85 & n150;
  assign n279 = ~n277 & ~n278;
  assign n64 = n61 & n63;
  assign n1075 = ~n64 & ~n166;
  assign n1076 = n279 & n1075;
  assign n1077 = n1074 & n1076;
  assign n156 = n147 & n150;
  assign n1078 = ~n156 & ~n946;
  assign n298 = n137 & n198;
  assign n351 = n85 & n198;
  assign n1079 = ~n298 & ~n351;
  assign n1080 = n1078 & n1079;
  assign n1081 = n1077 & n1080;
  assign n1082 = n1071 & n1081;
  assign n163 = n76 & n121;
  assign n164 = n82 & n150;
  assign n165 = ~n163 & ~n164;
  assign n1084 = n165 & n1083;
  assign n249 = n198 & n232;
  assign n1085 = ~n249 & ~n323;
  assign n1086 = n1084 & n1085;
  assign n202 = n61 & n82;
  assign n1087 = ~n79 & ~n202;
  assign n1088 = n1086 & n1087;
  assign n642 = n52 & n108;
  assign n826 = n67 & n642;
  assign n535 = n63 & n81;
  assign n1089 = ~n69 & ~n535;
  assign n1090 = ~n826 & n1089;
  assign n133 = n50 & n94;
  assign n373 = n68 & n108;
  assign n1091 = ~n133 & ~n373;
  assign n1092 = n1090 & n1091;
  assign n231 = n76 & n94;
  assign n540 = n150 & n232;
  assign n1093 = ~n231 & ~n540;
  assign n1094 = n1092 & n1093;
  assign n1095 = n1088 & n1094;
  assign n1096 = n1082 & n1095;
  assign n1266 = n147 & n198;
  assign n141 = n50 & n61;
  assign n334 = n108 & n147;
  assign n2692 = ~n87 & ~n334;
  assign n2693 = ~n141 & n2692;
  assign n303 = n63 & n116;
  assign n503 = n97 & n108;
  assign n2307 = ~n303 & ~n503;
  assign n301 = n116 & n142;
  assign n527 = n72 & n150;
  assign n2694 = ~n301 & ~n527;
  assign n2695 = n2307 & n2694;
  assign n2696 = n2693 & n2695;
  assign n404 = ~n402 & ~n403;
  assign n128 = n81 & n119;
  assign n183 = n92 & n182;
  assign n2595 = ~n128 & ~n183;
  assign n2697 = n404 & n2595;
  assign n2698 = n2696 & n2697;
  assign n2699 = ~n1266 & n2698;
  assign n146 = n94 & n142;
  assign n253 = n92 & n147;
  assign n11379 = ~n146 & ~n253;
  assign n11380 = ~n262 & n11379;
  assign n192 = n50 & n108;
  assign n476 = n108 & n137;
  assign n868 = ~n192 & ~n476;
  assign n234 = n121 & n182;
  assign n2968 = ~n234 & ~n439;
  assign n11381 = n868 & n2968;
  assign n11382 = n11380 & n11381;
  assign n385 = n76 & n108;
  assign n627 = n137 & n158;
  assign n4048 = ~n385 & ~n627;
  assign n378 = n63 & n108;
  assign n557 = n92 & n232;
  assign n4065 = ~n378 & ~n557;
  assign n11383 = n4048 & n4065;
  assign n190 = n82 & n94;
  assign n250 = n85 & n116;
  assign n884 = ~n190 & ~n250;
  assign n369 = n108 & n232;
  assign n630 = n63 & n150;
  assign n3473 = ~n369 & ~n630;
  assign n11384 = n884 & n3473;
  assign n11385 = n11383 & n11384;
  assign n11386 = n11382 & n11385;
  assign n218 = n61 & n119;
  assign n272 = n61 & n114;
  assign n949 = ~n272 & ~n948;
  assign n3005 = ~n218 & n949;
  assign n281 = n76 & n86;
  assign n709 = n114 & n198;
  assign n2385 = ~n281 & ~n709;
  assign n3828 = ~n640 & n2385;
  assign n11387 = n3005 & n3828;
  assign n319 = n82 & n121;
  assign n2104 = ~n319 & ~n509;
  assign n5534 = n2104 & n2654;
  assign n478 = n82 & n198;
  assign n584 = ~n111 & ~n478;
  assign n11388 = ~n370 & n584;
  assign n11389 = n5534 & n11388;
  assign n11390 = n11387 & n11389;
  assign n11391 = n11386 & n11390;
  assign n621 = ~x25 & n52;
  assign n623 = n621 & n622;
  assign n675 = n47 & n114;
  assign n915 = ~n623 & ~n675;
  assign n4054 = ~n228 & ~n755;
  assign n424 = n97 & n158;
  assign n4055 = ~n424 & ~n975;
  assign n4056 = n4054 & n4055;
  assign n4057 = n915 & n4056;
  assign n1155 = ~n269 & ~n350;
  assign n1156 = ~n296 & n1155;
  assign n4386 = ~n151 & n1156;
  assign n11392 = n4057 & n4386;
  assign n928 = n142 & n150;
  assign n136 = n61 & n97;
  assign n358 = n82 & n158;
  assign n2130 = ~n136 & ~n358;
  assign n2131 = ~n928 & n2130;
  assign n375 = n114 & n150;
  assign n2132 = ~n375 & ~n497;
  assign n2133 = n2131 & n2132;
  assign n109 = n102 & n108;
  assign n233 = n61 & n232;
  assign n4098 = ~n109 & ~n233;
  assign n189 = n108 & n182;
  assign n11393 = ~n189 & ~n475;
  assign n11394 = n4098 & n11393;
  assign n11395 = ~n199 & n11394;
  assign n11396 = n2133 & n11395;
  assign n11397 = n11392 & n11396;
  assign n11398 = n11391 & n11397;
  assign n11399 = n2699 & n11398;
  assign n170 = n85 & n94;
  assign n171 = n66 & n72;
  assign n172 = ~n170 & ~n171;
  assign n221 = n61 & n72;
  assign n4174 = ~n221 & ~n558;
  assign n4175 = n172 & n4174;
  assign n312 = n116 & n232;
  assign n429 = n63 & n92;
  assign n5130 = ~n312 & ~n429;
  assign n280 = n72 & n108;
  assign n11400 = ~n280 & ~n920;
  assign n11401 = n5130 & n11400;
  assign n304 = n72 & n158;
  assign n11402 = ~n304 & ~n409;
  assign n244 = n61 & n147;
  assign n11403 = ~n244 & ~n787;
  assign n11404 = n11402 & n11403;
  assign n11405 = n11401 & n11404;
  assign n148 = n94 & n147;
  assign n257 = n82 & n116;
  assign n473 = ~n148 & ~n257;
  assign n1240 = ~n308 & ~n353;
  assign n1241 = ~n588 & n1240;
  assign n11406 = n473 & n1241;
  assign n11407 = n11405 & n11406;
  assign n11408 = n4175 & n11407;
  assign n314 = n94 & n232;
  assign n346 = n92 & n142;
  assign n362 = n142 & n198;
  assign n11409 = ~n346 & ~n362;
  assign n11410 = ~n314 & n11409;
  assign n11411 = n11408 & n11410;
  assign n11412 = n11399 & n11411;
  assign n11413 = n1096 & n11412;
  assign n11836 = n11413 ^ x29;
  assign n412 = n47 & n63;
  assign n828 = ~n347 & ~n412;
  assign n714 = n47 & n147;
  assign n829 = ~n689 & ~n714;
  assign n830 = n828 & n829;
  assign n216 = n214 & n215;
  assign n3290 = ~n148 & ~n216;
  assign n3291 = ~n640 & n3290;
  assign n3247 = ~n103 & ~n549;
  assign n95 = n68 & n94;
  assign n570 = ~n95 & ~n323;
  assign n432 = n92 & n97;
  assign n676 = ~n432 & ~n675;
  assign n3292 = n570 & n676;
  assign n3293 = n3247 & n3292;
  assign n3294 = n3291 & n3293;
  assign n3295 = n830 & n3294;
  assign n359 = n158 & n232;
  assign n360 = ~n358 & ~n359;
  assign n1153 = ~n151 & ~n402;
  assign n1154 = ~n133 & n1153;
  assign n2038 = ~n146 & ~n314;
  assign n2267 = ~n429 & ~n666;
  assign n3296 = n2038 & n2267;
  assign n3297 = n1154 & n3296;
  assign n3298 = n360 & n3297;
  assign n3299 = n3295 & n3298;
  assign n3304 = ~n928 & n3303;
  assign n790 = n94 & n119;
  assign n1608 = ~n557 & ~n790;
  assign n126 = n72 & n94;
  assign n2121 = ~n126 & ~n322;
  assign n2122 = n1608 & n2121;
  assign n410 = n94 & n97;
  assign n2123 = ~n199 & ~n410;
  assign n2124 = n2122 & n2123;
  assign n3305 = ~n509 & n2124;
  assign n3306 = n3304 & n3305;
  assign n458 = n92 & n119;
  assign n173 = n63 & n158;
  assign n381 = ~n173 & ~n293;
  assign n390 = n142 & n158;
  assign n612 = n63 & n94;
  assign n3307 = ~n390 & ~n612;
  assign n3308 = n381 & n3307;
  assign n3309 = ~n458 & n3308;
  assign n418 = n94 & n137;
  assign n931 = ~n409 & ~n418;
  assign n3310 = ~n452 & ~n948;
  assign n3311 = n931 & n3310;
  assign n51 = n47 & n50;
  assign n354 = n47 & n72;
  assign n445 = ~n51 & ~n354;
  assign n2239 = ~n111 & ~n492;
  assign n3312 = n445 & n2239;
  assign n3313 = n3311 & n3312;
  assign n3314 = n3309 & n3313;
  assign n185 = n50 & n158;
  assign n437 = ~n134 & ~n185;
  assign n3199 = n437 & ~n552;
  assign n671 = n147 & n158;
  assign n237 = n47 & n142;
  assign n567 = n94 & n102;
  assign n3315 = ~n237 & ~n567;
  assign n3316 = ~n671 & n3315;
  assign n3317 = n3199 & n3316;
  assign n3319 = n3317 & n3318;
  assign n3320 = n3314 & n3319;
  assign n3321 = n3306 & n3320;
  assign n3322 = n3299 & n3321;
  assign n680 = n92 & n102;
  assign n4019 = ~n281 & ~n680;
  assign n226 = n72 & n92;
  assign n2623 = ~n170 & ~n226;
  assign n5623 = ~n298 & n2623;
  assign n11741 = n4019 & n5623;
  assign n11742 = n3322 & n11741;
  assign n2625 = ~n253 & ~n346;
  assign n11745 = n2625 & n11744;
  assign n270 = n94 & n182;
  assign n699 = n68 & n77;
  assign n1536 = n91 & n699;
  assign n1650 = ~n270 & ~n1536;
  assign n1866 = ~n475 & ~n920;
  assign n3347 = ~n403 & n1866;
  assign n11746 = n1650 & n3347;
  assign n11747 = n3081 & ~n3381;
  assign n11748 = n11746 & n11747;
  assign n11749 = ~n63 & ~n67;
  assign n11750 = n66 & ~n11749;
  assign n817 = ~x24 & ~x25;
  assign n11751 = n817 ^ x26;
  assign n11752 = n121 & ~n11751;
  assign n11753 = ~n11750 & ~n11752;
  assign n11754 = ~n115 & ~n190;
  assign n11755 = n11753 & n11754;
  assign n11756 = n3334 & n11755;
  assign n11757 = n11748 & n11756;
  assign n11758 = n11745 & n11757;
  assign n11759 = n11742 & n11758;
  assign n11837 = n11759 ^ n11413;
  assign n11838 = n11836 & ~n11837;
  assign n11839 = n11838 ^ x29;
  assign n11851 = n11850 ^ n11839;
  assign n3426 = ~x26 & n92;
  assign n3427 = ~n3300 & n3426;
  assign n3428 = ~n121 & ~n3427;
  assign n634 = n50 & n198;
  assign n635 = ~n416 & ~n634;
  assign n1299 = ~n199 & ~n582;
  assign n3863 = n158 & ~n3856;
  assign n3864 = n1299 & ~n3863;
  assign n3865 = n635 & n3864;
  assign n3866 = ~n67 & ~n646;
  assign n3867 = n3856 & n3866;
  assign n3868 = n198 & ~n3867;
  assign n3869 = n2625 & ~n3868;
  assign n3870 = n3865 & n3869;
  assign n3871 = n3862 & n3870;
  assign n3872 = ~n709 & n3871;
  assign n3398 = n48 & ~n52;
  assign n3399 = ~n215 & ~n3398;
  assign n3400 = n92 & ~n3399;
  assign n3873 = ~n226 & ~n3400;
  assign n3874 = n3872 & n3873;
  assign n3875 = n3428 & n3874;
  assign n41 = x30 ^ x29;
  assign n3325 = ~n929 & n2625;
  assign n652 = n86 & n137;
  assign n1183 = ~n456 & ~n652;
  assign n3175 = ~n170 & ~n281;
  assign n3252 = n1183 & n3175;
  assign n1302 = ~n186 & ~n627;
  assign n1005 = n76 & n158;
  assign n2401 = ~n93 & ~n1005;
  assign n3253 = n1302 & n2401;
  assign n3254 = n3252 & n3253;
  assign n723 = n86 & n102;
  assign n3255 = ~n723 & n3085;
  assign n3256 = n3254 & n3255;
  assign n536 = ~n304 & ~n314;
  assign n781 = ~n424 & ~n660;
  assign n3386 = n781 & ~n975;
  assign n3387 = n536 & n3386;
  assign n1500 = x24 & x25;
  assign n1507 = x26 & n198;
  assign n1508 = n1500 & n1507;
  assign n3388 = ~n94 & ~n1508;
  assign n3389 = n3387 & n3388;
  assign n3390 = n3256 & n3389;
  assign n3391 = n3325 & n3390;
  assign n3392 = n297 & n3081;
  assign n1501 = x26 & ~n1500;
  assign n3393 = n86 & n1501;
  assign n3394 = ~n610 & ~n3393;
  assign n3395 = ~n228 & n3394;
  assign n3396 = n3392 & n3395;
  assign n3397 = ~n500 & n3396;
  assign n617 = n119 & n158;
  assign n3401 = ~n617 & ~n3400;
  assign n3402 = n3397 & n3401;
  assign n3403 = n3391 & n3402;
  assign n3404 = n3385 & n3403;
  assign n3324 = ~n163 & n3323;
  assign n3326 = ~n87 & ~n1135;
  assign n3327 = ~n919 & n3326;
  assign n3328 = n3325 & n3327;
  assign n3329 = n3324 & n3328;
  assign n441 = ~n439 & ~n440;
  assign n518 = n85 & n121;
  assign n3330 = ~n234 & ~n518;
  assign n3331 = n441 & n3330;
  assign n3335 = n1240 & n3334;
  assign n3336 = n3331 & n3335;
  assign n893 = ~n270 & ~n351;
  assign n3337 = n1063 & n1197;
  assign n3338 = n893 & n3337;
  assign n3339 = n3336 & n3338;
  assign n3340 = n3329 & n3339;
  assign n309 = n121 & n205;
  assign n592 = n114 & n121;
  assign n3341 = ~n478 & ~n592;
  assign n3342 = ~n309 & n3341;
  assign n254 = n121 & n142;
  assign n3343 = ~n231 & ~n254;
  assign n3344 = n3342 & n3343;
  assign n3348 = n3346 & n3347;
  assign n3349 = n3344 & n3348;
  assign n3350 = n3340 & n3349;
  assign n3351 = n3322 & n3350;
  assign n3200 = n78 & n499;
  assign n3201 = ~n1345 & ~n3200;
  assign n463 = n50 & n78;
  assign n3202 = ~n250 & ~n463;
  assign n3203 = n3201 & n3202;
  assign n3204 = n3199 & n3203;
  assign n386 = ~n350 & ~n385;
  assign n238 = n50 & n66;
  assign n1611 = ~n87 & ~n238;
  assign n3205 = n386 & n1611;
  assign n3206 = n3204 & n3205;
  assign n797 = n621 & n796;
  assign n3207 = ~n206 & ~n303;
  assign n3208 = n893 & n3207;
  assign n3209 = ~n797 & n3208;
  assign n3210 = n3206 & n3209;
  assign n1335 = ~n152 & ~n576;
  assign n3211 = ~n710 & ~n841;
  assign n3212 = n1335 & n3211;
  assign n405 = n61 & n76;
  assign n406 = n76 & n150;
  assign n407 = ~n405 & ~n406;
  assign n3213 = ~n257 & ~n787;
  assign n3214 = n407 & n3213;
  assign n3215 = n3212 & n3214;
  assign n326 = n78 & n114;
  assign n217 = n68 & n78;
  assign n2137 = ~n217 & ~n409;
  assign n3216 = ~n326 & n2137;
  assign n292 = n78 & n102;
  assign n482 = ~n292 & ~n361;
  assign n2391 = ~n312 & ~n403;
  assign n3217 = n482 & n2391;
  assign n3218 = n3216 & n3217;
  assign n3219 = n3215 & n3218;
  assign n3220 = n3210 & n3219;
  assign n2731 = ~n429 & ~n750;
  assign n1227 = n116 & n147;
  assign n2732 = ~n83 & ~n1227;
  assign n2733 = n2731 & n2732;
  assign n392 = n66 & n82;
  assign n553 = n78 & n232;
  assign n727 = ~n392 & ~n553;
  assign n560 = n66 & n232;
  assign n2734 = ~n560 & ~n567;
  assign n2735 = n727 & n2734;
  assign n2736 = n2733 & n2735;
  assign n2738 = n2736 & n2737;
  assign n2159 = ~n151 & ~n758;
  assign n245 = n66 & n114;
  assign n313 = n78 & n142;
  assign n3221 = ~n245 & ~n313;
  assign n3222 = n2159 & n3221;
  assign n3223 = ~n458 & n3222;
  assign n3224 = n2738 & n3223;
  assign n3225 = n3220 & n3224;
  assign n897 = ~x27 & n54;
  assign n898 = n50 & n897;
  assign n899 = ~x28 & n898;
  assign n900 = ~n525 & ~n899;
  assign n901 = n63 & n78;
  assign n902 = ~n478 & ~n901;
  assign n903 = ~n189 & ~n432;
  assign n904 = n902 & n903;
  assign n905 = n900 & n904;
  assign n531 = n121 & n232;
  assign n859 = ~n418 & ~n531;
  assign n3226 = ~n919 & n1058;
  assign n3227 = n859 & n3226;
  assign n3228 = n905 & n3227;
  assign n273 = n78 & n97;
  assign n2771 = ~n273 & ~n301;
  assign n2772 = ~n201 & ~n689;
  assign n2773 = n2771 & n2772;
  assign n3229 = ~n439 & ~n558;
  assign n3230 = n2773 & n3229;
  assign n3231 = n3228 & n3230;
  assign n256 = n66 & n85;
  assign n327 = n66 & n142;
  assign n2165 = ~n256 & ~n327;
  assign n1520 = ~n117 & ~n197;
  assign n3232 = ~n173 & ~n476;
  assign n3233 = n1520 & n3232;
  assign n3234 = n2165 & n3233;
  assign n344 = n78 & n147;
  assign n2634 = ~n69 & ~n166;
  assign n3235 = ~n344 & n2634;
  assign n3236 = n3234 & n3235;
  assign n628 = n78 & n85;
  assign n1670 = ~n300 & ~n628;
  assign n1671 = ~n227 & n1670;
  assign n1109 = ~x26 & n62;
  assign n3237 = n94 & n1109;
  assign n3238 = ~n390 & ~n3237;
  assign n3239 = ~n1060 & n3238;
  assign n193 = n150 & n182;
  assign n683 = n78 & n82;
  assign n3240 = ~n193 & ~n683;
  assign n3241 = n3239 & n3240;
  assign n3242 = n1671 & n3241;
  assign n3243 = n3236 & n3242;
  assign n3244 = n3231 & n3243;
  assign n3245 = n3225 & n3244;
  assign n331 = n72 & n198;
  assign n1765 = ~n331 & ~n354;
  assign n687 = n61 & n182;
  assign n3246 = ~n492 & ~n687;
  assign n3248 = n3246 & n3247;
  assign n3249 = n1765 & n3248;
  assign n283 = n97 & n198;
  assign n657 = ~n109 & ~n283;
  assign n3250 = ~n412 & n657;
  assign n3251 = n3249 & n3250;
  assign n3257 = n3251 & n3256;
  assign n3258 = ~n216 & ~n504;
  assign n374 = ~n190 & ~n373;
  assign n3259 = n374 & n1240;
  assign n3260 = n3258 & n3259;
  assign n3261 = ~n319 & ~n517;
  assign n3262 = ~n183 & n3261;
  assign n494 = n119 & n198;
  assign n3263 = ~n298 & ~n494;
  assign n3264 = n3262 & n3263;
  assign n3265 = n3260 & n3264;
  assign n471 = n121 & n470;
  assign n544 = n68 & n198;
  assign n843 = n102 & n198;
  assign n844 = ~n544 & ~n843;
  assign n3266 = n602 & n844;
  assign n3267 = ~n471 & n3266;
  assign n3268 = n3265 & n3267;
  assign n3269 = n3257 & n3268;
  assign n3270 = n3245 & n3269;
  assign n333 = n61 & n68;
  assign n1771 = ~n333 & ~n458;
  assign n3108 = n602 & ~n901;
  assign n3109 = n1771 & n3108;
  assign n3110 = ~n197 & ~n514;
  assign n3111 = ~n51 & ~n540;
  assign n3112 = n3110 & n3111;
  assign n3113 = ~n69 & ~n612;
  assign n3114 = n3112 & n3113;
  assign n3115 = n3109 & n3114;
  assign n155 = n61 & n102;
  assign n3116 = ~n155 & ~n529;
  assign n3117 = ~n163 & ~n588;
  assign n3118 = n3116 & n3117;
  assign n222 = n108 & n119;
  assign n223 = ~n221 & ~n222;
  assign n2453 = ~n503 & ~n948;
  assign n3119 = n223 & n2453;
  assign n3120 = n3118 & n3119;
  assign n174 = n108 & n114;
  assign n175 = ~n173 & ~n174;
  assign n3121 = n175 & ~n478;
  assign n3123 = ~n630 & n3122;
  assign n3124 = n3121 & n3123;
  assign n3125 = n3120 & n3124;
  assign n3126 = n3115 & n3125;
  assign n3127 = ~n334 & ~n558;
  assign n3128 = ~n208 & ~n843;
  assign n3129 = n3127 & n3128;
  assign n1103 = ~n295 & ~n416;
  assign n506 = n85 & n108;
  assign n3130 = ~n463 & ~n506;
  assign n3131 = n1103 & n3130;
  assign n3132 = n3129 & n3131;
  assign n3133 = ~n469 & n3132;
  assign n3134 = n3126 & n3133;
  assign n2298 = ~n136 & ~n378;
  assign n3137 = ~n152 & ~n369;
  assign n3138 = n2298 & n3137;
  assign n1047 = n78 & n119;
  assign n1678 = ~n544 & ~n1047;
  assign n3139 = n1075 & n1678;
  assign n3140 = n3138 & n3139;
  assign n3141 = n3136 & n3140;
  assign n219 = ~n217 & ~n218;
  assign n2618 = ~n156 & n219;
  assign n791 = n61 & n137;
  assign n1332 = ~n298 & ~n791;
  assign n2760 = ~n432 & n1332;
  assign n3142 = n2618 & n2760;
  assign n3143 = n3141 & n3142;
  assign n3144 = ~n319 & ~n610;
  assign n3145 = ~n812 & n3144;
  assign n99 = n72 & n78;
  assign n376 = ~n99 & ~n375;
  assign n442 = n108 & n142;
  assign n3146 = ~n442 & ~n928;
  assign n3147 = n376 & n3146;
  assign n3148 = n3145 & n3147;
  assign n229 = ~n227 & ~n228;
  assign n3149 = n229 & ~n273;
  assign n3150 = n3148 & n3149;
  assign n1158 = ~n280 & ~n330;
  assign n3151 = n893 & n1158;
  assign n3152 = ~n192 & ~n500;
  assign n3153 = n2401 & n3152;
  assign n3154 = n3151 & n3153;
  assign n294 = ~n292 & ~n293;
  assign n3155 = n294 & n437;
  assign n3156 = ~n171 & ~n231;
  assign n3157 = n3155 & n3156;
  assign n3158 = n3154 & n3157;
  assign n3159 = n3150 & n3158;
  assign n3160 = n3143 & n3159;
  assign n3161 = n3134 & n3160;
  assign n255 = ~n253 & ~n254;
  assign n3162 = n255 & n2654;
  assign n955 = ~n504 & ~n680;
  assign n138 = n55 & n137;
  assign n3163 = ~n138 & ~n660;
  assign n3164 = n955 & n3163;
  assign n3165 = n3162 & n3164;
  assign n411 = ~n409 & ~n410;
  assign n799 = n55 & n102;
  assign n1021 = ~n557 & ~n799;
  assign n3166 = n411 & n1021;
  assign n889 = ~n237 & ~n439;
  assign n396 = n55 & n76;
  assign n1305 = ~n396 & ~n787;
  assign n3167 = n889 & n1305;
  assign n3168 = n3166 & n3167;
  assign n3169 = n3165 & n3168;
  assign n3170 = ~n417 & n1611;
  assign n656 = n84 & n655;
  assign n593 = n121 & n147;
  assign n3171 = ~n201 & ~n593;
  assign n3172 = ~n656 & n3171;
  assign n3173 = n3170 & n3172;
  assign n3174 = ~n689 & n1240;
  assign n3176 = ~n249 & n3175;
  assign n3177 = n3174 & n3176;
  assign n3178 = n3173 & n3177;
  assign n3179 = n3169 & n3178;
  assign n3180 = ~n322 & ~n666;
  assign n127 = n102 & n121;
  assign n740 = n55 & n182;
  assign n3181 = ~n127 & ~n740;
  assign n3182 = n3180 & n3181;
  assign n104 = n55 & n68;
  assign n336 = n63 & n198;
  assign n2806 = ~n104 & ~n336;
  assign n3183 = ~n527 & ~n919;
  assign n3184 = n2806 & n3183;
  assign n3185 = n3182 & n3184;
  assign n597 = ~n209 & ~n452;
  assign n263 = n82 & n108;
  assign n800 = n55 & n72;
  assign n2240 = ~n263 & ~n800;
  assign n3186 = n597 & n2240;
  assign n3187 = n404 & n3186;
  assign n3188 = n3185 & n3187;
  assign n2187 = ~n509 & ~n675;
  assign n3189 = ~n560 & ~n634;
  assign n3190 = n2187 & n3189;
  assign n976 = ~n126 & ~n975;
  assign n690 = x25 & n52;
  assign n691 = n94 & n690;
  assign n3191 = ~n691 & ~n714;
  assign n3192 = n976 & n3191;
  assign n3193 = n3190 & n3192;
  assign n3194 = n3188 & n3193;
  assign n3195 = n3179 & n3194;
  assign n3196 = n3161 & n3195;
  assign n1352 = ~n369 & ~n442;
  assign n1353 = ~n164 & ~n1227;
  assign n1354 = n1352 & n1353;
  assign n210 = ~n208 & ~n209;
  assign n2067 = ~n797 & ~n826;
  assign n2068 = n210 & n2067;
  assign n2069 = n1354 & n2068;
  assign n2070 = ~n652 & ~n1266;
  assign n2071 = ~n899 & n2070;
  assign n2072 = n2069 & n2071;
  assign n1825 = ~n628 & ~n841;
  assign n1826 = ~n244 & ~n634;
  assign n1827 = n1825 & n1826;
  assign n3038 = ~n201 & ~n920;
  assign n1166 = n55 & n232;
  assign n3039 = ~n531 & ~n1166;
  assign n3040 = n3038 & n3039;
  assign n3041 = ~n192 & ~n410;
  assign n3042 = ~n155 & ~n277;
  assign n3043 = n3041 & n3042;
  assign n3044 = n3040 & n3043;
  assign n3045 = n1827 & n3044;
  assign n3046 = ~n133 & ~n370;
  assign n3047 = ~n126 & n3046;
  assign n860 = ~n567 & ~n640;
  assign n2035 = ~n245 & ~n478;
  assign n3048 = n860 & n2035;
  assign n3049 = n3047 & n3048;
  assign n3050 = n294 & ~n630;
  assign n461 = n55 & n119;
  assign n2986 = ~n83 & ~n461;
  assign n3051 = ~n417 & ~n557;
  assign n3052 = n2986 & n3051;
  assign n3053 = n3050 & n3052;
  assign n3054 = n3049 & n3053;
  assign n3055 = n3045 & n3054;
  assign n443 = n50 & n55;
  assign n2813 = ~n443 & ~n843;
  assign n3056 = ~n141 & ~n553;
  assign n659 = n72 & n86;
  assign n3057 = ~n378 & ~n659;
  assign n3058 = n3056 & n3057;
  assign n3059 = ~n170 & ~n217;
  assign n3060 = n3058 & n3059;
  assign n3061 = n2813 & n3060;
  assign n3062 = n3055 & n3061;
  assign n3063 = n2072 & n3062;
  assign n1728 = ~n656 & ~n975;
  assign n1729 = ~n432 & ~n710;
  assign n1730 = ~n503 & n1729;
  assign n1731 = n1728 & n1730;
  assign n1834 = ~n233 & ~n452;
  assign n243 = n55 & n63;
  assign n3064 = ~n243 & ~n1060;
  assign n3065 = n1834 & n3064;
  assign n3066 = n2267 & n3065;
  assign n3067 = n1731 & n3066;
  assign n2808 = ~n51 & ~n173;
  assign n3068 = ~n592 & ~n791;
  assign n3069 = n2808 & n3068;
  assign n3070 = ~n418 & n3069;
  assign n3071 = n3067 & n3070;
  assign n526 = ~n524 & ~n525;
  assign n528 = n526 & ~n527;
  assign n143 = n61 & n142;
  assign n3072 = ~n758 & ~n787;
  assign n3073 = ~n143 & n3072;
  assign n3074 = ~n280 & ~n714;
  assign n98 = n55 & n97;
  assign n3075 = ~n98 & ~n115;
  assign n3076 = n3074 & n3075;
  assign n3077 = n3073 & n3076;
  assign n3078 = n528 & n3077;
  assign n3079 = n3071 & n3078;
  assign n3080 = n3063 & n3079;
  assign n299 = n297 & ~n298;
  assign n302 = ~n300 & ~n301;
  assign n305 = ~n303 & ~n304;
  assign n306 = n302 & n305;
  assign n307 = n299 & n306;
  assign n310 = x23 & n309;
  assign n311 = ~n308 & ~n310;
  assign n315 = ~n313 & ~n314;
  assign n316 = ~n312 & n315;
  assign n317 = n311 & n316;
  assign n318 = n307 & n317;
  assign n320 = n68 & n92;
  assign n321 = ~n319 & ~n320;
  assign n324 = ~n322 & ~n323;
  assign n325 = n321 & n324;
  assign n328 = ~n326 & ~n327;
  assign n329 = n325 & n328;
  assign n332 = ~n330 & ~n331;
  assign n335 = ~n333 & ~n334;
  assign n337 = n55 & n147;
  assign n338 = ~n336 & ~n337;
  assign n339 = n335 & n338;
  assign n340 = n332 & n339;
  assign n341 = n329 & n340;
  assign n342 = n318 & n341;
  assign n343 = n55 & n114;
  assign n345 = ~n343 & ~n344;
  assign n348 = ~n346 & ~n347;
  assign n349 = n345 & n348;
  assign n352 = ~n350 & ~n351;
  assign n355 = ~n353 & ~n354;
  assign n356 = n352 & n355;
  assign n357 = n349 & n356;
  assign n363 = ~n361 & ~n362;
  assign n364 = n360 & n363;
  assign n365 = n357 & n364;
  assign n366 = n342 & n365;
  assign n3097 = n366 & n3096;
  assign n3098 = n3080 & n3097;
  assign n57 = n52 & n56;
  assign n58 = ~n51 & ~n57;
  assign n70 = ~n64 & ~n69;
  assign n71 = n58 & n70;
  assign n80 = ~n74 & ~n79;
  assign n88 = ~n83 & ~n87;
  assign n89 = n80 & n88;
  assign n90 = n71 & n89;
  assign n96 = ~n93 & ~n95;
  assign n100 = ~n98 & ~n99;
  assign n101 = n96 & n100;
  assign n105 = ~n103 & ~n104;
  assign n106 = n101 & n105;
  assign n107 = n90 & n106;
  assign n110 = n68 & n81;
  assign n112 = ~n110 & ~n111;
  assign n113 = ~n109 & n112;
  assign n118 = ~n115 & ~n117;
  assign n120 = n86 & n119;
  assign n123 = ~n120 & ~n122;
  assign n124 = n118 & n123;
  assign n125 = n113 & n124;
  assign n129 = ~n127 & ~n128;
  assign n130 = ~n126 & n129;
  assign n131 = n125 & n130;
  assign n132 = n107 & n131;
  assign n135 = ~n133 & ~n134;
  assign n139 = ~n136 & ~n138;
  assign n140 = n135 & n139;
  assign n144 = ~n141 & ~n143;
  assign n145 = n140 & n144;
  assign n149 = ~n146 & ~n148;
  assign n153 = ~n151 & ~n152;
  assign n154 = n149 & n153;
  assign n157 = ~n155 & ~n156;
  assign n159 = n75 & n158;
  assign n160 = x23 & n159;
  assign n161 = n157 & ~n160;
  assign n162 = n154 & n161;
  assign n167 = n76 & n81;
  assign n168 = ~n166 & ~n167;
  assign n169 = n165 & n168;
  assign n176 = n172 & n175;
  assign n177 = n169 & n176;
  assign n178 = n162 & n177;
  assign n179 = n145 & n178;
  assign n180 = n132 & n179;
  assign n181 = n72 & n81;
  assign n184 = ~n181 & ~n183;
  assign n187 = ~n185 & ~n186;
  assign n188 = n184 & n187;
  assign n191 = ~n189 & ~n190;
  assign n194 = ~n192 & ~n193;
  assign n195 = n191 & n194;
  assign n196 = n188 & n195;
  assign n200 = ~n197 & ~n199;
  assign n203 = ~n201 & ~n202;
  assign n204 = n200 & n203;
  assign n207 = x23 & n206;
  assign n211 = ~n207 & n210;
  assign n212 = n204 & n211;
  assign n213 = n196 & n212;
  assign n220 = ~n216 & n219;
  assign n224 = n220 & n223;
  assign n225 = n213 & n224;
  assign n230 = ~n226 & n229;
  assign n235 = ~n233 & ~n234;
  assign n236 = ~n231 & n235;
  assign n239 = ~n237 & ~n238;
  assign n240 = n236 & n239;
  assign n241 = n230 & n240;
  assign n242 = n225 & n241;
  assign n246 = ~n244 & ~n245;
  assign n247 = ~n243 & n246;
  assign n251 = ~n249 & ~n250;
  assign n252 = ~n248 & n251;
  assign n258 = ~n256 & ~n257;
  assign n259 = n255 & n258;
  assign n260 = n252 & n259;
  assign n261 = n247 & n260;
  assign n264 = ~n262 & ~n263;
  assign n265 = n63 & n73;
  assign n266 = n81 & n137;
  assign n267 = ~n265 & ~n266;
  assign n268 = n264 & n267;
  assign n271 = ~n269 & ~n270;
  assign n274 = ~n272 & ~n273;
  assign n275 = n271 & n274;
  assign n276 = n268 & n275;
  assign n282 = ~n280 & ~n281;
  assign n284 = n61 & n85;
  assign n285 = ~n283 & ~n284;
  assign n286 = n282 & n285;
  assign n287 = n279 & n286;
  assign n288 = n276 & n287;
  assign n289 = n261 & n288;
  assign n290 = n242 & n289;
  assign n291 = n180 & n290;
  assign n367 = n294 & n366;
  assign n368 = n291 & n367;
  assign n371 = ~n57 & ~n370;
  assign n372 = ~n369 & n371;
  assign n377 = n374 & n376;
  assign n379 = ~n95 & ~n378;
  assign n380 = n377 & n379;
  assign n382 = n81 & n102;
  assign n383 = ~n227 & ~n382;
  assign n384 = n381 & n383;
  assign n387 = n384 & n386;
  assign n388 = n380 & n387;
  assign n389 = n372 & n388;
  assign n391 = ~n333 & ~n390;
  assign n393 = ~n262 & ~n392;
  assign n394 = ~n280 & n393;
  assign n395 = n391 & n394;
  assign n397 = ~n209 & ~n319;
  assign n398 = ~n396 & n397;
  assign n399 = ~n216 & ~n283;
  assign n400 = n398 & n399;
  assign n401 = n395 & n400;
  assign n408 = n404 & n407;
  assign n413 = ~n320 & ~n412;
  assign n414 = n411 & n413;
  assign n415 = n408 & n414;
  assign n419 = ~n417 & ~n418;
  assign n420 = ~n416 & n419;
  assign n421 = n415 & n420;
  assign n422 = n401 & n421;
  assign n423 = n389 & n422;
  assign n425 = ~n245 & ~n424;
  assign n426 = ~n248 & ~n326;
  assign n427 = n425 & n426;
  assign n430 = ~n428 & ~n429;
  assign n431 = n427 & n430;
  assign n433 = ~n346 & ~n432;
  assign n434 = ~n222 & n433;
  assign n435 = n431 & n434;
  assign n436 = n423 & n435;
  assign n438 = ~n199 & n437;
  assign n444 = ~n442 & ~n443;
  assign n446 = n444 & n445;
  assign n447 = n441 & n446;
  assign n448 = n438 & n447;
  assign n450 = ~n155 & ~n449;
  assign n451 = ~n87 & n450;
  assign n453 = ~n103 & ~n452;
  assign n454 = ~n303 & n453;
  assign n455 = n451 & n454;
  assign n459 = ~n133 & ~n458;
  assign n460 = n457 & n459;
  assign n462 = ~n166 & ~n461;
  assign n464 = ~n254 & ~n463;
  assign n465 = n462 & n464;
  assign n466 = n460 & n465;
  assign n467 = n455 & n466;
  assign n468 = n448 & n467;
  assign n472 = ~n469 & ~n471;
  assign n474 = n472 & n473;
  assign n477 = ~n475 & ~n476;
  assign n479 = ~n174 & ~n478;
  assign n480 = n477 & n479;
  assign n481 = n474 & n480;
  assign n483 = ~n186 & ~n263;
  assign n484 = n482 & n483;
  assign n485 = ~n98 & ~n197;
  assign n486 = ~n110 & ~n192;
  assign n487 = n485 & n486;
  assign n488 = n484 & n487;
  assign n489 = n481 & n488;
  assign n490 = n468 & n489;
  assign n491 = n436 & n490;
  assign n493 = ~n327 & ~n492;
  assign n495 = ~n243 & ~n494;
  assign n496 = n493 & n495;
  assign n498 = ~n231 & ~n497;
  assign n501 = n498 & ~n500;
  assign n502 = n496 & n501;
  assign n505 = ~n503 & ~n504;
  assign n507 = ~n234 & ~n506;
  assign n508 = n505 & n507;
  assign n510 = ~n273 & ~n509;
  assign n511 = ~n69 & n510;
  assign n512 = n508 & n511;
  assign n513 = n502 & n512;
  assign n515 = ~n189 & ~n514;
  assign n516 = ~n183 & n515;
  assign n519 = ~n517 & ~n518;
  assign n520 = ~n221 & ~n281;
  assign n521 = n519 & n520;
  assign n522 = n516 & n521;
  assign n523 = n513 & n522;
  assign n530 = ~n164 & ~n529;
  assign n532 = ~n334 & ~n531;
  assign n533 = n530 & n532;
  assign n534 = n528 & n533;
  assign n537 = ~n535 & n536;
  assign n538 = n534 & n537;
  assign n539 = n523 & n538;
  assign n542 = ~n111 & ~n541;
  assign n543 = ~n540 & n542;
  assign n545 = ~n217 & ~n544;
  assign n546 = ~n109 & ~n322;
  assign n547 = n545 & n546;
  assign n548 = n543 & n547;
  assign n551 = ~n549 & ~n550;
  assign n554 = ~n552 & ~n553;
  assign n555 = n551 & n554;
  assign n556 = n548 & n555;
  assign n559 = ~n557 & ~n558;
  assign n561 = ~n296 & ~n560;
  assign n562 = n559 & n561;
  assign n563 = ~n298 & n562;
  assign n564 = n556 & n563;
  assign n565 = n539 & n564;
  assign n566 = n491 & n565;
  assign n568 = ~n185 & ~n567;
  assign n569 = ~n192 & n568;
  assign n571 = ~n152 & ~n504;
  assign n572 = n570 & n571;
  assign n573 = n569 & n572;
  assign n577 = ~n201 & ~n576;
  assign n578 = ~n254 & ~n354;
  assign n579 = n577 & n578;
  assign n580 = n573 & n579;
  assign n581 = ~n245 & ~n304;
  assign n583 = ~n262 & ~n582;
  assign n585 = n583 & n584;
  assign n586 = n581 & n585;
  assign n587 = n580 & n586;
  assign n589 = ~n167 & ~n424;
  assign n590 = ~n588 & n589;
  assign n591 = ~n218 & ~n303;
  assign n594 = ~n592 & ~n593;
  assign n595 = n591 & n594;
  assign n596 = n590 & n595;
  assign n598 = ~n133 & ~n440;
  assign n599 = n597 & n598;
  assign n600 = n596 & n599;
  assign n601 = ~n57 & ~n418;
  assign n603 = ~n79 & n602;
  assign n604 = n601 & n603;
  assign n605 = n81 & n182;
  assign n606 = ~n284 & ~n605;
  assign n607 = n604 & n606;
  assign n608 = n600 & n607;
  assign n609 = n587 & n608;
  assign n613 = ~n492 & ~n612;
  assign n614 = ~n544 & n613;
  assign n615 = n611 & n614;
  assign n616 = n50 & n73;
  assign n618 = ~n616 & ~n617;
  assign n619 = n53 & n108;
  assign n620 = n49 & n619;
  assign n624 = ~n620 & ~n623;
  assign n625 = n618 & n624;
  assign n626 = n615 & n625;
  assign n629 = ~n627 & ~n628;
  assign n631 = ~n557 & ~n630;
  assign n632 = n251 & n631;
  assign n633 = n629 & n632;
  assign n636 = ~n343 & n635;
  assign n637 = n633 & n636;
  assign n638 = n626 & n637;
  assign n639 = n609 & n638;
  assign n641 = ~n503 & ~n640;
  assign n643 = x26 ^ x25;
  assign n644 = n642 & n643;
  assign n645 = n641 & ~n644;
  assign n648 = ~n313 & ~n647;
  assign n649 = n645 & n648;
  assign n650 = ~n308 & ~n405;
  assign n651 = ~n461 & n650;
  assign n653 = n651 & ~n652;
  assign n654 = n649 & n653;
  assign n658 = ~n656 & n657;
  assign n661 = ~n266 & ~n660;
  assign n662 = ~n659 & n661;
  assign n663 = n658 & n662;
  assign n664 = n654 & n663;
  assign n665 = ~n51 & ~n244;
  assign n667 = n665 & ~n666;
  assign n668 = ~n181 & ~n361;
  assign n669 = ~n265 & n668;
  assign n670 = n667 & n669;
  assign n672 = ~n300 & ~n671;
  assign n673 = ~n171 & ~n406;
  assign n674 = n672 & n673;
  assign n677 = n674 & n676;
  assign n678 = n670 & n677;
  assign n679 = ~n527 & ~n558;
  assign n681 = ~n475 & ~n680;
  assign n682 = n679 & n681;
  assign n684 = ~n369 & ~n683;
  assign n685 = ~n443 & n684;
  assign n686 = n682 & n685;
  assign n688 = n332 & ~n687;
  assign n692 = ~n689 & ~n691;
  assign n693 = n688 & n692;
  assign n694 = n686 & n693;
  assign n695 = n678 & n694;
  assign n696 = n664 & n695;
  assign n697 = ~n189 & ~n403;
  assign n698 = ~n143 & n697;
  assign n700 = ~x29 & n699;
  assign n701 = n698 & ~n700;
  assign n702 = ~n351 & ~n535;
  assign n703 = ~n197 & ~n353;
  assign n704 = n702 & n703;
  assign n705 = n701 & n704;
  assign n706 = ~n136 & ~n301;
  assign n707 = n279 & n706;
  assign n708 = n705 & n707;
  assign n711 = ~n709 & ~n710;
  assign n712 = ~n69 & n711;
  assign n713 = ~n410 & ~n552;
  assign n715 = ~n525 & ~n714;
  assign n716 = n713 & n715;
  assign n717 = n712 & n716;
  assign n718 = ~n93 & ~n269;
  assign n719 = ~n346 & n718;
  assign n720 = n717 & n719;
  assign n721 = ~n104 & n551;
  assign n722 = ~n134 & ~n327;
  assign n724 = ~n208 & ~n723;
  assign n725 = n722 & n724;
  assign n726 = n721 & n725;
  assign n728 = ~n110 & ~n248;
  assign n729 = n727 & n728;
  assign n730 = n726 & n729;
  assign n731 = n720 & n730;
  assign n732 = n708 & n731;
  assign n733 = n696 & n732;
  assign n734 = n639 & n733;
  assign n735 = x24 ^ x23;
  assign n736 = n159 & ~n735;
  assign n737 = ~n263 & ~n736;
  assign n738 = ~n199 & ~n527;
  assign n739 = n737 & n738;
  assign n741 = ~n233 & ~n740;
  assign n742 = ~n277 & n741;
  assign n743 = n116 & n690;
  assign n744 = ~n497 & ~n743;
  assign n745 = ~n248 & n744;
  assign n746 = n742 & n745;
  assign n747 = n739 & n746;
  assign n748 = ~n331 & ~n659;
  assign n749 = n629 & n748;
  assign n752 = ~n750 & ~n751;
  assign n753 = n749 & n752;
  assign n754 = n747 & n753;
  assign n756 = ~n417 & ~n440;
  assign n757 = ~n755 & n756;
  assign n759 = ~n249 & ~n758;
  assign n760 = n757 & n759;
  assign n764 = ~n163 & ~n336;
  assign n765 = ~n763 & n764;
  assign n766 = ~n231 & ~n303;
  assign n767 = n765 & n766;
  assign n768 = n760 & n767;
  assign n769 = ~n127 & n302;
  assign n770 = n651 & n769;
  assign n771 = ~n115 & ~n593;
  assign n772 = n770 & n771;
  assign n773 = n768 & n772;
  assign n774 = n754 & n773;
  assign n775 = ~n506 & ~n723;
  assign n776 = ~n243 & n775;
  assign n777 = n372 & n776;
  assign n778 = ~n189 & ~n612;
  assign n779 = ~n558 & ~n671;
  assign n780 = n778 & n779;
  assign n782 = ~n122 & ~n514;
  assign n783 = n781 & n782;
  assign n784 = n780 & n783;
  assign n785 = n777 & n784;
  assign n786 = ~n442 & ~n552;
  assign n788 = ~n87 & ~n787;
  assign n789 = n786 & n788;
  assign n792 = ~n790 & ~n791;
  assign n793 = n184 & n792;
  assign n794 = n789 & n793;
  assign n795 = n785 & n794;
  assign n798 = ~n298 & ~n797;
  assign n801 = ~n799 & ~n800;
  assign n802 = ~n228 & ~n322;
  assign n803 = n801 & n802;
  assign n804 = n798 & n803;
  assign n805 = ~n69 & ~n323;
  assign n806 = ~n333 & n805;
  assign n807 = ~n409 & ~n575;
  assign n808 = ~n244 & n807;
  assign n809 = n806 & n808;
  assign n810 = n804 & n809;
  assign n811 = ~n208 & ~n592;
  assign n813 = n811 & ~n812;
  assign n814 = ~n158 & ~n262;
  assign n815 = ~x26 & n49;
  assign n816 = ~n814 & n815;
  assign n818 = x23 & n817;
  assign n819 = n121 & n818;
  assign n820 = ~n452 & ~n819;
  assign n821 = ~n816 & n820;
  assign n822 = n813 & n821;
  assign n823 = n810 & n822;
  assign n824 = n795 & n823;
  assign n825 = n774 & n824;
  assign n827 = ~n656 & ~n826;
  assign n831 = n827 & n830;
  assign n832 = n145 & n831;
  assign n833 = ~n362 & ~n518;
  assign n834 = ~n64 & ~n492;
  assign n835 = n833 & n834;
  assign n836 = ~n151 & ~n295;
  assign n837 = n835 & n836;
  assign n838 = ~n353 & ~n529;
  assign n839 = ~n186 & ~n463;
  assign n840 = n838 & n839;
  assign n845 = n842 & n844;
  assign n846 = n840 & n845;
  assign n847 = n837 & n846;
  assign n848 = n832 & n847;
  assign n849 = ~n560 & n848;
  assign n851 = ~n541 & ~n850;
  assign n852 = ~n167 & ~n504;
  assign n853 = n851 & n852;
  assign n854 = ~n269 & ~n313;
  assign n855 = n853 & n854;
  assign n856 = ~n126 & ~n666;
  assign n857 = ~n120 & ~n164;
  assign n858 = n856 & n857;
  assign n861 = n859 & n860;
  assign n862 = n858 & n861;
  assign n863 = n855 & n862;
  assign n864 = ~n402 & ~n709;
  assign n865 = ~n382 & n864;
  assign n866 = ~n326 & ~n361;
  assign n867 = n865 & n866;
  assign n869 = ~n292 & ~n320;
  assign n870 = n868 & n869;
  assign n871 = n867 & n870;
  assign n872 = n863 & n871;
  assign n873 = ~n509 & ~n549;
  assign n874 = ~n256 & n873;
  assign n875 = ~n358 & ~n680;
  assign n876 = n874 & n875;
  assign n877 = ~n312 & ~n330;
  assign n878 = ~n683 & n877;
  assign n879 = n876 & n878;
  assign n880 = n872 & n879;
  assign n881 = n849 & n880;
  assign n882 = n825 & n881;
  assign n883 = ~n358 & ~n616;
  assign n885 = n883 & n884;
  assign n886 = ~n280 & ~n416;
  assign n887 = ~n592 & n886;
  assign n888 = n885 & n887;
  assign n890 = ~n326 & ~n529;
  assign n891 = n889 & n890;
  assign n892 = ~n346 & ~n557;
  assign n894 = n892 & n893;
  assign n895 = n891 & n894;
  assign n896 = n888 & n895;
  assign n906 = n246 & ~n791;
  assign n907 = n219 & n906;
  assign n908 = n905 & n907;
  assign n909 = n896 & n908;
  assign n910 = n107 & n909;
  assign n911 = ~n283 & ~n723;
  assign n912 = ~n330 & ~n503;
  assign n913 = ~n354 & n912;
  assign n914 = n911 & n913;
  assign n916 = n914 & n915;
  assign n917 = ~n541 & n916;
  assign n918 = n910 & n917;
  assign n921 = ~n919 & ~n920;
  assign n922 = ~n443 & ~n799;
  assign n923 = n921 & n922;
  assign n924 = n230 & n923;
  assign n925 = ~n687 & ~n850;
  assign n926 = n713 & n925;
  assign n927 = n924 & n926;
  assign n930 = ~n928 & ~n929;
  assign n932 = n930 & n931;
  assign n933 = ~n128 & n932;
  assign n934 = ~n284 & ~n456;
  assign n935 = ~n152 & ~n164;
  assign n936 = n934 & n935;
  assign n938 = n172 & n937;
  assign n939 = n936 & n938;
  assign n940 = n933 & n939;
  assign n941 = n927 & n940;
  assign n942 = n918 & n941;
  assign n943 = ~n234 & ~n314;
  assign n944 = ~n120 & ~n378;
  assign n945 = n943 & n944;
  assign n947 = ~n475 & ~n946;
  assign n950 = n947 & n949;
  assign n951 = n945 & n950;
  assign n952 = n611 & ~n826;
  assign n953 = n951 & n952;
  assign n954 = ~n109 & n157;
  assign n956 = n954 & n955;
  assign n957 = ~n143 & ~n428;
  assign n958 = n956 & n957;
  assign n959 = n953 & n958;
  assign n960 = n297 & ~n402;
  assign n961 = ~n424 & ~n843;
  assign n962 = ~n269 & n961;
  assign n963 = n960 & n962;
  assign n964 = ~n192 & ~n514;
  assign n965 = ~n494 & n964;
  assign n966 = n321 & n965;
  assign n967 = n963 & n966;
  assign n968 = n959 & n967;
  assign n969 = n774 & n968;
  assign n970 = n942 & n969;
  assign n971 = ~n269 & ~n281;
  assign n972 = ~n610 & n971;
  assign n973 = ~n155 & ~n333;
  assign n974 = n972 & n973;
  assign n977 = n974 & n976;
  assign n978 = ~n167 & ~n671;
  assign n979 = ~n263 & n978;
  assign n980 = ~n57 & n979;
  assign n981 = n977 & n980;
  assign n982 = ~n418 & ~n797;
  assign n983 = ~n396 & ~n680;
  assign n984 = n982 & n983;
  assign n985 = ~n750 & n833;
  assign n986 = ~n549 & ~n617;
  assign n987 = n985 & n986;
  assign n988 = n984 & n987;
  assign n989 = ~n456 & ~n630;
  assign n990 = ~n98 & ~n250;
  assign n991 = n989 & n990;
  assign n992 = ~n375 & ~n841;
  assign n993 = n991 & n992;
  assign n994 = ~n337 & ~n506;
  assign n995 = ~n620 & n994;
  assign n996 = n993 & n995;
  assign n997 = n988 & n996;
  assign n998 = n981 & n997;
  assign n1000 = ~n181 & n999;
  assign n1001 = ~n248 & ~n458;
  assign n1002 = n1000 & n1001;
  assign n1003 = ~n185 & ~n850;
  assign n1004 = ~n272 & n1003;
  assign n1006 = n302 & ~n1005;
  assign n1007 = n1004 & n1006;
  assign n1008 = n1002 & n1007;
  assign n1009 = n581 & ~n623;
  assign n1010 = ~n111 & ~n370;
  assign n1011 = n1009 & n1010;
  assign n1012 = n1008 & n1011;
  assign n1013 = n998 & n1012;
  assign n1014 = ~n120 & ~n675;
  assign n1015 = ~n266 & ~n361;
  assign n1016 = n1014 & n1015;
  assign n1017 = ~n233 & ~n313;
  assign n1018 = n1016 & n1017;
  assign n1019 = ~n312 & ~n529;
  assign n1020 = ~n392 & n1019;
  assign n1022 = ~n283 & ~n687;
  assign n1023 = n1021 & n1022;
  assign n1024 = n1020 & n1023;
  assign n1025 = n1018 & n1024;
  assign n1026 = ~n790 & ~n901;
  assign n1027 = ~n787 & n1026;
  assign n1028 = n1025 & n1027;
  assign n1029 = ~n226 & ~n531;
  assign n1030 = ~n173 & ~n432;
  assign n1031 = n1029 & n1030;
  assign n1032 = ~n238 & ~n452;
  assign n1033 = ~n217 & ~n478;
  assign n1034 = n1032 & n1033;
  assign n1035 = n1031 & n1034;
  assign n1036 = ~n428 & ~n443;
  assign n1037 = ~n405 & n1036;
  assign n1038 = n1035 & n1037;
  assign n1039 = ~n253 & ~n525;
  assign n1040 = ~n647 & n1039;
  assign n1041 = ~n152 & ~n755;
  assign n1042 = n1040 & n1041;
  assign n1043 = ~n83 & ~n463;
  assign n1044 = ~n273 & ~n494;
  assign n1045 = n1043 & n1044;
  assign n1046 = ~n243 & ~n449;
  assign n1048 = ~n440 & ~n1047;
  assign n1049 = n1046 & n1048;
  assign n1050 = n1045 & n1049;
  assign n1051 = n1042 & n1050;
  assign n1052 = n1038 & n1051;
  assign n1053 = n1028 & n1052;
  assign n1054 = n1013 & n1053;
  assign n1097 = n1054 & n1096;
  assign n1098 = n882 & n1097;
  assign n1099 = ~n970 & ~n1098;
  assign n1100 = ~n170 & ~n758;
  assign n1101 = ~n475 & ~n531;
  assign n1102 = n1100 & n1101;
  assign n1104 = ~n262 & n1103;
  assign n1105 = n1102 & n1104;
  assign n1106 = n651 & n1069;
  assign n1107 = n1105 & n1106;
  assign n1110 = ~n1108 & ~n1109;
  assign n1111 = n55 & ~n1110;
  assign n1112 = ~n263 & ~n799;
  assign n1113 = ~n1111 & n1112;
  assign n1114 = n667 & n1113;
  assign n1115 = n1107 & n1114;
  assign n1116 = ~n277 & ~n503;
  assign n1117 = ~n517 & n1116;
  assign n1118 = n1004 & n1117;
  assign n1119 = ~n201 & ~n478;
  assign n1120 = ~n141 & ~n249;
  assign n1121 = n1119 & n1120;
  assign n1122 = n1118 & n1121;
  assign n1123 = n1115 & n1122;
  assign n1124 = ~n237 & ~n385;
  assign n1125 = ~n544 & n1124;
  assign n1126 = ~n117 & ~n630;
  assign n1127 = ~n390 & n1126;
  assign n1128 = n1125 & n1127;
  assign n1129 = ~n428 & ~n689;
  assign n1130 = ~n343 & ~n567;
  assign n1131 = n1129 & n1130;
  assign n1132 = n1128 & n1131;
  assign n1133 = ~n238 & n883;
  assign n1134 = ~n588 & ~n709;
  assign n1136 = n1134 & ~n1135;
  assign n1137 = n1133 & n1136;
  assign n1138 = n1132 & n1137;
  assign n1139 = n1123 & n1138;
  assign n1140 = ~n605 & ~n797;
  assign n1141 = ~n659 & ~n710;
  assign n1142 = ~n202 & n1141;
  assign n1143 = n1140 & n1142;
  assign n1144 = ~n83 & ~n620;
  assign n1145 = n1143 & n1144;
  assign n1146 = ~n409 & ~n675;
  assign n1147 = ~n336 & n1146;
  assign n1148 = n121 & n499;
  assign n1149 = ~n841 & ~n1148;
  assign n1150 = ~n231 & n1149;
  assign n1151 = n1147 & n1150;
  assign n1152 = n1145 & n1151;
  assign n1157 = n1154 & n1156;
  assign n1159 = ~n278 & n1158;
  assign n1160 = ~n233 & ~n392;
  assign n1161 = ~n110 & n1160;
  assign n1162 = n1159 & n1161;
  assign n1163 = n1157 & n1162;
  assign n1165 = ~n518 & n1164;
  assign n1167 = ~n375 & ~n1166;
  assign n1168 = ~n313 & ~n946;
  assign n1169 = n1167 & n1168;
  assign n1170 = n1165 & n1169;
  assign n1171 = ~n549 & ~n1005;
  assign n1172 = ~n283 & ~n750;
  assign n1173 = n1171 & n1172;
  assign n1174 = n892 & n1173;
  assign n1175 = n1170 & n1174;
  assign n1176 = n1163 & n1175;
  assign n1177 = n1152 & n1176;
  assign n1178 = n1139 & n1177;
  assign n1179 = n828 & n1075;
  assign n1180 = ~n181 & ~n256;
  assign n1181 = n482 & n1180;
  assign n1182 = n1179 & n1181;
  assign n1184 = ~n378 & n1183;
  assign n1185 = n1182 & n1184;
  assign n1186 = ~n660 & ~n671;
  assign n1187 = n149 & n1186;
  assign n1188 = ~n250 & ~n253;
  assign n1189 = n1187 & n1188;
  assign n1190 = n1185 & n1189;
  assign n1191 = ~n592 & ~n1047;
  assign n1192 = ~n74 & ~n163;
  assign n1193 = n1191 & n1192;
  assign n1194 = ~n126 & ~n612;
  assign n1195 = ~n442 & n1194;
  assign n1196 = n1193 & n1195;
  assign n1198 = ~n627 & n1197;
  assign n1199 = ~n136 & ~n740;
  assign n1200 = ~n687 & n1199;
  assign n1201 = n1198 & n1200;
  assign n1202 = n1196 & n1201;
  assign n1203 = n705 & n1202;
  assign n1204 = n1190 & n1203;
  assign n1205 = ~n326 & ~n751;
  assign n1206 = n1072 & n1205;
  assign n1207 = n1204 & n1206;
  assign n1208 = n1178 & n1207;
  assign n1209 = ~n346 & ~n424;
  assign n1210 = ~n227 & ~n403;
  assign n1211 = n1209 & n1210;
  assign n1212 = ~n127 & ~n920;
  assign n1213 = n1211 & n1212;
  assign n1214 = ~n79 & ~n273;
  assign n1216 = n1214 & ~n1215;
  assign n1217 = ~n417 & ~n552;
  assign n1218 = n462 & n1217;
  assign n1219 = n1216 & n1218;
  assign n1220 = n1213 & n1219;
  assign n1221 = ~n117 & ~n948;
  assign n1222 = n391 & n1221;
  assign n1223 = ~n378 & n1222;
  assign n1224 = n1220 & n1223;
  assign n1225 = ~n167 & ~n458;
  assign n1226 = n441 & n1225;
  assign n1228 = ~n549 & ~n1227;
  assign n1229 = n911 & n1228;
  assign n1230 = n1226 & n1229;
  assign n1231 = ~n370 & ~n385;
  assign n1232 = ~n456 & n1231;
  assign n1233 = n813 & n1232;
  assign n1234 = n1230 & n1233;
  assign n1235 = n1224 & n1234;
  assign n1236 = ~n98 & ~n141;
  assign n1237 = n801 & n1236;
  assign n1238 = ~n612 & ~n714;
  assign n1239 = n1237 & n1238;
  assign n1242 = n1239 & n1241;
  assign n1243 = ~n155 & ~n541;
  assign n1244 = ~n257 & n1243;
  assign n1245 = ~n269 & ~n605;
  assign n1246 = n1043 & n1245;
  assign n1247 = n1244 & n1246;
  assign n1248 = n1242 & n1247;
  assign n1249 = n1235 & n1248;
  assign n1250 = ~n111 & ~n675;
  assign n1251 = ~n192 & ~n373;
  assign n1252 = n1250 & n1251;
  assign n1253 = ~n666 & ~n1135;
  assign n1254 = ~n755 & n1253;
  assign n1255 = n1252 & n1254;
  assign n1256 = ~n336 & ~n412;
  assign n1257 = n727 & n1256;
  assign n1258 = ~n126 & ~n790;
  assign n1259 = ~n109 & ~n416;
  assign n1260 = n1258 & n1259;
  assign n1261 = n1257 & n1260;
  assign n1262 = n1255 & n1261;
  assign n1263 = ~n544 & ~n797;
  assign n1264 = ~n410 & ~n535;
  assign n1265 = n1263 & n1264;
  assign n1267 = ~n254 & ~n1266;
  assign n1268 = n728 & n1267;
  assign n1269 = n1265 & n1268;
  assign n1270 = n1262 & n1269;
  assign n1271 = ~n337 & n437;
  assign n1272 = n960 & n1271;
  assign n1273 = ~n284 & ~n375;
  assign n1274 = ~n209 & ~n628;
  assign n1275 = n1273 & n1274;
  assign n1276 = ~n432 & n530;
  assign n1277 = n1275 & n1276;
  assign n1278 = n1272 & n1277;
  assign n1279 = n1270 & n1278;
  assign n1280 = ~n449 & ~n928;
  assign n1281 = ~n148 & ~n303;
  assign n1282 = n1280 & n1281;
  assign n1283 = ~n193 & ~n751;
  assign n1284 = ~n975 & n1283;
  assign n1285 = n1282 & n1284;
  assign n1286 = ~n143 & ~n354;
  assign n1287 = n947 & n1286;
  assign n1288 = ~n146 & ~n151;
  assign n1289 = n672 & n1288;
  assign n1290 = n1287 & n1289;
  assign n1291 = n1285 & n1290;
  assign n1292 = ~n216 & n1141;
  assign n1293 = n96 & ~n567;
  assign n1294 = n1292 & n1293;
  assign n1295 = ~n469 & ~n494;
  assign n1296 = ~n233 & n1295;
  assign n1297 = n1294 & n1296;
  assign n1298 = n1291 & n1297;
  assign n1300 = ~n351 & n1299;
  assign n1303 = n1301 & n1302;
  assign n1304 = n1300 & n1303;
  assign n1306 = ~n322 & ~n1166;
  assign n1307 = n1305 & n1306;
  assign n1308 = n453 & n526;
  assign n1309 = n1307 & n1308;
  assign n1310 = n1304 & n1309;
  assign n1311 = ~n280 & ~n334;
  assign n1312 = ~n163 & ~n190;
  assign n1313 = n1311 & n1312;
  assign n1314 = ~n429 & ~n709;
  assign n1315 = n1313 & n1314;
  assign n1316 = n1310 & n1315;
  assign n1317 = n1298 & n1316;
  assign n1318 = n1279 & n1317;
  assign n1319 = n1249 & n1318;
  assign n1320 = ~n1208 & ~n1319;
  assign n1321 = ~n882 & ~n1097;
  assign n1322 = n1320 & n1321;
  assign n1323 = ~n1099 & ~n1322;
  assign n1324 = ~n390 & ~n560;
  assign n1325 = ~n166 & n1324;
  assign n1326 = ~n249 & ~n627;
  assign n1327 = n1325 & n1326;
  assign n1328 = ~n155 & ~n723;
  assign n1329 = ~n254 & n1328;
  assign n1330 = ~n898 & n1329;
  assign n1331 = n1327 & n1330;
  assign n1333 = ~n126 & n1332;
  assign n1334 = n1331 & n1333;
  assign n1336 = ~n281 & ~n452;
  assign n1337 = ~n292 & n1336;
  assign n1338 = n1335 & n1337;
  assign n1339 = n618 & n1338;
  assign n1340 = n1334 & n1339;
  assign n1341 = ~n506 & n851;
  assign n1342 = ~n138 & ~n449;
  assign n1343 = n1341 & n1342;
  assign n1344 = ~n475 & ~n787;
  assign n1346 = ~n344 & ~n1345;
  assign n1347 = n1344 & n1346;
  assign n1348 = ~n117 & ~n361;
  assign n1349 = ~n634 & n1348;
  assign n1350 = n1347 & n1349;
  assign n1351 = n1343 & n1350;
  assign n1355 = n1351 & n1354;
  assign n1356 = ~n343 & ~n417;
  assign n1357 = n47 & n621;
  assign n1358 = n1356 & ~n1357;
  assign n1359 = ~n257 & ~n640;
  assign n1360 = ~n370 & ~n509;
  assign n1361 = n1359 & n1360;
  assign n1362 = n1358 & n1361;
  assign n1363 = ~n593 & ~n901;
  assign n1364 = n1362 & n1363;
  assign n1365 = ~n331 & ~n544;
  assign n1366 = ~n99 & n1365;
  assign n1367 = n1286 & n1366;
  assign n1368 = ~n478 & ~n656;
  assign n1369 = n1367 & n1368;
  assign n1370 = n1364 & n1369;
  assign n1371 = n1355 & n1370;
  assign n1372 = n1340 & n1371;
  assign n1373 = ~n173 & ~n265;
  assign n1374 = ~n463 & n1373;
  assign n1375 = ~n128 & ~n975;
  assign n1376 = n1374 & n1375;
  assign n1377 = ~n134 & ~n406;
  assign n1378 = ~n812 & ~n1266;
  assign n1379 = n1377 & n1378;
  assign n1380 = ~n322 & ~n418;
  assign n1381 = ~n79 & ~n248;
  assign n1382 = n1380 & n1381;
  assign n1383 = n1379 & n1382;
  assign n1384 = n1376 & n1383;
  assign n1385 = ~n120 & ~n319;
  assign n1386 = n78 & n215;
  assign n1387 = ~n266 & ~n1386;
  assign n1388 = n1385 & n1387;
  assign n1389 = ~n234 & ~n540;
  assign n1390 = ~n410 & ~n948;
  assign n1391 = n1389 & n1390;
  assign n1392 = n1388 & n1391;
  assign n1393 = n1384 & n1392;
  assign n1394 = ~n476 & ~n525;
  assign n1395 = ~n527 & ~n683;
  assign n1396 = n1394 & n1395;
  assign n1397 = n220 & n1396;
  assign n1398 = ~n111 & n1225;
  assign n1399 = n1397 & n1398;
  assign n1400 = n425 & n930;
  assign n1401 = ~n327 & ~n440;
  assign n1402 = n828 & n1401;
  assign n1403 = n1400 & n1402;
  assign n1404 = ~n97 & ~n182;
  assign n1405 = n61 & ~n1404;
  assign n1406 = ~n95 & ~n612;
  assign n1407 = ~n1405 & n1406;
  assign n1408 = n536 & n893;
  assign n1409 = n1407 & n1408;
  assign n1410 = n1403 & n1409;
  assign n1411 = n1399 & n1410;
  assign n1412 = n1393 & n1411;
  assign n1413 = n1177 & n1412;
  assign n1414 = n1372 & n1413;
  assign n1415 = ~n970 & ~n1208;
  assign n1416 = ~n1321 & ~n1415;
  assign n1417 = ~n1414 & ~n1416;
  assign n1418 = n1323 & ~n1417;
  assign n1419 = ~n882 & ~n1418;
  assign n1420 = n734 & ~n1419;
  assign n1421 = ~n207 & ~n461;
  assign n1422 = ~n183 & ~n331;
  assign n1423 = n1421 & n1422;
  assign n1424 = ~n122 & ~n257;
  assign n1425 = n1423 & n1424;
  assign n1426 = ~n588 & ~n1047;
  assign n1427 = ~n254 & ~n334;
  assign n1428 = n1426 & n1427;
  assign n1429 = ~n109 & ~n143;
  assign n1430 = ~n69 & ~n1227;
  assign n1431 = n1429 & n1430;
  assign n1432 = n1428 & n1431;
  assign n1433 = n1425 & n1432;
  assign n1434 = ~n524 & ~n1135;
  assign n1435 = n1231 & n1434;
  assign n1436 = ~n346 & n1435;
  assign n1437 = n1433 & n1436;
  assign n1438 = ~n138 & ~n901;
  assign n1439 = n697 & n1438;
  assign n1440 = ~n358 & ~n527;
  assign n1441 = n1274 & n1440;
  assign n1442 = n1439 & n1441;
  assign n1443 = n1031 & n1442;
  assign n1444 = ~n322 & ~n755;
  assign n1445 = ~n850 & n1444;
  assign n1446 = n995 & n1445;
  assign n1447 = n1443 & n1446;
  assign n1448 = ~n390 & ~n841;
  assign n1449 = n890 & n1448;
  assign n1450 = ~n160 & n1449;
  assign n1451 = ~n128 & n1061;
  assign n1452 = n1117 & n1451;
  assign n1453 = n1450 & n1452;
  assign n1454 = ~n416 & ~n642;
  assign n1455 = n844 & n1454;
  assign n1456 = ~n284 & n294;
  assign n1457 = n1455 & n1456;
  assign n1458 = ~n378 & ~n791;
  assign n1459 = ~n156 & n1458;
  assign n1460 = ~n458 & ~n525;
  assign n1461 = n1459 & n1460;
  assign n1462 = n1457 & n1461;
  assign n1463 = n1453 & n1462;
  assign n1464 = n1447 & n1463;
  assign n1465 = n1437 & n1464;
  assign n1466 = x23 & ~n817;
  assign n1468 = ~x26 & ~n1467;
  assign n1469 = ~n1466 & n1468;
  assign n1473 = ~n1469 & ~n1472;
  assign n1474 = n86 & ~n1473;
  assign n1476 = ~x24 & ~x26;
  assign n1477 = ~n1475 & ~n1476;
  assign n1478 = n47 & ~n1477;
  assign n1479 = n214 & ~n643;
  assign n1480 = ~n1478 & ~n1479;
  assign n1481 = ~n1474 & n1480;
  assign n1483 = ~n141 & ~n449;
  assign n1484 = ~n1482 & n1483;
  assign n1485 = ~n272 & ~n314;
  assign n1486 = n973 & n1485;
  assign n1487 = n1484 & n1486;
  assign n1488 = n1481 & n1487;
  assign n1489 = ~n250 & ~n560;
  assign n1490 = ~n442 & n1489;
  assign n1491 = ~n353 & ~n948;
  assign n1492 = ~n494 & ~n689;
  assign n1493 = n1491 & n1492;
  assign n1494 = n1490 & n1493;
  assign n1495 = n1488 & n1494;
  assign n1496 = ~n666 & ~n799;
  assign n1497 = ~n281 & n1496;
  assign n1498 = ~n164 & n1314;
  assign n1499 = n1497 & n1498;
  assign n1502 = x23 & ~n1501;
  assign n1503 = ~n817 & ~n1502;
  assign n1504 = ~x23 & x26;
  assign n1505 = n94 & ~n1504;
  assign n1506 = ~n1503 & n1505;
  assign n1509 = ~n134 & ~n687;
  assign n1510 = ~n1508 & n1509;
  assign n1511 = ~n1506 & n1510;
  assign n1512 = n1499 & n1511;
  assign n1513 = ~n359 & ~n656;
  assign n1514 = ~n248 & ~n283;
  assign n1515 = ~n170 & ~n929;
  assign n1516 = n1514 & n1515;
  assign n1517 = n1513 & n1516;
  assign n1518 = n1512 & n1517;
  assign n1519 = n1495 & n1518;
  assign n1521 = ~n298 & ~n1166;
  assign n1522 = n1520 & n1521;
  assign n1523 = ~n152 & ~n928;
  assign n1524 = ~n202 & ~n323;
  assign n1525 = n1523 & n1524;
  assign n1526 = n1522 & n1525;
  assign n1527 = ~n193 & ~n347;
  assign n1528 = ~n304 & n1527;
  assign n1529 = n1526 & n1528;
  assign n1530 = ~n199 & ~n406;
  assign n1531 = n1301 & n1530;
  assign n1532 = n684 & n1531;
  assign n1533 = n1529 & n1532;
  assign n1534 = ~n266 & n727;
  assign n1535 = n591 & n1534;
  assign n1537 = ~n405 & ~n1536;
  assign n1538 = ~n610 & ~n1266;
  assign n1539 = n983 & n1538;
  assign n1540 = n1537 & n1539;
  assign n1541 = n1535 & n1540;
  assign n1542 = n1533 & n1541;
  assign n1543 = n1519 & n1542;
  assign n1544 = n1465 & n1543;
  assign n1545 = ~n1420 & ~n1544;
  assign n1546 = ~n560 & ~n920;
  assign n1547 = n1283 & n1546;
  assign n1548 = ~n362 & ~n416;
  assign n1549 = n1547 & n1548;
  assign n1550 = ~n346 & ~n476;
  assign n1551 = ~n245 & ~n428;
  assign n1552 = n1550 & n1551;
  assign n1553 = n1549 & n1552;
  assign n1554 = ~n350 & ~n535;
  assign n1555 = ~n110 & n1554;
  assign n1556 = ~n270 & ~n843;
  assign n1557 = n1003 & n1556;
  assign n1558 = n1555 & n1557;
  assign n1559 = n1553 & n1558;
  assign n1560 = ~n69 & ~n740;
  assign n1561 = ~n529 & ~n640;
  assign n1562 = n1560 & n1561;
  assign n1563 = ~n126 & ~n901;
  assign n1564 = ~n524 & ~n683;
  assign n1565 = n1563 & n1564;
  assign n1566 = n1562 & n1565;
  assign n1567 = ~n189 & ~n331;
  assign n1568 = n781 & n1567;
  assign n1569 = ~n221 & ~n347;
  assign n1570 = n1273 & n1569;
  assign n1571 = n1568 & n1570;
  assign n1572 = n1566 & n1571;
  assign n1573 = ~n396 & ~n755;
  assign n1574 = n713 & n1573;
  assign n1575 = ~n266 & ~n1135;
  assign n1576 = ~n382 & n1575;
  assign n1577 = n1574 & n1576;
  assign n1578 = n648 & n1577;
  assign n1579 = n1572 & n1578;
  assign n1580 = n1559 & n1579;
  assign n1581 = n519 & n1580;
  assign n1582 = ~n928 & n1238;
  assign n1583 = ~n134 & ~n593;
  assign n1584 = ~n231 & n1583;
  assign n1585 = n1582 & n1584;
  assign n1586 = ~n456 & n1301;
  assign n1587 = n1585 & n1586;
  assign n1588 = ~n799 & ~n1060;
  assign n1589 = ~n202 & ~n254;
  assign n1590 = n1588 & n1589;
  assign n1591 = ~n148 & ~n689;
  assign n1592 = ~n234 & n1591;
  assign n1593 = n1590 & n1592;
  assign n1594 = ~n616 & ~n1047;
  assign n1595 = n1126 & n1594;
  assign n1596 = n1593 & n1595;
  assign n1597 = n1587 & n1596;
  assign n1598 = ~n659 & ~n723;
  assign n1599 = ~n304 & ~n558;
  assign n1600 = n1598 & n1599;
  assign n1601 = n756 & n1600;
  assign n1602 = ~n322 & ~n550;
  assign n1603 = n105 & n1602;
  assign n1604 = n1601 & n1603;
  assign n1605 = n1597 & n1604;
  assign n1606 = ~n439 & ~n710;
  assign n1607 = ~n218 & n1606;
  assign n1609 = n1607 & n1608;
  assign n1610 = n1058 & n1085;
  assign n1612 = n1610 & n1611;
  assign n1613 = n1609 & n1612;
  assign n1614 = ~n181 & ~n296;
  assign n1615 = ~n156 & ~n228;
  assign n1616 = n1614 & n1615;
  assign n1617 = n302 & ~n343;
  assign n1618 = n1616 & n1617;
  assign n1619 = n1613 & n1618;
  assign n1620 = ~n283 & ~n432;
  assign n1621 = ~n503 & n1620;
  assign n1622 = ~n443 & ~n791;
  assign n1623 = n1621 & n1622;
  assign n1624 = n485 & n999;
  assign n1625 = n144 & n1624;
  assign n1626 = n1623 & n1625;
  assign n1627 = ~n201 & ~n409;
  assign n1628 = ~n278 & n1627;
  assign n1629 = n321 & n1628;
  assign n1630 = n532 & n852;
  assign n1631 = ~n475 & ~n758;
  assign n1632 = n738 & n1631;
  assign n1633 = n1630 & n1632;
  assign n1634 = n1629 & n1633;
  assign n1635 = n1626 & n1634;
  assign n1636 = n1619 & n1635;
  assign n1637 = n1605 & n1636;
  assign n1638 = n1581 & n1637;
  assign n1639 = ~n1545 & n1638;
  assign n1640 = ~n550 & ~n1135;
  assign n1641 = ~n103 & n1640;
  assign n1642 = n144 & n493;
  assign n1643 = n1641 & n1642;
  assign n1644 = ~n308 & ~n946;
  assign n1645 = n118 & n1644;
  assign n1646 = ~n83 & ~n301;
  assign n1647 = ~n975 & n1646;
  assign n1648 = n1645 & n1647;
  assign n1649 = n1643 & n1648;
  assign n1651 = n210 & ~n634;
  assign n1652 = n1650 & n1651;
  assign n1653 = ~n403 & ~n476;
  assign n1654 = ~n375 & n1653;
  assign n1655 = ~n254 & n788;
  assign n1656 = n1654 & n1655;
  assign n1657 = n1652 & n1656;
  assign n1658 = n1649 & n1657;
  assign n1659 = ~n127 & ~n506;
  assign n1660 = ~n440 & ~n442;
  assign n1661 = n1659 & n1660;
  assign n1662 = n1658 & n1661;
  assign n1663 = ~n272 & ~n410;
  assign n1664 = ~n221 & n1663;
  assign n1665 = ~n138 & ~n1166;
  assign n1666 = n584 & n1665;
  assign n1667 = n1664 & n1666;
  assign n1668 = ~n263 & ~n405;
  assign n1669 = n1667 & n1668;
  assign n1672 = ~n248 & ~n920;
  assign n1673 = ~n99 & n1672;
  assign n1674 = n1671 & n1673;
  assign n1675 = n1184 & n1674;
  assign n1676 = n1669 & n1675;
  assign n1677 = n1019 & n1301;
  assign n1679 = n332 & n1678;
  assign n1680 = n1677 & n1679;
  assign n1681 = ~n524 & ~n709;
  assign n1682 = n438 & n1681;
  assign n1683 = n1680 & n1682;
  assign n1684 = n810 & n1683;
  assign n1685 = n1676 & n1684;
  assign n1686 = n1662 & n1685;
  assign n1687 = ~n449 & n833;
  assign n1688 = ~n181 & ~n337;
  assign n1689 = n1311 & n1688;
  assign n1690 = n1687 & n1689;
  assign n1691 = n875 & n1622;
  assign n1692 = n1690 & n1691;
  assign n1693 = ~n540 & ~n671;
  assign n1694 = ~n104 & ~n812;
  assign n1695 = n1693 & n1694;
  assign n1696 = n1582 & n1695;
  assign n1697 = n1692 & n1696;
  assign n1698 = ~n385 & ~n675;
  assign n1699 = n1555 & n1698;
  assign n1700 = n624 & n1699;
  assign n1701 = ~n265 & ~n553;
  assign n1702 = ~n292 & ~n359;
  assign n1703 = n1701 & n1702;
  assign n1704 = ~n98 & ~n683;
  assign n1705 = ~n253 & ~n710;
  assign n1706 = n1704 & n1705;
  assign n1707 = n1703 & n1706;
  assign n1708 = n1700 & n1707;
  assign n1709 = n1697 & n1708;
  assign n1710 = ~n64 & ~n461;
  assign n1711 = n1424 & n1710;
  assign n1712 = ~n346 & ~n402;
  assign n1713 = ~n351 & n1712;
  assign n1714 = n1711 & n1713;
  assign n1715 = ~n164 & n679;
  assign n1716 = ~n475 & ~n1060;
  assign n1717 = ~n163 & ~n313;
  assign n1718 = n1716 & n1717;
  assign n1719 = n1715 & n1718;
  assign n1720 = n1714 & n1719;
  assign n1721 = n673 & n1363;
  assign n1722 = n1720 & n1721;
  assign n1723 = ~n418 & ~n740;
  assign n1724 = n1722 & n1723;
  assign n1725 = n1709 & n1724;
  assign n1726 = n1686 & n1725;
  assign n1727 = ~n1639 & ~n1726;
  assign n1732 = n100 & ~n1405;
  assign n1733 = ~n163 & n1732;
  assign n1734 = n1731 & n1733;
  assign n1735 = ~n103 & ~n249;
  assign n1736 = ~n1135 & n1735;
  assign n1737 = ~n362 & ~n517;
  assign n1738 = n1736 & n1737;
  assign n1739 = ~n439 & ~n652;
  assign n1740 = n1483 & n1739;
  assign n1741 = ~n138 & ~n303;
  assign n1742 = n1072 & n1741;
  assign n1743 = n1740 & n1742;
  assign n1744 = n1738 & n1743;
  assign n1745 = n1734 & n1744;
  assign n1746 = ~n337 & ~n544;
  assign n1747 = n893 & n1746;
  assign n1748 = ~n111 & ~n222;
  assign n1749 = ~n406 & ~n443;
  assign n1750 = n1748 & n1749;
  assign n1751 = n1747 & n1750;
  assign n1752 = n1161 & n1751;
  assign n1753 = n1745 & n1752;
  assign n1754 = ~n628 & ~n714;
  assign n1755 = ~n344 & ~n617;
  assign n1756 = ~n226 & ~n237;
  assign n1757 = n1755 & n1756;
  assign n1758 = n1754 & n1757;
  assign n1759 = ~n314 & ~n410;
  assign n1760 = ~n190 & ~n588;
  assign n1761 = n1759 & n1760;
  assign n1762 = n397 & n1167;
  assign n1763 = n1761 & n1762;
  assign n1764 = n1758 & n1763;
  assign n1766 = n464 & n1765;
  assign n1767 = n1764 & n1766;
  assign n1768 = n1753 & n1767;
  assign n1769 = n880 & n1768;
  assign n1770 = n247 & n1165;
  assign n1772 = n1332 & n1771;
  assign n1773 = n1770 & n1772;
  assign n1774 = ~n170 & ~n948;
  assign n1775 = ~n627 & n1774;
  assign n1776 = ~n186 & ~n197;
  assign n1777 = n1775 & n1776;
  assign n1778 = n1773 & n1777;
  assign n1779 = ~n659 & n1778;
  assign n1780 = ~n199 & ~n353;
  assign n1781 = n902 & n1780;
  assign n1782 = ~n723 & ~n758;
  assign n1783 = n302 & n1782;
  assign n1784 = n1781 & n1783;
  assign n1785 = ~n593 & ~n1266;
  assign n1786 = n1784 & n1785;
  assign n1787 = ~n336 & ~n396;
  assign n1788 = ~n560 & n1787;
  assign n1790 = n1788 & n1789;
  assign n1791 = n118 & n1283;
  assign n1792 = ~n273 & ~n843;
  assign n1793 = n1614 & n1792;
  assign n1794 = n1791 & n1793;
  assign n1795 = n1790 & n1794;
  assign n1796 = n1786 & n1795;
  assign n1797 = n1779 & n1796;
  assign n1798 = n1769 & n1797;
  assign n1799 = ~n1727 & n1798;
  assign n1800 = ~n553 & n1514;
  assign n1801 = ~n163 & ~n506;
  assign n1802 = n1800 & n1801;
  assign n1803 = ~n95 & ~n671;
  assign n1804 = ~n216 & n1803;
  assign n1805 = ~n231 & ~n504;
  assign n1806 = ~n443 & n1805;
  assign n1807 = n1804 & n1806;
  assign n1808 = n1802 & n1807;
  assign n1809 = ~n104 & n1283;
  assign n1810 = ~n186 & ~n277;
  assign n1811 = ~n901 & n1810;
  assign n1812 = n1809 & n1811;
  assign n1813 = n1808 & n1812;
  assign n1814 = ~n227 & ~n592;
  assign n1815 = ~n975 & n1814;
  assign n1816 = n1451 & n1815;
  assign n1817 = ~n117 & ~n919;
  assign n1818 = ~n471 & ~n652;
  assign n1819 = n1817 & n1818;
  assign n1820 = n1816 & n1819;
  assign n1821 = ~n256 & n986;
  assign n1822 = n1327 & n1821;
  assign n1823 = n1820 & n1822;
  assign n1824 = n1813 & n1823;
  assign n1828 = ~n234 & n1827;
  assign n1829 = n1824 & n1828;
  assign n1830 = n366 & n1829;
  assign n1831 = ~n406 & ~n787;
  assign n1832 = ~n226 & n1831;
  assign n1833 = n545 & n1832;
  assign n1835 = n1665 & n1834;
  assign n1836 = ~n456 & ~n458;
  assign n1837 = n1835 & n1836;
  assign n1838 = n1833 & n1837;
  assign n1839 = ~n126 & ~n723;
  assign n1840 = ~n535 & n1839;
  assign n1841 = ~n152 & ~n476;
  assign n1842 = n437 & n1841;
  assign n1843 = n1840 & n1842;
  assign n1844 = n1838 & n1843;
  assign n1845 = ~n209 & ~n582;
  assign n1846 = ~n680 & n1845;
  assign n1847 = ~n269 & ~n928;
  assign n1848 = n1846 & n1847;
  assign n1849 = ~n201 & ~n791;
  assign n1850 = ~n64 & ~n799;
  assign n1851 = n1849 & n1850;
  assign n1852 = n1848 & n1851;
  assign n1853 = ~n74 & ~n605;
  assign n1854 = ~n424 & n1853;
  assign n1855 = ~n284 & n530;
  assign n1856 = n1854 & n1855;
  assign n1857 = ~n518 & n884;
  assign n1858 = n796 & n818;
  assign n1859 = ~n396 & ~n1858;
  assign n1860 = n1857 & n1859;
  assign n1861 = n1856 & n1860;
  assign n1862 = n1852 & n1861;
  assign n1863 = n1844 & n1862;
  assign n1864 = ~n263 & ~n948;
  assign n1865 = ~n527 & n1864;
  assign n1867 = ~n115 & ~n514;
  assign n1868 = n1866 & n1867;
  assign n1869 = n1865 & n1868;
  assign n1870 = ~n463 & ~n758;
  assign n1871 = ~n109 & n1870;
  assign n1872 = n1869 & n1871;
  assign n1873 = n713 & n1072;
  assign n1874 = ~n133 & ~n382;
  assign n1875 = n1873 & n1874;
  assign n1876 = n1872 & n1875;
  assign n1877 = n1863 & n1876;
  assign n1878 = n1830 & n1877;
  assign n1879 = ~n1799 & ~n1878;
  assign n1880 = ~n103 & ~n929;
  assign n1881 = ~n266 & n1880;
  assign n1882 = ~n95 & ~n588;
  assign n1883 = ~n476 & ~n627;
  assign n1884 = n1882 & n1883;
  assign n1885 = n1881 & n1884;
  assign n1886 = n601 & n1885;
  assign n1887 = ~n217 & ~n710;
  assign n1888 = n1616 & n1887;
  assign n1889 = ~n303 & ~n1227;
  assign n1890 = n1888 & n1889;
  assign n1891 = n1886 & n1890;
  assign n1892 = ~n221 & ~n740;
  assign n1893 = n833 & n1892;
  assign n1894 = n738 & n1893;
  assign n1895 = ~n122 & ~n370;
  assign n1896 = ~n812 & n1895;
  assign n1897 = n1894 & n1896;
  assign n1898 = n1593 & n1897;
  assign n1899 = n1891 & n1898;
  assign n1900 = ~n127 & ~n628;
  assign n1901 = ~n244 & n1900;
  assign n1902 = ~n277 & ~n350;
  assign n1903 = ~n524 & n1902;
  assign n1904 = n1901 & n1903;
  assign n1905 = ~n171 & ~n463;
  assign n1906 = ~n51 & ~n301;
  assign n1907 = n1905 & n1906;
  assign n1908 = n1904 & n1907;
  assign n1909 = ~n314 & ~n605;
  assign n1910 = n1491 & n1909;
  assign n1911 = ~n190 & ~n751;
  assign n1912 = n1910 & n1911;
  assign n1913 = n1908 & n1912;
  assign n1914 = n1899 & n1913;
  assign n1915 = ~n173 & n672;
  assign n1916 = n1058 & n1915;
  assign n1917 = n1800 & n1916;
  assign n1918 = ~n313 & ~n373;
  assign n1919 = ~n309 & n1918;
  assign n1920 = ~n369 & ~n535;
  assign n1921 = n1919 & n1920;
  assign n1922 = n1917 & n1921;
  assign n1923 = n1640 & n1698;
  assign n1924 = ~n736 & n1923;
  assign n1925 = ~n412 & ~n787;
  assign n1926 = ~n540 & ~n919;
  assign n1927 = n1925 & n1926;
  assign n1928 = n1924 & n1927;
  assign n1929 = ~n262 & ~n323;
  assign n1930 = ~n284 & n1929;
  assign n1931 = ~n243 & ~n409;
  assign n1932 = n1930 & n1931;
  assign n1933 = ~n557 & ~n1047;
  assign n1934 = ~n298 & n1933;
  assign n1935 = ~n151 & n271;
  assign n1936 = n1934 & n1935;
  assign n1937 = n1932 & n1936;
  assign n1938 = n1928 & n1937;
  assign n1939 = n1922 & n1938;
  assign n1940 = ~n312 & ~n666;
  assign n1941 = ~n295 & ~n354;
  assign n1942 = n1940 & n1941;
  assign n1943 = ~n280 & ~n292;
  assign n1944 = ~n99 & ~n278;
  assign n1945 = n1943 & n1944;
  assign n1946 = n1942 & n1945;
  assign n1947 = ~n250 & ~n683;
  assign n1948 = ~n218 & ~n227;
  assign n1949 = n1947 & n1948;
  assign n1950 = n860 & n1787;
  assign n1951 = n1949 & n1950;
  assign n1952 = n1946 & n1951;
  assign n1953 = n1601 & n1952;
  assign n1954 = ~n74 & ~n201;
  assign n1955 = ~n69 & ~n1266;
  assign n1956 = n1954 & n1955;
  assign n1957 = ~n104 & ~n432;
  assign n1958 = ~n378 & ~n514;
  assign n1959 = n1957 & n1958;
  assign n1960 = n1956 & n1959;
  assign n1961 = ~n334 & ~n390;
  assign n1962 = n1567 & n1961;
  assign n1963 = n1960 & n1962;
  assign n1964 = ~n222 & ~n843;
  assign n1965 = ~n382 & ~n850;
  assign n1966 = n1964 & n1965;
  assign n1967 = ~n93 & ~n517;
  assign n1968 = ~n238 & ~n630;
  assign n1969 = n1967 & n1968;
  assign n1970 = n1966 & n1969;
  assign n1971 = n1963 & n1970;
  assign n1972 = n1953 & n1971;
  assign n1973 = n1939 & n1972;
  assign n1974 = n1914 & n1973;
  assign n1975 = ~n1879 & n1974;
  assign n1976 = ~n201 & ~n405;
  assign n1977 = ~n181 & ~n333;
  assign n1978 = n1976 & n1977;
  assign n1979 = ~n109 & n1087;
  assign n1980 = n1978 & n1979;
  assign n1981 = ~n492 & ~n691;
  assign n1982 = ~n265 & ~n270;
  assign n1983 = n1981 & n1982;
  assign n1984 = n219 & n1983;
  assign n1985 = n1980 & n1984;
  assign n1986 = ~n527 & ~n588;
  assign n1987 = ~n337 & n1986;
  assign n1988 = ~n192 & ~n901;
  assign n1989 = ~n231 & n1988;
  assign n1990 = n1987 & n1989;
  assign n1991 = n1985 & n1990;
  assign n1992 = ~n755 & ~n946;
  assign n1993 = n371 & n1992;
  assign n1994 = ~n250 & n453;
  assign n1995 = n1993 & n1994;
  assign n1996 = ~n416 & n485;
  assign n1997 = ~n126 & ~n652;
  assign n1998 = n519 & n1997;
  assign n1999 = n1996 & n1998;
  assign n2000 = n1995 & n1999;
  assign n2001 = n1991 & n2000;
  assign n2002 = ~n243 & n1205;
  assign n2003 = ~n461 & ~n503;
  assign n2004 = ~n93 & ~n843;
  assign n2005 = n2003 & n2004;
  assign n2006 = n2002 & n2005;
  assign n2007 = n1671 & n2006;
  assign n2008 = ~n358 & ~n841;
  assign n2009 = n1883 & n2008;
  assign n2010 = n713 & n2009;
  assign n2011 = n2007 & n2010;
  assign n2012 = n2001 & n2011;
  assign n2013 = ~n163 & ~n353;
  assign n2014 = ~n174 & ~n226;
  assign n2015 = n2013 & n2014;
  assign n2016 = n321 & n1209;
  assign n2017 = n2015 & n2016;
  assign n2018 = n438 & n2017;
  assign n2019 = ~n138 & ~n257;
  assign n2020 = n444 & n2019;
  assign n2021 = ~n171 & n2020;
  assign n2022 = ~n327 & ~n567;
  assign n2023 = n851 & n2022;
  assign n2024 = ~n156 & ~n529;
  assign n2025 = ~n99 & ~n605;
  assign n2026 = n2024 & n2025;
  assign n2027 = n2023 & n2026;
  assign n2028 = n2021 & n2027;
  assign n2029 = n2018 & n2028;
  assign n2030 = n1928 & n2029;
  assign n2031 = n2012 & n2030;
  assign n2032 = ~n640 & ~n1047;
  assign n2033 = ~n396 & n2032;
  assign n2034 = n1785 & n2033;
  assign n2036 = ~n295 & n2035;
  assign n2037 = n2034 & n2036;
  assign n2039 = n441 & n2038;
  assign n2040 = ~n64 & ~n525;
  assign n2041 = n2039 & n2040;
  assign n2042 = ~n253 & ~n428;
  assign n2043 = n684 & n2042;
  assign n2044 = n2041 & n2043;
  assign n2045 = n2037 & n2044;
  assign n2046 = ~n69 & ~n1166;
  assign n2047 = ~n280 & n2046;
  assign n2048 = n1723 & n1748;
  assign n2049 = n2047 & n2048;
  assign n2050 = n583 & n1492;
  assign n2051 = ~n322 & ~n409;
  assign n2052 = n1836 & n2051;
  assign n2053 = n2050 & n2052;
  assign n2054 = n2049 & n2053;
  assign n2055 = ~n313 & ~n610;
  assign n2056 = n1335 & n2055;
  assign n2057 = ~n524 & ~n660;
  assign n2058 = ~n141 & ~n375;
  assign n2059 = n2057 & n2058;
  assign n2060 = n2056 & n2059;
  assign n2061 = n2054 & n2060;
  assign n2062 = n2045 & n2061;
  assign n2063 = ~n432 & ~n758;
  assign n2064 = n2062 & n2063;
  assign n2065 = n2031 & n2064;
  assign n2066 = ~n1975 & ~n2065;
  assign n2074 = ~n163 & ~n344;
  assign n2075 = n2073 & n2074;
  assign n2076 = ~n440 & ~n560;
  assign n2077 = n2075 & n2076;
  assign n2078 = n867 & n2077;
  assign n2079 = ~n301 & ~n689;
  assign n2080 = ~n127 & n2079;
  assign n2081 = ~n263 & ~n1482;
  assign n2082 = n2080 & n2081;
  assign n2083 = ~n181 & ~n492;
  assign n2084 = n583 & n2083;
  assign n2085 = ~n156 & ~n227;
  assign n2086 = n2084 & n2085;
  assign n2087 = n2082 & n2086;
  assign n2088 = n2078 & n2087;
  assign n2089 = n2072 & n2088;
  assign n2090 = ~n293 & ~n552;
  assign n2091 = ~n406 & ~n558;
  assign n2092 = n2090 & n2091;
  assign n2093 = n1359 & n2092;
  assign n2094 = ~n170 & ~n680;
  assign n2095 = n2093 & n2094;
  assign n2096 = ~n417 & n1389;
  assign n2097 = ~n456 & n2096;
  assign n2098 = ~n763 & n1171;
  assign n2099 = n425 & n852;
  assign n2100 = n2098 & n2099;
  assign n2101 = n2097 & n2100;
  assign n2102 = n2095 & n2101;
  assign n2103 = n2089 & n2102;
  assign n2105 = n335 & n2104;
  assign n2106 = n1909 & n2105;
  assign n2107 = ~n221 & ~n254;
  assign n2108 = n1295 & n2107;
  assign n2109 = n878 & n2108;
  assign n2110 = n2106 & n2109;
  assign n2111 = n2103 & n2110;
  assign n2112 = ~n253 & ~n812;
  assign n2113 = ~n461 & n2112;
  assign n2114 = ~n270 & ~n350;
  assign n2115 = ~n74 & ~n553;
  assign n2116 = n2114 & n2115;
  assign n2117 = n2113 & n2116;
  assign n2118 = ~n323 & ~n353;
  assign n2119 = ~n403 & n2118;
  assign n2120 = n2117 & n2119;
  assign n2125 = n282 & n1172;
  assign n2126 = ~n343 & ~n1166;
  assign n2127 = n2125 & n2126;
  assign n2128 = n2124 & n2127;
  assign n2129 = n2120 & n2128;
  assign n2134 = ~n192 & ~n612;
  assign n2135 = ~n115 & ~n428;
  assign n2136 = n2134 & n2135;
  assign n2138 = ~n174 & ~n266;
  assign n2139 = n2137 & n2138;
  assign n2140 = n2136 & n2139;
  assign n2141 = n2133 & n2140;
  assign n2142 = n2129 & n2141;
  assign n2143 = ~n202 & ~n478;
  assign n2144 = n1792 & n2143;
  assign n2145 = ~n336 & ~n351;
  assign n2146 = n2144 & n2145;
  assign n2147 = ~n284 & n1075;
  assign n2148 = n1091 & n1882;
  assign n2149 = n2147 & n2148;
  assign n2150 = n2146 & n2149;
  assign n2151 = ~n841 & ~n946;
  assign n2152 = ~n592 & ~n675;
  assign n2153 = n2151 & n2152;
  assign n2154 = ~n243 & ~n298;
  assign n2155 = n2153 & n2154;
  assign n2156 = n2150 & n2155;
  assign n2157 = ~n439 & ~n518;
  assign n2158 = ~n616 & n2157;
  assign n2160 = ~n141 & ~n173;
  assign n2161 = n2159 & n2160;
  assign n2162 = n2158 & n2161;
  assign n2163 = ~n295 & ~n671;
  assign n2164 = n2162 & n2163;
  assign n2166 = ~n544 & n2165;
  assign n2167 = ~n155 & ~n527;
  assign n2168 = ~n244 & n2167;
  assign n2169 = n2166 & n2168;
  assign n2170 = ~n385 & ~n416;
  assign n2171 = n2169 & n2170;
  assign n2172 = n2164 & n2171;
  assign n2173 = n2156 & n2172;
  assign n2174 = n2142 & n2173;
  assign n2175 = n2111 & n2174;
  assign n2176 = ~n2066 & n2175;
  assign n2177 = ~n253 & ~n323;
  assign n2178 = ~n110 & ~n429;
  assign n2179 = n2177 & n2178;
  assign n2180 = ~n217 & ~n385;
  assign n2181 = n2179 & n2180;
  assign n2182 = ~n660 & ~n1135;
  assign n2183 = n191 & n2182;
  assign n2184 = n2181 & n2183;
  assign n2185 = ~n167 & ~n208;
  assign n2186 = ~n216 & n2185;
  assign n2188 = n1286 & n2187;
  assign n2189 = n2186 & n2188;
  assign n2190 = ~n293 & ~n709;
  assign n2191 = n1264 & n2190;
  assign n2192 = n1659 & n1831;
  assign n2193 = n2191 & n2192;
  assign n2194 = n2189 & n2193;
  assign n2195 = n2184 & n2194;
  assign n2196 = n1778 & n2195;
  assign n2197 = ~n497 & ~n929;
  assign n2198 = n70 & n2197;
  assign n2199 = ~n687 & n2198;
  assign n2200 = ~n541 & ~n750;
  assign n2201 = ~n616 & n2200;
  assign n2202 = ~n432 & ~n919;
  assign n2203 = ~n57 & n2202;
  assign n2204 = n2201 & n2203;
  assign n2205 = n2199 & n2204;
  assign n2206 = n2196 & n2205;
  assign n2207 = ~n272 & ~n392;
  assign n2208 = ~n403 & n2207;
  assign n2209 = ~n93 & ~n652;
  assign n2210 = n2208 & n2209;
  assign n2211 = n1835 & n2210;
  assign n2212 = ~n266 & ~n689;
  assign n2213 = n532 & n2212;
  assign n2214 = ~n183 & ~n308;
  assign n2215 = n2213 & n2214;
  assign n2216 = ~n83 & ~n417;
  assign n2217 = ~n231 & n2216;
  assign n2218 = n135 & n1902;
  assign n2219 = n2217 & n2218;
  assign n2220 = n2215 & n2219;
  assign n2221 = n2211 & n2220;
  assign n2222 = ~n270 & ~n544;
  assign n2223 = ~n202 & ~n850;
  assign n2224 = n2222 & n2223;
  assign n2225 = ~n128 & ~n630;
  assign n2226 = n2224 & n2225;
  assign n2227 = ~n79 & ~n359;
  assign n2228 = ~n257 & n2227;
  assign n2229 = n1695 & n2228;
  assign n2230 = n2226 & n2229;
  assign n2231 = n2221 & n2230;
  assign n2232 = ~n126 & ~n469;
  assign n2233 = ~n248 & ~n314;
  assign n2234 = n2232 & n2233;
  assign n2235 = ~n439 & ~n517;
  assign n2236 = ~n192 & ~n390;
  assign n2237 = n2235 & n2236;
  assign n2238 = n2234 & n2237;
  assign n2241 = n2239 & n2240;
  assign n2242 = ~n1482 & n1569;
  assign n2243 = n2241 & n2242;
  assign n2244 = n2238 & n2243;
  assign n2245 = n1796 & n2244;
  assign n2246 = n2231 & n2245;
  assign n2247 = n2206 & n2246;
  assign n2248 = ~n2176 & ~n2247;
  assign n2249 = ~n390 & ~n582;
  assign n2250 = n1909 & n2249;
  assign n2251 = n271 & n2250;
  assign n2252 = ~n233 & ~n919;
  assign n2253 = ~n659 & n2252;
  assign n2254 = n2251 & n2253;
  assign n2255 = ~n143 & ~n226;
  assign n2256 = ~n265 & ~n617;
  assign n2257 = n2255 & n2256;
  assign n2258 = n834 & n2257;
  assign n2259 = n2254 & n2258;
  assign n2260 = ~n128 & ~n418;
  assign n2261 = ~n301 & ~n535;
  assign n2262 = n2260 & n2261;
  assign n2263 = ~n262 & ~n347;
  assign n2264 = ~n683 & ~n799;
  assign n2265 = n2263 & n2264;
  assign n2266 = n2262 & n2265;
  assign n2268 = n2151 & n2267;
  assign n2269 = n2266 & n2268;
  assign n2270 = ~n382 & ~n723;
  assign n2271 = ~n98 & ~n238;
  assign n2272 = n2270 & n2271;
  assign n2273 = n786 & n2272;
  assign n2274 = n2269 & n2273;
  assign n2275 = n2259 & n2274;
  assign n2276 = ~n148 & ~n1060;
  assign n2277 = ~n93 & ~n174;
  assign n2278 = n2276 & n2277;
  assign n2279 = n1640 & n2278;
  assign n2280 = ~n237 & ~n304;
  assign n2281 = ~n359 & n2280;
  assign n2282 = n2279 & n2281;
  assign n2283 = n2275 & n2282;
  assign n2284 = ~n576 & ~n797;
  assign n2285 = ~n323 & ~n709;
  assign n2286 = ~n207 & n2285;
  assign n2287 = n2284 & n2286;
  assign n2288 = ~n146 & ~n173;
  assign n2289 = ~n319 & ~n800;
  assign n2290 = n2288 & n2289;
  assign n2291 = n2287 & n2290;
  assign n2293 = ~n449 & ~n758;
  assign n2294 = n2292 & n2293;
  assign n2295 = n135 & ~n506;
  assign n2296 = n2294 & n2295;
  assign n2297 = n2291 & n2296;
  assign n2299 = ~n83 & ~n497;
  assign n2300 = n2298 & n2299;
  assign n2301 = n1809 & n2300;
  assign n2302 = ~n185 & ~n458;
  assign n2303 = n542 & n2302;
  assign n2304 = n682 & n2303;
  assign n2305 = n2301 & n2304;
  assign n2306 = n2297 & n2305;
  assign n2308 = ~n257 & ~n278;
  assign n2309 = n2307 & n2308;
  assign n2310 = ~n228 & ~n312;
  assign n2311 = ~n691 & n2310;
  assign n2312 = n2309 & n2311;
  assign n2313 = n860 & n2165;
  assign n2314 = ~n201 & ~n392;
  assign n2315 = n1739 & n2314;
  assign n2316 = n2313 & n2315;
  assign n2317 = n2312 & n2316;
  assign n2318 = ~n334 & ~n346;
  assign n2319 = ~n410 & ~n660;
  assign n2320 = n2318 & n2319;
  assign n2321 = ~n428 & n2320;
  assign n2322 = n2317 & n2321;
  assign n2323 = n2306 & n2322;
  assign n2324 = n2283 & n2323;
  assign n2325 = ~n263 & ~n351;
  assign n2326 = ~n313 & ~n787;
  assign n2327 = n2325 & n2326;
  assign n2328 = ~n170 & ~n452;
  assign n2329 = n973 & n2328;
  assign n2330 = n2327 & n2329;
  assign n2331 = ~n99 & n2330;
  assign n2332 = n445 & n1728;
  assign n2333 = ~n273 & ~n293;
  assign n2334 = ~n249 & n2333;
  assign n2335 = ~n151 & n184;
  assign n2336 = n2334 & n2335;
  assign n2337 = n2332 & n2336;
  assign n2338 = n2331 & n2337;
  assign n2339 = ~n517 & ~n929;
  assign n2340 = n1530 & n2339;
  assign n2341 = n297 & n2340;
  assign n2342 = n220 & n2341;
  assign n2343 = n2338 & n2342;
  assign n2344 = ~n244 & ~n630;
  assign n2345 = n1776 & n2344;
  assign n2346 = n1546 & n2345;
  assign n2347 = ~n544 & ~n791;
  assign n2348 = ~n755 & n2347;
  assign n2349 = ~n331 & ~n350;
  assign n2350 = n857 & n2349;
  assign n2351 = n2348 & n2350;
  assign n2352 = n2346 & n2351;
  assign n2353 = ~n57 & n1805;
  assign n2354 = n2097 & n2353;
  assign n2355 = n2352 & n2354;
  assign n2356 = n2343 & n2355;
  assign n2357 = n2324 & n2356;
  assign n2358 = ~n2248 & n2357;
  assign n2359 = ~n1208 & ~n1414;
  assign n2360 = n1097 & ~n2359;
  assign n2361 = ~n970 & ~n2360;
  assign n2362 = n882 & ~n2361;
  assign n2363 = ~n734 & ~n2362;
  assign n2364 = n1544 & ~n2363;
  assign n2365 = ~n1638 & ~n2364;
  assign n2366 = n1726 & ~n2365;
  assign n2367 = ~n1798 & ~n2366;
  assign n2368 = n1878 & ~n2367;
  assign n2369 = ~n1974 & ~n2368;
  assign n2370 = n2065 & ~n2369;
  assign n2371 = ~n2175 & ~n2370;
  assign n2372 = n2247 & ~n2371;
  assign n2373 = ~n2357 & ~n2372;
  assign n2374 = ~n206 & ~n293;
  assign n2375 = ~n1060 & n2374;
  assign n2376 = n2113 & n2375;
  assign n2377 = ~n192 & n1741;
  assign n2378 = ~n186 & n397;
  assign n2379 = n2377 & n2378;
  assign n2380 = n2376 & n2379;
  assign n2381 = n1152 & n2380;
  assign n2382 = ~n167 & ~n351;
  assign n2383 = n2293 & n2382;
  assign n2384 = ~n373 & ~n582;
  assign n2386 = n2384 & n2385;
  assign n2387 = n2383 & n2386;
  assign n2388 = ~n354 & ~n689;
  assign n2389 = ~n333 & ~n406;
  assign n2390 = n2388 & n2389;
  assign n2392 = ~n497 & ~n540;
  assign n2393 = n2391 & n2392;
  assign n2394 = n2390 & n2393;
  assign n2395 = n2387 & n2394;
  assign n2396 = ~n109 & ~n170;
  assign n2397 = ~n429 & ~n634;
  assign n2398 = n2396 & n2397;
  assign n2399 = n2395 & n2398;
  assign n2400 = n2381 & n2399;
  assign n2402 = ~n369 & ~n628;
  assign n2403 = n2401 & n2402;
  assign n2404 = ~n197 & ~n787;
  assign n2405 = ~n257 & ~n439;
  assign n2406 = n2404 & n2405;
  assign n2407 = n2403 & n2406;
  assign n2408 = ~n244 & ~n504;
  assign n2409 = ~n173 & n2408;
  assign n2410 = n1193 & n2409;
  assign n2411 = n2407 & n2410;
  assign n2412 = n118 & n989;
  assign n2413 = n1328 & n2412;
  assign n2414 = n2258 & n2413;
  assign n2415 = n2411 & n2414;
  assign n2416 = ~n326 & n1288;
  assign n2417 = ~n295 & n1238;
  assign n2418 = n2416 & n2417;
  assign n2419 = ~n687 & n994;
  assign n2420 = n2418 & n2419;
  assign n2421 = n2415 & n2420;
  assign n2422 = n2400 & n2421;
  assign n2423 = n1581 & n2422;
  assign n2424 = ~n2373 & n2423;
  assign n2425 = ~n2358 & ~n2424;
  assign n2426 = ~n385 & ~n456;
  assign n2427 = ~n750 & n2426;
  assign n2428 = ~n120 & ~n509;
  assign n2429 = n1273 & n2428;
  assign n2430 = n2427 & n2429;
  assign n2431 = n603 & n2430;
  assign n2432 = ~n406 & ~n1047;
  assign n2433 = ~n117 & ~n143;
  assign n2434 = n2432 & n2433;
  assign n2435 = ~n343 & ~n531;
  assign n2436 = n546 & n2435;
  assign n2437 = n2434 & n2436;
  assign n2438 = n1042 & n2437;
  assign n2439 = n2431 & n2438;
  assign n2440 = ~n216 & ~n429;
  assign n2441 = ~n373 & n2440;
  assign n2442 = ~n192 & ~n529;
  assign n2443 = ~n128 & ~n313;
  assign n2444 = n2442 & n2443;
  assign n2445 = n2166 & n2444;
  assign n2446 = n2441 & n2445;
  assign n2447 = n2439 & n2446;
  assign n2448 = n2297 & n2447;
  assign n2449 = n1972 & n2448;
  assign n2450 = ~n418 & ~n1005;
  assign n2451 = ~n326 & ~n1060;
  assign n2452 = n2450 & n2451;
  assign n2454 = ~n443 & n2453;
  assign n2455 = n2452 & n2454;
  assign n2456 = ~n64 & ~n181;
  assign n2457 = ~n616 & n2456;
  assign n2458 = n247 & n2457;
  assign n2459 = n2455 & n2458;
  assign n2460 = n235 & n2392;
  assign n2461 = ~n494 & ~n628;
  assign n2462 = n2460 & n2461;
  assign n2463 = n1652 & n2462;
  assign n2464 = n2459 & n2463;
  assign n2465 = ~n370 & n453;
  assign n2466 = ~n553 & n738;
  assign n2467 = n2465 & n2466;
  assign n2468 = ~n300 & n1665;
  assign n2469 = n2467 & n2468;
  assign n2470 = n1517 & n2469;
  assign n2471 = n2464 & n2470;
  assign n2472 = ~n314 & ~n439;
  assign n2473 = n584 & n2472;
  assign n2474 = n1027 & n2473;
  assign n2475 = n2208 & n2474;
  assign n2476 = n1212 & n2263;
  assign n2477 = ~n226 & ~n428;
  assign n2478 = ~n1148 & n2477;
  assign n2479 = n2476 & n2478;
  assign n2480 = n2475 & n2479;
  assign n2481 = n2471 & n2480;
  assign n2482 = n2449 & n2481;
  assign n2483 = ~n227 & ~n634;
  assign n2484 = ~n390 & ~n553;
  assign n2485 = n2483 & n2484;
  assign n2486 = n1567 & n1611;
  assign n2487 = n2485 & n2486;
  assign n2488 = ~n193 & ~n409;
  assign n2489 = ~n152 & ~n790;
  assign n2490 = n2488 & n2489;
  assign n2491 = n651 & n2490;
  assign n2492 = n2487 & n2491;
  assign n2493 = ~n412 & ~n750;
  assign n2494 = ~n109 & ~n358;
  assign n2495 = n2493 & n2494;
  assign n2496 = ~n197 & n1678;
  assign n2497 = n2495 & n2496;
  assign n2498 = n679 & n1288;
  assign n2499 = n1238 & n2498;
  assign n2500 = n2497 & n2499;
  assign n2501 = n2492 & n2500;
  assign n2502 = n247 & n519;
  assign n2503 = ~n593 & n1171;
  assign n2504 = n2502 & n2503;
  assign n2505 = n2501 & n2504;
  assign n2506 = x24 & n1148;
  assign n2507 = n713 & ~n2506;
  assign n2508 = n2104 & n2507;
  assign n2509 = ~n190 & ~n1266;
  assign n2510 = ~n202 & n2509;
  assign n2511 = n2508 & n2510;
  assign n2512 = ~n428 & n2453;
  assign n2513 = n1069 & n2512;
  assign n2514 = n2511 & n2513;
  assign n2515 = ~n582 & ~n946;
  assign n2516 = ~n1405 & n2515;
  assign n2517 = n1085 & n2516;
  assign n2518 = ~n51 & ~n671;
  assign n2519 = n1188 & n2518;
  assign n2520 = ~n298 & ~n373;
  assign n2521 = ~n296 & ~n680;
  assign n2522 = n2520 & n2521;
  assign n2523 = n2519 & n2522;
  assign n2524 = n2517 & n2523;
  assign n2525 = n2514 & n2524;
  assign n2527 = ~n382 & ~n841;
  assign n2528 = n2526 & n2527;
  assign n2529 = ~n148 & ~n504;
  assign n2530 = n2528 & n2529;
  assign n2531 = ~n660 & ~n920;
  assign n2532 = ~n899 & n2531;
  assign n2533 = n2461 & n2532;
  assign n2534 = n2530 & n2533;
  assign n2535 = n1167 & n1739;
  assign n2536 = ~n156 & ~n812;
  assign n2537 = n2535 & n2536;
  assign n2538 = n2534 & n2537;
  assign n2539 = n2525 & n2538;
  assign n2540 = n2505 & n2539;
  assign n2541 = ~n208 & ~n301;
  assign n2542 = ~n347 & ~n901;
  assign n2543 = n2541 & n2542;
  assign n2544 = ~n278 & ~n362;
  assign n2545 = n1847 & n2544;
  assign n2546 = n2543 & n2545;
  assign n2547 = ~n312 & ~n449;
  assign n2548 = ~n620 & n2547;
  assign n2549 = n2546 & n2548;
  assign n2552 = ~n231 & ~n617;
  assign n2553 = n1554 & n2552;
  assign n2554 = n2551 & n2553;
  assign n2555 = n2549 & n2554;
  assign n2556 = ~n326 & ~n514;
  assign n2557 = ~n656 & n2556;
  assign n2558 = n1029 & n2557;
  assign n2559 = n1436 & n2558;
  assign n2560 = n419 & ~n740;
  assign n2561 = ~n199 & ~n292;
  assign n2562 = ~n120 & n2561;
  assign n2563 = n2560 & n2562;
  assign n2564 = n457 & n536;
  assign n2565 = n274 & n2564;
  assign n2566 = n2563 & n2565;
  assign n2567 = n2559 & n2566;
  assign n2568 = n2555 & n2567;
  assign n2569 = ~n192 & ~n819;
  assign n2570 = ~n79 & ~n218;
  assign n2571 = n2569 & n2570;
  assign n2572 = n2314 & n2571;
  assign n2573 = n2568 & n2572;
  assign n2574 = n2540 & n2573;
  assign n2575 = ~n2482 & ~n2574;
  assign n2576 = n2425 & n2575;
  assign n2577 = ~n343 & ~n475;
  assign n2578 = ~n170 & n2577;
  assign n2579 = n1292 & n2578;
  assign n2580 = n578 & n2579;
  assign n2581 = ~n350 & ~n424;
  assign n2582 = ~n378 & ~n497;
  assign n2583 = n2581 & n2582;
  assign n2584 = ~n344 & ~n592;
  assign n2585 = n1352 & n2584;
  assign n2586 = n2583 & n2585;
  assign n2587 = n2580 & n2586;
  assign n2588 = ~n93 & ~n273;
  assign n2589 = ~n763 & n2588;
  assign n2590 = ~n110 & ~n300;
  assign n2591 = ~n385 & n2590;
  assign n2592 = n2589 & n2591;
  assign n2593 = ~n270 & ~n709;
  assign n2594 = n1771 & n2593;
  assign n2596 = n1103 & n2595;
  assign n2597 = n2594 & n2596;
  assign n2598 = n2592 & n2597;
  assign n2599 = n1886 & n2598;
  assign n2600 = n2587 & n2599;
  assign n2601 = n1096 & n2600;
  assign n2602 = ~n185 & ~n237;
  assign n2603 = ~n346 & ~n440;
  assign n2604 = n2602 & n2603;
  assign n2605 = ~n337 & ~n531;
  assign n2606 = n2604 & n2605;
  assign n2607 = ~n120 & n1328;
  assign n2608 = ~n256 & ~n800;
  assign n2609 = n2607 & n2608;
  assign n2610 = n2606 & n2609;
  assign n2611 = n2505 & n2610;
  assign n2612 = n2601 & n2611;
  assign n2613 = ~n358 & ~n552;
  assign n2614 = ~n304 & n2613;
  assign n2615 = ~n461 & ~n683;
  assign n2616 = n1324 & n2615;
  assign n2617 = n2614 & n2616;
  assign n2619 = n2617 & n2618;
  assign n2620 = ~n333 & n2526;
  assign n2621 = n419 & n1976;
  assign n2622 = n2620 & n2621;
  assign n2624 = n2577 & n2623;
  assign n2626 = n2624 & n2625;
  assign n2627 = n2622 & n2626;
  assign n2628 = n2619 & n2627;
  assign n2629 = ~n110 & ~n1060;
  assign n2630 = ~n375 & n2629;
  assign n2631 = n2334 & n2630;
  assign n2632 = ~n138 & ~n610;
  assign n2633 = n2631 & n2632;
  assign n2635 = ~n193 & ~n612;
  assign n2636 = n2634 & n2635;
  assign n2637 = ~n362 & ~n442;
  assign n2638 = n2636 & n2637;
  assign n2639 = ~n227 & ~n410;
  assign n2640 = ~n456 & ~n592;
  assign n2641 = n2639 & n2640;
  assign n2642 = n2638 & n2641;
  assign n2643 = n2633 & n2642;
  assign n2644 = n2628 & n2643;
  assign n2645 = n1939 & n2644;
  assign n2646 = n279 & ~n1405;
  assign n2647 = n191 & n530;
  assign n2648 = n2646 & n2647;
  assign n2649 = ~n755 & ~n948;
  assign n2650 = n1940 & n2649;
  assign n2651 = n352 & n961;
  assign n2652 = n2650 & n2651;
  assign n2653 = n2648 & n2652;
  assign n2655 = n282 & n2654;
  assign n2656 = ~n146 & ~n494;
  assign n2657 = n986 & n2656;
  assign n2658 = n2655 & n2657;
  assign n2659 = n451 & n2658;
  assign n2660 = n2653 & n2659;
  assign n2661 = ~n104 & ~n320;
  assign n2662 = ~n117 & ~n183;
  assign n2663 = n2661 & n2662;
  assign n2664 = n1271 & n2663;
  assign n2665 = ~n120 & ~n929;
  assign n2666 = ~n347 & n2665;
  assign n2667 = n2664 & n2666;
  assign n2668 = n2660 & n2667;
  assign n2669 = n2645 & n2668;
  assign n2670 = n2612 & n2669;
  assign n2671 = ~n2574 & ~n2670;
  assign n2672 = ~n2612 & ~n2669;
  assign n2673 = ~n2482 & n2672;
  assign n2674 = ~n2671 & ~n2673;
  assign n2675 = ~n2423 & n2575;
  assign n2676 = n2674 & ~n2675;
  assign n2677 = ~n2576 & n2676;
  assign n2678 = ~n2358 & ~n2423;
  assign n2679 = n2672 & n2678;
  assign n2680 = n2677 & ~n2679;
  assign n2681 = n956 & n1059;
  assign n2682 = n1629 & n2681;
  assign n2683 = ~n605 & n893;
  assign n2684 = ~n337 & n1548;
  assign n2685 = n2683 & n2684;
  assign n2686 = ~n300 & ~n841;
  assign n2687 = n282 & n2686;
  assign n2688 = n1788 & n2687;
  assign n2689 = n2685 & n2688;
  assign n2690 = n2244 & n2689;
  assign n2691 = n2682 & n2690;
  assign n2700 = n2691 & n2699;
  assign n2701 = ~n327 & ~n429;
  assign n2702 = ~n791 & n2701;
  assign n2703 = n311 & n2702;
  assign n2704 = n118 & ~n509;
  assign n2705 = n2416 & n2704;
  assign n2706 = n2703 & n2705;
  assign n2707 = ~n406 & ~n948;
  assign n2708 = ~n136 & n2707;
  assign n2709 = n1359 & n2708;
  assign n2710 = n1164 & n2639;
  assign n2711 = ~n758 & ~n812;
  assign n2712 = n2710 & n2711;
  assign n2713 = n2709 & n2712;
  assign n2714 = n2706 & n2713;
  assign n2715 = n2587 & n2714;
  assign n2716 = n1053 & n2715;
  assign n2717 = n2700 & n2716;
  assign n2718 = n1095 & n2717;
  assign n2719 = n566 & n2718;
  assign n2720 = n2669 & n2719;
  assign n2722 = n371 & n2721;
  assign n2723 = ~n93 & ~n265;
  assign n2724 = n2623 & n2723;
  assign n2725 = n2722 & n2724;
  assign n2726 = n956 & n2725;
  assign n2727 = n149 & ~n402;
  assign n2728 = n462 & n2727;
  assign n2729 = n2709 & n2728;
  assign n2730 = n2726 & n2729;
  assign n2739 = ~n143 & ~n1060;
  assign n2740 = n419 & n2739;
  assign n2741 = ~n540 & ~n850;
  assign n2742 = ~n612 & n2741;
  assign n2743 = n2740 & n2742;
  assign n2744 = n472 & n1574;
  assign n2745 = n2743 & n2744;
  assign n2746 = n2738 & n2745;
  assign n2747 = n2730 & n2746;
  assign n2748 = ~n336 & ~n797;
  assign n2749 = n2114 & n2748;
  assign n2750 = ~n79 & ~n382;
  assign n2751 = ~n799 & n2750;
  assign n2752 = n2749 & n2751;
  assign n2753 = ~n272 & ~n343;
  assign n2754 = n1073 & n2753;
  assign n2755 = ~n326 & ~n506;
  assign n2756 = ~n762 & n2755;
  assign n2757 = n2754 & n2756;
  assign n2758 = n2752 & n2757;
  assign n2759 = n1673 & n2758;
  assign n2761 = ~n314 & ~n666;
  assign n2762 = ~n128 & ~n141;
  assign n2763 = n2761 & n2762;
  assign n2764 = n2760 & n2763;
  assign n2765 = ~n218 & ~n787;
  assign n2766 = n285 & n2765;
  assign n2767 = n493 & n1124;
  assign n2768 = n2766 & n2767;
  assign n2769 = n2764 & n2768;
  assign n2770 = n2504 & n2769;
  assign n2774 = n1810 & n2773;
  assign n2775 = n532 & n1741;
  assign n2776 = n602 & n2775;
  assign n2777 = n2774 & n2776;
  assign n2778 = ~n331 & ~n683;
  assign n2779 = n1882 & n2778;
  assign n2780 = ~n208 & ~n442;
  assign n2781 = n1853 & n2780;
  assign n2782 = n2779 & n2781;
  assign n2783 = n2777 & n2782;
  assign n2784 = n2770 & n2783;
  assign n2785 = n2759 & n2784;
  assign n2786 = n2747 & n2785;
  assign n2787 = ~n57 & ~n308;
  assign n2788 = n2165 & n2787;
  assign n2789 = ~n128 & n2723;
  assign n2790 = n2788 & n2789;
  assign n2791 = ~n83 & n297;
  assign n2792 = n2790 & n2791;
  assign n2793 = ~n133 & ~n283;
  assign n2794 = ~n659 & n2793;
  assign n2795 = ~n186 & ~n402;
  assign n2796 = ~n103 & ~n683;
  assign n2797 = n2795 & n2796;
  assign n2798 = n2794 & n2797;
  assign n2799 = ~n134 & ~n174;
  assign n2800 = ~n709 & n2799;
  assign n2801 = ~n227 & n781;
  assign n2802 = n2800 & n2801;
  assign n2803 = n2798 & n2802;
  assign n2804 = n2792 & n2803;
  assign n2805 = ~n509 & ~n763;
  assign n2807 = n2805 & n2806;
  assign n2809 = n2040 & n2808;
  assign n2810 = n2807 & n2809;
  assign n2811 = ~n273 & ~n469;
  assign n2812 = n2051 & n2811;
  assign n2814 = ~n323 & n2813;
  assign n2815 = n2812 & n2814;
  assign n2816 = n2810 & n2815;
  assign n2817 = ~n156 & ~n266;
  assign n2818 = n2349 & n2817;
  assign n2819 = ~n751 & ~n1227;
  assign n2820 = ~n115 & ~n390;
  assign n2821 = n2819 & n2820;
  assign n2822 = n2818 & n2821;
  assign n2823 = n2816 & n2822;
  assign n2824 = n2804 & n2823;
  assign n2825 = ~n257 & ~n312;
  assign n2826 = ~n396 & n2825;
  assign n2827 = ~n750 & ~n901;
  assign n2828 = n2590 & n2827;
  assign n2829 = n2826 & n2828;
  assign n2830 = n1001 & n1231;
  assign n2831 = n2829 & n2830;
  assign n2832 = n1263 & n2577;
  assign n2833 = n1491 & n2063;
  assign n2834 = n925 & n2833;
  assign n2835 = n2832 & n2834;
  assign n2836 = n2831 & n2835;
  assign n2837 = n2331 & n2836;
  assign n2838 = ~n189 & ~n553;
  assign n2839 = ~n136 & n2838;
  assign n2840 = ~n518 & ~n946;
  assign n2841 = n2839 & n2840;
  assign n2842 = ~n723 & ~n800;
  assign n2843 = ~n540 & n2842;
  assign n2844 = n2841 & n2843;
  assign n2845 = ~n74 & ~n531;
  assign n2846 = ~n417 & ~n819;
  assign n2847 = n2845 & n2846;
  assign n2848 = ~n634 & ~n675;
  assign n2849 = n2847 & n2848;
  assign n2850 = ~n359 & ~n524;
  assign n2851 = n1288 & n2850;
  assign n2852 = n2849 & n2851;
  assign n2853 = n2844 & n2852;
  assign n2854 = ~n392 & n498;
  assign n2855 = ~n476 & ~n506;
  assign n2856 = ~n298 & n2855;
  assign n2857 = n2854 & n2856;
  assign n2858 = n1609 & n2857;
  assign n2859 = n2853 & n2858;
  assign n2860 = n2837 & n2859;
  assign n2861 = n2824 & n2860;
  assign n2862 = n2786 & n2861;
  assign n2863 = ~n2720 & ~n2862;
  assign n2864 = n2680 & ~n2863;
  assign n2865 = ~n566 & ~n2718;
  assign n2866 = n2861 & ~n2865;
  assign n2867 = n2669 & n2862;
  assign n2868 = ~n2866 & ~n2867;
  assign n2869 = n2719 & n2786;
  assign n2870 = n2868 & ~n2869;
  assign n2871 = ~n2864 & n2870;
  assign n2872 = ~n566 & n2871;
  assign n2873 = n368 & ~n2872;
  assign n2874 = ~n948 & ~n2506;
  assign n2875 = ~n237 & ~n656;
  assign n2876 = n2874 & n2875;
  assign n2877 = ~n120 & ~n284;
  assign n2878 = ~n524 & n2877;
  assign n2879 = n2876 & n2878;
  assign n2880 = n305 & n2392;
  assign n2881 = n223 & n2880;
  assign n2882 = n2879 & n2881;
  assign n2883 = ~n233 & ~n385;
  assign n2884 = ~n99 & n2883;
  assign n2885 = n1483 & n2884;
  assign n2886 = n692 & n1159;
  assign n2887 = n2885 & n2886;
  assign n2888 = n2882 & n2887;
  assign n2889 = ~n262 & n875;
  assign n2890 = ~n396 & ~n432;
  assign n2891 = n1421 & n2890;
  assign n2892 = n2889 & n2891;
  assign n2893 = n2803 & n2892;
  assign n2894 = n2888 & n2893;
  assign n2895 = ~n552 & ~n740;
  assign n2896 = ~n263 & ~n553;
  assign n2897 = n2895 & n2896;
  assign n2898 = ~n359 & ~n610;
  assign n2899 = ~n254 & ~n605;
  assign n2900 = n2898 & n2899;
  assign n2901 = n2897 & n2900;
  assign n2902 = n856 & n2526;
  assign n2903 = n2634 & n2902;
  assign n2904 = n2901 & n2903;
  assign n2905 = n2894 & n2904;
  assign n2906 = n1902 & n2527;
  assign n2907 = n2787 & n2906;
  assign n2908 = ~n74 & ~n797;
  assign n2909 = n420 & n2908;
  assign n2910 = n2907 & n2909;
  assign n2911 = ~n492 & ~n527;
  assign n2912 = n530 & n2911;
  assign n2913 = n551 & n1785;
  assign n2914 = n2912 & n2913;
  assign n2915 = n2910 & n2914;
  assign n2916 = ~n475 & ~n929;
  assign n2917 = ~n1166 & n2916;
  assign n2918 = ~n1482 & n2584;
  assign n2919 = n2917 & n2918;
  assign n2920 = n1832 & n2919;
  assign n2921 = n2915 & n2920;
  assign n2922 = ~n209 & ~n243;
  assign n2923 = ~n250 & ~n300;
  assign n2924 = n2922 & n2923;
  assign n2925 = ~n266 & ~n751;
  assign n2926 = n2924 & n2925;
  assign n2927 = ~n351 & n2625;
  assign n2928 = n2926 & n2927;
  assign n2929 = n1622 & n1967;
  assign n2930 = n2928 & n2929;
  assign n2931 = n2921 & n2930;
  assign n2932 = n1422 & n1782;
  assign n2933 = n473 & n2051;
  assign n2934 = n2932 & n2933;
  assign n2935 = ~n87 & ~n152;
  assign n2936 = ~n98 & ~n336;
  assign n2937 = n2935 & n2936;
  assign n2938 = ~n51 & ~n256;
  assign n2939 = n2298 & n2938;
  assign n2940 = n2937 & n2939;
  assign n2941 = n2934 & n2940;
  assign n2943 = ~n231 & ~n429;
  assign n2944 = n2942 & n2943;
  assign n2945 = ~n115 & n2811;
  assign n2946 = n2944 & n2945;
  assign n2947 = n2941 & n2946;
  assign n2948 = n1398 & n1934;
  assign n2949 = ~n320 & n2207;
  assign n2950 = n508 & n2949;
  assign n2951 = n2948 & n2950;
  assign n2952 = n2947 & n2951;
  assign n2953 = n2931 & n2952;
  assign n2954 = n2905 & n2953;
  assign n2955 = n2873 & n2954;
  assign n2956 = n566 & ~n2871;
  assign n2957 = ~n405 & ~n928;
  assign n2958 = n2827 & n2957;
  assign n2959 = n66 & n1109;
  assign n2960 = ~n185 & ~n2959;
  assign n2961 = ~n553 & n2960;
  assign n2962 = n2958 & n2961;
  assign n2963 = ~n330 & ~n946;
  assign n2964 = n2187 & n2963;
  assign n2965 = ~n57 & ~n310;
  assign n2966 = n2964 & n2965;
  assign n2967 = n2962 & n2966;
  assign n2969 = ~n93 & ~n919;
  assign n2970 = n2968 & n2969;
  assign n2971 = n486 & n2013;
  assign n2972 = n2970 & n2971;
  assign n2973 = n780 & n2972;
  assign n2974 = n2967 & n2973;
  assign n2976 = ~n370 & n2975;
  assign n2977 = n994 & n1514;
  assign n2978 = n2976 & n2977;
  assign n2979 = n1999 & n2978;
  assign n2980 = n2974 & n2979;
  assign n2981 = n1342 & n1943;
  assign n2982 = ~n156 & ~n627;
  assign n2983 = ~n111 & ~n295;
  assign n2984 = n2982 & n2983;
  assign n2985 = n2981 & n2984;
  assign n2987 = n2165 & n2986;
  assign n2988 = n2799 & n2987;
  assign n2989 = n2985 & n2988;
  assign n2990 = ~n221 & ~n456;
  assign n2991 = n854 & n2990;
  assign n2992 = n1263 & n2991;
  assign n2993 = ~n87 & n526;
  assign n2994 = n2992 & n2993;
  assign n2995 = n2989 & n2994;
  assign n2996 = n2980 & n2995;
  assign n2997 = ~n403 & ~n929;
  assign n2998 = ~n504 & ~n549;
  assign n2999 = n2997 & n2998;
  assign n3000 = n1496 & n2999;
  assign n3001 = n2889 & n3000;
  assign n3002 = n684 & n792;
  assign n3003 = n3001 & n3002;
  assign n3004 = ~n476 & ~n1227;
  assign n3006 = n3004 & n3005;
  assign n3007 = ~n751 & ~n1858;
  assign n3008 = n3006 & n3007;
  assign n3009 = ~n244 & ~n440;
  assign n3010 = n2382 & n3009;
  assign n3011 = n1116 & n2143;
  assign n3012 = n3010 & n3011;
  assign n3013 = ~n410 & ~n659;
  assign n3014 = n184 & n3013;
  assign n3015 = n1994 & n3014;
  assign n3016 = n3012 & n3015;
  assign n3017 = n3008 & n3016;
  assign n3018 = n3003 & n3017;
  assign n3019 = ~n199 & ~n494;
  assign n3020 = ~n99 & ~n1266;
  assign n3021 = n3019 & n3020;
  assign n3022 = ~n141 & ~n193;
  assign n3023 = n3021 & n3022;
  assign n3024 = n1445 & n3023;
  assign n3025 = ~n312 & ~n417;
  assign n3026 = n123 & n3025;
  assign n3027 = ~n975 & n3026;
  assign n3028 = n3024 & n3027;
  assign n3029 = ~n95 & ~n424;
  assign n3030 = ~n208 & n3029;
  assign n3031 = n759 & n1328;
  assign n3032 = n3030 & n3031;
  assign n3033 = ~n216 & ~n605;
  assign n3034 = n3032 & n3033;
  assign n3035 = n3028 & n3034;
  assign n3036 = n3018 & n3035;
  assign n3037 = n2996 & n3036;
  assign n3099 = n3037 & n3098;
  assign n3100 = n2956 & n3099;
  assign n3101 = ~n3037 & ~n3098;
  assign n3102 = n2954 & ~n3101;
  assign n3103 = n368 & n3099;
  assign n3104 = ~n3102 & ~n3103;
  assign n3105 = ~n3100 & n3104;
  assign n3106 = ~n2955 & n3105;
  assign n3406 = n3098 & ~n3106;
  assign n3407 = ~n3196 & ~n3406;
  assign n3408 = n3270 & ~n3407;
  assign n3409 = ~n3351 & ~n3408;
  assign n3410 = n3404 & ~n3409;
  assign n3420 = ~n281 & n3388;
  assign n3421 = n1481 & n3420;
  assign n3422 = n3419 & n3421;
  assign n3423 = n66 & ~n76;
  assign n3424 = ~n61 & ~n3423;
  assign n3425 = n3422 & n3424;
  assign n3429 = ~n79 & ~n226;
  assign n3430 = n3428 & n3429;
  assign n3431 = n3425 & n3430;
  assign n3877 = ~n3410 & ~n3431;
  assign n3286 = ~n3098 & n3106;
  assign n3287 = ~n3270 & n3286;
  assign n3288 = ~n3196 & ~n3270;
  assign n3289 = ~n3287 & ~n3288;
  assign n3352 = n3289 & n3351;
  assign n3405 = ~n3352 & ~n3404;
  assign n3876 = ~n3405 & n3431;
  assign n5756 = n3877 ^ n3876;
  assign n5757 = n3875 & n5756;
  assign n5758 = n5757 ^ n3876;
  assign n11852 = n41 & n5758;
  assign n11853 = n3875 & ~n11852;
  assign n11854 = x31 & ~n11853;
  assign n11878 = n11854 ^ n11839;
  assign n11879 = n11851 & ~n11878;
  assign n11880 = n11879 ^ n11854;
  assign n11760 = n11759 ^ x29;
  assign n11761 = n11760 ^ n11413;
  assign n11855 = n11854 ^ n11851;
  assign n4519 = ~n152 & ~n687;
  assign n4520 = ~n333 & n4519;
  assign n4521 = n2874 & n4520;
  assign n4522 = ~n298 & ~n326;
  assign n4523 = n1273 & n4522;
  assign n4524 = n4521 & n4523;
  assign n3824 = ~n308 & ~n424;
  assign n4525 = n282 & n2615;
  assign n4526 = n3824 & n4525;
  assign n3596 = ~n476 & ~n714;
  assign n4527 = ~n126 & n3596;
  assign n4528 = n4526 & n4527;
  assign n4529 = n4524 & n4528;
  assign n4530 = ~n1005 & n1905;
  assign n4531 = n2817 & n3110;
  assign n4532 = n4530 & n4531;
  assign n4533 = n4529 & n4532;
  assign n4534 = ~n344 & ~n610;
  assign n4535 = n2233 & n4534;
  assign n4536 = n2570 & n4535;
  assign n4537 = ~n148 & ~n557;
  assign n4538 = ~n164 & n4537;
  assign n4539 = ~n170 & ~n1060;
  assign n4540 = n1688 & n4539;
  assign n4541 = n4538 & n4540;
  assign n4542 = n4536 & n4541;
  assign n4543 = n4533 & n4542;
  assign n10887 = n118 & n3033;
  assign n10888 = ~n244 & ~n402;
  assign n10889 = n2590 & n10888;
  assign n10890 = n10887 & n10889;
  assign n10891 = n597 & n1406;
  assign n10892 = n833 & n1302;
  assign n10893 = n10891 & n10892;
  assign n10894 = n10890 & n10893;
  assign n10895 = ~n390 & ~n1047;
  assign n10896 = ~n361 & ~n723;
  assign n10897 = n10895 & n10896;
  assign n10898 = ~n354 & ~n524;
  assign n10899 = n1306 & n10898;
  assign n10900 = n10897 & n10899;
  assign n10901 = n10894 & n10900;
  assign n5116 = n495 & n2895;
  assign n5117 = ~n283 & ~n525;
  assign n5118 = ~n320 & ~n535;
  assign n5119 = n5117 & n5118;
  assign n5120 = n5116 & n5119;
  assign n5121 = ~n529 & ~n1266;
  assign n5122 = n2202 & n5121;
  assign n5123 = n2170 & n5122;
  assign n5124 = n5120 & n5123;
  assign n4739 = ~n99 & ~n109;
  assign n5033 = ~n296 & n4739;
  assign n10902 = n144 & n294;
  assign n10903 = n5033 & n10902;
  assign n10904 = n1133 & n10903;
  assign n10905 = n5124 & n10904;
  assign n10906 = n10901 & n10905;
  assign n10907 = n4543 & n10906;
  assign n10908 = n2323 & n10907;
  assign n11241 = n10908 ^ x26;
  assign n4566 = ~n110 & ~n190;
  assign n5032 = n937 & n4566;
  assign n4565 = ~n202 & ~n216;
  assign n11242 = ~n358 & n4565;
  assign n11243 = n5032 & n11242;
  assign n11244 = ~n244 & ~n336;
  assign n11245 = n782 & n11244;
  assign n11246 = n2353 & n11245;
  assign n11247 = n11243 & n11246;
  assign n11248 = ~n146 & ~n558;
  assign n11249 = n2165 & n11248;
  assign n11250 = ~n120 & n11249;
  assign n11251 = ~n362 & ~n582;
  assign n11252 = n1363 & n11251;
  assign n11253 = n302 & n860;
  assign n11254 = n11252 & n11253;
  assign n11255 = n11250 & n11254;
  assign n11256 = n11247 & n11255;
  assign n3912 = ~n185 & n635;
  assign n3913 = ~n222 & ~n518;
  assign n3914 = n3912 & n3913;
  assign n4232 = ~n197 & ~n262;
  assign n11257 = n2632 & n4232;
  assign n11258 = n530 & n2035;
  assign n11259 = n11257 & n11258;
  assign n11260 = ~n95 & ~n497;
  assign n11261 = ~n298 & ~n331;
  assign n11262 = n11260 & n11261;
  assign n11263 = n11259 & n11262;
  assign n11264 = n3914 & n11263;
  assign n11265 = n11256 & n11264;
  assign n11266 = n235 & n3064;
  assign n4198 = ~n181 & ~n409;
  assign n11267 = n2432 & n4198;
  assign n11268 = n11266 & n11267;
  assign n3500 = ~n148 & n2385;
  assign n11269 = ~n253 & ~n334;
  assign n11270 = ~n630 & n11269;
  assign n11271 = n3500 & n11270;
  assign n11272 = n11268 & n11271;
  assign n11273 = n3002 & n11272;
  assign n5047 = ~n323 & ~n750;
  assign n5048 = ~n250 & n5047;
  assign n5049 = ~n192 & ~n919;
  assign n5050 = n2212 & n5049;
  assign n5051 = n5048 & n5050;
  assign n5052 = n1284 & n5051;
  assign n5381 = ~n64 & ~n382;
  assign n5382 = ~n104 & n5381;
  assign n11274 = ~n277 & ~n1536;
  assign n11275 = n5382 & n11274;
  assign n11276 = ~n237 & ~n628;
  assign n11277 = n11275 & n11276;
  assign n11278 = n5052 & n11277;
  assign n11279 = n11273 & n11278;
  assign n11280 = n11265 & n11279;
  assign n11281 = n1249 & n11280;
  assign n11282 = n11281 ^ n10908;
  assign n11283 = n11241 & ~n11282;
  assign n11284 = n11283 ^ x26;
  assign n10091 = n649 & n1656;
  assign n10092 = ~n812 & n2623;
  assign n10093 = n10091 & n10092;
  assign n10094 = ~n156 & n282;
  assign n10095 = n371 & n10094;
  assign n5442 = ~n452 & ~n710;
  assign n5443 = ~n326 & n5442;
  assign n10096 = n1754 & n5443;
  assign n10097 = n10095 & n10096;
  assign n3453 = ~n337 & ~n592;
  assign n4380 = ~n277 & ~n588;
  assign n10098 = n3453 & n4380;
  assign n10099 = n4065 & n10098;
  assign n10100 = n1036 & n10099;
  assign n10101 = n10097 & n10100;
  assign n10102 = n10093 & n10101;
  assign n10103 = n1533 & n10102;
  assign n11285 = ~n514 & ~n517;
  assign n11286 = ~n432 & ~n478;
  assign n11287 = n11285 & n11286;
  assign n11288 = n1209 & n2207;
  assign n11289 = n11287 & n11288;
  assign n11290 = n3235 & n11289;
  assign n5618 = ~n576 & n2145;
  assign n11291 = ~n691 & n5618;
  assign n4100 = ~n155 & ~n359;
  assign n11292 = n606 & n4100;
  assign n5520 = ~n333 & ~n1005;
  assign n11293 = ~n171 & ~n417;
  assign n11294 = n5520 & n11293;
  assign n11295 = n11292 & n11294;
  assign n11296 = n11291 & n11295;
  assign n11297 = n11290 & n11296;
  assign n3529 = ~n791 & n925;
  assign n11298 = ~n79 & ~n167;
  assign n11299 = ~n231 & ~n295;
  assign n11300 = n11298 & n11299;
  assign n11301 = n3529 & n11300;
  assign n11302 = ~n115 & ~n308;
  assign n11303 = n2515 & n11302;
  assign n11304 = ~n109 & ~n529;
  assign n11305 = n1039 & n11304;
  assign n11306 = n11303 & n11305;
  assign n11307 = n11301 & n11306;
  assign n11308 = n2973 & n11307;
  assign n11309 = n11297 & n11308;
  assign n3712 = ~n410 & ~n518;
  assign n11310 = n2527 & n3712;
  assign n11311 = ~n500 & n3111;
  assign n11312 = n11310 & n11311;
  assign n5091 = ~n126 & ~n494;
  assign n5092 = ~n343 & n5091;
  assign n11313 = ~n266 & ~n458;
  assign n11314 = ~n143 & ~n164;
  assign n11315 = n11313 & n11314;
  assign n11316 = n5092 & n11315;
  assign n11317 = n11312 & n11316;
  assign n4014 = ~n373 & n1976;
  assign n11318 = n184 & ~n610;
  assign n11319 = n2485 & n11318;
  assign n11320 = n4014 & n11319;
  assign n11321 = n11317 & n11320;
  assign n11322 = n11309 & n11321;
  assign n11323 = n10103 & n11322;
  assign n5769 = ~n3352 & ~n3409;
  assign n5770 = n5769 ^ n3404;
  assign n11325 = n41 & ~n5770;
  assign n11326 = n54 & ~n3270;
  assign n11327 = n91 & ~n3351;
  assign n11328 = ~n11326 & ~n11327;
  assign n11329 = ~n11325 & n11328;
  assign n11330 = x31 & ~n11329;
  assign n3671 = ~x31 & n54;
  assign n11331 = ~n3351 & n3671;
  assign n3676 = ~x31 & n41;
  assign n11332 = ~n3404 & n3676;
  assign n11333 = ~n11331 & ~n11332;
  assign n11334 = ~n11330 & n11333;
  assign n11414 = n11323 & n11334;
  assign n11415 = n11284 & n11414;
  assign n11416 = ~n11323 & ~n11334;
  assign n11417 = ~n11284 & n11416;
  assign n11418 = ~n11415 & ~n11417;
  assign n11419 = n11418 ^ n11413;
  assign n3411 = ~n3405 & ~n3410;
  assign n11371 = x31 & n3411;
  assign n11372 = n11371 ^ n3431;
  assign n11373 = n41 & ~n11372;
  assign n3669 = x31 & n54;
  assign n11374 = ~n3351 & n3669;
  assign n3672 = x31 & n91;
  assign n3673 = ~n3671 & ~n3672;
  assign n11375 = ~n3404 & ~n3673;
  assign n11376 = ~n11374 & ~n11375;
  assign n11377 = ~n11373 & n11376;
  assign n42 = x27 ^ x26;
  assign n43 = x29 ^ x28;
  assign n3273 = x28 ^ x27;
  assign n3274 = n43 & ~n3273;
  assign n3275 = ~n42 & n3274;
  assign n11369 = n3275 & ~n3875;
  assign n11370 = ~x29 & ~n11369;
  assign n11378 = n11377 ^ n11370;
  assign n11420 = n11419 ^ n11378;
  assign n44 = n42 & n43;
  assign n11336 = n44 & n5758;
  assign n3277 = ~n42 & n3273;
  assign n11337 = n3277 & ~n3875;
  assign n11338 = n3275 & ~n3431;
  assign n11339 = ~n11337 & ~n11338;
  assign n11340 = ~n11336 & n11339;
  assign n11341 = n11340 ^ x29;
  assign n11324 = n11323 ^ n11284;
  assign n11335 = n11334 ^ n11324;
  assign n11342 = n11341 ^ n11335;
  assign n11109 = n3287 ^ x30;
  assign n11110 = n41 & n11109;
  assign n11111 = n11110 ^ x29;
  assign n11112 = n3196 & ~n11111;
  assign n11113 = ~n91 & n3098;
  assign n11114 = n41 & ~n3196;
  assign n11115 = ~n11113 & ~n11114;
  assign n11116 = n3106 & n11115;
  assign n11117 = n3270 & ~n11116;
  assign n11118 = n41 & ~n3098;
  assign n11119 = ~n54 & n3196;
  assign n11120 = ~n11118 & ~n11119;
  assign n11121 = ~n3106 & n11120;
  assign n11122 = n11117 & ~n11121;
  assign n11123 = ~n3106 & n3288;
  assign n11124 = ~n54 & ~n11123;
  assign n11125 = n11113 & ~n11124;
  assign n11126 = ~n11122 & ~n11125;
  assign n11127 = ~n11112 & n11126;
  assign n11106 = n41 & ~n3270;
  assign n11107 = n54 & ~n3196;
  assign n11108 = ~n11106 & ~n11107;
  assign n11128 = n11127 ^ n11108;
  assign n11129 = ~x31 & ~n11128;
  assign n11130 = n11129 ^ n11127;
  assign n11131 = n194 & n1378;
  assign n4552 = ~n245 & ~n503;
  assign n11132 = n1406 & n4552;
  assign n11133 = n11131 & n11132;
  assign n3553 = ~n281 & ~n671;
  assign n11134 = ~n1005 & ~n1345;
  assign n11135 = ~n284 & n11134;
  assign n11136 = n3553 & n11135;
  assign n11137 = n11133 & n11136;
  assign n11138 = n2837 & n11137;
  assign n4731 = ~n326 & ~n354;
  assign n4732 = ~n375 & ~n463;
  assign n4733 = n4731 & n4732;
  assign n4734 = ~n243 & ~n928;
  assign n4735 = n4733 & n4734;
  assign n4736 = ~n173 & ~n201;
  assign n4737 = n1126 & n4736;
  assign n4738 = n4735 & n4737;
  assign n4788 = ~n283 & n2943;
  assign n11139 = n297 & ~n666;
  assign n11140 = n4788 & n11139;
  assign n11141 = ~n183 & n419;
  assign n11142 = n2084 & n11141;
  assign n11143 = n11140 & n11142;
  assign n4141 = ~n373 & ~n560;
  assign n11144 = ~n233 & ~n272;
  assign n11145 = n4141 & n11144;
  assign n11146 = n397 & n536;
  assign n11147 = n11145 & n11146;
  assign n3737 = ~n541 & ~n550;
  assign n11148 = ~n269 & ~n382;
  assign n11149 = n3737 & n11148;
  assign n11150 = n990 & n3137;
  assign n11151 = n11149 & n11150;
  assign n11152 = n11147 & n11151;
  assign n11153 = n11143 & n11152;
  assign n11154 = n4738 & n11153;
  assign n11155 = ~n256 & n738;
  assign n4555 = ~n74 & ~n497;
  assign n11156 = n665 & n4555;
  assign n11157 = n11155 & n11156;
  assign n11158 = ~n634 & n2634;
  assign n11159 = n220 & n11158;
  assign n11160 = n11157 & n11159;
  assign n11161 = n407 & n999;
  assign n11162 = n1158 & n1183;
  assign n11163 = n11161 & n11162;
  assign n11164 = n11160 & n11163;
  assign n11165 = ~n504 & ~n740;
  assign n11166 = ~n146 & ~n308;
  assign n11167 = n11165 & n11166;
  assign n11168 = ~n514 & ~n710;
  assign n11169 = n11167 & n11168;
  assign n11016 = ~n461 & ~n709;
  assign n11170 = ~n323 & ~n518;
  assign n11171 = n11016 & n11170;
  assign n11172 = n889 & n11171;
  assign n11173 = n11169 & n11172;
  assign n11174 = n2321 & n11173;
  assign n11175 = n11164 & n11174;
  assign n11176 = n11154 & n11175;
  assign n11177 = n11138 & n11176;
  assign n11343 = ~n11130 & n11177;
  assign n3988 = n3289 & ~n3408;
  assign n3989 = n3988 ^ n3351;
  assign n11344 = n41 & ~n3989;
  assign n11345 = n91 & ~n3270;
  assign n11346 = x31 & ~n11107;
  assign n11347 = ~n11345 & n11346;
  assign n11348 = ~n11344 & n11347;
  assign n11349 = n41 & ~n3351;
  assign n11350 = ~x31 & ~n11349;
  assign n11351 = ~n11326 & n11350;
  assign n11352 = ~n11348 & ~n11351;
  assign n11353 = n11281 ^ x26;
  assign n11354 = n11352 & n11353;
  assign n11355 = n11343 & ~n11354;
  assign n11356 = ~n11352 & ~n11353;
  assign n11357 = n10908 & ~n11356;
  assign n11358 = ~n11355 & n11357;
  assign n11359 = n11130 & ~n11177;
  assign n11360 = n11359 ^ n11352;
  assign n11361 = ~n10908 & ~n11353;
  assign n11362 = n11361 ^ n11352;
  assign n11363 = n11360 & ~n11362;
  assign n11364 = n11363 ^ n11359;
  assign n11365 = ~n11358 & ~n11364;
  assign n11366 = n11365 ^ n11335;
  assign n11367 = ~n11342 & n11366;
  assign n11368 = n11367 ^ n11341;
  assign n11421 = n11420 ^ n11368;
  assign n4352 = ~n301 & ~n841;
  assign n4353 = n559 & n4352;
  assign n4354 = n264 & n1918;
  assign n4355 = n4353 & n4354;
  assign n4356 = ~n524 & ~n544;
  assign n4357 = n2635 & n4356;
  assign n4358 = ~n359 & ~n369;
  assign n4359 = n4357 & n4358;
  assign n4360 = ~n202 & ~n652;
  assign n4361 = n1180 & n4360;
  assign n4362 = n486 & n4361;
  assign n4363 = n4359 & n4362;
  assign n4364 = n4355 & n4363;
  assign n4365 = ~n292 & n1085;
  assign n4366 = ~n227 & ~n334;
  assign n4367 = n4365 & n4366;
  assign n4368 = ~n736 & n1305;
  assign n4369 = n1273 & n2983;
  assign n4370 = n4368 & n4369;
  assign n4371 = n4367 & n4370;
  assign n4372 = n4364 & n4371;
  assign n4373 = ~n310 & ~n901;
  assign n4374 = ~n126 & ~n497;
  assign n4375 = n1324 & n4374;
  assign n4376 = n4373 & n4375;
  assign n4377 = n3095 & n4376;
  assign n4378 = n907 & n4377;
  assign n4379 = n4372 & n4378;
  assign n3836 = ~n265 & n2625;
  assign n4381 = ~n312 & ~n412;
  assign n4382 = n4380 & n4381;
  assign n4383 = ~n207 & n883;
  assign n4384 = n4382 & n4383;
  assign n4385 = n3836 & n4384;
  assign n4387 = ~n122 & ~n304;
  assign n4388 = ~n74 & ~n659;
  assign n4389 = n4387 & n4388;
  assign n4390 = n4386 & n4389;
  assign n4391 = n4385 & n4390;
  assign n4392 = ~n133 & ~n330;
  assign n4393 = ~n406 & ~n478;
  assign n4394 = n4392 & n4393;
  assign n4395 = n3596 & n4394;
  assign n4396 = ~n87 & ~n128;
  assign n4397 = ~n104 & n4396;
  assign n4398 = n4395 & n4397;
  assign n4399 = n2946 & n4398;
  assign n4400 = n4391 & n4399;
  assign n4401 = ~n327 & n676;
  assign n4402 = n1240 & n1520;
  assign n4403 = n4401 & n4402;
  assign n4404 = n635 & n2813;
  assign n4405 = n4403 & n4404;
  assign n4406 = ~n1536 & n1931;
  assign n4407 = ~n410 & ~n449;
  assign n4408 = n4406 & n4407;
  assign n4409 = n4405 & n4408;
  assign n4077 = ~n79 & ~n463;
  assign n4078 = ~n199 & ~n553;
  assign n4079 = n4077 & n4078;
  assign n4080 = n1301 & n2842;
  assign n4081 = n4079 & n4080;
  assign n4082 = n982 & n4081;
  assign n4410 = n2578 & n3033;
  assign n4411 = ~n103 & n1075;
  assign n4412 = n4410 & n4411;
  assign n4413 = n4082 & n4412;
  assign n4414 = n4409 & n4413;
  assign n4415 = n4400 & n4414;
  assign n4416 = n4379 & n4415;
  assign n3685 = ~n300 & ~n592;
  assign n4417 = ~n228 & ~n237;
  assign n4418 = n3685 & n4417;
  assign n3813 = ~n552 & ~n850;
  assign n4419 = n1889 & n3813;
  assign n4420 = n4418 & n4419;
  assign n4421 = ~n83 & ~n152;
  assign n4422 = ~n155 & n4421;
  assign n4423 = n4420 & n4422;
  assign n4424 = ~n378 & ~n689;
  assign n4425 = n1286 & n4424;
  assign n4426 = n3330 & n4425;
  assign n4427 = n4423 & n4426;
  assign n4428 = n4416 & n4427;
  assign n4433 = ~n2424 & ~n2678;
  assign n4434 = n4433 ^ n2482;
  assign n4435 = n41 & ~n4434;
  assign n4296 = n54 & ~n2357;
  assign n4436 = n91 & ~n2423;
  assign n4437 = ~n4296 & ~n4436;
  assign n4438 = x31 & n4437;
  assign n4439 = ~n4435 & n4438;
  assign n4440 = n41 & ~n2482;
  assign n4441 = n54 & ~n2423;
  assign n4442 = ~n4440 & ~n4441;
  assign n4443 = ~x31 & n4442;
  assign n4444 = ~n4439 & ~n4443;
  assign n4309 = ~n2424 & ~n2482;
  assign n4310 = n2612 & ~n4309;
  assign n4307 = n2482 & ~n2678;
  assign n4308 = ~n2612 & ~n4307;
  assign n4450 = n4310 ^ n4308;
  assign n4451 = ~n2574 & n4450;
  assign n4452 = n4451 ^ n4308;
  assign n4453 = n4452 ^ n2669;
  assign n4454 = n44 & ~n4453;
  assign n4455 = ~n2574 & n3277;
  assign n3280 = n42 & ~n43;
  assign n4456 = ~n2669 & n3280;
  assign n4457 = ~n4455 & ~n4456;
  assign n4458 = ~n2612 & n3275;
  assign n4459 = n4457 & ~n4458;
  assign n4460 = ~n4454 & n4459;
  assign n4461 = n4460 ^ x29;
  assign n3667 = x31 & n41;
  assign n4292 = ~n2358 & ~n2373;
  assign n4293 = n4292 ^ n2423;
  assign n4294 = n3667 & ~n4293;
  assign n4295 = n41 & ~n2423;
  assign n4297 = ~n4295 & ~n4296;
  assign n4298 = ~x31 & ~n4297;
  assign n4299 = ~n2357 & n3672;
  assign n4300 = n54 & ~n2247;
  assign n4301 = x31 & n4300;
  assign n4302 = ~n4299 & ~n4301;
  assign n4303 = ~n4298 & n4302;
  assign n4304 = ~n4294 & n4303;
  assign n4252 = ~n2176 & ~n2371;
  assign n4253 = n4252 ^ n2247;
  assign n4254 = n41 & n4253;
  assign n4255 = n54 & n2065;
  assign n4256 = n91 & n2175;
  assign n4257 = ~n4255 & ~n4256;
  assign n4258 = x31 & n4257;
  assign n4259 = ~n4254 & n4258;
  assign n4260 = n54 & n2175;
  assign n3640 = ~x31 & ~n91;
  assign n4261 = ~n54 & n2247;
  assign n4262 = n3640 & ~n4261;
  assign n4263 = ~n4260 & n4262;
  assign n4264 = ~n4259 & ~n4263;
  assign n4109 = ~n347 & ~n503;
  assign n4110 = n3330 & n4109;
  assign n4111 = n3116 & n4110;
  assign n4112 = ~n293 & n2925;
  assign n4113 = n4111 & n4112;
  assign n4114 = n1932 & n4113;
  assign n4115 = ~n610 & ~n634;
  assign n4116 = n1460 & n4115;
  assign n4117 = n3163 & n4116;
  assign n4118 = ~n83 & ~n567;
  assign n4119 = ~n120 & ~n358;
  assign n4120 = n4118 & n4119;
  assign n4121 = n4117 & n4120;
  assign n4122 = n4114 & n4121;
  assign n3904 = ~n265 & ~n517;
  assign n3905 = ~n497 & n3904;
  assign n4123 = ~n277 & ~n343;
  assign n4124 = ~n283 & ~n541;
  assign n4125 = n4123 & n4124;
  assign n4126 = ~n163 & ~n666;
  assign n4127 = n1168 & n4126;
  assign n4128 = n4125 & n4127;
  assign n4129 = n3905 & n4128;
  assign n4130 = ~n418 & ~n787;
  assign n4131 = n2318 & n4130;
  assign n4132 = n3246 & n4131;
  assign n4133 = n653 & n4132;
  assign n4134 = n4129 & n4133;
  assign n4135 = n4122 & n4134;
  assign n4136 = n792 & n1263;
  assign n4137 = ~n300 & ~n640;
  assign n4138 = ~n69 & ~n683;
  assign n4139 = n4137 & n4138;
  assign n4140 = n4136 & n4139;
  assign n4072 = ~n296 & ~n1166;
  assign n4142 = n4072 & n4141;
  assign n4143 = n2180 & n2806;
  assign n4144 = n4142 & n4143;
  assign n4145 = n4140 & n4144;
  assign n4146 = ~n183 & ~n361;
  assign n4147 = n3089 & n4146;
  assign n4148 = ~n57 & n771;
  assign n4149 = n4147 & n4148;
  assign n4150 = n1990 & n4149;
  assign n4151 = n4145 & n4150;
  assign n3726 = ~n227 & ~n476;
  assign n4161 = n1199 & n1485;
  assign n4162 = n3726 & n4161;
  assign n4163 = ~n244 & n3146;
  assign n4164 = n4162 & n4163;
  assign n4165 = n4160 & n4164;
  assign n4166 = n4151 & n4165;
  assign n3935 = ~n134 & ~n396;
  assign n4167 = n3935 & n4077;
  assign n4168 = n483 & n1314;
  assign n4169 = n4167 & n4168;
  assign n3471 = ~n87 & ~n540;
  assign n3576 = ~n344 & ~n552;
  assign n4170 = n3471 & n3576;
  assign n4171 = n1288 & n1977;
  assign n4172 = n4170 & n4171;
  assign n4173 = n4169 & n4172;
  assign n3606 = ~n392 & ~n616;
  assign n4176 = ~n424 & ~n506;
  assign n4177 = n3606 & n4176;
  assign n4178 = n4175 & n4177;
  assign n4179 = n4173 & n4178;
  assign n4180 = ~n237 & ~n929;
  assign n4181 = ~n758 & n4180;
  assign n4182 = ~n280 & ~n378;
  assign n4183 = n144 & n4182;
  assign n4184 = n4181 & n4183;
  assign n4185 = n2417 & n4184;
  assign n4186 = n4179 & n4185;
  assign n4187 = n4166 & n4186;
  assign n4188 = n4135 & n4187;
  assign n4189 = n4188 ^ x8;
  assign n3707 = ~n256 & ~n514;
  assign n3708 = n2267 & n3707;
  assign n3709 = n1225 & n3708;
  assign n3710 = ~n245 & n1787;
  assign n3711 = n3709 & n3710;
  assign n3713 = ~n331 & ~n382;
  assign n3714 = n3712 & n3713;
  assign n3715 = n532 & n2310;
  assign n3716 = n3714 & n3715;
  assign n3717 = n2728 & n3716;
  assign n3718 = n3711 & n3717;
  assign n3719 = ~n593 & ~n610;
  assign n3720 = ~n217 & n3719;
  assign n3721 = ~n456 & ~n1005;
  assign n3722 = n3720 & n3721;
  assign n3723 = n2683 & n3722;
  assign n3724 = ~n405 & n1631;
  assign n3725 = n2271 & n3724;
  assign n3727 = n1594 & n3726;
  assign n3728 = n3725 & n3727;
  assign n3729 = n3723 & n3728;
  assign n3730 = n3718 & n3729;
  assign n4190 = ~n126 & n3365;
  assign n4191 = n1302 & n3020;
  assign n4192 = n4141 & n4191;
  assign n4193 = n4190 & n4192;
  assign n4194 = ~n406 & n2787;
  assign n4195 = n4193 & n4194;
  assign n4196 = ~n151 & ~n525;
  assign n4197 = ~n216 & n4196;
  assign n4199 = n2461 & n4198;
  assign n4200 = n4197 & n4199;
  assign n4201 = n2182 & n2569;
  assign n4202 = n3121 & n4201;
  assign n4203 = n4200 & n4202;
  assign n4204 = n4195 & n4203;
  assign n4205 = ~n133 & ~n412;
  assign n4206 = ~n812 & n4205;
  assign n4207 = ~n87 & ~n710;
  assign n4208 = ~n202 & ~n617;
  assign n4209 = n4207 & n4208;
  assign n4210 = n4206 & n4209;
  assign n4211 = n2468 & n4210;
  assign n3699 = n472 & ~n790;
  assign n3700 = ~n1065 & n3699;
  assign n4212 = ~n226 & ~n322;
  assign n4213 = n255 & n4212;
  assign n4214 = n2949 & n4213;
  assign n4215 = n3700 & n4214;
  assign n4216 = n4211 & n4215;
  assign n4217 = n4204 & n4216;
  assign n4218 = n3730 & n4217;
  assign n4219 = n786 & n2925;
  assign n4220 = n2227 & n4219;
  assign n4221 = n1332 & n1554;
  assign n4222 = ~n630 & n4221;
  assign n4223 = n4220 & n4222;
  assign n4224 = n3230 & n4223;
  assign n4225 = ~n304 & n1238;
  assign n4226 = ~n281 & n297;
  assign n4227 = n4225 & n4226;
  assign n4228 = n3912 & n4227;
  assign n4229 = n4224 & n4228;
  assign n4230 = ~n249 & ~n327;
  assign n4231 = n602 & n4230;
  assign n4233 = n4231 & n4232;
  assign n4234 = n1263 & n4233;
  assign n4235 = ~n233 & n925;
  assign n4236 = n4234 & n4235;
  assign n4237 = ~n497 & ~n1060;
  assign n4238 = ~n164 & ~n292;
  assign n4239 = n4237 & n4238;
  assign n4240 = ~n743 & n875;
  assign n4241 = n4239 & n4240;
  assign n4242 = ~n141 & ~n333;
  assign n4243 = ~n652 & n4242;
  assign n4244 = n3262 & n4243;
  assign n4245 = n4241 & n4244;
  assign n4246 = n4236 & n4245;
  assign n4247 = n4229 & n4246;
  assign n4248 = n4218 & n4247;
  assign n4249 = n4248 ^ n4188;
  assign n4250 = n4189 & ~n4249;
  assign n4251 = n4250 ^ x8;
  assign n4265 = n4264 ^ n4251;
  assign n4064 = n782 & ~n1405;
  assign n4066 = ~n104 & ~n234;
  assign n4067 = n4065 & n4066;
  assign n4068 = n4064 & n4067;
  assign n4069 = ~n370 & n2314;
  assign n4070 = n4068 & n4069;
  assign n4071 = ~n270 & ~n841;
  assign n4073 = n4071 & n4072;
  assign n4074 = n1019 & n3146;
  assign n4075 = n4073 & n4074;
  assign n4076 = n4070 & n4075;
  assign n4083 = n2184 & n4082;
  assign n4084 = n4076 & n4083;
  assign n4035 = n1273 & n2805;
  assign n4036 = n526 & n1001;
  assign n4037 = n4035 & n4036;
  assign n4038 = ~n630 & ~n634;
  assign n4039 = n3290 & n4038;
  assign n4040 = ~n390 & ~n740;
  assign n4041 = n2134 & n4040;
  assign n4042 = ~n209 & ~n249;
  assign n4043 = ~n170 & ~n304;
  assign n4044 = n4042 & n4043;
  assign n4045 = n4041 & n4044;
  assign n4046 = n4039 & n4045;
  assign n4047 = n4037 & n4046;
  assign n4085 = ~n278 & n860;
  assign n4086 = n81 & n215;
  assign n4087 = ~n439 & ~n4086;
  assign n4088 = n4085 & n4087;
  assign n3577 = ~n492 & n3576;
  assign n4089 = ~n245 & ~n265;
  assign n4090 = n1964 & n4089;
  assign n4091 = n3577 & n4090;
  assign n4092 = n4088 & n4091;
  assign n4093 = ~n531 & ~n975;
  assign n4094 = n935 & n4093;
  assign n4095 = ~n95 & ~n314;
  assign n4096 = n1295 & n4095;
  assign n4097 = n4094 & n4096;
  assign n4099 = n1918 & n4098;
  assign n4101 = n1670 & n4100;
  assign n4102 = n4099 & n4101;
  assign n4103 = n4097 & n4102;
  assign n4104 = n4092 & n4103;
  assign n4105 = n4047 & n4104;
  assign n4106 = n4084 & n4105;
  assign n4107 = n3018 & n4106;
  assign n4266 = n4251 ^ n4107;
  assign n3805 = ~n283 & n2130;
  assign n3806 = ~n418 & ~n582;
  assign n3807 = n3805 & n3806;
  assign n3808 = ~n343 & ~n405;
  assign n3809 = n297 & n3808;
  assign n3810 = n3807 & n3809;
  assign n4267 = n892 & n2067;
  assign n4268 = n860 & n934;
  assign n4269 = n4267 & n4268;
  assign n4270 = ~n558 & n2310;
  assign n4271 = ~n238 & n4270;
  assign n4272 = n4269 & n4271;
  assign n4273 = ~n174 & ~n412;
  assign n4274 = ~n292 & ~n331;
  assign n4275 = n4273 & n4274;
  assign n4276 = n1072 & n4275;
  assign n4277 = ~n95 & ~n634;
  assign n4278 = n1847 & n4277;
  assign n4279 = n4276 & n4278;
  assign n4280 = n4272 & n4279;
  assign n4281 = n1728 & n1755;
  assign n4282 = ~n443 & n1444;
  assign n4283 = n4281 & n4282;
  assign n4284 = n4280 & n4283;
  assign n4285 = n3810 & n4284;
  assign n4286 = n2206 & n2700;
  assign n4287 = n4285 & n4286;
  assign n4288 = n4287 ^ n4107;
  assign n4289 = ~n4266 & ~n4288;
  assign n4290 = ~n4265 & n4289;
  assign n4291 = n4290 ^ n4107;
  assign n4305 = n4304 ^ n4291;
  assign n3788 = n130 & n1140;
  assign n3789 = ~n333 & ~n370;
  assign n3790 = ~n244 & n3789;
  assign n3791 = n2799 & n3790;
  assign n3792 = n3788 & n3791;
  assign n3738 = ~n280 & ~n347;
  assign n3793 = n355 & n1210;
  assign n3794 = n3738 & n3793;
  assign n3795 = n2929 & n3794;
  assign n3796 = n3792 & n3795;
  assign n3446 = ~n133 & ~n452;
  assign n3447 = ~n155 & ~n616;
  assign n3448 = n3446 & n3447;
  assign n3449 = ~n826 & n3448;
  assign n3451 = n2787 & n3450;
  assign n3452 = n3449 & n3451;
  assign n3454 = ~n310 & n2307;
  assign n3455 = n3453 & n3454;
  assign n3456 = n3452 & n3455;
  assign n3925 = ~n544 & n1017;
  assign n4002 = n1624 & n3925;
  assign n4003 = ~n183 & n1739;
  assign n4004 = n1142 & n4003;
  assign n4005 = n4002 & n4004;
  assign n4006 = n3456 & n4005;
  assign n4007 = n3796 & n4006;
  assign n4008 = ~n64 & ~n640;
  assign n4009 = ~n217 & ~n314;
  assign n4010 = n4008 & n4009;
  assign n4011 = ~n173 & ~n270;
  assign n4012 = n583 & n4011;
  assign n4013 = n4010 & n4012;
  assign n4015 = n144 & ~n320;
  assign n4016 = n4014 & n4015;
  assign n4017 = n4013 & n4016;
  assign n4018 = n852 & ~n3200;
  assign n4020 = ~n361 & ~n948;
  assign n4021 = n4019 & n4020;
  assign n4022 = n4018 & n4021;
  assign n4023 = n4017 & n4022;
  assign n4024 = ~n323 & ~n478;
  assign n4025 = n1920 & n4024;
  assign n4026 = ~n234 & ~n666;
  assign n4027 = ~n392 & ~n463;
  assign n4028 = n4026 & n4027;
  assign n4029 = n4025 & n4028;
  assign n4030 = n926 & n2856;
  assign n4031 = n4029 & n4030;
  assign n4032 = n2844 & n4031;
  assign n4033 = n4023 & n4032;
  assign n4034 = n4007 & n4033;
  assign n4049 = n1546 & n4048;
  assign n4050 = ~n1005 & n2073;
  assign n4051 = n4049 & n4050;
  assign n4052 = n294 & n530;
  assign n4053 = n4051 & n4052;
  assign n4058 = ~n461 & ~n660;
  assign n4059 = n4057 & n4058;
  assign n4060 = n4053 & n4059;
  assign n4061 = n4047 & n4060;
  assign n4062 = n4034 & n4061;
  assign n4063 = n4062 ^ x11;
  assign n4108 = n4107 ^ n4063;
  assign n4447 = n4304 ^ n4108;
  assign n4448 = ~n4305 & ~n4447;
  assign n4449 = n4448 ^ n4291;
  assign n4462 = n4461 ^ n4449;
  assign n4429 = n4107 ^ x11;
  assign n4430 = n4107 ^ n4062;
  assign n4431 = n4429 & ~n4430;
  assign n4432 = n4431 ^ x11;
  assign n4827 = n4449 ^ n4432;
  assign n4828 = ~n4462 & n4827;
  assign n4829 = n4828 ^ n4461;
  assign n4830 = ~n4444 & n4829;
  assign n4831 = ~n4449 & n4461;
  assign n4832 = n4432 & n4831;
  assign n4833 = ~n4830 & ~n4832;
  assign n4802 = ~n91 & n2423;
  assign n4803 = ~n4440 & ~n4802;
  assign n4804 = n2425 & n4803;
  assign n4805 = n2612 & ~n4804;
  assign n4806 = ~n54 & n2482;
  assign n4807 = ~n4295 & ~n4806;
  assign n4808 = ~n2425 & n4807;
  assign n4809 = n4805 & ~n4808;
  assign n4810 = ~n2612 & n4806;
  assign n4811 = n2678 & n4810;
  assign n4812 = n91 & n2482;
  assign n4813 = x31 & ~n4812;
  assign n4814 = ~n4811 & n4813;
  assign n4815 = ~n4809 & n4814;
  assign n4816 = ~n2482 & ~n2612;
  assign n4817 = ~n2425 & n4816;
  assign n4818 = ~n54 & ~n4817;
  assign n4819 = n4802 & ~n4818;
  assign n4820 = n4815 & ~n4819;
  assign n4821 = n54 & n2482;
  assign n4822 = n3640 & ~n4821;
  assign n4823 = ~n54 & n2612;
  assign n4824 = n4822 & ~n4823;
  assign n4825 = ~n4820 & ~n4824;
  assign n4723 = ~n605 & n844;
  assign n4724 = ~n535 & n4566;
  assign n4725 = n4723 & n4724;
  assign n4726 = n1756 & n4725;
  assign n4727 = ~n319 & n1445;
  assign n4728 = n3240 & n4232;
  assign n4729 = n4727 & n4728;
  assign n4730 = n4726 & n4729;
  assign n4740 = n2055 & n4739;
  assign n4741 = ~n405 & ~n592;
  assign n4742 = ~n527 & n4741;
  assign n4743 = n4740 & n4742;
  assign n3482 = n105 & n542;
  assign n4744 = ~n331 & n1171;
  assign n4745 = n3482 & n4744;
  assign n4746 = n4743 & n4745;
  assign n4747 = n4738 & n4746;
  assign n4748 = n4730 & n4747;
  assign n4749 = ~n278 & n4748;
  assign n4750 = ~n382 & ~n1227;
  assign n4751 = n4146 & n4750;
  assign n4752 = n597 & n1771;
  assign n4753 = n4751 & n4752;
  assign n4754 = n162 & n4753;
  assign n4755 = ~n51 & ~n93;
  assign n4756 = ~n497 & n4755;
  assign n4757 = n994 & n4756;
  assign n4758 = n4754 & n4757;
  assign n4759 = ~n396 & ~n567;
  assign n4760 = ~n304 & ~n412;
  assign n4761 = n4759 & n4760;
  assign n4762 = n1197 & n2634;
  assign n4763 = n4761 & n4762;
  assign n4764 = n1492 & n3738;
  assign n4765 = ~n269 & ~n617;
  assign n4766 = n1810 & n4765;
  assign n4767 = n4764 & n4766;
  assign n4768 = n4763 & n4767;
  assign n4769 = n4758 & n4768;
  assign n4770 = n1360 & n2753;
  assign n4771 = n1575 & n4770;
  assign n4772 = ~n295 & ~n675;
  assign n4773 = ~n406 & n4772;
  assign n4774 = ~n351 & ~n656;
  assign n4775 = n4773 & n4774;
  assign n4776 = n4771 & n4775;
  assign n4777 = ~n253 & ~n402;
  assign n4778 = ~n170 & ~n222;
  assign n4779 = n4777 & n4778;
  assign n4780 = n420 & n4779;
  assign n4781 = n4776 & n4780;
  assign n4782 = n533 & n2232;
  assign n4783 = ~n167 & n1665;
  assign n4784 = n4782 & n4783;
  assign n4785 = ~n710 & ~n1060;
  assign n4786 = n964 & n4785;
  assign n4787 = n1785 & n4786;
  assign n4789 = n4787 & n4788;
  assign n4790 = n4784 & n4789;
  assign n4791 = n4781 & n4790;
  assign n4792 = n4769 & n4791;
  assign n4793 = n4749 & n4792;
  assign n4794 = ~n323 & ~n390;
  assign n4795 = ~n79 & ~n300;
  assign n4796 = n4794 & n4795;
  assign n4797 = ~n476 & ~n948;
  assign n4798 = n1026 & n4797;
  assign n4799 = n4796 & n4798;
  assign n4800 = n1828 & n4799;
  assign n4801 = n4793 & n4800;
  assign n4826 = n4825 ^ n4801;
  assign n4834 = n4449 & ~n4461;
  assign n4835 = ~n4432 & n4834;
  assign n4836 = n4444 & n4835;
  assign n4945 = ~n4826 & ~n4836;
  assign n4946 = n4833 & ~n4945;
  assign n4947 = ~n4428 & ~n4946;
  assign n4948 = n4428 & n4826;
  assign n4949 = ~n4832 & ~n4948;
  assign n4950 = ~n4444 & ~n4949;
  assign n4951 = ~n4835 & n4950;
  assign n4952 = n4829 & n4948;
  assign n4953 = ~n4951 & ~n4952;
  assign n4954 = ~n4947 & n4953;
  assign n3657 = ~n2669 & ~n2680;
  assign n3658 = n2786 & ~n3657;
  assign n3660 = n2669 & n2680;
  assign n3661 = ~n2786 & ~n3660;
  assign n4494 = ~n3658 & ~n3661;
  assign n4495 = n4494 ^ n2718;
  assign n4936 = n44 & ~n4495;
  assign n4937 = ~n2718 & n3280;
  assign n4938 = ~n2669 & n3275;
  assign n4939 = ~n2786 & n3277;
  assign n4940 = ~n4938 & ~n4939;
  assign n4941 = ~n4937 & n4940;
  assign n4942 = ~n4936 & n4941;
  assign n4943 = n4942 ^ x29;
  assign n4311 = ~n4308 & ~n4310;
  assign n4312 = n4311 ^ n2574;
  assign n4924 = n41 & n4312;
  assign n4925 = x31 & ~n4821;
  assign n4926 = n91 & n2612;
  assign n4927 = n4925 & ~n4926;
  assign n4928 = ~n4924 & n4927;
  assign n4929 = ~n54 & n2574;
  assign n4930 = n3640 & ~n4929;
  assign n4931 = n54 & n2612;
  assign n4932 = n4930 & ~n4931;
  assign n4933 = ~n4928 & ~n4932;
  assign n4567 = n4565 & n4566;
  assign n4568 = n570 & n4567;
  assign n4569 = ~n303 & ~n320;
  assign n4570 = n2780 & n4569;
  assign n4571 = ~n361 & ~n617;
  assign n4572 = n2249 & n4571;
  assign n4573 = n4570 & n4572;
  assign n4574 = n4568 & n4573;
  assign n4575 = n1641 & n4574;
  assign n4576 = ~n226 & ~n296;
  assign n4577 = n1530 & n4576;
  assign n4578 = ~n262 & ~n612;
  assign n4579 = ~n334 & n4578;
  assign n4580 = n4577 & n4579;
  assign n4581 = n543 & n4580;
  assign n4582 = n2813 & n2943;
  assign n4583 = n2665 & n3122;
  assign n4584 = n4582 & n4583;
  assign n4585 = n4581 & n4584;
  assign n4586 = n3188 & n4585;
  assign n4587 = n4575 & n4586;
  assign n4887 = ~n647 & ~n709;
  assign n4888 = ~n354 & ~n750;
  assign n4889 = n4887 & n4888;
  assign n4890 = n464 & n4889;
  assign n4891 = n624 & n4890;
  assign n4892 = n4207 & n4242;
  assign n4893 = n860 & n2654;
  assign n4894 = n4892 & n4893;
  assign n4895 = n2788 & n4894;
  assign n4896 = n4891 & n4895;
  assign n4897 = n663 & n3723;
  assign n4898 = n4896 & n4897;
  assign n4899 = ~n312 & ~n358;
  assign n4900 = n376 & n4899;
  assign n4901 = n3155 & n4900;
  assign n4902 = ~n627 & n1091;
  assign n4903 = n2433 & n4902;
  assign n4904 = n4901 & n4903;
  assign n3521 = ~n277 & n2649;
  assign n4905 = n235 & n1548;
  assign n4906 = ~n249 & ~n410;
  assign n4907 = n1101 & n4906;
  assign n4908 = n4905 & n4907;
  assign n4909 = n3521 & n4908;
  assign n4910 = n4904 & n4909;
  assign n4911 = n4178 & n4910;
  assign n3609 = ~n163 & ~n337;
  assign n4912 = ~n250 & ~n272;
  assign n4913 = n3609 & n4912;
  assign n4914 = n719 & n4913;
  assign n4915 = n2490 & n4914;
  assign n4916 = ~n634 & ~n799;
  assign n4917 = n2344 & n4916;
  assign n4918 = n1976 & n4917;
  assign n4919 = n4915 & n4918;
  assign n4920 = n4911 & n4919;
  assign n4921 = n4898 & n4920;
  assign n4922 = n4587 & n4921;
  assign n4923 = n4922 ^ x14;
  assign n4934 = n4933 ^ n4923;
  assign n4885 = n4825 ^ n4428;
  assign n4886 = ~n4826 & ~n4885;
  assign n4935 = n4934 ^ n4886;
  assign n4944 = n4943 ^ n4935;
  assign n4955 = n4954 ^ n4944;
  assign n3285 = n643 & n735;
  assign n3748 = n2871 ^ n566;
  assign n3749 = n3748 ^ n368;
  assign n4877 = n3285 & n3749;
  assign n3434 = ~n817 & ~n1467;
  assign n3435 = ~n3300 & n3434;
  assign n4878 = ~n566 & n3435;
  assign n3437 = ~n643 & n735;
  assign n4879 = ~n368 & n3437;
  assign n4880 = ~n4878 & ~n4879;
  assign n3440 = ~n63 & ~n119;
  assign n4881 = ~n2861 & ~n3440;
  assign n4882 = n4880 & ~n4881;
  assign n4883 = ~n4877 & n4882;
  assign n4884 = n4883 ^ x26;
  assign n4956 = n4955 ^ n4884;
  assign n3662 = n2718 & ~n3661;
  assign n3659 = ~n2718 & ~n3658;
  assign n3663 = n3662 ^ n3659;
  assign n3664 = n2861 & n3663;
  assign n3665 = n3664 ^ n3662;
  assign n3666 = n3665 ^ n566;
  assign n4714 = n3285 & ~n3666;
  assign n4715 = ~n566 & n3437;
  assign n4716 = ~n2861 & n3435;
  assign n4717 = ~n4715 & ~n4716;
  assign n4718 = ~n2718 & ~n3440;
  assign n4719 = n4717 & ~n4718;
  assign n4720 = ~n4714 & n4719;
  assign n4721 = n4720 ^ x26;
  assign n4652 = n2680 ^ n2669;
  assign n4653 = n4652 ^ n2786;
  assign n4706 = n44 & ~n4653;
  assign n4707 = ~n2574 & n3275;
  assign n4708 = ~n2669 & n3277;
  assign n4709 = ~n2786 & n3280;
  assign n4710 = ~n4708 & ~n4709;
  assign n4711 = ~n4707 & n4710;
  assign n4712 = ~n4706 & n4711;
  assign n4713 = n4712 ^ x29;
  assign n4722 = n4721 ^ n4713;
  assign n4837 = ~n4428 & ~n4836;
  assign n4838 = n4833 & n4837;
  assign n4445 = n4444 ^ n4432;
  assign n4839 = ~n4445 & ~n4834;
  assign n4840 = n4428 & ~n4839;
  assign n4841 = n4831 ^ n4432;
  assign n4842 = ~n4831 & n4841;
  assign n4843 = n4444 & n4842;
  assign n4844 = n4843 ^ n4841;
  assign n4845 = n4840 & ~n4844;
  assign n4846 = ~n4838 & ~n4845;
  assign n4847 = n4846 ^ n4826;
  assign n4874 = n4847 ^ n4721;
  assign n4875 = ~n4722 & n4874;
  assign n4876 = n4875 ^ n4847;
  assign n4957 = n4956 ^ n4876;
  assign n3775 = ~n2873 & ~n3037;
  assign n3630 = ~n368 & ~n2956;
  assign n3774 = n3037 & ~n3630;
  assign n3971 = n3775 ^ n3774;
  assign n3972 = n2954 & n3971;
  assign n3973 = n3972 ^ n3774;
  assign n3974 = n3973 ^ n3098;
  assign n4476 = x21 ^ x20;
  assign n4477 = x23 ^ x22;
  assign n4478 = n4476 & n4477;
  assign n4865 = ~n3974 & n4478;
  assign n4487 = n4476 & ~n4477;
  assign n4866 = ~n3098 & n4487;
  assign n36 = x20 & x21;
  assign n34 = ~x20 & ~x21;
  assign n4482 = n36 ^ n34;
  assign n4483 = x22 & n4482;
  assign n4484 = n4483 ^ n36;
  assign n4867 = ~n2954 & n4484;
  assign n4868 = ~n4866 & ~n4867;
  assign n35 = ~x22 & n34;
  assign n37 = x22 & n36;
  assign n38 = ~n35 & ~n37;
  assign n4480 = ~n38 & n4477;
  assign n4869 = ~n3037 & n4480;
  assign n4870 = n4868 & ~n4869;
  assign n4871 = ~n4865 & n4870;
  assign n4872 = n4871 ^ x23;
  assign n3776 = ~n3774 & ~n3775;
  assign n3777 = n3776 ^ n2954;
  assign n4697 = ~n3777 & n4478;
  assign n4698 = ~n368 & n4480;
  assign n4699 = ~n3037 & n4484;
  assign n4700 = ~n4698 & ~n4699;
  assign n4701 = ~n2954 & n4487;
  assign n4702 = n4700 & ~n4701;
  assign n4703 = ~n4697 & n4702;
  assign n4704 = n4703 ^ x23;
  assign n4446 = n4445 ^ n4428;
  assign n4463 = n4462 ^ n4446;
  assign n4313 = n44 & ~n4312;
  assign n4314 = ~n2612 & n3277;
  assign n4315 = ~n2482 & n3275;
  assign n4316 = ~n4314 & ~n4315;
  assign n4317 = ~n2574 & n3280;
  assign n4318 = n4316 & ~n4317;
  assign n4319 = ~n4313 & n4318;
  assign n4320 = n4319 ^ x29;
  assign n4306 = n4305 ^ n4108;
  assign n4321 = n4320 ^ n4306;
  assign n4333 = ~n4307 & ~n4309;
  assign n4334 = n4333 ^ n2612;
  assign n4335 = n44 & ~n4334;
  assign n4336 = ~n2482 & n3277;
  assign n4337 = ~n2423 & n3275;
  assign n4338 = ~n4336 & ~n4337;
  assign n4339 = ~n2612 & n3280;
  assign n4340 = n4338 & ~n4339;
  assign n4341 = ~n4335 & n4340;
  assign n4342 = n4341 ^ x29;
  assign n4322 = ~n2248 & ~n2372;
  assign n4323 = n4322 ^ n2357;
  assign n4324 = n41 & n4323;
  assign n4325 = n91 & n2247;
  assign n4326 = x31 & ~n4325;
  assign n4327 = ~n4260 & n4326;
  assign n4328 = ~n4324 & n4327;
  assign n4329 = ~x31 & n4300;
  assign n4330 = ~n2357 & n3676;
  assign n4331 = ~n4329 & ~n4330;
  assign n4332 = ~n4328 & n4331;
  assign n4343 = n4342 ^ n4332;
  assign n4344 = ~n4265 & ~n4266;
  assign n4345 = n4344 ^ n4287;
  assign n4346 = n4345 ^ n4332;
  assign n4347 = n4343 & ~n4346;
  assign n4348 = n4347 ^ n4342;
  assign n4349 = n4348 ^ n4320;
  assign n4350 = n4321 & n4349;
  assign n4351 = n4350 ^ n4348;
  assign n4464 = n4463 ^ n4351;
  assign n4465 = ~n3659 & ~n3662;
  assign n4466 = n4465 ^ n2861;
  assign n4467 = n3285 & ~n4466;
  assign n4468 = ~n2718 & n3435;
  assign n4469 = ~n2861 & n3437;
  assign n4470 = ~n2786 & ~n3440;
  assign n4471 = ~n4469 & ~n4470;
  assign n4472 = ~n4468 & n4471;
  assign n4473 = ~n4467 & n4472;
  assign n4474 = n4473 ^ x26;
  assign n4694 = n4474 ^ n4463;
  assign n4695 = n4464 & ~n4694;
  assign n4696 = n4695 ^ n4474;
  assign n4705 = n4704 ^ n4696;
  assign n4848 = n4847 ^ n4722;
  assign n4862 = n4848 ^ n4704;
  assign n4863 = ~n4705 & n4862;
  assign n4864 = n4863 ^ n4848;
  assign n4873 = n4872 ^ n4864;
  assign n4958 = n4957 ^ n4873;
  assign n4671 = x18 ^ x17;
  assign n4672 = x20 ^ x19;
  assign n4673 = n4671 & n4672;
  assign n4853 = ~n3989 & n4673;
  assign n4678 = x17 & x18;
  assign n4675 = ~x17 & ~x18;
  assign n4683 = n4678 ^ n4675;
  assign n4684 = x19 & n4683;
  assign n4685 = n4684 ^ n4678;
  assign n4854 = ~n3270 & n4685;
  assign n4676 = ~x19 & n4675;
  assign n4677 = x20 & n4676;
  assign n4679 = x19 & ~x20;
  assign n4680 = n4678 & n4679;
  assign n4681 = ~n4677 & ~n4680;
  assign n4855 = ~n3196 & ~n4681;
  assign n4688 = n4671 & ~n4672;
  assign n4856 = ~n3351 & n4688;
  assign n4857 = ~n4855 & ~n4856;
  assign n4858 = ~n4854 & n4857;
  assign n4859 = ~n4853 & n4858;
  assign n4860 = n4859 ^ x20;
  assign n3107 = n3106 ^ n3098;
  assign n3197 = n3196 ^ n3106;
  assign n3198 = n3107 & ~n3197;
  assign n3271 = n3270 ^ n3198;
  assign n4674 = ~n3271 & n4673;
  assign n4682 = ~n3098 & ~n4681;
  assign n4686 = ~n3196 & n4685;
  assign n4687 = ~n4682 & ~n4686;
  assign n4689 = ~n3270 & n4688;
  assign n4690 = n4687 & ~n4689;
  assign n4691 = ~n4674 & n4690;
  assign n4692 = n4691 ^ x20;
  assign n3631 = ~n2873 & ~n3630;
  assign n3632 = n3631 ^ n3037;
  assign n4479 = ~n3632 & n4478;
  assign n4481 = ~n566 & n4480;
  assign n4485 = ~n368 & n4484;
  assign n4486 = ~n4481 & ~n4485;
  assign n4488 = ~n3037 & n4487;
  assign n4489 = n4486 & ~n4488;
  assign n4490 = ~n4479 & n4489;
  assign n4491 = n4490 ^ x23;
  assign n4475 = n4474 ^ n4464;
  assign n4492 = n4491 ^ n4475;
  assign n4496 = n3285 & ~n4495;
  assign n4497 = ~n2718 & n3437;
  assign n4498 = ~n2669 & ~n3440;
  assign n4499 = ~n2786 & n3435;
  assign n4500 = ~n4498 & ~n4499;
  assign n4501 = ~n4497 & n4500;
  assign n4502 = ~n4496 & n4501;
  assign n4503 = n4502 ^ x26;
  assign n4493 = n4348 ^ n4321;
  assign n4504 = n4503 ^ n4493;
  assign n4650 = n4345 ^ n4343;
  assign n4637 = n4266 ^ n4264;
  assign n4506 = ~n2066 & ~n2370;
  assign n4507 = n4506 ^ n2175;
  assign n4508 = n3667 & ~n4507;
  assign n4509 = n3640 & ~n4255;
  assign n4510 = ~n54 & n2175;
  assign n4511 = n4509 & ~n4510;
  assign n4512 = ~n2065 & n3672;
  assign n4513 = ~n1974 & n3669;
  assign n4514 = ~n4512 & ~n4513;
  assign n4515 = ~n4511 & n4514;
  assign n4516 = ~n4508 & n4515;
  assign n4505 = n4248 ^ n4189;
  assign n4517 = n4516 ^ n4505;
  assign n4592 = ~n1879 & ~n2368;
  assign n4593 = x31 & n4592;
  assign n4594 = n4593 ^ n1974;
  assign n4595 = n41 & ~n4594;
  assign n4596 = ~n1798 & n3669;
  assign n4597 = ~n1878 & ~n3673;
  assign n4598 = ~n4596 & ~n4597;
  assign n4599 = ~n4595 & n4598;
  assign n4518 = x5 ^ x2;
  assign n4544 = ~n790 & ~n799;
  assign n4545 = n1368 & n4544;
  assign n4546 = n1422 & n1906;
  assign n4547 = n4545 & n4546;
  assign n4548 = ~n277 & n4547;
  assign n4549 = ~n253 & ~n787;
  assign n4550 = ~n166 & n4549;
  assign n4551 = n2789 & n4550;
  assign n4553 = n2526 & n4552;
  assign n4554 = ~n173 & ~n256;
  assign n4556 = n4554 & n4555;
  assign n4557 = n4553 & n4556;
  assign n4558 = n4551 & n4557;
  assign n4559 = n1226 & n2992;
  assign n4560 = n4558 & n4559;
  assign n4561 = n4548 & n4560;
  assign n4562 = ~n791 & n2967;
  assign n4563 = n4561 & n4562;
  assign n4564 = n4543 & n4563;
  assign n4588 = n4564 & n4587;
  assign n4589 = n4588 ^ x5;
  assign n4590 = n4518 & ~n4589;
  assign n4591 = n4590 ^ x2;
  assign n4600 = n4599 ^ n4591;
  assign n4601 = n4591 ^ n4188;
  assign n3537 = n2382 & ~n2506;
  assign n3538 = n462 & ~n1135;
  assign n3539 = n3537 & n3538;
  assign n3540 = n685 & n2965;
  assign n3541 = n3539 & n3540;
  assign n3542 = ~n74 & n1787;
  assign n3543 = ~n193 & ~n333;
  assign n3544 = n584 & n3543;
  assign n3545 = n3542 & n3544;
  assign n3546 = n3541 & n3545;
  assign n3547 = ~n127 & ~n358;
  assign n3548 = ~n337 & n3547;
  assign n3549 = n450 & n1944;
  assign n3550 = n3548 & n3549;
  assign n3551 = n239 & n321;
  assign n3552 = ~n293 & ~n385;
  assign n3554 = n3552 & n3553;
  assign n3555 = n3551 & n3554;
  assign n3556 = n3550 & n3555;
  assign n3557 = n2342 & n3556;
  assign n3558 = n3546 & n3557;
  assign n4602 = ~n110 & ~n723;
  assign n4603 = n1153 & n4602;
  assign n4604 = ~n143 & n3330;
  assign n4605 = n4603 & n4604;
  assign n4606 = n420 & n4605;
  assign n3458 = ~n181 & ~n350;
  assign n4607 = n1569 & n3458;
  assign n4608 = n4238 & n4607;
  assign n4609 = n2800 & n4608;
  assign n4610 = n4606 & n4609;
  assign n4611 = n4164 & n4234;
  assign n4612 = n4610 & n4611;
  assign n3560 = ~n95 & ~n1047;
  assign n4613 = ~n362 & ~n946;
  assign n4614 = n3560 & n4613;
  assign n4615 = ~n424 & ~n627;
  assign n4616 = ~n656 & n4615;
  assign n4617 = n4614 & n4616;
  assign n4618 = n834 & n2227;
  assign n4619 = n3058 & n4618;
  assign n4620 = n4617 & n4619;
  assign n4621 = n453 & n2051;
  assign n4622 = n2477 & n4621;
  assign n4623 = n1324 & n3183;
  assign n4624 = n4237 & n4623;
  assign n4625 = n4622 & n4624;
  assign n4626 = n4620 & n4625;
  assign n4627 = n1028 & n4626;
  assign n4628 = n4612 & n4627;
  assign n4629 = n3558 & n4628;
  assign n4630 = n4629 ^ n4188;
  assign n4631 = ~n4601 & ~n4630;
  assign n4632 = ~n4600 & n4631;
  assign n4633 = n4632 ^ n4188;
  assign n4634 = n4633 ^ n4516;
  assign n4635 = ~n4517 & ~n4634;
  assign n4636 = n4635 ^ n4633;
  assign n4638 = n4637 ^ n4636;
  assign n4639 = n44 & ~n4434;
  assign n4640 = ~n2482 & n3280;
  assign n4641 = ~n2357 & n3275;
  assign n4642 = ~n4640 & ~n4641;
  assign n4643 = ~n2423 & n3277;
  assign n4644 = n4642 & ~n4643;
  assign n4645 = ~n4639 & n4644;
  assign n4646 = n4645 ^ x29;
  assign n4647 = n4646 ^ n4636;
  assign n4648 = ~n4638 & ~n4647;
  assign n4649 = n4648 ^ n4646;
  assign n4651 = n4650 ^ n4649;
  assign n4654 = n3285 & ~n4653;
  assign n4655 = ~n2574 & ~n3440;
  assign n4656 = ~n2669 & n3435;
  assign n4657 = ~n2786 & n3437;
  assign n4658 = ~n4656 & ~n4657;
  assign n4659 = ~n4655 & n4658;
  assign n4660 = ~n4654 & n4659;
  assign n4661 = n4660 ^ x26;
  assign n4662 = n4661 ^ n4649;
  assign n4663 = n4651 & ~n4662;
  assign n4664 = n4663 ^ n4650;
  assign n4665 = n4664 ^ n4503;
  assign n4666 = n4504 & n4665;
  assign n4667 = n4666 ^ n4664;
  assign n4668 = n4667 ^ n4491;
  assign n4669 = n4492 & n4668;
  assign n4670 = n4669 ^ n4667;
  assign n4693 = n4692 ^ n4670;
  assign n4849 = n4848 ^ n4705;
  assign n4850 = n4849 ^ n4692;
  assign n4851 = ~n4693 & n4850;
  assign n4852 = n4851 ^ n4849;
  assign n4861 = n4860 ^ n4852;
  assign n4959 = n4958 ^ n4861;
  assign n3432 = n3431 ^ n3411;
  assign n4961 = x15 ^ x14;
  assign n4962 = x17 ^ x16;
  assign n4963 = n4961 & n4962;
  assign n4964 = ~n3432 & n4963;
  assign n4965 = ~x14 & ~x15;
  assign n4966 = ~x16 & n4965;
  assign n4967 = x14 & x15;
  assign n4968 = x16 & n4967;
  assign n4969 = ~n4966 & ~n4968;
  assign n4970 = n4962 & ~n4969;
  assign n4971 = ~n3351 & n4970;
  assign n4972 = n4961 & ~n4962;
  assign n4973 = ~n3431 & n4972;
  assign n4974 = ~n4971 & ~n4973;
  assign n4975 = x16 ^ x15;
  assign n4976 = ~n4961 & n4975;
  assign n4977 = ~n3404 & n4976;
  assign n4978 = n4974 & ~n4977;
  assign n4979 = ~n4964 & n4978;
  assign n4980 = n4979 ^ x17;
  assign n4960 = n4849 ^ n4693;
  assign n4981 = n4980 ^ n4960;
  assign n3647 = n3196 ^ n3107;
  assign n5193 = n3647 & n4673;
  assign n5194 = ~n3098 & n4685;
  assign n5195 = ~n3196 & n4688;
  assign n5196 = ~n5194 & ~n5195;
  assign n5197 = ~n2954 & ~n4681;
  assign n5198 = n5196 & ~n5197;
  assign n5199 = ~n5193 & n5198;
  assign n5200 = n5199 ^ x20;
  assign n4990 = n4664 ^ n4504;
  assign n4982 = n3749 & n4478;
  assign n4983 = ~n368 & n4487;
  assign n4984 = ~n2861 & n4480;
  assign n4985 = ~n4983 & ~n4984;
  assign n4986 = ~n566 & n4484;
  assign n4987 = n4985 & ~n4986;
  assign n4988 = ~n4982 & n4987;
  assign n4989 = n4988 ^ x23;
  assign n4991 = n4990 ^ n4989;
  assign n4993 = ~n3666 & n4478;
  assign n4994 = ~n2718 & n4480;
  assign n4995 = ~n2861 & n4484;
  assign n4996 = ~n4994 & ~n4995;
  assign n4997 = ~n566 & n4487;
  assign n4998 = n4996 & ~n4997;
  assign n4999 = ~n4993 & n4998;
  assign n5000 = n4999 ^ x23;
  assign n4992 = n4661 ^ n4651;
  assign n5001 = n5000 ^ n4992;
  assign n5003 = n3285 & ~n4453;
  assign n5004 = ~n2612 & ~n3440;
  assign n5005 = ~n2574 & n3435;
  assign n5006 = ~n5004 & ~n5005;
  assign n5007 = ~n2669 & n3437;
  assign n5008 = n5006 & ~n5007;
  assign n5009 = ~n5003 & n5008;
  assign n5010 = n5009 ^ x26;
  assign n5002 = n4646 ^ n4638;
  assign n5011 = n5010 ^ n5002;
  assign n5013 = n44 & ~n4293;
  assign n5014 = ~n2423 & n3280;
  assign n5015 = ~n2247 & n3275;
  assign n5016 = ~n5014 & ~n5015;
  assign n5017 = ~n2357 & n3277;
  assign n5018 = n5016 & ~n5017;
  assign n5019 = ~n5013 & n5018;
  assign n5020 = n5019 ^ x29;
  assign n5012 = n4633 ^ n4517;
  assign n5021 = n5020 ^ n5012;
  assign n5166 = ~n1975 & ~n2369;
  assign n5167 = n5166 ^ n2065;
  assign n5168 = n3667 & ~n5167;
  assign n5169 = ~n2065 & n3676;
  assign n5170 = ~n1974 & ~n3673;
  assign n5171 = ~n5169 & ~n5170;
  assign n5172 = ~n1878 & n3669;
  assign n5173 = n5171 & ~n5172;
  assign n5174 = ~n5168 & n5173;
  assign n5153 = n44 & ~n4253;
  assign n5154 = ~n2065 & n3275;
  assign n5155 = ~n2175 & n3277;
  assign n5156 = ~n5154 & ~n5155;
  assign n5157 = ~n2247 & n3280;
  assign n5158 = n5156 & ~n5157;
  assign n5159 = ~n5153 & n5158;
  assign n5160 = n5159 ^ x29;
  assign n5023 = ~n1799 & ~n2367;
  assign n5024 = x31 & n5023;
  assign n5025 = n5024 ^ n1878;
  assign n5026 = n41 & ~n5025;
  assign n5027 = ~n1726 & n3669;
  assign n5028 = ~n1798 & ~n3673;
  assign n5029 = ~n5027 & ~n5028;
  assign n5030 = ~n5026 & n5029;
  assign n5022 = n4588 ^ n4518;
  assign n5031 = n5030 ^ n5022;
  assign n5068 = ~n1545 & ~n2364;
  assign n5069 = n5068 ^ n1638;
  assign n5070 = n3667 & ~n5069;
  assign n5071 = n54 & n1544;
  assign n5072 = n3640 & ~n5071;
  assign n5073 = ~n54 & n1638;
  assign n5074 = n5072 & ~n5073;
  assign n5075 = ~n1544 & n3672;
  assign n5076 = ~n734 & n3669;
  assign n5077 = ~n5075 & ~n5076;
  assign n5078 = ~n5074 & n5077;
  assign n5079 = ~n5070 & n5078;
  assign n5034 = n5032 & n5033;
  assign n5035 = n1293 & n5034;
  assign n5036 = ~n330 & ~n928;
  assign n5037 = ~n843 & n5036;
  assign n5038 = ~n492 & ~n1266;
  assign n5039 = n2165 & n5038;
  assign n5040 = n5037 & n5039;
  assign n5041 = ~n313 & ~n410;
  assign n5042 = n4273 & n5041;
  assign n5043 = n1906 & n3085;
  assign n5044 = n5042 & n5043;
  assign n5045 = n5040 & n5044;
  assign n5046 = n5035 & n5045;
  assign n5053 = n5046 & n5052;
  assign n5054 = n1248 & n5053;
  assign n5055 = ~n280 & n3110;
  assign n5056 = n2906 & n5055;
  assign n5057 = n239 & n1934;
  assign n5058 = n5056 & n5057;
  assign n5059 = ~n284 & n519;
  assign n5060 = n1326 & n5059;
  assign n5061 = n5058 & n5060;
  assign n5062 = n1200 & n2107;
  assign n5063 = n4270 & n5062;
  assign n5064 = n4149 & n5063;
  assign n5065 = n5061 & n5064;
  assign n5066 = n5054 & n5065;
  assign n5067 = n2481 & n5066;
  assign n5080 = n5079 ^ n5067;
  assign n5139 = n5079 ^ x2;
  assign n5109 = n781 & n4237;
  assign n5110 = n989 & n5109;
  assign n5111 = n4355 & n5110;
  assign n3472 = ~n323 & ~n843;
  assign n5112 = n1491 & n3738;
  assign n5113 = n3472 & n5112;
  assign n5114 = n3000 & n5113;
  assign n5115 = n5111 & n5114;
  assign n5125 = n519 & n1787;
  assign n5126 = ~n253 & ~n751;
  assign n5127 = ~n567 & n5126;
  assign n5128 = n5125 & n5127;
  assign n5129 = n297 & n532;
  assign n5131 = n3453 & n5130;
  assign n5132 = n5129 & n5131;
  assign n5133 = n5128 & n5132;
  assign n5134 = n5124 & n5133;
  assign n5135 = n5115 & n5134;
  assign n5136 = n242 & n5135;
  assign n5137 = n1372 & n5136;
  assign n5081 = ~n166 & ~n439;
  assign n5082 = n860 & n2025;
  assign n5083 = n5081 & n5082;
  assign n5084 = n391 & n3163;
  assign n5085 = n61 & n815;
  assign n5086 = ~n323 & ~n5085;
  assign n5087 = n5084 & n5086;
  assign n5088 = n5083 & n5087;
  assign n5089 = n2558 & n5088;
  assign n5090 = n2070 & n2908;
  assign n5093 = ~n250 & ~n790;
  assign n5094 = n239 & n5093;
  assign n5095 = n5092 & n5094;
  assign n5096 = n5090 & n5095;
  assign n5097 = ~n148 & ~n269;
  assign n5098 = ~n243 & ~n344;
  assign n5099 = n5097 & n5098;
  assign n5100 = n1934 & n5099;
  assign n5101 = n657 & n1491;
  assign n5102 = n4028 & n5101;
  assign n5103 = n5100 & n5102;
  assign n5104 = n5096 & n5103;
  assign n5105 = n5089 & n5104;
  assign n5106 = n1709 & n5105;
  assign n5107 = n774 & n3096;
  assign n5108 = n5106 & n5107;
  assign n5138 = n5137 ^ n5108;
  assign n5140 = n5139 ^ n5138;
  assign n5141 = ~n5080 & n5140;
  assign n5142 = n5141 ^ n5080;
  assign n5143 = n5137 ^ n5067;
  assign n5144 = n5143 ^ n5141;
  assign n5145 = ~n5138 & ~n5144;
  assign n5146 = n5145 ^ n5138;
  assign n5147 = n5146 ^ n5139;
  assign n5148 = ~n5142 & n5147;
  assign n5149 = n5148 ^ x2;
  assign n5150 = n5149 ^ n5030;
  assign n5151 = ~n5031 & ~n5150;
  assign n5152 = n5151 ^ n5149;
  assign n5161 = n5160 ^ n5152;
  assign n5162 = n4601 ^ n4599;
  assign n5163 = n5162 ^ n5152;
  assign n5164 = ~n5161 & ~n5163;
  assign n5165 = n5164 ^ n5160;
  assign n5175 = n5174 ^ n5165;
  assign n5176 = ~n4600 & ~n4601;
  assign n5177 = n5176 ^ n4629;
  assign n5178 = n5177 ^ n5174;
  assign n5179 = n5175 & ~n5178;
  assign n5180 = n5179 ^ n5165;
  assign n5181 = n5180 ^ n5020;
  assign n5182 = n5021 & n5181;
  assign n5183 = n5182 ^ n5180;
  assign n5184 = n5183 ^ n5010;
  assign n5185 = ~n5011 & n5184;
  assign n5186 = n5185 ^ n5183;
  assign n5187 = n5186 ^ n5000;
  assign n5188 = ~n5001 & n5187;
  assign n5189 = n5188 ^ n5186;
  assign n5190 = n5189 ^ n4990;
  assign n5191 = n4991 & ~n5190;
  assign n5192 = n5191 ^ n5189;
  assign n5201 = n5200 ^ n5192;
  assign n5202 = n4667 ^ n4492;
  assign n5203 = n5202 ^ n5200;
  assign n5204 = n5201 & n5203;
  assign n5205 = n5204 ^ n5192;
  assign n5206 = n5205 ^ n4980;
  assign n5207 = ~n4981 & n5206;
  assign n5208 = n5207 ^ n5205;
  assign n5209 = n4959 & n5208;
  assign n3878 = ~n3876 & ~n3877;
  assign n3879 = n3878 ^ n3875;
  assign n5748 = x12 ^ x11;
  assign n5796 = x13 & n5748;
  assign n5797 = ~n3879 & n5796;
  assign n5749 = x14 ^ x13;
  assign n5750 = x13 ^ x12;
  assign n5751 = n5749 & ~n5750;
  assign n5752 = ~n5748 & n5751;
  assign n5798 = ~n3404 & n5752;
  assign n5742 = x11 & x12;
  assign n5743 = ~x13 & n5742;
  assign n5744 = ~x11 & ~x12;
  assign n5745 = x13 & n5744;
  assign n5746 = ~n5743 & ~n5745;
  assign n5799 = ~n3431 & ~n5746;
  assign n5800 = ~n5798 & ~n5799;
  assign n5801 = ~x13 & n5748;
  assign n5802 = ~n3875 & n5801;
  assign n5803 = n5800 & ~n5802;
  assign n5804 = ~n5797 & n5803;
  assign n5805 = ~x14 & ~n5804;
  assign n5806 = ~n3879 & n5801;
  assign n5807 = x14 & n5800;
  assign n5808 = ~n3875 & n5796;
  assign n5809 = n5807 & ~n5808;
  assign n5810 = ~n5806 & n5809;
  assign n5811 = ~n5805 & ~n5810;
  assign n6285 = ~n3875 & ~n3876;
  assign n6286 = n5814 & n6285;
  assign n5819 = ~x8 & ~x9;
  assign n5820 = ~x10 & n5819;
  assign n5821 = x8 & x9;
  assign n5822 = x10 & n5821;
  assign n5823 = ~n5820 & ~n5822;
  assign n5824 = n5813 & ~n5823;
  assign n6287 = ~n3875 & n5824;
  assign n6288 = ~n6286 & ~n6287;
  assign n6289 = n6288 ^ x11;
  assign n6000 = ~n5770 & n5801;
  assign n6001 = ~n3270 & n5752;
  assign n6002 = ~n3351 & ~n5746;
  assign n6003 = ~n6001 & ~n6002;
  assign n6004 = ~n3404 & n5796;
  assign n6005 = n6003 & ~n6004;
  assign n6006 = ~n6000 & n6005;
  assign n6007 = x14 & ~n6006;
  assign n6008 = ~n5770 & n5796;
  assign n6009 = ~n3404 & n5801;
  assign n6010 = ~x14 & ~n6009;
  assign n6011 = n6003 & n6010;
  assign n6012 = ~n6008 & n6011;
  assign n6013 = ~n6007 & ~n6012;
  assign n5331 = n643 & n4433;
  assign n5332 = n5331 ^ n2482;
  assign n5333 = n735 & ~n5332;
  assign n5334 = ~n2357 & ~n3440;
  assign n5335 = ~n2423 & n3435;
  assign n5336 = ~n5334 & ~n5335;
  assign n5337 = ~n5333 & n5336;
  assign n5338 = n5337 ^ x26;
  assign n5330 = n5162 ^ n5161;
  assign n5339 = n5338 ^ n5330;
  assign n5341 = n44 & ~n4507;
  assign n5342 = ~n2065 & n3277;
  assign n5343 = ~n1974 & n3275;
  assign n5344 = ~n5342 & ~n5343;
  assign n5345 = ~n2175 & n3280;
  assign n5346 = n5344 & ~n5345;
  assign n5347 = ~n5341 & n5346;
  assign n5348 = n5347 ^ x29;
  assign n5340 = n5149 ^ n5031;
  assign n5349 = n5348 ^ n5340;
  assign n5364 = n5137 ^ n5079;
  assign n5365 = ~n5080 & ~n5139;
  assign n5366 = ~n5364 & n5365;
  assign n5367 = n5366 ^ n5108;
  assign n5350 = ~n1727 & ~n2366;
  assign n5351 = n5350 ^ n1798;
  assign n5352 = n3667 & ~n5351;
  assign n5353 = n54 & ~n1638;
  assign n5354 = ~n91 & ~n3671;
  assign n5355 = ~n1726 & ~n5354;
  assign n5356 = ~n5353 & ~n5355;
  assign n5357 = ~x31 & n1726;
  assign n5358 = ~x31 & ~n54;
  assign n5359 = ~n5357 & ~n5358;
  assign n5360 = ~n5356 & n5359;
  assign n5361 = ~n1798 & n3676;
  assign n5362 = ~n5360 & ~n5361;
  assign n5363 = ~n5352 & n5362;
  assign n5368 = n5367 ^ n5363;
  assign n5702 = ~n1639 & ~n2365;
  assign n5703 = n5702 ^ n1726;
  assign n5704 = n41 & n5703;
  assign n5705 = x31 & ~n5071;
  assign n5706 = n91 & n1638;
  assign n5707 = n5705 & ~n5706;
  assign n5708 = ~n5704 & n5707;
  assign n5709 = ~x31 & n5353;
  assign n5710 = ~n1726 & n3676;
  assign n5711 = ~n5709 & ~n5710;
  assign n5712 = ~n5708 & n5711;
  assign n5371 = n5023 ^ n1878;
  assign n5372 = n44 & ~n5371;
  assign n5373 = ~n1726 & n3275;
  assign n5374 = ~n1878 & n3280;
  assign n5375 = ~n5373 & ~n5374;
  assign n5376 = ~n1798 & n3277;
  assign n5377 = n5375 & ~n5376;
  assign n5378 = ~n5372 & n5377;
  assign n5379 = n5378 ^ x29;
  assign n5369 = n5067 ^ x2;
  assign n5370 = n5369 ^ n5079;
  assign n5380 = n5379 ^ n5370;
  assign n5415 = ~n1420 & ~n2363;
  assign n5416 = n5415 ^ n1544;
  assign n5417 = n3667 & ~n5416;
  assign n5418 = ~n882 & n3669;
  assign n5419 = ~n1544 & n3676;
  assign n5420 = ~n5418 & ~n5419;
  assign n5421 = ~n734 & ~n3673;
  assign n5422 = n5420 & ~n5421;
  assign n5423 = ~n5417 & n5422;
  assign n5383 = ~n238 & ~n304;
  assign n5384 = n3354 & n5383;
  assign n5385 = n5382 & n5384;
  assign n5386 = ~n535 & ~n549;
  assign n5387 = n2595 & n5386;
  assign n5388 = n1615 & n2518;
  assign n5389 = n5387 & n5388;
  assign n5390 = n5385 & n5389;
  assign n5391 = ~n791 & n2126;
  assign n5392 = n2963 & n5391;
  assign n5393 = n5390 & n5392;
  assign n5394 = ~n263 & n1295;
  assign n5395 = n5125 & n5394;
  assign n5396 = n4538 & n5395;
  assign n5397 = n5393 & n5396;
  assign n5398 = n4575 & n5397;
  assign n5399 = ~n429 & ~n1060;
  assign n5400 = ~n273 & ~n506;
  assign n5401 = n5399 & n5400;
  assign n5402 = n3050 & n5401;
  assign n5403 = ~n127 & ~n478;
  assign n5404 = n2707 & n5403;
  assign n5405 = n1567 & n2975;
  assign n5406 = n5404 & n5405;
  assign n5407 = n5402 & n5406;
  assign n5408 = n1810 & n4916;
  assign n5409 = n1191 & n5408;
  assign n5410 = n4359 & n5409;
  assign n5411 = n5407 & n5410;
  assign n5412 = n2011 & n5411;
  assign n5413 = n4898 & n5412;
  assign n5414 = n5398 & n5413;
  assign n5424 = n5423 ^ n5414;
  assign n5463 = n54 & ~n970;
  assign n5464 = n1418 ^ n882;
  assign n5465 = n5464 ^ n734;
  assign n5466 = n41 & ~n5465;
  assign n5467 = ~n5463 & ~n5466;
  assign n5468 = x31 & ~n5467;
  assign n5469 = ~n882 & ~n3673;
  assign n5470 = ~n734 & n3676;
  assign n5471 = ~n5469 & ~n5470;
  assign n5472 = ~n5468 & n5471;
  assign n5425 = ~n228 & ~n740;
  assign n5426 = n1716 & n5425;
  assign n5427 = n532 & n5426;
  assign n5428 = n2417 & n5427;
  assign n5429 = n1296 & n2135;
  assign n5430 = n5428 & n5429;
  assign n5431 = n498 & n1421;
  assign n5432 = n1854 & n5431;
  assign n5433 = n4109 & n4566;
  assign n5434 = n844 & n2076;
  assign n5435 = n5433 & n5434;
  assign n5436 = ~n197 & n3353;
  assign n5437 = n3155 & n5436;
  assign n5438 = n5435 & n5437;
  assign n5439 = n5432 & n5438;
  assign n5440 = n5430 & n5439;
  assign n5441 = n4031 & n5440;
  assign n5444 = n4190 & n5443;
  assign n5445 = ~n202 & ~n901;
  assign n5446 = n1782 & n5445;
  assign n5447 = n1198 & n5446;
  assign n5448 = n5444 & n5447;
  assign n5449 = ~n170 & ~n382;
  assign n5450 = ~n301 & n5449;
  assign n5452 = n158 & n5451;
  assign n5453 = ~n362 & ~n5452;
  assign n5454 = n930 & n5453;
  assign n5455 = n5450 & n5454;
  assign n5456 = n4273 & n5081;
  assign n5457 = n360 & n4424;
  assign n5458 = n5456 & n5457;
  assign n5459 = n5455 & n5458;
  assign n5460 = n5448 & n5459;
  assign n5461 = n289 & n5460;
  assign n5462 = n5441 & n5461;
  assign n5473 = n5472 ^ n5462;
  assign n5490 = ~n281 & ~n353;
  assign n5491 = ~n319 & ~n799;
  assign n5492 = n5490 & n5491;
  assign n5493 = ~n109 & ~n549;
  assign n5494 = n5492 & n5493;
  assign n5495 = ~n359 & ~n755;
  assign n5496 = n706 & n5495;
  assign n5497 = n5494 & n5496;
  assign n5498 = n3236 & n5497;
  assign n5499 = ~n57 & ~n475;
  assign n5500 = n1749 & n1957;
  assign n5501 = n5499 & n5500;
  assign n5502 = n600 & n5501;
  assign n5503 = n5498 & n5502;
  assign n5504 = n4387 & n4565;
  assign n5505 = ~n221 & ~n253;
  assign n5506 = n5091 & n5505;
  assign n5507 = n5504 & n5506;
  assign n5508 = ~n193 & ~n675;
  assign n5509 = ~n1047 & n5508;
  assign n5510 = n1673 & n5509;
  assign n5511 = n5507 & n5510;
  assign n5512 = n5503 & n5511;
  assign n5513 = ~n186 & ~n351;
  assign n5514 = ~n362 & ~n812;
  assign n5515 = n5513 & n5514;
  assign n5516 = n1360 & n2038;
  assign n5517 = n5515 & n5516;
  assign n5518 = n438 & n2521;
  assign n5519 = n5517 & n5518;
  assign n5521 = n5403 & n5520;
  assign n5522 = n4071 & n4424;
  assign n5523 = n5521 & n5522;
  assign n5524 = n1265 & n5523;
  assign n5525 = n5519 & n5524;
  assign n5526 = ~n79 & n957;
  assign n5527 = n4276 & n5526;
  assign n5528 = n5525 & n5527;
  assign n5529 = n5512 & n5528;
  assign n5530 = n4135 & n5529;
  assign n5476 = ~n1320 & n1414;
  assign n5477 = ~n1097 & ~n5476;
  assign n5478 = n5477 ^ n2360;
  assign n5479 = ~n970 & n5478;
  assign n5480 = n5479 ^ n5477;
  assign n5481 = n5480 ^ n882;
  assign n5482 = n41 & n5481;
  assign n5483 = n54 & n1097;
  assign n5484 = n91 & n970;
  assign n5485 = ~n5483 & ~n5484;
  assign n5486 = ~n5482 & n5485;
  assign n5474 = n41 & ~n882;
  assign n5475 = ~n5463 & ~n5474;
  assign n5487 = n5486 ^ n5475;
  assign n5488 = ~x31 & ~n5487;
  assign n5489 = n5488 ^ n5486;
  assign n5531 = n5530 ^ n5489;
  assign n5563 = ~n2360 & ~n5477;
  assign n5564 = n5563 ^ n970;
  assign n5565 = n41 & ~n5564;
  assign n5566 = n54 & ~n1414;
  assign n5567 = n91 & ~n1097;
  assign n5568 = ~n5566 & ~n5567;
  assign n5569 = ~n5565 & n5568;
  assign n5570 = x31 & ~n5569;
  assign n5571 = n3640 & ~n5483;
  assign n5572 = ~n54 & n970;
  assign n5573 = n5571 & ~n5572;
  assign n5574 = ~n5570 & ~n5573;
  assign n3906 = ~n354 & ~n456;
  assign n3907 = ~n201 & ~n256;
  assign n3908 = n3906 & n3907;
  assign n5532 = n1165 & n3908;
  assign n5533 = ~n51 & ~n691;
  assign n5535 = n5533 & n5534;
  assign n5536 = n5532 & n5535;
  assign n5537 = ~n351 & n2326;
  assign n5538 = n706 & n1406;
  assign n5539 = n5537 & n5538;
  assign n5540 = n2137 & n2801;
  assign n5541 = n5539 & n5540;
  assign n5542 = n5536 & n5541;
  assign n5543 = ~n314 & ~n647;
  assign n5544 = n598 & n5543;
  assign n5545 = ~n185 & ~n558;
  assign n5546 = n5544 & n5545;
  assign n5547 = n1036 & n3170;
  assign n5548 = n5546 & n5547;
  assign n5549 = n5542 & n5548;
  assign n5550 = ~n151 & ~n557;
  assign n5551 = n376 & n5550;
  assign n5552 = n1214 & n5551;
  assign n5553 = ~n373 & ~n540;
  assign n5554 = ~n64 & n5553;
  assign n5555 = n3074 & n5554;
  assign n5556 = n5552 & n5555;
  assign n5557 = ~n103 & n2310;
  assign n5558 = n1739 & n3737;
  assign n5559 = n5557 & n5558;
  assign n5560 = n5556 & n5559;
  assign n5561 = n5549 & n5560;
  assign n5562 = n1465 & n5561;
  assign n5575 = n5574 ^ n5562;
  assign n5588 = n282 & n1039;
  assign n5589 = ~n492 & ~n1005;
  assign n5590 = ~n1166 & n5589;
  assign n5591 = n5588 & n5590;
  assign n5592 = n1537 & n1715;
  assign n5593 = n5591 & n5592;
  assign n5594 = n820 & n3009;
  assign n5595 = n3471 & n5594;
  assign n5596 = n5593 & n5595;
  assign n5597 = ~n296 & ~n582;
  assign n5598 = n3056 & n5597;
  assign n5599 = n771 & n5533;
  assign n5600 = n5598 & n5599;
  assign n5601 = n5596 & n5600;
  assign n5602 = ~n163 & n1153;
  assign n5603 = n3290 & n5602;
  assign n5604 = n1140 & n5603;
  assign n5605 = n1014 & n2298;
  assign n5606 = n2190 & n5605;
  assign n5607 = n5604 & n5606;
  assign n5608 = n5601 & n5607;
  assign n3812 = ~n531 & ~n946;
  assign n5609 = n2608 & n3812;
  assign n5610 = n875 & n2209;
  assign n5611 = n5609 & n5610;
  assign n5612 = n2204 & n5611;
  assign n5613 = ~n83 & ~n628;
  assign n5614 = ~n208 & n5613;
  assign n5615 = n229 & n1688;
  assign n5616 = n5614 & n5615;
  assign n5617 = n5612 & n5616;
  assign n5619 = ~n243 & ~n392;
  assign n5620 = ~n186 & ~n514;
  assign n5621 = n5619 & n5620;
  assign n5622 = n5618 & n5621;
  assign n5624 = n5622 & n5623;
  assign n5625 = n1384 & n5624;
  assign n5626 = n5617 & n5625;
  assign n5627 = n1580 & n5626;
  assign n5628 = n5608 & n5627;
  assign n5578 = ~n2359 & ~n5476;
  assign n5579 = n5578 ^ n1097;
  assign n5580 = n41 & n5579;
  assign n5581 = n54 & n1208;
  assign n5582 = n91 & n1414;
  assign n5583 = ~n5581 & ~n5582;
  assign n5584 = ~n5580 & n5583;
  assign n5576 = n41 & ~n1097;
  assign n5577 = ~n5566 & ~n5576;
  assign n5585 = n5584 ^ n5577;
  assign n5586 = ~x31 & ~n5585;
  assign n5587 = n5586 ^ n5584;
  assign n5629 = n5628 ^ n5587;
  assign n5630 = ~n1208 & n1319;
  assign n5631 = x31 & n5630;
  assign n5632 = n41 & ~n1414;
  assign n5633 = ~n5631 & n5632;
  assign n5634 = n1319 & n1414;
  assign n5635 = n41 & ~n5634;
  assign n5636 = n54 ^ x31;
  assign n5637 = ~n1208 & n5636;
  assign n5638 = ~n5635 & n5637;
  assign n5639 = ~n1319 & n3669;
  assign n5640 = ~n5638 & ~n5639;
  assign n5641 = ~n5633 & n5640;
  assign n5642 = n852 & n2842;
  assign n5643 = n949 & n5505;
  assign n5644 = n5642 & n5643;
  assign n5645 = ~n273 & ~n689;
  assign n5646 = ~n277 & n5645;
  assign n5647 = n184 & n1021;
  assign n5648 = n5646 & n5647;
  assign n5649 = n5644 & n5648;
  assign n5650 = ~n797 & ~n850;
  assign n5651 = n3191 & n5650;
  assign n5652 = n5649 & n5651;
  assign n5653 = n2190 & n2550;
  assign n5654 = n229 & n5653;
  assign n5655 = ~n93 & ~n416;
  assign n5656 = n2225 & n5655;
  assign n5657 = n5654 & n5656;
  assign n5658 = n285 & n1871;
  assign n5659 = ~n337 & ~n576;
  assign n5660 = n5658 & n5659;
  assign n5661 = n5657 & n5660;
  assign n5662 = n5652 & n5661;
  assign n5663 = n1722 & n5662;
  assign n5664 = n411 & n3004;
  assign n5665 = n5455 & n5664;
  assign n5666 = ~n652 & n2076;
  assign n5667 = n2618 & n5666;
  assign n5668 = ~n98 & ~n843;
  assign n5669 = ~n1166 & n5668;
  assign n5670 = n2486 & n5669;
  assign n5671 = n5667 & n5670;
  assign n5672 = n5665 & n5671;
  assign n5673 = n836 & n1652;
  assign n3499 = ~n248 & n1992;
  assign n5674 = n1020 & n3499;
  assign n5675 = ~n373 & ~n535;
  assign n5676 = n1771 & n5675;
  assign n5677 = n5674 & n5676;
  assign n5678 = n5673 & n5677;
  assign n5679 = n5672 & n5678;
  assign n5680 = n5663 & n5679;
  assign n3892 = n495 & n1087;
  assign n3893 = ~n616 & ~n683;
  assign n3894 = n2435 & n3893;
  assign n3895 = n3892 & n3894;
  assign n3896 = n1301 & n2038;
  assign n3897 = ~n680 & n3307;
  assign n3898 = n3896 & n3897;
  assign n3899 = n3895 & n3898;
  assign n3900 = n1731 & n3899;
  assign n3901 = ~n308 & ~n660;
  assign n3902 = ~n326 & n3901;
  assign n3903 = n1332 & n3902;
  assign n3909 = n3905 & n3908;
  assign n3910 = n3903 & n3909;
  assign n3911 = n3900 & n3910;
  assign n5681 = n450 & n3911;
  assign n5682 = n5680 & n5681;
  assign n5683 = ~n5641 & ~n5682;
  assign n5684 = n5683 ^ n5587;
  assign n5685 = n5629 & n5684;
  assign n5686 = n5685 ^ n5683;
  assign n5687 = n5686 ^ n5574;
  assign n5688 = ~n5575 & ~n5687;
  assign n5689 = n5688 ^ n5686;
  assign n5690 = n5689 ^ n5489;
  assign n5691 = n5531 & n5690;
  assign n5692 = n5691 ^ n5689;
  assign n5693 = n5692 ^ n5472;
  assign n5694 = ~n5473 & ~n5693;
  assign n5695 = n5694 ^ n5692;
  assign n5696 = n5695 ^ n5423;
  assign n5697 = ~n5424 & ~n5696;
  assign n5698 = n5697 ^ n5695;
  assign n5699 = n5698 ^ n5379;
  assign n5700 = n5380 & ~n5699;
  assign n5701 = n5700 ^ n5698;
  assign n5713 = n5712 ^ n5701;
  assign n5714 = n5365 ^ n5137;
  assign n5715 = n5714 ^ n5712;
  assign n5716 = ~n5713 & ~n5715;
  assign n5717 = n5716 ^ n5701;
  assign n5718 = n5717 ^ n5367;
  assign n5719 = ~n5368 & ~n5718;
  assign n5720 = n5719 ^ n5717;
  assign n5721 = n5720 ^ n5348;
  assign n5722 = n5349 & ~n5721;
  assign n5723 = n5722 ^ n5720;
  assign n5724 = n5723 ^ n5338;
  assign n5725 = ~n5339 & ~n5724;
  assign n5726 = n5725 ^ n5723;
  assign n5238 = n3285 & ~n4334;
  assign n5239 = ~n2482 & n3435;
  assign n5240 = ~n2423 & ~n3440;
  assign n5241 = ~n5239 & ~n5240;
  assign n5242 = ~n2612 & n3437;
  assign n5243 = n5241 & ~n5242;
  assign n5244 = ~n5238 & n5243;
  assign n5245 = n5244 ^ x26;
  assign n5236 = n5177 ^ n5175;
  assign n5228 = n44 & ~n4323;
  assign n5229 = ~n2357 & n3280;
  assign n5230 = ~n2175 & n3275;
  assign n5231 = ~n5229 & ~n5230;
  assign n5232 = ~n2247 & n3277;
  assign n5233 = n5231 & ~n5232;
  assign n5234 = ~n5228 & n5233;
  assign n5235 = n5234 ^ x29;
  assign n5237 = n5236 ^ n5235;
  assign n5328 = n5245 ^ n5237;
  assign n5320 = n4478 & ~n4653;
  assign n5321 = ~n2574 & n4480;
  assign n5322 = ~n2669 & n4484;
  assign n5323 = ~n2786 & n4487;
  assign n5324 = ~n5322 & ~n5323;
  assign n5325 = ~n5321 & n5324;
  assign n5326 = ~n5320 & n5325;
  assign n5327 = n5326 ^ x23;
  assign n5329 = n5328 ^ n5327;
  assign n5847 = n5726 ^ n5329;
  assign n5839 = ~n3666 & n4673;
  assign n5840 = ~n2718 & ~n4681;
  assign n5841 = ~n2861 & n4685;
  assign n5842 = ~n5840 & ~n5841;
  assign n5843 = ~n566 & n4688;
  assign n5844 = n5842 & ~n5843;
  assign n5845 = ~n5839 & n5844;
  assign n5846 = n5845 ^ x20;
  assign n5848 = n5847 ^ n5846;
  assign n5883 = n5723 ^ n5339;
  assign n5870 = n5720 ^ n5349;
  assign n5857 = n3285 & ~n4323;
  assign n5858 = ~n2357 & n3437;
  assign n5859 = ~n2247 & n3435;
  assign n5860 = ~n5858 & ~n5859;
  assign n5861 = ~n2175 & ~n3440;
  assign n5862 = n5860 & ~n5861;
  assign n5863 = ~n5857 & n5862;
  assign n5864 = n5863 ^ x26;
  assign n5849 = n44 & ~n5167;
  assign n5850 = ~n1878 & n3275;
  assign n5851 = ~n1974 & n3277;
  assign n5852 = ~n5850 & ~n5851;
  assign n5853 = ~n2065 & n3280;
  assign n5854 = n5852 & ~n5853;
  assign n5855 = ~n5849 & n5854;
  assign n5856 = n5855 ^ x29;
  assign n5865 = n5864 ^ n5856;
  assign n5866 = n5717 ^ n5368;
  assign n5867 = n5866 ^ n5864;
  assign n5868 = ~n5865 & ~n5867;
  assign n5869 = n5868 ^ n5866;
  assign n5871 = n5870 ^ n5869;
  assign n5872 = n3285 & ~n4293;
  assign n5873 = ~n2423 & n3437;
  assign n5874 = ~n2247 & ~n3440;
  assign n5875 = ~n5873 & ~n5874;
  assign n5876 = ~n2357 & n3435;
  assign n5877 = n5875 & ~n5876;
  assign n5878 = ~n5872 & n5877;
  assign n5879 = n5878 ^ x26;
  assign n5880 = n5879 ^ n5869;
  assign n5881 = ~n5871 & n5880;
  assign n5882 = n5881 ^ n5870;
  assign n5884 = n5883 ^ n5882;
  assign n5885 = ~n4453 & n4478;
  assign n5886 = ~n2612 & n4480;
  assign n5887 = ~n2669 & n4487;
  assign n5888 = ~n5886 & ~n5887;
  assign n5889 = ~n2574 & n4484;
  assign n5890 = n5888 & ~n5889;
  assign n5891 = ~n5885 & n5890;
  assign n5892 = n5891 ^ x23;
  assign n5893 = n5892 ^ n5882;
  assign n5894 = ~n5884 & ~n5893;
  assign n5895 = n5894 ^ n5883;
  assign n5896 = n5895 ^ n5847;
  assign n5897 = n5848 & n5896;
  assign n5898 = n5897 ^ n5895;
  assign n5727 = n5726 ^ n5328;
  assign n5728 = ~n5329 & ~n5727;
  assign n5729 = n5728 ^ n5726;
  assign n5246 = n5245 ^ n5235;
  assign n5247 = n5237 & ~n5246;
  assign n5248 = n5247 ^ n5236;
  assign n5226 = n5180 ^ n5021;
  assign n5218 = n3285 & ~n4312;
  assign n5219 = ~n2612 & n3435;
  assign n5220 = ~n2574 & n3437;
  assign n5221 = ~n5219 & ~n5220;
  assign n5222 = ~n2482 & ~n3440;
  assign n5223 = n5221 & ~n5222;
  assign n5224 = ~n5218 & n5223;
  assign n5225 = n5224 ^ x26;
  assign n5227 = n5226 ^ n5225;
  assign n5318 = n5248 ^ n5227;
  assign n5310 = n4478 & ~n4495;
  assign n5311 = ~n2718 & n4487;
  assign n5312 = ~n2669 & n4480;
  assign n5313 = ~n2786 & n4484;
  assign n5314 = ~n5312 & ~n5313;
  assign n5315 = ~n5311 & n5314;
  assign n5316 = ~n5310 & n5315;
  assign n5317 = n5316 ^ x23;
  assign n5319 = n5318 ^ n5317;
  assign n5837 = n5729 ^ n5319;
  assign n5829 = n3749 & n4673;
  assign n5830 = ~n368 & n4688;
  assign n5831 = ~n2861 & ~n4681;
  assign n5832 = ~n5830 & ~n5831;
  assign n5833 = ~n566 & n4685;
  assign n5834 = n5832 & ~n5833;
  assign n5835 = ~n5829 & n5834;
  assign n5836 = n5835 ^ x20;
  assign n5838 = n5837 ^ n5836;
  assign n5987 = n5898 ^ n5838;
  assign n5921 = n5895 ^ n5848;
  assign n5913 = ~n3777 & n4963;
  assign n5914 = ~n2954 & n4972;
  assign n5915 = ~n368 & n4970;
  assign n5916 = ~n5914 & ~n5915;
  assign n5917 = ~n3037 & n4976;
  assign n5918 = n5916 & ~n5917;
  assign n5919 = ~n5913 & n5918;
  assign n5920 = n5919 ^ x17;
  assign n5922 = n5921 ^ n5920;
  assign n5971 = n5892 ^ n5884;
  assign n5958 = ~n4312 & n4478;
  assign n5959 = ~n2612 & n4484;
  assign n5960 = ~n2482 & n4480;
  assign n5961 = ~n5959 & ~n5960;
  assign n5962 = ~n2574 & n4487;
  assign n5963 = n5961 & ~n5962;
  assign n5964 = ~n5958 & n5963;
  assign n5965 = n5964 ^ x23;
  assign n5945 = ~n4334 & n4478;
  assign n5946 = ~n2482 & n4484;
  assign n5947 = ~n2423 & n4480;
  assign n5948 = ~n5946 & ~n5947;
  assign n5949 = ~n2612 & n4487;
  assign n5950 = n5948 & ~n5949;
  assign n5951 = ~n5945 & n5950;
  assign n5952 = n5951 ^ x23;
  assign n5932 = n3285 & ~n4253;
  assign n5933 = ~n2175 & n3435;
  assign n5934 = ~n2247 & n3437;
  assign n5935 = ~n5933 & ~n5934;
  assign n5936 = ~n2065 & ~n3440;
  assign n5937 = n5935 & ~n5936;
  assign n5938 = ~n5932 & n5937;
  assign n5939 = n5938 ^ x26;
  assign n5923 = n4592 ^ n1974;
  assign n5924 = n44 & ~n5923;
  assign n5925 = ~n1878 & n3277;
  assign n5926 = ~n1974 & n3280;
  assign n5927 = ~n5925 & ~n5926;
  assign n5928 = ~n1798 & n3275;
  assign n5929 = n5927 & ~n5928;
  assign n5930 = ~n5924 & n5929;
  assign n5931 = n5930 ^ x29;
  assign n5940 = n5939 ^ n5931;
  assign n5941 = n5714 ^ n5713;
  assign n5942 = n5941 ^ n5939;
  assign n5943 = ~n5940 & ~n5942;
  assign n5944 = n5943 ^ n5941;
  assign n5953 = n5952 ^ n5944;
  assign n5954 = n5866 ^ n5865;
  assign n5955 = n5954 ^ n5944;
  assign n5956 = n5953 & n5955;
  assign n5957 = n5956 ^ n5954;
  assign n5966 = n5965 ^ n5957;
  assign n5967 = n5879 ^ n5871;
  assign n5968 = n5967 ^ n5957;
  assign n5969 = n5966 & n5968;
  assign n5970 = n5969 ^ n5967;
  assign n5972 = n5971 ^ n5970;
  assign n5973 = ~n4466 & n4673;
  assign n5974 = ~n2718 & n4685;
  assign n5975 = ~n2786 & ~n4681;
  assign n5976 = ~n2861 & n4688;
  assign n5977 = ~n5975 & ~n5976;
  assign n5978 = ~n5974 & n5977;
  assign n5979 = ~n5973 & n5978;
  assign n5980 = n5979 ^ x20;
  assign n5981 = n5980 ^ n5970;
  assign n5982 = n5972 & n5981;
  assign n5983 = n5982 ^ n5971;
  assign n5984 = n5983 ^ n5921;
  assign n5985 = ~n5922 & ~n5984;
  assign n5986 = n5985 ^ n5983;
  assign n5988 = n5987 ^ n5986;
  assign n5989 = ~n3974 & n4963;
  assign n5990 = ~n2954 & n4976;
  assign n5991 = ~n3037 & n4970;
  assign n5992 = ~n5990 & ~n5991;
  assign n5993 = ~n3098 & n4972;
  assign n5994 = n5992 & ~n5993;
  assign n5995 = ~n5989 & n5994;
  assign n5996 = n5995 ^ x17;
  assign n5997 = n5996 ^ n5986;
  assign n5998 = n5988 & n5997;
  assign n5999 = n5998 ^ n5987;
  assign n6014 = n6013 ^ n5999;
  assign n5730 = n5729 ^ n5318;
  assign n5731 = n5319 & n5730;
  assign n5732 = n5731 ^ n5729;
  assign n5261 = n5183 ^ n5011;
  assign n5252 = ~n4466 & n4478;
  assign n5253 = ~n2718 & n4484;
  assign n5254 = ~n2786 & n4480;
  assign n5255 = ~n2861 & n4487;
  assign n5256 = ~n5254 & ~n5255;
  assign n5257 = ~n5253 & n5256;
  assign n5258 = ~n5252 & n5257;
  assign n5259 = n5258 ^ x23;
  assign n5249 = n5248 ^ n5226;
  assign n5250 = n5227 & ~n5249;
  assign n5251 = n5250 ^ n5248;
  assign n5260 = n5259 ^ n5251;
  assign n5308 = n5261 ^ n5260;
  assign n5300 = ~n3632 & n4673;
  assign n5301 = ~n368 & n4685;
  assign n5302 = ~n3037 & n4688;
  assign n5303 = ~n5301 & ~n5302;
  assign n5304 = ~n566 & ~n4681;
  assign n5305 = n5303 & ~n5304;
  assign n5306 = ~n5300 & n5305;
  assign n5307 = n5306 ^ x20;
  assign n5309 = n5308 ^ n5307;
  assign n5910 = n5732 ^ n5309;
  assign n5902 = n3647 & n4963;
  assign n5903 = ~n2954 & n4970;
  assign n5904 = ~n3098 & n4976;
  assign n5905 = ~n5903 & ~n5904;
  assign n5906 = ~n3196 & n4972;
  assign n5907 = n5905 & ~n5906;
  assign n5908 = ~n5902 & n5907;
  assign n5909 = n5908 ^ x17;
  assign n5911 = n5910 ^ n5909;
  assign n5899 = n5898 ^ n5837;
  assign n5900 = ~n5838 & ~n5899;
  assign n5901 = n5900 ^ n5898;
  assign n5912 = n5911 ^ n5901;
  assign n6282 = n6013 ^ n5912;
  assign n6283 = n6014 & n6282;
  assign n6284 = n6283 ^ n5999;
  assign n6290 = n6289 ^ n6284;
  assign n5733 = n5732 ^ n5308;
  assign n5734 = ~n5309 & ~n5733;
  assign n5735 = n5734 ^ n5732;
  assign n5267 = ~n3777 & n4673;
  assign n5268 = ~n2954 & n4688;
  assign n5269 = ~n368 & ~n4681;
  assign n5270 = ~n5268 & ~n5269;
  assign n5271 = ~n3037 & n4685;
  assign n5272 = n5270 & ~n5271;
  assign n5273 = ~n5267 & n5272;
  assign n5274 = n5273 ^ x20;
  assign n5265 = n5186 ^ n5001;
  assign n5262 = n5261 ^ n5259;
  assign n5263 = n5260 & ~n5262;
  assign n5264 = n5263 ^ n5251;
  assign n5266 = n5265 ^ n5264;
  assign n5298 = n5274 ^ n5266;
  assign n5290 = ~n3271 & n4963;
  assign n5291 = ~n3098 & n4970;
  assign n5292 = ~n3196 & n4976;
  assign n5293 = ~n5291 & ~n5292;
  assign n5294 = ~n3270 & n4972;
  assign n5295 = n5293 & ~n5294;
  assign n5296 = ~n5290 & n5295;
  assign n5297 = n5296 ^ x17;
  assign n5299 = n5298 ^ n5297;
  assign n6279 = n5735 ^ n5299;
  assign n6265 = ~n3432 & n5801;
  assign n6266 = ~n3404 & ~n5746;
  assign n6267 = ~n3351 & n5752;
  assign n6268 = ~n6266 & ~n6267;
  assign n6269 = ~n3431 & n5796;
  assign n6270 = n6268 & ~n6269;
  assign n6271 = ~n6265 & n6270;
  assign n6272 = x14 & ~n6271;
  assign n6273 = ~n3432 & n5796;
  assign n6274 = ~n3431 & n5801;
  assign n6275 = ~x14 & ~n6274;
  assign n6276 = n6268 & n6275;
  assign n6277 = ~n6273 & n6276;
  assign n6278 = ~n6272 & ~n6277;
  assign n6280 = n6279 ^ n6278;
  assign n6262 = n5910 ^ n5901;
  assign n6263 = n5911 & n6262;
  assign n6264 = n6263 ^ n5901;
  assign n6281 = n6280 ^ n6264;
  assign n6291 = n6290 ^ n6281;
  assign n6015 = n6014 ^ n5912;
  assign n5815 = n5758 & n5814;
  assign n5816 = x10 ^ x9;
  assign n5817 = ~n5812 & n5816;
  assign n5818 = ~n3875 & n5817;
  assign n5825 = ~n3431 & n5824;
  assign n5826 = ~n5818 & ~n5825;
  assign n5827 = ~n5815 & n5826;
  assign n5828 = n5827 ^ x11;
  assign n6016 = n6015 ^ n5828;
  assign n6031 = n5996 ^ n5988;
  assign n6017 = ~n3989 & n5801;
  assign n6018 = ~n3270 & ~n5746;
  assign n6019 = ~n3196 & n5752;
  assign n6020 = ~n6018 & ~n6019;
  assign n6021 = ~n3351 & n5796;
  assign n6022 = n6020 & ~n6021;
  assign n6023 = ~n6017 & n6022;
  assign n6024 = x14 & ~n6023;
  assign n6025 = ~n3989 & n5796;
  assign n6026 = ~n3351 & n5801;
  assign n6027 = ~x14 & ~n6026;
  assign n6028 = n6020 & n6027;
  assign n6029 = ~n6025 & n6028;
  assign n6030 = ~n6024 & ~n6029;
  assign n6032 = n6031 ^ n6030;
  assign n6053 = n5983 ^ n5922;
  assign n6033 = ~x14 & n5748;
  assign n6034 = n6033 ^ x13;
  assign n6035 = ~n3198 & ~n6034;
  assign n6036 = n6035 ^ x13;
  assign n6037 = ~n3270 & ~n6036;
  assign n6038 = n5748 & ~n6037;
  assign n6039 = ~x13 & n3198;
  assign n6040 = n3270 & ~n6039;
  assign n6041 = ~n3098 & n5752;
  assign n6042 = ~n3196 & ~n5746;
  assign n6043 = ~n6041 & ~n6042;
  assign n6044 = x14 & n6043;
  assign n6045 = ~n3198 & ~n6044;
  assign n6046 = n6040 & ~n6045;
  assign n6047 = n6038 & ~n6046;
  assign n6048 = ~x14 & ~n5748;
  assign n6049 = n6043 & ~n6048;
  assign n6050 = ~n6047 & n6049;
  assign n6051 = ~x14 & ~n6043;
  assign n6052 = ~n6050 & ~n6051;
  assign n6054 = n6053 ^ n6052;
  assign n6063 = n5980 ^ n5972;
  assign n6055 = ~n3632 & n4963;
  assign n6056 = ~n566 & n4970;
  assign n6057 = ~n3037 & n4972;
  assign n6058 = ~n6056 & ~n6057;
  assign n6059 = ~n368 & n4976;
  assign n6060 = n6058 & ~n6059;
  assign n6061 = ~n6055 & n6060;
  assign n6062 = n6061 ^ x17;
  assign n6064 = n6063 ^ n6062;
  assign n6073 = n5967 ^ n5966;
  assign n6065 = ~n4495 & n4673;
  assign n6066 = ~n2718 & n4688;
  assign n6067 = ~n2669 & ~n4681;
  assign n6068 = ~n2786 & n4685;
  assign n6069 = ~n6067 & ~n6068;
  assign n6070 = ~n6066 & n6069;
  assign n6071 = ~n6065 & n6070;
  assign n6072 = n6071 ^ x20;
  assign n6074 = n6073 ^ n6072;
  assign n6083 = n5954 ^ n5953;
  assign n6075 = ~n4653 & n4673;
  assign n6076 = ~n2574 & ~n4681;
  assign n6077 = ~n2669 & n4685;
  assign n6078 = ~n2786 & n4688;
  assign n6079 = ~n6077 & ~n6078;
  assign n6080 = ~n6076 & n6079;
  assign n6081 = ~n6075 & n6080;
  assign n6082 = n6081 ^ x20;
  assign n6084 = n6083 ^ n6082;
  assign n6093 = n5941 ^ n5940;
  assign n6085 = ~n4434 & n4478;
  assign n6086 = ~n2423 & n4484;
  assign n6087 = ~n2482 & n4487;
  assign n6088 = ~n6086 & ~n6087;
  assign n6089 = ~n2357 & n4480;
  assign n6090 = n6088 & ~n6089;
  assign n6091 = ~n6085 & n6090;
  assign n6092 = n6091 ^ x23;
  assign n6094 = n6093 ^ n6092;
  assign n6103 = n5698 ^ n5380;
  assign n6095 = n3285 & ~n4507;
  assign n6096 = ~n2065 & n3435;
  assign n6097 = ~n1974 & ~n3440;
  assign n6098 = ~n6096 & ~n6097;
  assign n6099 = ~n2175 & n3437;
  assign n6100 = n6098 & ~n6099;
  assign n6101 = ~n6095 & n6100;
  assign n6102 = n6101 ^ x26;
  assign n6104 = n6103 ^ n6102;
  assign n6113 = n5695 ^ n5424;
  assign n6105 = n44 & ~n5351;
  assign n6106 = ~n1726 & n3277;
  assign n6107 = ~n1638 & n3275;
  assign n6108 = ~n6106 & ~n6107;
  assign n6109 = ~n1798 & n3280;
  assign n6110 = n6108 & ~n6109;
  assign n6111 = ~n6105 & n6110;
  assign n6112 = n6111 ^ x29;
  assign n6114 = n6113 ^ n6112;
  assign n6123 = n5692 ^ n5473;
  assign n6115 = n44 & ~n5703;
  assign n6116 = ~n1726 & n3280;
  assign n6117 = ~n1638 & n3277;
  assign n6118 = ~n1544 & n3275;
  assign n6119 = ~n6117 & ~n6118;
  assign n6120 = ~n6116 & n6119;
  assign n6121 = ~n6115 & n6120;
  assign n6122 = n6121 ^ x29;
  assign n6124 = n6123 ^ n6122;
  assign n6133 = n5689 ^ n5531;
  assign n6125 = n44 & ~n5069;
  assign n6126 = ~n734 & n3275;
  assign n6127 = ~n1638 & n3280;
  assign n6128 = ~n6126 & ~n6127;
  assign n6129 = ~n1544 & n3277;
  assign n6130 = n6128 & ~n6129;
  assign n6131 = ~n6125 & n6130;
  assign n6132 = n6131 ^ x29;
  assign n6134 = n6133 ^ n6132;
  assign n6143 = n5686 ^ n5575;
  assign n6135 = n44 & ~n5416;
  assign n6136 = ~n882 & n3275;
  assign n6137 = ~n734 & n3277;
  assign n6138 = ~n1544 & n3280;
  assign n6139 = ~n6137 & ~n6138;
  assign n6140 = ~n6136 & n6139;
  assign n6141 = ~n6135 & n6140;
  assign n6142 = n6141 ^ x29;
  assign n6144 = n6143 ^ n6142;
  assign n6192 = n44 & ~n5481;
  assign n6193 = ~n882 & n3280;
  assign n6194 = ~n1097 & n3275;
  assign n6195 = ~n6193 & ~n6194;
  assign n6196 = ~n970 & n3277;
  assign n6197 = n6195 & ~n6196;
  assign n6198 = ~n6192 & n6197;
  assign n6199 = n6198 ^ x29;
  assign n6151 = n44 & ~n5564;
  assign n6152 = ~n1097 & n3277;
  assign n6153 = ~n1414 & n3275;
  assign n6154 = ~n6152 & ~n6153;
  assign n6155 = ~n970 & n3280;
  assign n6156 = n6154 & ~n6155;
  assign n6157 = ~n6151 & n6156;
  assign n6158 = n6157 ^ x29;
  assign n6145 = ~n91 & ~n1208;
  assign n6146 = n6145 ^ n1319;
  assign n6148 = n6146 ^ n6145;
  assign n6149 = ~x31 & ~n6148;
  assign n6147 = ~n54 & ~n6146;
  assign n6150 = n6149 ^ n6147;
  assign n6159 = n6158 ^ n6150;
  assign n6160 = n44 & ~n5579;
  assign n6161 = ~n1208 & n3275;
  assign n6162 = ~n1414 & n3277;
  assign n6163 = ~n6161 & ~n6162;
  assign n6164 = ~n1097 & n3280;
  assign n6165 = n6163 & ~n6164;
  assign n6166 = ~n6160 & n6165;
  assign n6168 = n43 & n5630;
  assign n6169 = n6168 ^ n1414;
  assign n6170 = n42 & ~n6169;
  assign n6171 = ~n1208 & n3277;
  assign n6172 = ~n1319 & n3275;
  assign n6173 = ~n6171 & ~n6172;
  assign n6174 = ~n6170 & n6173;
  assign n6175 = n42 & ~n1208;
  assign n6176 = x26 & n65;
  assign n6177 = ~x26 & ~x27;
  assign n6178 = ~x28 & n6177;
  assign n6179 = ~n6176 & ~n6178;
  assign n6180 = ~n1319 & n6179;
  assign n6181 = ~n6175 & ~n6180;
  assign n6182 = n6174 & n6181;
  assign n6183 = ~x30 & ~n1319;
  assign n6184 = ~n6182 & ~n6183;
  assign n6185 = x29 & ~n6184;
  assign n6167 = n60 & ~n1319;
  assign n6186 = n6185 ^ n6167;
  assign n6187 = ~n6166 & n6186;
  assign n6188 = n6187 ^ n6185;
  assign n6189 = n6188 ^ n6158;
  assign n6190 = n6159 & ~n6189;
  assign n6191 = n6190 ^ n6188;
  assign n6200 = n6199 ^ n6191;
  assign n6201 = n5641 & n5682;
  assign n6202 = n6201 ^ n6199;
  assign n6203 = ~n6200 & ~n6202;
  assign n6204 = n6203 ^ n6191;
  assign n6205 = n44 & ~n5465;
  assign n6206 = ~n882 & n3277;
  assign n6207 = ~n734 & n3280;
  assign n6208 = ~n6206 & ~n6207;
  assign n6209 = ~n970 & n3275;
  assign n6210 = n6208 & ~n6209;
  assign n6211 = ~n6205 & n6210;
  assign n6212 = n6211 ^ x29;
  assign n6213 = n5629 & ~n6212;
  assign n6214 = ~n5683 & n6213;
  assign n6215 = n6214 ^ n6212;
  assign n6216 = ~n6204 & n6215;
  assign n6217 = n6191 & ~n6199;
  assign n6218 = n5683 & n6217;
  assign n6219 = ~n5629 & n6212;
  assign n6220 = n6218 & ~n6219;
  assign n6221 = n6212 ^ n5683;
  assign n6222 = n5629 & n6221;
  assign n6223 = n6222 ^ n5683;
  assign n6224 = ~n6220 & n6223;
  assign n6225 = ~n6216 & ~n6224;
  assign n6226 = n6225 ^ n6143;
  assign n6227 = n6144 & n6226;
  assign n6228 = n6227 ^ n6225;
  assign n6229 = n6228 ^ n6133;
  assign n6230 = ~n6134 & ~n6229;
  assign n6231 = n6230 ^ n6228;
  assign n6232 = n6231 ^ n6123;
  assign n6233 = n6124 & n6232;
  assign n6234 = n6233 ^ n6231;
  assign n6235 = n6234 ^ n6113;
  assign n6236 = n6114 & n6235;
  assign n6237 = n6236 ^ n6234;
  assign n6238 = n6237 ^ n6103;
  assign n6239 = ~n6104 & ~n6238;
  assign n6240 = n6239 ^ n6237;
  assign n6241 = n6240 ^ n6093;
  assign n6242 = n6094 & n6241;
  assign n6243 = n6242 ^ n6240;
  assign n6244 = n6243 ^ n6083;
  assign n6245 = ~n6084 & ~n6244;
  assign n6246 = n6245 ^ n6243;
  assign n6247 = n6246 ^ n6073;
  assign n6248 = ~n6074 & ~n6247;
  assign n6249 = n6248 ^ n6246;
  assign n6250 = n6249 ^ n6063;
  assign n6251 = ~n6064 & ~n6250;
  assign n6252 = n6251 ^ n6249;
  assign n6253 = n6252 ^ n6053;
  assign n6254 = n6054 & n6253;
  assign n6255 = n6254 ^ n6252;
  assign n6256 = n6255 ^ n6031;
  assign n6257 = n6032 & ~n6256;
  assign n6258 = n6257 ^ n6255;
  assign n6259 = n6258 ^ n6015;
  assign n6260 = ~n6016 & ~n6259;
  assign n6261 = n6260 ^ n6258;
  assign n6292 = n6291 ^ n6261;
  assign n6293 = n6255 ^ n6032;
  assign n6294 = ~n3879 & n5814;
  assign n6295 = n5812 & ~n5813;
  assign n6296 = ~n3875 & n6295;
  assign n6297 = ~n3431 & n5817;
  assign n6298 = ~n6296 & ~n6297;
  assign n6299 = ~n3404 & n5824;
  assign n6300 = n6298 & ~n6299;
  assign n6301 = ~n6294 & n6300;
  assign n6302 = n6301 ^ x11;
  assign n6303 = ~n6293 & ~n6302;
  assign n7157 = n6252 ^ n6054;
  assign n7149 = ~n3432 & n5814;
  assign n7150 = ~n3351 & n5824;
  assign n7151 = ~n3431 & n6295;
  assign n7152 = ~n7150 & ~n7151;
  assign n7153 = ~n3404 & n5817;
  assign n7154 = n7152 & ~n7153;
  assign n7155 = ~n7149 & n7154;
  assign n7156 = n7155 ^ x11;
  assign n7158 = n7157 ^ n7156;
  assign n6836 = n6249 ^ n6064;
  assign n6820 = n3107 & n3196;
  assign n6821 = n5748 & ~n6820;
  assign n6822 = ~x14 & ~n6821;
  assign n6823 = n3196 ^ x13;
  assign n6824 = ~n3107 & n6823;
  assign n6825 = n5748 & n6824;
  assign n6826 = ~n6822 & ~n6825;
  assign n6827 = ~n2954 & n5752;
  assign n6828 = ~n3098 & ~n5746;
  assign n6829 = ~n6827 & ~n6828;
  assign n6830 = ~n6826 & n6829;
  assign n6831 = ~n3196 & n5748;
  assign n6832 = n3107 & n6831;
  assign n6833 = n6829 & ~n6832;
  assign n6834 = x14 & ~n6833;
  assign n6835 = ~n6830 & ~n6834;
  assign n6837 = n6836 ^ n6835;
  assign n6564 = n6246 ^ n6074;
  assign n6556 = n3749 & n4963;
  assign n6557 = ~n368 & n4972;
  assign n6558 = ~n2861 & n4970;
  assign n6559 = ~n6557 & ~n6558;
  assign n6560 = ~n566 & n4976;
  assign n6561 = n6559 & ~n6560;
  assign n6562 = ~n6556 & n6561;
  assign n6563 = n6562 ^ x17;
  assign n6565 = n6564 ^ n6563;
  assign n6351 = n6243 ^ n6084;
  assign n6343 = ~n3666 & n4963;
  assign n6344 = ~n2718 & n4970;
  assign n6345 = ~n2861 & n4976;
  assign n6346 = ~n6344 & ~n6345;
  assign n6347 = ~n566 & n4972;
  assign n6348 = n6346 & ~n6347;
  assign n6349 = ~n6343 & n6348;
  assign n6350 = n6349 ^ x17;
  assign n6352 = n6351 ^ n6350;
  assign n6361 = n6240 ^ n6094;
  assign n6353 = ~n4453 & n4673;
  assign n6354 = ~n2612 & ~n4681;
  assign n6355 = ~n2574 & n4685;
  assign n6356 = ~n6354 & ~n6355;
  assign n6357 = ~n2669 & n4688;
  assign n6358 = n6356 & ~n6357;
  assign n6359 = ~n6353 & n6358;
  assign n6360 = n6359 ^ x20;
  assign n6362 = n6361 ^ n6360;
  assign n6371 = n6237 ^ n6104;
  assign n6363 = ~n4293 & n4478;
  assign n6364 = ~n2423 & n4487;
  assign n6365 = ~n2247 & n4480;
  assign n6366 = ~n6364 & ~n6365;
  assign n6367 = ~n2357 & n4484;
  assign n6368 = n6366 & ~n6367;
  assign n6369 = ~n6363 & n6368;
  assign n6370 = n6369 ^ x23;
  assign n6372 = n6371 ^ n6370;
  assign n6381 = n6234 ^ n6114;
  assign n6373 = n3285 & ~n5167;
  assign n6374 = ~n1878 & ~n3440;
  assign n6375 = ~n1974 & n3435;
  assign n6376 = ~n6374 & ~n6375;
  assign n6377 = ~n2065 & n3437;
  assign n6378 = n6376 & ~n6377;
  assign n6379 = ~n6373 & n6378;
  assign n6380 = n6379 ^ x26;
  assign n6382 = n6381 ^ n6380;
  assign n6391 = n6231 ^ n6124;
  assign n6383 = n3285 & ~n5923;
  assign n6384 = ~n1798 & ~n3440;
  assign n6385 = ~n1878 & n3435;
  assign n6386 = ~n6384 & ~n6385;
  assign n6387 = ~n1974 & n3437;
  assign n6388 = n6386 & ~n6387;
  assign n6389 = ~n6383 & n6388;
  assign n6390 = n6389 ^ x26;
  assign n6392 = n6391 ^ n6390;
  assign n6401 = n6228 ^ n6134;
  assign n6393 = n3285 & ~n5371;
  assign n6394 = ~n1798 & n3435;
  assign n6395 = ~n1878 & n3437;
  assign n6396 = ~n6394 & ~n6395;
  assign n6397 = ~n1726 & ~n3440;
  assign n6398 = n6396 & ~n6397;
  assign n6399 = ~n6393 & n6398;
  assign n6400 = n6399 ^ x26;
  assign n6402 = n6401 ^ n6400;
  assign n6411 = n6225 ^ n6144;
  assign n6403 = n3285 & ~n5351;
  assign n6404 = ~n1798 & n3437;
  assign n6405 = ~n1726 & n3435;
  assign n6406 = ~n6404 & ~n6405;
  assign n6407 = ~n1638 & ~n3440;
  assign n6408 = n6406 & ~n6407;
  assign n6409 = ~n6403 & n6408;
  assign n6410 = n6409 ^ x26;
  assign n6412 = n6411 ^ n6410;
  assign n6424 = n6212 ^ n5629;
  assign n6421 = n6217 ^ n6204;
  assign n6422 = ~n5683 & ~n6421;
  assign n6423 = n6422 ^ n6217;
  assign n6425 = n6424 ^ n6423;
  assign n6413 = n3285 & ~n5703;
  assign n6414 = ~n1726 & n3437;
  assign n6415 = ~n1638 & n3435;
  assign n6416 = ~n1544 & ~n3440;
  assign n6417 = ~n6415 & ~n6416;
  assign n6418 = ~n6414 & n6417;
  assign n6419 = ~n6413 & n6418;
  assign n6420 = n6419 ^ x26;
  assign n6426 = n6425 ^ n6420;
  assign n6435 = n6199 ^ n5641;
  assign n6436 = n6435 ^ n5682;
  assign n6437 = n6436 ^ n6191;
  assign n6427 = n3285 & ~n5069;
  assign n6428 = ~n734 & ~n3440;
  assign n6429 = ~n1638 & n3437;
  assign n6430 = ~n6428 & ~n6429;
  assign n6431 = ~n1544 & n3435;
  assign n6432 = n6430 & ~n6431;
  assign n6433 = ~n6427 & n6432;
  assign n6434 = n6433 ^ x26;
  assign n6438 = n6437 ^ n6434;
  assign n6447 = n6188 ^ n6159;
  assign n6439 = n3285 & ~n5416;
  assign n6440 = ~n882 & ~n3440;
  assign n6441 = ~n734 & n3435;
  assign n6442 = ~n6440 & ~n6441;
  assign n6443 = ~n1544 & n3437;
  assign n6444 = n6442 & ~n6443;
  assign n6445 = ~n6439 & n6444;
  assign n6446 = n6445 ^ x26;
  assign n6448 = n6447 ^ n6446;
  assign n6455 = n3285 & ~n5465;
  assign n6456 = ~n882 & n3435;
  assign n6457 = ~n970 & ~n3440;
  assign n6458 = ~n6456 & ~n6457;
  assign n6459 = ~n734 & n3437;
  assign n6460 = n6458 & ~n6459;
  assign n6461 = ~n6455 & n6460;
  assign n6462 = n6461 ^ x26;
  assign n6453 = n6166 ^ x29;
  assign n6450 = n6182 ^ n1319;
  assign n6451 = x29 & ~n6450;
  assign n6449 = x30 & ~n1319;
  assign n6452 = n6451 ^ n6449;
  assign n6454 = n6453 ^ n6452;
  assign n6463 = n6462 ^ n6454;
  assign n6466 = n3285 & ~n5481;
  assign n6467 = ~n882 & n3437;
  assign n6468 = ~n970 & n3435;
  assign n6469 = ~n6467 & ~n6468;
  assign n6470 = ~n1097 & ~n3440;
  assign n6471 = n6469 & ~n6470;
  assign n6472 = ~n6466 & n6471;
  assign n6473 = n6472 ^ x26;
  assign n6464 = x29 & ~n6181;
  assign n6465 = n6464 ^ n6174;
  assign n6474 = n6473 ^ n6465;
  assign n6482 = n3285 & ~n5564;
  assign n6483 = ~n1097 & n3435;
  assign n6484 = ~n1414 & ~n3440;
  assign n6485 = ~n6483 & ~n6484;
  assign n6486 = ~n970 & n3437;
  assign n6487 = n6485 & ~n6486;
  assign n6488 = ~n6482 & n6487;
  assign n6489 = n6488 ^ x26;
  assign n6478 = x28 & ~n1319;
  assign n6475 = x26 & x27;
  assign n6476 = n6475 ^ x28;
  assign n6477 = ~n1319 & n6476;
  assign n6479 = n6478 ^ n6477;
  assign n6480 = ~n6175 & ~n6479;
  assign n6481 = n6480 ^ n6478;
  assign n6490 = n6489 ^ n6481;
  assign n6491 = n3285 & ~n5579;
  assign n6492 = ~n1097 & n3437;
  assign n6493 = ~n1414 & n3435;
  assign n6494 = ~n6492 & ~n6493;
  assign n6495 = ~n1208 & ~n3440;
  assign n6496 = n6494 & ~n6495;
  assign n6497 = ~n6491 & n6496;
  assign n6498 = n6497 ^ x26;
  assign n6499 = n643 & n5630;
  assign n6500 = n735 & ~n1414;
  assign n6501 = ~n6499 & n6500;
  assign n6502 = ~n1319 & ~n3440;
  assign n6503 = ~n6501 & ~n6502;
  assign n6504 = n3285 & n5634;
  assign n6505 = ~n3435 & ~n6504;
  assign n6506 = ~n1208 & ~n6505;
  assign n6507 = n6503 & ~n6506;
  assign n6508 = n735 & ~n1208;
  assign n6509 = ~n735 & ~n3435;
  assign n6510 = ~n1319 & ~n6509;
  assign n6511 = ~n6508 & ~n6510;
  assign n6512 = x26 & n6511;
  assign n6513 = n6507 & n6512;
  assign n6514 = n42 & ~n1319;
  assign n6515 = ~n6513 & ~n6514;
  assign n6516 = ~n6498 & ~n6515;
  assign n6517 = n6516 ^ n6481;
  assign n6518 = n6490 & n6517;
  assign n6519 = n6518 ^ n6489;
  assign n6520 = n6519 ^ n6473;
  assign n6521 = ~n6474 & n6520;
  assign n6522 = n6521 ^ n6519;
  assign n6523 = n6522 ^ n6454;
  assign n6524 = ~n6463 & n6523;
  assign n6525 = n6524 ^ n6522;
  assign n6526 = n6525 ^ n6447;
  assign n6527 = ~n6448 & n6526;
  assign n6528 = n6527 ^ n6525;
  assign n6529 = n6528 ^ n6437;
  assign n6530 = ~n6438 & n6529;
  assign n6531 = n6530 ^ n6528;
  assign n6532 = n6531 ^ n6425;
  assign n6533 = ~n6426 & n6532;
  assign n6534 = n6533 ^ n6531;
  assign n6535 = n6534 ^ n6411;
  assign n6536 = ~n6412 & n6535;
  assign n6537 = n6536 ^ n6534;
  assign n6538 = n6537 ^ n6401;
  assign n6539 = n6402 & ~n6538;
  assign n6540 = n6539 ^ n6537;
  assign n6541 = n6540 ^ n6391;
  assign n6542 = ~n6392 & n6541;
  assign n6543 = n6542 ^ n6540;
  assign n6544 = n6543 ^ n6381;
  assign n6545 = ~n6382 & n6544;
  assign n6546 = n6545 ^ n6543;
  assign n6547 = n6546 ^ n6371;
  assign n6548 = n6372 & ~n6547;
  assign n6549 = n6548 ^ n6546;
  assign n6550 = n6549 ^ n6361;
  assign n6551 = ~n6362 & n6550;
  assign n6552 = n6551 ^ n6549;
  assign n6553 = n6552 ^ n6351;
  assign n6554 = n6352 & ~n6553;
  assign n6555 = n6554 ^ n6552;
  assign n6817 = n6564 ^ n6555;
  assign n6818 = n6565 & ~n6817;
  assign n6819 = n6818 ^ n6555;
  assign n7146 = n6836 ^ n6819;
  assign n7147 = ~n6837 & ~n7146;
  assign n7148 = n7147 ^ n6819;
  assign n7159 = n7158 ^ n7148;
  assign n6838 = n6837 ^ n6819;
  assign n6566 = n6565 ^ n6555;
  assign n6329 = ~n3974 & n5796;
  assign n6330 = ~n2954 & ~n5746;
  assign n6331 = ~n3037 & n5752;
  assign n6332 = ~n6330 & ~n6331;
  assign n6333 = ~n3098 & n5801;
  assign n6334 = n6332 & ~n6333;
  assign n6335 = ~n6329 & n6334;
  assign n6336 = ~x14 & ~n6335;
  assign n6337 = ~n3974 & n5801;
  assign n6338 = ~n3098 & n5796;
  assign n6339 = x14 & ~n6338;
  assign n6340 = n6332 & n6339;
  assign n6341 = ~n6337 & n6340;
  assign n6342 = ~n6336 & ~n6341;
  assign n6567 = n6566 ^ n6342;
  assign n6582 = n6552 ^ n6352;
  assign n6568 = ~n3777 & n5796;
  assign n6569 = ~n368 & n5752;
  assign n6570 = ~n3037 & ~n5746;
  assign n6571 = ~n6569 & ~n6570;
  assign n6572 = ~n2954 & n5801;
  assign n6573 = n6571 & ~n6572;
  assign n6574 = ~n6568 & n6573;
  assign n6575 = ~x14 & ~n6574;
  assign n6576 = ~n3777 & n5801;
  assign n6577 = ~n2954 & n5796;
  assign n6578 = x14 & ~n6577;
  assign n6579 = n6571 & n6578;
  assign n6580 = ~n6576 & n6579;
  assign n6581 = ~n6575 & ~n6580;
  assign n6583 = n6582 ^ n6581;
  assign n6592 = n6549 ^ n6362;
  assign n6584 = ~n4466 & n4963;
  assign n6585 = ~n2718 & n4976;
  assign n6586 = ~n2786 & n4970;
  assign n6587 = ~n2861 & n4972;
  assign n6588 = ~n6586 & ~n6587;
  assign n6589 = ~n6585 & n6588;
  assign n6590 = ~n6584 & n6589;
  assign n6591 = n6590 ^ x17;
  assign n6593 = n6592 ^ n6591;
  assign n6602 = n6546 ^ n6372;
  assign n6594 = ~n4312 & n4673;
  assign n6595 = ~n2482 & ~n4681;
  assign n6596 = ~n2574 & n4688;
  assign n6597 = ~n6595 & ~n6596;
  assign n6598 = ~n2612 & n4685;
  assign n6599 = n6597 & ~n6598;
  assign n6600 = ~n6594 & n6599;
  assign n6601 = n6600 ^ x20;
  assign n6603 = n6602 ^ n6601;
  assign n6612 = n6543 ^ n6382;
  assign n6604 = ~n4323 & n4478;
  assign n6605 = ~n2357 & n4487;
  assign n6606 = ~n2247 & n4484;
  assign n6607 = ~n6605 & ~n6606;
  assign n6608 = ~n2175 & n4480;
  assign n6609 = n6607 & ~n6608;
  assign n6610 = ~n6604 & n6609;
  assign n6611 = n6610 ^ x23;
  assign n6613 = n6612 ^ n6611;
  assign n6622 = n6540 ^ n6392;
  assign n6614 = ~n4253 & n4478;
  assign n6615 = ~n2065 & n4480;
  assign n6616 = ~n2175 & n4484;
  assign n6617 = ~n6615 & ~n6616;
  assign n6618 = ~n2247 & n4487;
  assign n6619 = n6617 & ~n6618;
  assign n6620 = ~n6614 & n6619;
  assign n6621 = n6620 ^ x23;
  assign n6623 = n6622 ^ n6621;
  assign n6632 = n6537 ^ n6402;
  assign n6624 = n4478 & ~n4507;
  assign n6625 = ~n2065 & n4484;
  assign n6626 = ~n1974 & n4480;
  assign n6627 = ~n6625 & ~n6626;
  assign n6628 = ~n2175 & n4487;
  assign n6629 = n6627 & ~n6628;
  assign n6630 = ~n6624 & n6629;
  assign n6631 = n6630 ^ x23;
  assign n6633 = n6632 ^ n6631;
  assign n6642 = n6534 ^ n6412;
  assign n6634 = n4478 & ~n5167;
  assign n6635 = ~n1878 & n4480;
  assign n6636 = ~n2065 & n4487;
  assign n6637 = ~n6635 & ~n6636;
  assign n6638 = ~n1974 & n4484;
  assign n6639 = n6637 & ~n6638;
  assign n6640 = ~n6634 & n6639;
  assign n6641 = n6640 ^ x23;
  assign n6643 = n6642 ^ n6641;
  assign n6652 = n6531 ^ n6426;
  assign n6644 = n4478 & ~n5923;
  assign n6645 = ~n1878 & n4484;
  assign n6646 = ~n1974 & n4487;
  assign n6647 = ~n6645 & ~n6646;
  assign n6648 = ~n1798 & n4480;
  assign n6649 = n6647 & ~n6648;
  assign n6650 = ~n6644 & n6649;
  assign n6651 = n6650 ^ x23;
  assign n6653 = n6652 ^ n6651;
  assign n6662 = n6528 ^ n6438;
  assign n6654 = n4478 & ~n5371;
  assign n6655 = ~n1798 & n4484;
  assign n6656 = ~n1726 & n4480;
  assign n6657 = ~n6655 & ~n6656;
  assign n6658 = ~n1878 & n4487;
  assign n6659 = n6657 & ~n6658;
  assign n6660 = ~n6654 & n6659;
  assign n6661 = n6660 ^ x23;
  assign n6663 = n6662 ^ n6661;
  assign n6672 = n6525 ^ n6448;
  assign n6664 = n4478 & ~n5351;
  assign n6665 = ~n1726 & n4484;
  assign n6666 = ~n1638 & n4480;
  assign n6667 = ~n6665 & ~n6666;
  assign n6668 = ~n1798 & n4487;
  assign n6669 = n6667 & ~n6668;
  assign n6670 = ~n6664 & n6669;
  assign n6671 = n6670 ^ x23;
  assign n6673 = n6672 ^ n6671;
  assign n6682 = n6522 ^ n6463;
  assign n6674 = n4478 & ~n5703;
  assign n6675 = ~n1726 & n4487;
  assign n6676 = ~n1638 & n4484;
  assign n6677 = ~n6675 & ~n6676;
  assign n6678 = ~n1544 & n4480;
  assign n6679 = n6677 & ~n6678;
  assign n6680 = ~n6674 & n6679;
  assign n6681 = n6680 ^ x23;
  assign n6683 = n6682 ^ n6681;
  assign n6692 = n6519 ^ n6474;
  assign n6684 = n4478 & ~n5069;
  assign n6685 = ~n734 & n4480;
  assign n6686 = ~n1544 & n4484;
  assign n6687 = ~n6685 & ~n6686;
  assign n6688 = ~n1638 & n4487;
  assign n6689 = n6687 & ~n6688;
  assign n6690 = ~n6684 & n6689;
  assign n6691 = n6690 ^ x23;
  assign n6693 = n6692 ^ n6691;
  assign n6695 = n4478 & ~n5416;
  assign n6696 = ~n882 & n4480;
  assign n6697 = ~n734 & n4484;
  assign n6698 = ~n1544 & n4487;
  assign n6699 = ~n6697 & ~n6698;
  assign n6700 = ~n6696 & n6699;
  assign n6701 = ~n6695 & n6700;
  assign n6702 = n6701 ^ x23;
  assign n6694 = n6516 ^ n6490;
  assign n6703 = n6702 ^ n6694;
  assign n6761 = n6514 ^ n6513;
  assign n6762 = n6761 ^ n6498;
  assign n6706 = n4478 & ~n5481;
  assign n6707 = ~n882 & n4487;
  assign n6708 = ~n970 & n4484;
  assign n6709 = ~n6707 & ~n6708;
  assign n6710 = ~n1097 & n4480;
  assign n6711 = n6709 & ~n6710;
  assign n6712 = ~n6706 & n6711;
  assign n6713 = n6712 ^ x23;
  assign n6704 = x26 & ~n6511;
  assign n6705 = n6704 ^ n6507;
  assign n6714 = n6713 ^ n6705;
  assign n6721 = n4478 & ~n5564;
  assign n6722 = ~n1097 & n4484;
  assign n6723 = ~n1414 & n4480;
  assign n6724 = ~n6722 & ~n6723;
  assign n6725 = ~n970 & n4487;
  assign n6726 = n6724 & ~n6725;
  assign n6727 = ~n6721 & n6726;
  assign n6728 = n6727 ^ x23;
  assign n6717 = x25 & ~n1319;
  assign n6715 = ~n690 & n3434;
  assign n6716 = ~n1319 & n6715;
  assign n6718 = n6717 ^ n6716;
  assign n6719 = ~n6508 & ~n6718;
  assign n6720 = n6719 ^ n6717;
  assign n6729 = n6728 ^ n6720;
  assign n6730 = n4478 & ~n5579;
  assign n6731 = ~n1097 & n4487;
  assign n6732 = ~n1414 & n4484;
  assign n6733 = ~n6731 & ~n6732;
  assign n6734 = ~n1208 & n4480;
  assign n6735 = n6733 & ~n6734;
  assign n6736 = ~n6730 & n6735;
  assign n6737 = n6736 ^ x23;
  assign n6738 = n4477 & n5630;
  assign n6739 = ~n1414 & n4476;
  assign n6740 = ~n6738 & n6739;
  assign n6741 = ~n1319 & n4480;
  assign n6742 = ~n6740 & ~n6741;
  assign n6743 = n4478 & n5634;
  assign n6744 = ~n4484 & ~n6743;
  assign n6745 = ~n1208 & ~n6744;
  assign n6746 = n6742 & ~n6745;
  assign n6747 = ~n1208 & n4476;
  assign n6748 = n38 & ~n1319;
  assign n6749 = ~n6747 & ~n6748;
  assign n6750 = x23 & n6749;
  assign n6751 = n6746 & n6750;
  assign n6752 = n735 & ~n1319;
  assign n6753 = ~n6751 & ~n6752;
  assign n6754 = ~n6737 & ~n6753;
  assign n6755 = n6754 ^ n6720;
  assign n6756 = n6729 & n6755;
  assign n6757 = n6756 ^ n6728;
  assign n6758 = n6757 ^ n6713;
  assign n6759 = ~n6714 & n6758;
  assign n6760 = n6759 ^ n6757;
  assign n6763 = n6762 ^ n6760;
  assign n6764 = n4478 & ~n5465;
  assign n6765 = ~n882 & n4484;
  assign n6766 = ~n734 & n4487;
  assign n6767 = ~n6765 & ~n6766;
  assign n6768 = ~n970 & n4480;
  assign n6769 = n6767 & ~n6768;
  assign n6770 = ~n6764 & n6769;
  assign n6771 = n6770 ^ x23;
  assign n6772 = n6771 ^ n6762;
  assign n6773 = n6763 & ~n6772;
  assign n6774 = n6773 ^ n6760;
  assign n6775 = n6774 ^ n6702;
  assign n6776 = n6703 & n6775;
  assign n6777 = n6776 ^ n6774;
  assign n6778 = n6777 ^ n6692;
  assign n6779 = ~n6693 & n6778;
  assign n6780 = n6779 ^ n6777;
  assign n6781 = n6780 ^ n6682;
  assign n6782 = ~n6683 & n6781;
  assign n6783 = n6782 ^ n6780;
  assign n6784 = n6783 ^ n6672;
  assign n6785 = ~n6673 & n6784;
  assign n6786 = n6785 ^ n6783;
  assign n6787 = n6786 ^ n6662;
  assign n6788 = ~n6663 & n6787;
  assign n6789 = n6788 ^ n6786;
  assign n6790 = n6789 ^ n6652;
  assign n6791 = ~n6653 & n6790;
  assign n6792 = n6791 ^ n6789;
  assign n6793 = n6792 ^ n6642;
  assign n6794 = ~n6643 & n6793;
  assign n6795 = n6794 ^ n6792;
  assign n6796 = n6795 ^ n6632;
  assign n6797 = n6633 & ~n6796;
  assign n6798 = n6797 ^ n6795;
  assign n6799 = n6798 ^ n6622;
  assign n6800 = ~n6623 & n6799;
  assign n6801 = n6800 ^ n6798;
  assign n6802 = n6801 ^ n6612;
  assign n6803 = ~n6613 & n6802;
  assign n6804 = n6803 ^ n6801;
  assign n6805 = n6804 ^ n6602;
  assign n6806 = n6603 & ~n6805;
  assign n6807 = n6806 ^ n6804;
  assign n6808 = n6807 ^ n6592;
  assign n6809 = ~n6593 & n6808;
  assign n6810 = n6809 ^ n6807;
  assign n6811 = n6810 ^ n6581;
  assign n6812 = ~n6583 & ~n6811;
  assign n6813 = n6812 ^ n6582;
  assign n6814 = n6813 ^ n6342;
  assign n6815 = ~n6567 & n6814;
  assign n6816 = n6815 ^ n6566;
  assign n6839 = n6838 ^ n6816;
  assign n6321 = ~n5770 & n5814;
  assign n6322 = ~n3270 & n5824;
  assign n6323 = ~n3351 & n5817;
  assign n6324 = ~n3404 & n6295;
  assign n6325 = ~n6323 & ~n6324;
  assign n6326 = ~n6322 & n6325;
  assign n6327 = ~n6321 & n6326;
  assign n6328 = n6327 ^ x11;
  assign n7143 = n6816 ^ n6328;
  assign n7144 = ~n6839 & n7143;
  assign n7145 = n7144 ^ n6838;
  assign n7160 = n7159 ^ n7145;
  assign n6304 = x8 ^ x7;
  assign n6305 = x6 ^ x5;
  assign n6306 = n6304 & n6305;
  assign n7139 = n6285 & n6306;
  assign n6311 = x5 & x6;
  assign n6312 = x7 & n6311;
  assign n6313 = ~x5 & ~x6;
  assign n6314 = ~x7 & n6313;
  assign n6315 = ~n6312 & ~n6314;
  assign n6316 = n6304 & ~n6315;
  assign n7140 = ~n3875 & n6316;
  assign n7141 = ~n7139 & ~n7140;
  assign n7142 = n7141 ^ x8;
  assign n7161 = n7160 ^ n7142;
  assign n6840 = n6839 ^ n6328;
  assign n6307 = n5758 & n6306;
  assign n6308 = x7 ^ x6;
  assign n6309 = ~n6305 & n6308;
  assign n6310 = ~n3875 & n6309;
  assign n6317 = ~n3431 & n6316;
  assign n6318 = ~n6310 & ~n6317;
  assign n6319 = ~n6307 & n6318;
  assign n6320 = n6319 ^ x8;
  assign n6841 = n6840 ^ n6320;
  assign n6850 = n6813 ^ n6567;
  assign n6842 = ~n3989 & n5814;
  assign n6843 = ~n3270 & n5817;
  assign n6844 = ~n3351 & n6295;
  assign n6845 = ~n3196 & n5824;
  assign n6846 = ~n6844 & ~n6845;
  assign n6847 = ~n6843 & n6846;
  assign n6848 = ~n6842 & n6847;
  assign n6849 = n6848 ^ x11;
  assign n6851 = n6850 ^ n6849;
  assign n6860 = n6810 ^ n6583;
  assign n6852 = ~n3271 & n5814;
  assign n6853 = ~n3098 & n5824;
  assign n6854 = ~n3196 & n5817;
  assign n6855 = ~n6853 & ~n6854;
  assign n6856 = ~n3270 & n6295;
  assign n6857 = n6855 & ~n6856;
  assign n6858 = ~n6852 & n6857;
  assign n6859 = n6858 ^ x11;
  assign n6861 = n6860 ^ n6859;
  assign n6876 = n6807 ^ n6593;
  assign n6862 = ~n3632 & n5796;
  assign n6863 = ~n566 & n5752;
  assign n6864 = ~n368 & ~n5746;
  assign n6865 = ~n6863 & ~n6864;
  assign n6866 = ~n3037 & n5801;
  assign n6867 = n6865 & ~n6866;
  assign n6868 = ~n6862 & n6867;
  assign n6869 = ~x14 & ~n6868;
  assign n6870 = ~n3632 & n5801;
  assign n6871 = ~n3037 & n5796;
  assign n6872 = x14 & ~n6871;
  assign n6873 = n6865 & n6872;
  assign n6874 = ~n6870 & n6873;
  assign n6875 = ~n6869 & ~n6874;
  assign n6877 = n6876 ^ n6875;
  assign n6886 = n6804 ^ n6603;
  assign n6878 = ~n4495 & n4963;
  assign n6879 = ~n2718 & n4972;
  assign n6880 = ~n2786 & n4976;
  assign n6881 = ~n2669 & n4970;
  assign n6882 = ~n6880 & ~n6881;
  assign n6883 = ~n6879 & n6882;
  assign n6884 = ~n6878 & n6883;
  assign n6885 = n6884 ^ x17;
  assign n6887 = n6886 ^ n6885;
  assign n6896 = n6801 ^ n6613;
  assign n6888 = n4333 & n4672;
  assign n6889 = n6888 ^ n2612;
  assign n6890 = n4671 & ~n6889;
  assign n6891 = ~n2482 & n4685;
  assign n6892 = ~n2423 & ~n4681;
  assign n6893 = ~n6891 & ~n6892;
  assign n6894 = ~n6890 & n6893;
  assign n6895 = n6894 ^ x20;
  assign n6897 = n6896 ^ n6895;
  assign n6906 = n6798 ^ n6623;
  assign n6898 = ~n4434 & n4673;
  assign n6899 = ~n2482 & n4688;
  assign n6900 = ~n2423 & n4685;
  assign n6901 = ~n6899 & ~n6900;
  assign n6902 = ~n2357 & ~n4681;
  assign n6903 = n6901 & ~n6902;
  assign n6904 = ~n6898 & n6903;
  assign n6905 = n6904 ^ x20;
  assign n6907 = n6906 ^ n6905;
  assign n6916 = n6795 ^ n6633;
  assign n6908 = ~n4293 & n4673;
  assign n6909 = ~n2357 & n4685;
  assign n6910 = ~n2247 & ~n4681;
  assign n6911 = ~n6909 & ~n6910;
  assign n6912 = ~n2423 & n4688;
  assign n6913 = n6911 & ~n6912;
  assign n6914 = ~n6908 & n6913;
  assign n6915 = n6914 ^ x20;
  assign n6917 = n6916 ^ n6915;
  assign n6926 = n6792 ^ n6643;
  assign n6918 = ~n4323 & n4673;
  assign n6919 = ~n2357 & n4688;
  assign n6920 = ~n2175 & ~n4681;
  assign n6921 = ~n6919 & ~n6920;
  assign n6922 = ~n2247 & n4685;
  assign n6923 = n6921 & ~n6922;
  assign n6924 = ~n6918 & n6923;
  assign n6925 = n6924 ^ x20;
  assign n6927 = n6926 ^ n6925;
  assign n6936 = n6789 ^ n6653;
  assign n6928 = ~n4253 & n4673;
  assign n6929 = ~n2065 & ~n4681;
  assign n6930 = ~n2175 & n4685;
  assign n6931 = ~n6929 & ~n6930;
  assign n6932 = ~n2247 & n4688;
  assign n6933 = n6931 & ~n6932;
  assign n6934 = ~n6928 & n6933;
  assign n6935 = n6934 ^ x20;
  assign n6937 = n6936 ^ n6935;
  assign n7096 = ~n4507 & n4673;
  assign n7097 = ~n2065 & n4685;
  assign n7098 = ~n2175 & n4688;
  assign n7099 = ~n7097 & ~n7098;
  assign n7100 = ~n1974 & ~n4681;
  assign n7101 = n7099 & ~n7100;
  assign n7102 = ~n7096 & n7101;
  assign n7103 = n7102 ^ x20;
  assign n6946 = n6783 ^ n6673;
  assign n6938 = n4673 & ~n5167;
  assign n6939 = ~n1878 & ~n4681;
  assign n6940 = ~n1974 & n4685;
  assign n6941 = ~n6939 & ~n6940;
  assign n6942 = ~n2065 & n4688;
  assign n6943 = n6941 & ~n6942;
  assign n6944 = ~n6938 & n6943;
  assign n6945 = n6944 ^ x20;
  assign n6947 = n6946 ^ n6945;
  assign n6956 = n6780 ^ n6683;
  assign n6948 = n4673 & ~n5923;
  assign n6949 = ~n1798 & ~n4681;
  assign n6950 = ~n1878 & n4685;
  assign n6951 = ~n6949 & ~n6950;
  assign n6952 = ~n1974 & n4688;
  assign n6953 = n6951 & ~n6952;
  assign n6954 = ~n6948 & n6953;
  assign n6955 = n6954 ^ x20;
  assign n6957 = n6956 ^ n6955;
  assign n6966 = n6777 ^ n6693;
  assign n6958 = n4673 & ~n5371;
  assign n6959 = ~n1798 & n4685;
  assign n6960 = ~n1726 & ~n4681;
  assign n6961 = ~n6959 & ~n6960;
  assign n6962 = ~n1878 & n4688;
  assign n6963 = n6961 & ~n6962;
  assign n6964 = ~n6958 & n6963;
  assign n6965 = n6964 ^ x20;
  assign n6967 = n6966 ^ n6965;
  assign n6976 = n6774 ^ n6703;
  assign n6968 = n4673 & ~n5351;
  assign n6969 = ~n1726 & n4685;
  assign n6970 = ~n1638 & ~n4681;
  assign n6971 = ~n6969 & ~n6970;
  assign n6972 = ~n1798 & n4688;
  assign n6973 = n6971 & ~n6972;
  assign n6974 = ~n6968 & n6973;
  assign n6975 = n6974 ^ x20;
  assign n6977 = n6976 ^ n6975;
  assign n6986 = n6771 ^ n6763;
  assign n6978 = n4673 & ~n5703;
  assign n6979 = ~n1726 & n4688;
  assign n6980 = ~n1638 & n4685;
  assign n6981 = ~n1544 & ~n4681;
  assign n6982 = ~n6980 & ~n6981;
  assign n6983 = ~n6979 & n6982;
  assign n6984 = ~n6978 & n6983;
  assign n6985 = n6984 ^ x20;
  assign n6987 = n6986 ^ n6985;
  assign n6989 = n4673 & ~n5069;
  assign n6990 = ~n734 & ~n4681;
  assign n6991 = ~n1544 & n4685;
  assign n6992 = ~n6990 & ~n6991;
  assign n6993 = ~n1638 & n4688;
  assign n6994 = n6992 & ~n6993;
  assign n6995 = ~n6989 & n6994;
  assign n6996 = n6995 ^ x20;
  assign n6988 = n6757 ^ n6714;
  assign n6997 = n6996 ^ n6988;
  assign n6999 = n4673 & ~n5416;
  assign n7000 = ~n882 & ~n4681;
  assign n7001 = ~n734 & n4685;
  assign n7002 = ~n1544 & n4688;
  assign n7003 = ~n7001 & ~n7002;
  assign n7004 = ~n7000 & n7003;
  assign n7005 = ~n6999 & n7004;
  assign n7006 = n7005 ^ x20;
  assign n6998 = n6754 ^ n6729;
  assign n7007 = n7006 ^ n6998;
  assign n7010 = n4673 & ~n5465;
  assign n7011 = ~n882 & n4685;
  assign n7012 = ~n970 & ~n4681;
  assign n7013 = ~n7011 & ~n7012;
  assign n7014 = ~n734 & n4688;
  assign n7015 = n7013 & ~n7014;
  assign n7016 = ~n7010 & n7015;
  assign n7017 = n7016 ^ x20;
  assign n7008 = n6752 ^ n6751;
  assign n7009 = n7008 ^ n6737;
  assign n7018 = n7017 ^ n7009;
  assign n7021 = n4673 & ~n5481;
  assign n7022 = ~n882 & n4688;
  assign n7023 = ~n970 & n4685;
  assign n7024 = ~n7022 & ~n7023;
  assign n7025 = ~n1097 & ~n4681;
  assign n7026 = n7024 & ~n7025;
  assign n7027 = ~n7021 & n7026;
  assign n7028 = n7027 ^ x20;
  assign n7019 = x23 & ~n6749;
  assign n7020 = n7019 ^ n6746;
  assign n7029 = n7028 ^ n7020;
  assign n7036 = n4673 & ~n5564;
  assign n7037 = ~n1097 & n4685;
  assign n7038 = ~n1414 & ~n4681;
  assign n7039 = ~n7037 & ~n7038;
  assign n7040 = ~n970 & n4688;
  assign n7041 = n7039 & ~n7040;
  assign n7042 = ~n7036 & n7041;
  assign n7043 = n7042 ^ x20;
  assign n7032 = x22 & ~n1319;
  assign n7030 = n36 ^ x22;
  assign n7031 = ~n1319 & n7030;
  assign n7033 = n7032 ^ n7031;
  assign n7034 = ~n6747 & ~n7033;
  assign n7035 = n7034 ^ n7032;
  assign n7044 = n7043 ^ n7035;
  assign n7045 = n4673 & ~n5579;
  assign n7046 = ~n1097 & n4688;
  assign n7047 = ~n1208 & ~n4681;
  assign n7048 = ~n7046 & ~n7047;
  assign n7049 = ~n1414 & n4685;
  assign n7050 = n7048 & ~n7049;
  assign n7051 = ~n7045 & n7050;
  assign n7052 = n7051 ^ x20;
  assign n7053 = n4672 & n5630;
  assign n7054 = ~n1414 & n4671;
  assign n7055 = ~n7053 & n7054;
  assign n7056 = ~n1319 & ~n4681;
  assign n7057 = ~n7055 & ~n7056;
  assign n7058 = n1208 & n1319;
  assign n7059 = ~n4671 & ~n4685;
  assign n7060 = ~n7058 & ~n7059;
  assign n7061 = x20 & ~n7060;
  assign n7062 = n7057 & n7061;
  assign n7063 = ~n1319 & n4476;
  assign n7064 = ~n7062 & ~n7063;
  assign n7065 = ~n7052 & ~n7064;
  assign n7066 = n7065 ^ n7035;
  assign n7067 = n7044 & n7066;
  assign n7068 = n7067 ^ n7043;
  assign n7069 = n7068 ^ n7028;
  assign n7070 = ~n7029 & n7069;
  assign n7071 = n7070 ^ n7068;
  assign n7072 = n7071 ^ n7017;
  assign n7073 = ~n7018 & n7072;
  assign n7074 = n7073 ^ n7071;
  assign n7075 = n7074 ^ n7006;
  assign n7076 = n7007 & n7075;
  assign n7077 = n7076 ^ n7074;
  assign n7078 = n7077 ^ n6996;
  assign n7079 = ~n6997 & n7078;
  assign n7080 = n7079 ^ n7077;
  assign n7081 = n7080 ^ n6986;
  assign n7082 = ~n6987 & n7081;
  assign n7083 = n7082 ^ n7080;
  assign n7084 = n7083 ^ n6976;
  assign n7085 = n6977 & ~n7084;
  assign n7086 = n7085 ^ n7083;
  assign n7087 = n7086 ^ n6966;
  assign n7088 = ~n6967 & n7087;
  assign n7089 = n7088 ^ n7086;
  assign n7090 = n7089 ^ n6956;
  assign n7091 = ~n6957 & n7090;
  assign n7092 = n7091 ^ n7089;
  assign n7093 = n7092 ^ n6946;
  assign n7094 = ~n6947 & n7093;
  assign n7095 = n7094 ^ n7092;
  assign n7104 = n7103 ^ n7095;
  assign n7105 = n6786 ^ n6663;
  assign n7106 = n7105 ^ n7103;
  assign n7107 = n7104 & ~n7106;
  assign n7108 = n7107 ^ n7095;
  assign n7109 = n7108 ^ n6936;
  assign n7110 = ~n6937 & n7109;
  assign n7111 = n7110 ^ n7108;
  assign n7112 = n7111 ^ n6926;
  assign n7113 = ~n6927 & n7112;
  assign n7114 = n7113 ^ n7111;
  assign n7115 = n7114 ^ n6916;
  assign n7116 = n6917 & ~n7115;
  assign n7117 = n7116 ^ n7114;
  assign n7118 = n7117 ^ n6906;
  assign n7119 = ~n6907 & n7118;
  assign n7120 = n7119 ^ n7117;
  assign n7121 = n7120 ^ n6896;
  assign n7122 = ~n6897 & n7121;
  assign n7123 = n7122 ^ n7120;
  assign n7124 = n7123 ^ n6886;
  assign n7125 = n6887 & ~n7124;
  assign n7126 = n7125 ^ n7123;
  assign n7127 = n7126 ^ n6876;
  assign n7128 = ~n6877 & n7127;
  assign n7129 = n7128 ^ n7126;
  assign n7130 = n7129 ^ n6860;
  assign n7131 = n6861 & ~n7130;
  assign n7132 = n7131 ^ n7129;
  assign n7133 = n7132 ^ n6850;
  assign n7134 = ~n6851 & n7133;
  assign n7135 = n7134 ^ n7132;
  assign n7136 = n7135 ^ n6840;
  assign n7137 = n6841 & ~n7136;
  assign n7138 = n7137 ^ n7135;
  assign n7162 = n7161 ^ n7138;
  assign n7163 = n7135 ^ n6841;
  assign n7164 = ~n3879 & n6306;
  assign n7165 = ~n3404 & n6316;
  assign n7166 = ~n3431 & n6309;
  assign n7167 = ~n7165 & ~n7166;
  assign n7168 = ~n6304 & n6305;
  assign n7169 = ~n3875 & n7168;
  assign n7170 = n7167 & ~n7169;
  assign n7171 = ~n7164 & n7170;
  assign n7172 = n7171 ^ x8;
  assign n7181 = n7129 ^ n6861;
  assign n7173 = ~n3432 & n6306;
  assign n7174 = ~n3404 & n6309;
  assign n7175 = ~n3351 & n6316;
  assign n7176 = ~n7174 & ~n7175;
  assign n7177 = ~n3431 & n7168;
  assign n7178 = n7176 & ~n7177;
  assign n7179 = ~n7173 & n7178;
  assign n7180 = n7179 ^ x8;
  assign n7182 = n7181 ^ n7180;
  assign n7191 = n7126 ^ n6877;
  assign n7183 = n3647 & n5814;
  assign n7184 = ~n2954 & n5824;
  assign n7185 = ~n3196 & n6295;
  assign n7186 = ~n7184 & ~n7185;
  assign n7187 = ~n3098 & n5817;
  assign n7188 = n7186 & ~n7187;
  assign n7189 = ~n7183 & n7188;
  assign n7190 = n7189 ^ x11;
  assign n7192 = n7191 ^ n7190;
  assign n7210 = n7123 ^ n6887;
  assign n7193 = n3748 & ~n6034;
  assign n7194 = n7193 ^ x13;
  assign n7195 = ~n368 & ~n7194;
  assign n7196 = n5748 & ~n7195;
  assign n7197 = ~x13 & ~n3748;
  assign n7198 = n368 & ~n7197;
  assign n7199 = ~n566 & ~n5746;
  assign n7200 = ~n2861 & n5752;
  assign n7201 = ~n7199 & ~n7200;
  assign n7202 = x14 & n7201;
  assign n7203 = n3748 & ~n7202;
  assign n7204 = n7198 & ~n7203;
  assign n7205 = n7196 & ~n7204;
  assign n7206 = ~n6048 & n7201;
  assign n7207 = ~n7205 & n7206;
  assign n7208 = ~x14 & ~n7201;
  assign n7209 = ~n7207 & ~n7208;
  assign n7211 = n7210 ^ n7209;
  assign n7220 = n7120 ^ n6897;
  assign n7212 = ~n4653 & n4963;
  assign n7213 = ~n2574 & n4970;
  assign n7214 = ~n2669 & n4976;
  assign n7215 = ~n2786 & n4972;
  assign n7216 = ~n7214 & ~n7215;
  assign n7217 = ~n7213 & n7216;
  assign n7218 = ~n7212 & n7217;
  assign n7219 = n7218 ^ x17;
  assign n7221 = n7220 ^ n7219;
  assign n7230 = n7117 ^ n6907;
  assign n7222 = ~n4453 & n4963;
  assign n7223 = ~n2574 & n4976;
  assign n7224 = ~n2669 & n4972;
  assign n7225 = ~n7223 & ~n7224;
  assign n7226 = ~n2612 & n4970;
  assign n7227 = n7225 & ~n7226;
  assign n7228 = ~n7222 & n7227;
  assign n7229 = n7228 ^ x17;
  assign n7231 = n7230 ^ n7229;
  assign n7240 = n7114 ^ n6917;
  assign n7232 = ~n4312 & n4963;
  assign n7233 = ~n2482 & n4970;
  assign n7234 = ~n2574 & n4972;
  assign n7235 = ~n7233 & ~n7234;
  assign n7236 = ~n2612 & n4976;
  assign n7237 = n7235 & ~n7236;
  assign n7238 = ~n7232 & n7237;
  assign n7239 = n7238 ^ x17;
  assign n7241 = n7240 ^ n7239;
  assign n7250 = n7111 ^ n6927;
  assign n7242 = ~n4334 & n4963;
  assign n7243 = ~n2482 & n4976;
  assign n7244 = ~n2423 & n4970;
  assign n7245 = ~n7243 & ~n7244;
  assign n7246 = ~n2612 & n4972;
  assign n7247 = n7245 & ~n7246;
  assign n7248 = ~n7242 & n7247;
  assign n7249 = n7248 ^ x17;
  assign n7251 = n7250 ^ n7249;
  assign n7260 = n7108 ^ n6937;
  assign n7252 = ~n4434 & n4963;
  assign n7253 = ~n2357 & n4970;
  assign n7254 = ~n2423 & n4976;
  assign n7255 = ~n7253 & ~n7254;
  assign n7256 = ~n2482 & n4972;
  assign n7257 = n7255 & ~n7256;
  assign n7258 = ~n7252 & n7257;
  assign n7259 = n7258 ^ x17;
  assign n7261 = n7260 ^ n7259;
  assign n7270 = n7105 ^ n7104;
  assign n7262 = ~n4293 & n4963;
  assign n7263 = ~n2357 & n4976;
  assign n7264 = ~n2423 & n4972;
  assign n7265 = ~n7263 & ~n7264;
  assign n7266 = ~n2247 & n4970;
  assign n7267 = n7265 & ~n7266;
  assign n7268 = ~n7262 & n7267;
  assign n7269 = n7268 ^ x17;
  assign n7271 = n7270 ^ n7269;
  assign n7272 = n7089 ^ n6957;
  assign n7281 = n7086 ^ n6967;
  assign n7273 = ~n4507 & n4963;
  assign n7274 = ~n2065 & n4976;
  assign n7275 = ~n1974 & n4970;
  assign n7276 = ~n7274 & ~n7275;
  assign n7277 = ~n2175 & n4972;
  assign n7278 = n7276 & ~n7277;
  assign n7279 = ~n7273 & n7278;
  assign n7280 = n7279 ^ x17;
  assign n7282 = n7281 ^ n7280;
  assign n7291 = n7083 ^ n6977;
  assign n7283 = n4963 & ~n5167;
  assign n7284 = ~n2065 & n4972;
  assign n7285 = ~n1878 & n4970;
  assign n7286 = ~n7284 & ~n7285;
  assign n7287 = ~n1974 & n4976;
  assign n7288 = n7286 & ~n7287;
  assign n7289 = ~n7283 & n7288;
  assign n7290 = n7289 ^ x17;
  assign n7292 = n7291 ^ n7290;
  assign n7301 = n7080 ^ n6987;
  assign n7293 = n4963 & ~n5923;
  assign n7294 = ~n1798 & n4970;
  assign n7295 = ~n1878 & n4976;
  assign n7296 = ~n7294 & ~n7295;
  assign n7297 = ~n1974 & n4972;
  assign n7298 = n7296 & ~n7297;
  assign n7299 = ~n7293 & n7298;
  assign n7300 = n7299 ^ x17;
  assign n7302 = n7301 ^ n7300;
  assign n7311 = n7077 ^ n6997;
  assign n7303 = n4963 & ~n5371;
  assign n7304 = ~n1798 & n4976;
  assign n7305 = ~n1726 & n4970;
  assign n7306 = ~n7304 & ~n7305;
  assign n7307 = ~n1878 & n4972;
  assign n7308 = n7306 & ~n7307;
  assign n7309 = ~n7303 & n7308;
  assign n7310 = n7309 ^ x17;
  assign n7312 = n7311 ^ n7310;
  assign n7321 = n7074 ^ n7007;
  assign n7313 = n4963 & ~n5351;
  assign n7314 = ~n1798 & n4972;
  assign n7315 = ~n1726 & n4976;
  assign n7316 = ~n7314 & ~n7315;
  assign n7317 = ~n1638 & n4970;
  assign n7318 = n7316 & ~n7317;
  assign n7319 = ~n7313 & n7318;
  assign n7320 = n7319 ^ x17;
  assign n7322 = n7321 ^ n7320;
  assign n7331 = n7071 ^ n7018;
  assign n7323 = n4963 & ~n5703;
  assign n7324 = ~n1726 & n4972;
  assign n7325 = ~n1638 & n4976;
  assign n7326 = ~n1544 & n4970;
  assign n7327 = ~n7325 & ~n7326;
  assign n7328 = ~n7324 & n7327;
  assign n7329 = ~n7323 & n7328;
  assign n7330 = n7329 ^ x17;
  assign n7332 = n7331 ^ n7330;
  assign n7341 = n7068 ^ n7029;
  assign n7333 = n4963 & ~n5069;
  assign n7334 = ~n1638 & n4972;
  assign n7335 = ~n1544 & n4976;
  assign n7336 = ~n7334 & ~n7335;
  assign n7337 = ~n734 & n4970;
  assign n7338 = n7336 & ~n7337;
  assign n7339 = ~n7333 & n7338;
  assign n7340 = n7339 ^ x17;
  assign n7342 = n7341 ^ n7340;
  assign n7344 = n4963 & ~n5416;
  assign n7345 = ~n882 & n4970;
  assign n7346 = ~n734 & n4976;
  assign n7347 = ~n1544 & n4972;
  assign n7348 = ~n7346 & ~n7347;
  assign n7349 = ~n7345 & n7348;
  assign n7350 = ~n7344 & n7349;
  assign n7351 = n7350 ^ x17;
  assign n7343 = n7065 ^ n7044;
  assign n7352 = n7351 ^ n7343;
  assign n7355 = n4963 & ~n5465;
  assign n7356 = ~n970 & n4970;
  assign n7357 = ~n734 & n4972;
  assign n7358 = ~n7356 & ~n7357;
  assign n7359 = ~n882 & n4976;
  assign n7360 = n7358 & ~n7359;
  assign n7361 = ~n7355 & n7360;
  assign n7362 = n7361 ^ x17;
  assign n7353 = n7063 ^ n7062;
  assign n7354 = n7353 ^ n7052;
  assign n7363 = n7362 ^ n7354;
  assign n7373 = n4963 & ~n5481;
  assign n7374 = ~n882 & n4972;
  assign n7375 = ~n1097 & n4970;
  assign n7376 = ~n7374 & ~n7375;
  assign n7377 = ~n970 & n4976;
  assign n7378 = n7376 & ~n7377;
  assign n7379 = ~n7373 & n7378;
  assign n7380 = n7379 ^ x17;
  assign n7368 = n4673 & n5634;
  assign n7369 = ~n4685 & ~n7368;
  assign n7370 = ~n1208 & ~n7369;
  assign n7371 = n7057 & ~n7370;
  assign n7364 = ~n1208 & n4671;
  assign n7365 = n1319 & ~n7364;
  assign n7366 = x20 & ~n7059;
  assign n7367 = ~n7365 & n7366;
  assign n7372 = n7371 ^ n7367;
  assign n7381 = n7380 ^ n7372;
  assign n7386 = n4963 & ~n5564;
  assign n7387 = ~n1097 & n4976;
  assign n7388 = ~n1414 & n4970;
  assign n7389 = ~n7387 & ~n7388;
  assign n7390 = ~n970 & n4972;
  assign n7391 = n7389 & ~n7390;
  assign n7392 = ~n7386 & n7391;
  assign n7393 = n7392 ^ x17;
  assign n7383 = ~n1319 & n4678;
  assign n7384 = ~n7364 & ~n7383;
  assign n7382 = x19 & ~n1319;
  assign n7385 = n7384 ^ n7382;
  assign n7394 = n7393 ^ n7385;
  assign n7395 = n4963 & ~n5579;
  assign n7396 = ~n1097 & n4972;
  assign n7397 = ~n1414 & n4976;
  assign n7398 = ~n7396 & ~n7397;
  assign n7399 = ~n1208 & n4970;
  assign n7400 = n7398 & ~n7399;
  assign n7401 = ~n7395 & n7400;
  assign n7402 = n7401 ^ x17;
  assign n7403 = n4963 & n5634;
  assign n7404 = ~n4976 & ~n7403;
  assign n7405 = ~n1208 & ~n7404;
  assign n7406 = ~n1414 & n4963;
  assign n7407 = ~n4970 & ~n7406;
  assign n7408 = ~n1319 & ~n7407;
  assign n7409 = ~n1208 & n4962;
  assign n7410 = ~n1414 & n4961;
  assign n7411 = ~n7409 & n7410;
  assign n7412 = ~n7408 & ~n7411;
  assign n7413 = ~n7405 & n7412;
  assign n7414 = ~n1208 & n4961;
  assign n7415 = ~n1319 & n4969;
  assign n7416 = ~n7414 & ~n7415;
  assign n7417 = x17 & n7416;
  assign n7418 = n7413 & n7417;
  assign n7419 = ~n1319 & n4671;
  assign n7420 = ~n7418 & ~n7419;
  assign n7421 = ~n7402 & ~n7420;
  assign n7422 = n7421 ^ n7385;
  assign n7423 = n7394 & n7422;
  assign n7424 = n7423 ^ n7393;
  assign n7425 = n7424 ^ n7380;
  assign n7426 = ~n7381 & n7425;
  assign n7427 = n7426 ^ n7424;
  assign n7428 = n7427 ^ n7362;
  assign n7429 = ~n7363 & n7428;
  assign n7430 = n7429 ^ n7427;
  assign n7431 = n7430 ^ n7351;
  assign n7432 = n7352 & n7431;
  assign n7433 = n7432 ^ n7430;
  assign n7434 = n7433 ^ n7341;
  assign n7435 = ~n7342 & n7434;
  assign n7436 = n7435 ^ n7433;
  assign n7437 = n7436 ^ n7331;
  assign n7438 = ~n7332 & n7437;
  assign n7439 = n7438 ^ n7436;
  assign n7440 = n7439 ^ n7321;
  assign n7441 = n7322 & ~n7440;
  assign n7442 = n7441 ^ n7439;
  assign n7443 = n7442 ^ n7311;
  assign n7444 = ~n7312 & n7443;
  assign n7445 = n7444 ^ n7442;
  assign n7446 = n7445 ^ n7301;
  assign n7447 = ~n7302 & n7446;
  assign n7448 = n7447 ^ n7445;
  assign n7449 = n7448 ^ n7291;
  assign n7450 = n7292 & ~n7449;
  assign n7451 = n7450 ^ n7448;
  assign n7452 = n7451 ^ n7281;
  assign n7453 = ~n7282 & n7452;
  assign n7454 = n7453 ^ n7451;
  assign n7455 = n7272 & n7454;
  assign n7456 = n7092 ^ n6947;
  assign n7457 = ~n7455 & ~n7456;
  assign n7458 = ~n4323 & n4963;
  assign n7459 = ~n2357 & n4972;
  assign n7460 = ~n2247 & n4976;
  assign n7461 = ~n7459 & ~n7460;
  assign n7462 = ~n2175 & n4970;
  assign n7463 = n7461 & ~n7462;
  assign n7464 = ~n7458 & n7463;
  assign n7465 = n7464 ^ x17;
  assign n7466 = ~n7457 & n7465;
  assign n7467 = ~n7272 & ~n7454;
  assign n7468 = ~n4253 & n4963;
  assign n7469 = ~n2065 & n4970;
  assign n7470 = ~n2247 & n4972;
  assign n7471 = ~n7469 & ~n7470;
  assign n7472 = ~n2175 & n4976;
  assign n7473 = n7471 & ~n7472;
  assign n7474 = ~n7468 & n7473;
  assign n7475 = n7474 ^ x17;
  assign n7476 = n7474 ^ n7464;
  assign n7477 = ~n7456 & n7476;
  assign n7478 = n7475 & n7477;
  assign n7479 = n7478 ^ n7475;
  assign n7480 = ~n7467 & n7479;
  assign n7481 = n7455 & n7456;
  assign n7482 = ~n7480 & ~n7481;
  assign n7483 = ~n7466 & n7482;
  assign n7484 = n7483 ^ n7270;
  assign n7485 = ~n7271 & ~n7484;
  assign n7486 = n7485 ^ n7483;
  assign n7487 = n7486 ^ n7260;
  assign n7488 = ~n7261 & ~n7487;
  assign n7489 = n7488 ^ n7486;
  assign n7490 = n7489 ^ n7250;
  assign n7491 = ~n7251 & ~n7490;
  assign n7492 = n7491 ^ n7489;
  assign n7493 = n7492 ^ n7240;
  assign n7494 = n7241 & n7493;
  assign n7495 = n7494 ^ n7492;
  assign n7496 = n7495 ^ n7230;
  assign n7497 = ~n7231 & ~n7496;
  assign n7498 = n7497 ^ n7495;
  assign n7499 = n7498 ^ n7220;
  assign n7500 = ~n7221 & ~n7499;
  assign n7501 = n7500 ^ n7498;
  assign n7502 = n7501 ^ n7210;
  assign n7503 = n7211 & n7502;
  assign n7504 = n7503 ^ n7501;
  assign n7505 = n7504 ^ n7191;
  assign n7506 = ~n7192 & ~n7505;
  assign n7507 = n7506 ^ n7504;
  assign n7508 = n7507 ^ n7180;
  assign n7509 = ~n7182 & n7508;
  assign n7510 = n7509 ^ n7181;
  assign n7511 = ~n7172 & n7510;
  assign n7512 = ~n7163 & ~n7511;
  assign n7574 = n7498 ^ n7221;
  assign n7557 = n566 & ~n3665;
  assign n7558 = x14 & n7557;
  assign n7559 = x14 & ~n5748;
  assign n7560 = n566 ^ x13;
  assign n7561 = n5748 & ~n7560;
  assign n7562 = n3665 & n7561;
  assign n7563 = ~n7559 & ~n7562;
  assign n7564 = ~n7558 & n7563;
  assign n7565 = ~n2718 & n5752;
  assign n7566 = ~n2861 & ~n5746;
  assign n7567 = ~n7565 & ~n7566;
  assign n7568 = ~n7564 & n7567;
  assign n7569 = ~n566 & n5748;
  assign n7570 = ~n3665 & n7569;
  assign n7571 = n7567 & ~n7570;
  assign n7572 = ~x14 & ~n7571;
  assign n7573 = ~n7568 & ~n7572;
  assign n7575 = n7574 ^ n7573;
  assign n7593 = n7495 ^ n7231;
  assign n7576 = ~n4466 & n6033;
  assign n7577 = ~n2718 & ~n5746;
  assign n7578 = ~n2786 & n5752;
  assign n7579 = ~n7577 & ~n7578;
  assign n7580 = x14 & n7579;
  assign n7581 = n2861 & n7580;
  assign n7582 = x13 & ~n7581;
  assign n7583 = ~n7576 & n7582;
  assign n7584 = n4466 & n7580;
  assign n7585 = ~n2861 & n6033;
  assign n7586 = ~x13 & ~n7585;
  assign n7587 = ~n7584 & n7586;
  assign n7588 = ~n7583 & ~n7587;
  assign n7589 = n7559 ^ x14;
  assign n7590 = n7579 & ~n7589;
  assign n7591 = n7590 ^ x14;
  assign n7592 = ~n7588 & n7591;
  assign n7594 = n7593 ^ n7592;
  assign n7609 = n7492 ^ n7241;
  assign n7595 = ~n4495 & n5796;
  assign n7596 = ~n2669 & n5752;
  assign n7597 = ~n2786 & ~n5746;
  assign n7598 = ~n7596 & ~n7597;
  assign n7599 = ~n2718 & n5801;
  assign n7600 = n7598 & ~n7599;
  assign n7601 = ~n7595 & n7600;
  assign n7602 = ~x14 & ~n7601;
  assign n7603 = ~n4495 & n5801;
  assign n7604 = x14 & n7598;
  assign n7605 = ~n2718 & n5796;
  assign n7606 = n7604 & ~n7605;
  assign n7607 = ~n7603 & n7606;
  assign n7608 = ~n7602 & ~n7607;
  assign n7610 = n7609 ^ n7608;
  assign n7620 = n7489 ^ n7251;
  assign n7611 = n4653 & n5749;
  assign n7612 = n2786 & ~n5749;
  assign n7613 = n5748 & ~n7612;
  assign n7614 = ~n7611 & n7613;
  assign n7615 = ~n2574 & n5752;
  assign n7616 = ~n2669 & ~n5746;
  assign n7617 = ~n7615 & ~n7616;
  assign n7618 = ~n7614 & n7617;
  assign n7619 = n7618 ^ x14;
  assign n7621 = n7620 ^ n7619;
  assign n7636 = n7486 ^ n7261;
  assign n7622 = ~n4453 & n5801;
  assign n7623 = ~n2612 & n5752;
  assign n7624 = ~n2574 & ~n5746;
  assign n7625 = ~n7623 & ~n7624;
  assign n7626 = ~n2669 & n5796;
  assign n7627 = n7625 & ~n7626;
  assign n7628 = ~n7622 & n7627;
  assign n7629 = x14 & ~n7628;
  assign n7630 = ~n4453 & n5796;
  assign n7631 = ~n2669 & n5801;
  assign n7632 = ~x14 & ~n7631;
  assign n7633 = n7625 & n7632;
  assign n7634 = ~n7630 & n7633;
  assign n7635 = ~n7629 & ~n7634;
  assign n7637 = n7636 ^ n7635;
  assign n7646 = n7483 ^ n7271;
  assign n7638 = n4311 & n5749;
  assign n7639 = n7638 ^ n2574;
  assign n7640 = n5748 & ~n7639;
  assign n7641 = ~n2482 & n5752;
  assign n7642 = ~n2612 & ~n5746;
  assign n7643 = ~n7641 & ~n7642;
  assign n7644 = ~n7640 & n7643;
  assign n7645 = n7644 ^ x14;
  assign n7647 = n7646 ^ n7645;
  assign n7669 = n7464 ^ n7456;
  assign n7664 = n7454 ^ n7272;
  assign n7665 = n7272 ^ x17;
  assign n7666 = n7665 ^ n7474;
  assign n7667 = ~n7664 & n7666;
  assign n7668 = n7667 ^ n7474;
  assign n7670 = n7669 ^ n7668;
  assign n7648 = n2612 & ~n4333;
  assign n7649 = ~x14 & n7648;
  assign n7650 = n2612 ^ x13;
  assign n7651 = n5748 & n7650;
  assign n7652 = n4333 & n7651;
  assign n7653 = ~n6048 & ~n7652;
  assign n7654 = ~n7649 & n7653;
  assign n7655 = ~n2423 & n5752;
  assign n7656 = ~n2482 & ~n5746;
  assign n7657 = ~n7655 & ~n7656;
  assign n7658 = ~n7654 & n7657;
  assign n7659 = ~n2612 & n5748;
  assign n7660 = ~n4333 & n7659;
  assign n7661 = n7657 & ~n7660;
  assign n7662 = x14 & ~n7661;
  assign n7663 = ~n7658 & ~n7662;
  assign n7671 = n7670 ^ n7663;
  assign n7686 = n7664 ^ n7475;
  assign n7672 = ~n4434 & n5796;
  assign n7673 = ~n2357 & n5752;
  assign n7674 = ~n2423 & ~n5746;
  assign n7675 = ~n7673 & ~n7674;
  assign n7676 = ~n2482 & n5801;
  assign n7677 = n7675 & ~n7676;
  assign n7678 = ~n7672 & n7677;
  assign n7679 = ~x14 & ~n7678;
  assign n7680 = ~n4434 & n5801;
  assign n7681 = ~n2482 & n5796;
  assign n7682 = x14 & ~n7681;
  assign n7683 = n7675 & n7682;
  assign n7684 = ~n7680 & n7683;
  assign n7685 = ~n7679 & ~n7684;
  assign n7687 = n7686 ^ n7685;
  assign n7702 = n7451 ^ n7282;
  assign n7688 = ~n4293 & n5796;
  assign n7689 = ~n2357 & ~n5746;
  assign n7690 = ~n2247 & n5752;
  assign n7691 = ~n7689 & ~n7690;
  assign n7692 = ~n2423 & n5801;
  assign n7693 = n7691 & ~n7692;
  assign n7694 = ~n7688 & n7693;
  assign n7695 = ~x14 & ~n7694;
  assign n7696 = ~n4293 & n5801;
  assign n7697 = ~n2423 & n5796;
  assign n7698 = x14 & ~n7697;
  assign n7699 = n7691 & n7698;
  assign n7700 = ~n7696 & n7699;
  assign n7701 = ~n7695 & ~n7700;
  assign n7703 = n7702 ^ n7701;
  assign n7720 = n7448 ^ n7292;
  assign n7704 = n2357 & ~n4322;
  assign n7705 = x14 & n7704;
  assign n7706 = n2357 ^ x13;
  assign n7707 = n5748 & ~n7706;
  assign n7708 = n4322 & n7707;
  assign n7709 = ~n7559 & ~n7708;
  assign n7710 = ~n7705 & n7709;
  assign n7711 = ~n2175 & n5752;
  assign n7712 = ~n2247 & ~n5746;
  assign n7713 = ~n7711 & ~n7712;
  assign n7714 = ~n7710 & n7713;
  assign n7715 = ~n2357 & n5748;
  assign n7716 = ~n4322 & n7715;
  assign n7717 = n7713 & ~n7716;
  assign n7718 = ~x14 & ~n7717;
  assign n7719 = ~n7714 & ~n7718;
  assign n7721 = n7720 ^ n7719;
  assign n7731 = n7445 ^ n7302;
  assign n7722 = n4253 & n5749;
  assign n7723 = n2247 & ~n5749;
  assign n7724 = n5748 & ~n7723;
  assign n7725 = ~n7722 & n7724;
  assign n7726 = ~n2175 & ~n5746;
  assign n7727 = ~n2065 & n5752;
  assign n7728 = ~n7726 & ~n7727;
  assign n7729 = ~n7725 & n7728;
  assign n7730 = n7729 ^ x14;
  assign n7732 = n7731 ^ n7730;
  assign n7750 = n7442 ^ n7312;
  assign n7733 = ~n4506 & ~n6034;
  assign n7734 = n7733 ^ x13;
  assign n7735 = ~n2175 & ~n7734;
  assign n7736 = n5748 & ~n7735;
  assign n7737 = ~x13 & n4506;
  assign n7738 = n2175 & ~n7737;
  assign n7739 = ~n2065 & ~n5746;
  assign n7740 = ~n1974 & n5752;
  assign n7741 = ~n7739 & ~n7740;
  assign n7742 = x14 & n7741;
  assign n7743 = ~n4506 & ~n7742;
  assign n7744 = n7738 & ~n7743;
  assign n7745 = n7736 & ~n7744;
  assign n7746 = ~n6048 & n7741;
  assign n7747 = ~n7745 & n7746;
  assign n7748 = ~x14 & ~n7741;
  assign n7749 = ~n7747 & ~n7748;
  assign n7751 = n7750 ^ n7749;
  assign n7766 = n7439 ^ n7322;
  assign n7752 = ~n5167 & n5801;
  assign n7753 = ~n1878 & n5752;
  assign n7754 = ~n1974 & ~n5746;
  assign n7755 = ~n7753 & ~n7754;
  assign n7756 = ~n2065 & n5796;
  assign n7757 = n7755 & ~n7756;
  assign n7758 = ~n7752 & n7757;
  assign n7759 = x14 & ~n7758;
  assign n7760 = ~n5167 & n5796;
  assign n7761 = ~n2065 & n5801;
  assign n7762 = ~x14 & ~n7761;
  assign n7763 = n7755 & n7762;
  assign n7764 = ~n7760 & n7763;
  assign n7765 = ~n7759 & ~n7764;
  assign n7767 = n7766 ^ n7765;
  assign n7782 = n7436 ^ n7332;
  assign n7768 = n5796 & ~n5923;
  assign n7769 = ~n1798 & n5752;
  assign n7770 = ~n1878 & ~n5746;
  assign n7771 = ~n7769 & ~n7770;
  assign n7772 = ~n1974 & n5801;
  assign n7773 = n7771 & ~n7772;
  assign n7774 = ~n7768 & n7773;
  assign n7775 = ~x14 & ~n7774;
  assign n7776 = n5801 & ~n5923;
  assign n7777 = ~n1974 & n5796;
  assign n7778 = x14 & ~n7777;
  assign n7779 = n7771 & n7778;
  assign n7780 = ~n7776 & n7779;
  assign n7781 = ~n7775 & ~n7780;
  assign n7783 = n7782 ^ n7781;
  assign n7801 = n7433 ^ n7342;
  assign n7784 = ~n1798 & ~n5746;
  assign n7785 = ~n1726 & n5752;
  assign n7786 = ~n7784 & ~n7785;
  assign n7788 = x13 & n5023;
  assign n7789 = n1878 & ~n7788;
  assign n7790 = x14 & n7786;
  assign n7791 = ~n5023 & n7790;
  assign n7792 = n7789 & ~n7791;
  assign n7793 = ~n5023 & ~n6034;
  assign n7794 = n7793 ^ x13;
  assign n7795 = ~n1878 & n7794;
  assign n7796 = ~n7792 & ~n7795;
  assign n7787 = n7786 ^ x14;
  assign n7797 = n7796 ^ n7787;
  assign n7798 = n7786 & ~n7797;
  assign n7799 = n5748 & n7798;
  assign n7800 = n7799 ^ n7787;
  assign n7802 = n7801 ^ n7800;
  assign n7811 = n7430 ^ n7352;
  assign n7803 = n5350 & n5749;
  assign n7804 = n7803 ^ n1798;
  assign n7805 = n5748 & ~n7804;
  assign n7806 = ~n1726 & ~n5746;
  assign n7807 = ~n1638 & n5752;
  assign n7808 = ~n7806 & ~n7807;
  assign n7809 = ~n7805 & n7808;
  assign n7810 = n7809 ^ x14;
  assign n7812 = n7811 ^ n7810;
  assign n7829 = n7427 ^ n7363;
  assign n7813 = ~n5703 & n6033;
  assign n7814 = ~n1544 & n5752;
  assign n7815 = ~n1638 & ~n5746;
  assign n7816 = ~n7814 & ~n7815;
  assign n7817 = x14 & n7816;
  assign n7818 = n1726 & n7817;
  assign n7819 = x13 & ~n7818;
  assign n7820 = ~n7813 & n7819;
  assign n7821 = n5703 & n7817;
  assign n7822 = ~n1726 & n6033;
  assign n7823 = ~x13 & ~n7822;
  assign n7824 = ~n7821 & n7823;
  assign n7825 = ~n7820 & ~n7824;
  assign n7826 = ~n7589 & n7816;
  assign n7827 = n7826 ^ x14;
  assign n7828 = ~n7825 & n7827;
  assign n7830 = n7829 ^ n7828;
  assign n7832 = ~n5069 & n5801;
  assign n7833 = ~n734 & n5752;
  assign n7834 = ~n1544 & ~n5746;
  assign n7835 = ~n7833 & ~n7834;
  assign n7836 = ~n1638 & n5796;
  assign n7837 = n7835 & ~n7836;
  assign n7838 = ~n7832 & n7837;
  assign n7839 = x14 & ~n7838;
  assign n7840 = ~n5069 & n5796;
  assign n7841 = ~n1638 & n5801;
  assign n7842 = ~x14 & ~n7841;
  assign n7843 = n7835 & n7842;
  assign n7844 = ~n7840 & n7843;
  assign n7845 = ~n7839 & ~n7844;
  assign n7831 = n7424 ^ n7381;
  assign n7846 = n7845 ^ n7831;
  assign n7848 = ~x14 & n1544;
  assign n7849 = ~n5415 & n7848;
  assign n7850 = ~n6048 & ~n7849;
  assign n7851 = n1544 ^ x13;
  assign n7852 = n5748 & n7851;
  assign n7853 = n5415 & n7852;
  assign n7854 = n7850 & ~n7853;
  assign n7855 = ~n882 & n5752;
  assign n7856 = ~n734 & ~n5746;
  assign n7857 = ~n7855 & ~n7856;
  assign n7858 = ~n7854 & n7857;
  assign n7859 = ~n1544 & ~n5415;
  assign n7860 = x14 & n5748;
  assign n7861 = n7859 & n7860;
  assign n7862 = x14 & ~n7857;
  assign n7863 = ~n7861 & ~n7862;
  assign n7864 = ~n7858 & n7863;
  assign n7847 = n7421 ^ n7394;
  assign n7865 = n7864 ^ n7847;
  assign n7868 = ~n5465 & n5796;
  assign n7869 = ~n970 & n5752;
  assign n7870 = ~n882 & ~n5746;
  assign n7871 = ~n7869 & ~n7870;
  assign n7872 = ~n734 & n5801;
  assign n7873 = n7871 & ~n7872;
  assign n7874 = ~n7868 & n7873;
  assign n7875 = ~x14 & ~n7874;
  assign n7876 = ~n5465 & n5801;
  assign n7877 = ~n734 & n5796;
  assign n7878 = x14 & ~n7877;
  assign n7879 = n7871 & n7878;
  assign n7880 = ~n7876 & n7879;
  assign n7881 = ~n7875 & ~n7880;
  assign n7866 = n7419 ^ n7418;
  assign n7867 = n7866 ^ n7402;
  assign n7882 = n7881 ^ n7867;
  assign n7885 = ~n5481 & n5796;
  assign n7886 = ~n1097 & n5752;
  assign n7887 = ~n970 & ~n5746;
  assign n7888 = ~n7886 & ~n7887;
  assign n7889 = ~n882 & n5801;
  assign n7890 = n7888 & ~n7889;
  assign n7891 = ~n7885 & n7890;
  assign n7892 = ~x14 & ~n7891;
  assign n7893 = ~n5481 & n5801;
  assign n7894 = ~n882 & n5796;
  assign n7895 = x14 & ~n7894;
  assign n7896 = n7888 & n7895;
  assign n7897 = ~n7893 & n7896;
  assign n7898 = ~n7892 & ~n7897;
  assign n7883 = x17 & ~n7416;
  assign n7884 = n7883 ^ n7413;
  assign n7899 = n7898 ^ n7884;
  assign n7900 = ~n5579 & n5801;
  assign n7901 = ~n1208 & n5752;
  assign n7902 = ~n1414 & ~n5746;
  assign n7903 = ~n7901 & ~n7902;
  assign n7904 = ~n1097 & n5796;
  assign n7905 = n7903 & ~n7904;
  assign n7906 = ~n7900 & n7905;
  assign n7907 = x14 & ~n7906;
  assign n7908 = ~n5579 & n5796;
  assign n7909 = ~n1097 & n5801;
  assign n7910 = ~x14 & ~n7909;
  assign n7911 = n7903 & n7910;
  assign n7912 = ~n7908 & n7911;
  assign n7913 = ~n7907 & ~n7912;
  assign n7914 = n5630 & n5749;
  assign n7915 = n7914 ^ n1414;
  assign n7916 = n5748 & ~n7915;
  assign n7917 = ~n1208 & ~n5746;
  assign n7918 = ~n1319 & n5752;
  assign n7919 = ~n7917 & ~n7918;
  assign n7920 = ~n7916 & n7919;
  assign n7921 = ~n1319 & ~n5746;
  assign n7922 = ~n5748 & ~n7921;
  assign n7923 = ~n7058 & ~n7922;
  assign n7924 = x14 & ~n7923;
  assign n7925 = n7920 & n7924;
  assign n7926 = ~n1319 & n4961;
  assign n7927 = ~n7925 & ~n7926;
  assign n7928 = n7913 & ~n7927;
  assign n7929 = n970 ^ x13;
  assign n7930 = n5748 & n7929;
  assign n7931 = n5563 & n7930;
  assign n7932 = ~n6048 & ~n7931;
  assign n7933 = ~x14 & n970;
  assign n7934 = ~n5563 & n7933;
  assign n7935 = n7932 & ~n7934;
  assign n7936 = ~n1097 & ~n5746;
  assign n7937 = ~n1414 & n5752;
  assign n7938 = ~n7936 & ~n7937;
  assign n7939 = ~n7935 & n7938;
  assign n7940 = ~n970 & n5748;
  assign n7941 = ~n5564 & n7940;
  assign n7942 = n7938 & ~n7941;
  assign n7943 = x14 & ~n7942;
  assign n7944 = ~n7939 & ~n7943;
  assign n7945 = ~n7928 & ~n7944;
  assign n7947 = ~n1319 & n4967;
  assign n7948 = ~n7414 & ~n7947;
  assign n7946 = x16 & ~n1319;
  assign n7949 = n7948 ^ n7946;
  assign n7950 = n7928 & n7944;
  assign n7951 = n7949 & ~n7950;
  assign n7952 = ~n7945 & ~n7951;
  assign n7953 = n7952 ^ n7884;
  assign n7954 = n7899 & n7953;
  assign n7955 = n7954 ^ n7898;
  assign n7956 = n7955 ^ n7881;
  assign n7957 = ~n7882 & n7956;
  assign n7958 = n7957 ^ n7955;
  assign n7959 = n7958 ^ n7864;
  assign n7960 = ~n7865 & ~n7959;
  assign n7961 = n7960 ^ n7958;
  assign n7962 = n7961 ^ n7845;
  assign n7963 = n7846 & ~n7962;
  assign n7964 = n7963 ^ n7961;
  assign n7965 = n7964 ^ n7829;
  assign n7966 = ~n7830 & n7965;
  assign n7967 = n7966 ^ n7964;
  assign n7968 = n7967 ^ n7811;
  assign n7969 = n7812 & ~n7968;
  assign n7970 = n7969 ^ n7967;
  assign n7971 = n7970 ^ n7801;
  assign n7972 = ~n7802 & n7971;
  assign n7973 = n7972 ^ n7970;
  assign n7974 = n7973 ^ n7782;
  assign n7975 = ~n7783 & n7974;
  assign n7976 = n7975 ^ n7973;
  assign n7977 = n7976 ^ n7766;
  assign n7978 = ~n7767 & ~n7977;
  assign n7979 = n7978 ^ n7976;
  assign n7980 = n7979 ^ n7750;
  assign n7981 = ~n7751 & n7980;
  assign n7982 = n7981 ^ n7979;
  assign n7983 = n7982 ^ n7731;
  assign n7984 = ~n7732 & n7983;
  assign n7985 = n7984 ^ n7982;
  assign n7986 = n7985 ^ n7720;
  assign n7987 = n7721 & ~n7986;
  assign n7988 = n7987 ^ n7985;
  assign n7989 = n7988 ^ n7702;
  assign n7990 = ~n7703 & n7989;
  assign n7991 = n7990 ^ n7988;
  assign n7992 = n7991 ^ n7686;
  assign n7993 = ~n7687 & n7992;
  assign n7994 = n7993 ^ n7991;
  assign n7995 = n7994 ^ n7670;
  assign n7996 = n7671 & n7995;
  assign n7997 = n7996 ^ n7994;
  assign n7998 = n7997 ^ n7646;
  assign n7999 = n7647 & ~n7998;
  assign n8000 = n7999 ^ n7997;
  assign n8001 = n8000 ^ n7636;
  assign n8002 = ~n7637 & ~n8001;
  assign n8003 = n8002 ^ n8000;
  assign n8004 = n8003 ^ n7620;
  assign n8005 = n7621 & ~n8004;
  assign n8006 = n8005 ^ n8003;
  assign n8007 = n8006 ^ n7609;
  assign n8008 = ~n7610 & n8007;
  assign n8009 = n8008 ^ n8006;
  assign n8010 = n8009 ^ n7593;
  assign n8011 = n7594 & ~n8010;
  assign n8012 = n8011 ^ n8009;
  assign n8013 = n8012 ^ n7574;
  assign n8014 = n7575 & ~n8013;
  assign n8015 = n8014 ^ n8012;
  assign n7555 = n7501 ^ n7211;
  assign n7536 = ~x11 & n5812;
  assign n7537 = ~n3974 & n7536;
  assign n7538 = ~n2954 & n5817;
  assign n7539 = ~n3037 & n5824;
  assign n7540 = ~n7538 & ~n7539;
  assign n7541 = x11 & n7540;
  assign n7542 = n3098 & n7541;
  assign n7543 = x10 & ~n7542;
  assign n7544 = ~n7537 & n7543;
  assign n7545 = n3974 & n7541;
  assign n7546 = ~n3098 & n7536;
  assign n7547 = ~x10 & ~n7546;
  assign n7548 = ~n7545 & n7547;
  assign n7549 = ~n7544 & ~n7548;
  assign n7550 = x11 & ~n5812;
  assign n7551 = n7550 ^ x11;
  assign n7552 = n7540 & ~n7551;
  assign n7553 = n7552 ^ x11;
  assign n7554 = ~n7549 & n7553;
  assign n7556 = n7555 ^ n7554;
  assign n8417 = n8015 ^ n7556;
  assign n8409 = ~n3989 & n6306;
  assign n8410 = ~n3270 & n6309;
  assign n8411 = ~n3196 & n6316;
  assign n8412 = ~n3351 & n7168;
  assign n8413 = ~n8411 & ~n8412;
  assign n8414 = ~n8410 & n8413;
  assign n8415 = ~n8409 & n8414;
  assign n8416 = n8415 ^ x8;
  assign n8418 = n8417 ^ n8416;
  assign n8042 = n8012 ^ n7575;
  assign n8034 = ~n3777 & n5814;
  assign n8035 = ~n368 & n5824;
  assign n8036 = ~n3037 & n5817;
  assign n8037 = ~n8035 & ~n8036;
  assign n8038 = ~n2954 & n6295;
  assign n8039 = n8037 & ~n8038;
  assign n8040 = ~n8034 & n8039;
  assign n8041 = n8040 ^ x11;
  assign n8043 = n8042 ^ n8041;
  assign n8052 = n8009 ^ n7594;
  assign n8044 = ~n3632 & n5814;
  assign n8045 = ~n566 & n5824;
  assign n8046 = ~n368 & n5817;
  assign n8047 = ~n8045 & ~n8046;
  assign n8048 = ~n3037 & n6295;
  assign n8049 = n8047 & ~n8048;
  assign n8050 = ~n8044 & n8049;
  assign n8051 = n8050 ^ x11;
  assign n8053 = n8052 ^ n8051;
  assign n8062 = n8006 ^ n7610;
  assign n8054 = n3749 & n5814;
  assign n8055 = ~n566 & n5817;
  assign n8056 = ~n2861 & n5824;
  assign n8057 = ~n8055 & ~n8056;
  assign n8058 = ~n368 & n6295;
  assign n8059 = n8057 & ~n8058;
  assign n8060 = ~n8054 & n8059;
  assign n8061 = n8060 ^ x11;
  assign n8063 = n8062 ^ n8061;
  assign n8072 = n8003 ^ n7621;
  assign n8064 = ~n3666 & n5814;
  assign n8065 = ~n2718 & n5824;
  assign n8066 = ~n2861 & n5817;
  assign n8067 = ~n8065 & ~n8066;
  assign n8068 = ~n566 & n6295;
  assign n8069 = n8067 & ~n8068;
  assign n8070 = ~n8064 & n8069;
  assign n8071 = n8070 ^ x11;
  assign n8073 = n8072 ^ n8071;
  assign n8082 = n8000 ^ n7637;
  assign n8074 = ~n4466 & n5814;
  assign n8075 = ~n2718 & n5817;
  assign n8076 = ~n2861 & n6295;
  assign n8077 = ~n2786 & n5824;
  assign n8078 = ~n8076 & ~n8077;
  assign n8079 = ~n8075 & n8078;
  assign n8080 = ~n8074 & n8079;
  assign n8081 = n8080 ^ x11;
  assign n8083 = n8082 ^ n8081;
  assign n8092 = n7997 ^ n7647;
  assign n8084 = ~n4495 & n5814;
  assign n8085 = ~n2718 & n6295;
  assign n8086 = ~n2786 & n5817;
  assign n8087 = ~n2669 & n5824;
  assign n8088 = ~n8086 & ~n8087;
  assign n8089 = ~n8085 & n8088;
  assign n8090 = ~n8084 & n8089;
  assign n8091 = n8090 ^ x11;
  assign n8093 = n8092 ^ n8091;
  assign n8102 = n7994 ^ n7671;
  assign n8094 = ~n4653 & n5814;
  assign n8095 = ~n2574 & n5824;
  assign n8096 = ~n2669 & n5817;
  assign n8097 = ~n2786 & n6295;
  assign n8098 = ~n8096 & ~n8097;
  assign n8099 = ~n8095 & n8098;
  assign n8100 = ~n8094 & n8099;
  assign n8101 = n8100 ^ x11;
  assign n8103 = n8102 ^ n8101;
  assign n8112 = n7991 ^ n7687;
  assign n8104 = ~n4453 & n5814;
  assign n8105 = ~n2574 & n5817;
  assign n8106 = ~n2669 & n6295;
  assign n8107 = ~n8105 & ~n8106;
  assign n8108 = ~n2612 & n5824;
  assign n8109 = n8107 & ~n8108;
  assign n8110 = ~n8104 & n8109;
  assign n8111 = n8110 ^ x11;
  assign n8113 = n8112 ^ n8111;
  assign n8122 = n7988 ^ n7703;
  assign n8114 = ~n4312 & n5814;
  assign n8115 = ~n2612 & n5817;
  assign n8116 = ~n2482 & n5824;
  assign n8117 = ~n8115 & ~n8116;
  assign n8118 = ~n2574 & n6295;
  assign n8119 = n8117 & ~n8118;
  assign n8120 = ~n8114 & n8119;
  assign n8121 = n8120 ^ x11;
  assign n8123 = n8122 ^ n8121;
  assign n8132 = n7985 ^ n7721;
  assign n8124 = ~n4334 & n5814;
  assign n8125 = ~n2482 & n5817;
  assign n8126 = ~n2423 & n5824;
  assign n8127 = ~n8125 & ~n8126;
  assign n8128 = ~n2612 & n6295;
  assign n8129 = n8127 & ~n8128;
  assign n8130 = ~n8124 & n8129;
  assign n8131 = n8130 ^ x11;
  assign n8133 = n8132 ^ n8131;
  assign n8142 = n7982 ^ n7732;
  assign n8134 = n4433 & n5813;
  assign n8135 = n8134 ^ n2482;
  assign n8136 = n5812 & ~n8135;
  assign n8137 = ~n2357 & n5824;
  assign n8138 = ~n2423 & n5817;
  assign n8139 = ~n8137 & ~n8138;
  assign n8140 = ~n8136 & n8139;
  assign n8141 = n8140 ^ x11;
  assign n8143 = n8142 ^ n8141;
  assign n8145 = n7973 ^ n7783;
  assign n8154 = n7970 ^ n7802;
  assign n8146 = ~n4507 & n5814;
  assign n8147 = ~n2065 & n5817;
  assign n8148 = ~n1974 & n5824;
  assign n8149 = ~n8147 & ~n8148;
  assign n8150 = ~n2175 & n6295;
  assign n8151 = n8149 & ~n8150;
  assign n8152 = ~n8146 & n8151;
  assign n8153 = n8152 ^ x11;
  assign n8155 = n8154 ^ n8153;
  assign n8314 = ~n5167 & n5814;
  assign n8315 = ~n1878 & n5824;
  assign n8316 = ~n1974 & n5817;
  assign n8317 = ~n8315 & ~n8316;
  assign n8318 = ~n2065 & n6295;
  assign n8319 = n8317 & ~n8318;
  assign n8320 = ~n8314 & n8319;
  assign n8321 = n8320 ^ x11;
  assign n8164 = n7964 ^ n7830;
  assign n8156 = n5814 & ~n5923;
  assign n8157 = ~n1878 & n5817;
  assign n8158 = ~n1974 & n6295;
  assign n8159 = ~n8157 & ~n8158;
  assign n8160 = ~n1798 & n5824;
  assign n8161 = n8159 & ~n8160;
  assign n8162 = ~n8156 & n8161;
  assign n8163 = n8162 ^ x11;
  assign n8165 = n8164 ^ n8163;
  assign n8174 = n7961 ^ n7846;
  assign n8166 = n5023 & n5813;
  assign n8167 = n8166 ^ n1878;
  assign n8168 = n5812 & ~n8167;
  assign n8169 = ~n1726 & n5824;
  assign n8170 = ~n1798 & n5817;
  assign n8171 = ~n8169 & ~n8170;
  assign n8172 = ~n8168 & n8171;
  assign n8173 = n8172 ^ x11;
  assign n8175 = n8174 ^ n8173;
  assign n8176 = ~n5416 & n5814;
  assign n8177 = ~n882 & n5824;
  assign n8178 = ~n1544 & n6295;
  assign n8179 = ~n734 & n5817;
  assign n8180 = ~n8178 & ~n8179;
  assign n8181 = ~n8177 & n8180;
  assign n8182 = ~n8176 & n8181;
  assign n8183 = n8182 ^ x11;
  assign n8184 = n7944 ^ n7928;
  assign n8185 = n8184 ^ n7949;
  assign n8186 = n8183 & n8185;
  assign n8195 = n7926 ^ n7925;
  assign n8196 = n8195 ^ n7913;
  assign n8187 = ~n5465 & n5814;
  assign n8188 = ~n970 & n5824;
  assign n8189 = ~n734 & n6295;
  assign n8190 = ~n8188 & ~n8189;
  assign n8191 = ~n882 & n5817;
  assign n8192 = n8190 & ~n8191;
  assign n8193 = ~n8187 & n8192;
  assign n8194 = n8193 ^ x11;
  assign n8197 = n8196 ^ n8194;
  assign n8200 = ~n5481 & n5814;
  assign n8201 = ~n882 & n6295;
  assign n8202 = ~n1097 & n5824;
  assign n8203 = ~n8201 & ~n8202;
  assign n8204 = ~n970 & n5817;
  assign n8205 = n8203 & ~n8204;
  assign n8206 = ~n8200 & n8205;
  assign n8207 = n8206 ^ x11;
  assign n8198 = x14 & n7923;
  assign n8199 = n8198 ^ n7920;
  assign n8208 = n8207 ^ n8199;
  assign n8218 = ~n5564 & n5814;
  assign n8219 = ~n970 & n6295;
  assign n8220 = ~n1414 & n5824;
  assign n8221 = ~n8219 & ~n8220;
  assign n8222 = ~n1097 & n5817;
  assign n8223 = n8221 & ~n8222;
  assign n8224 = ~n8218 & n8223;
  assign n8225 = n8224 ^ x11;
  assign n8209 = ~n1208 & ~n5744;
  assign n8210 = x13 & ~n5742;
  assign n8211 = ~n8209 & n8210;
  assign n8212 = ~n5743 & ~n8211;
  assign n8213 = ~n1319 & ~n8212;
  assign n8214 = x13 & ~n1319;
  assign n8215 = n5748 & ~n8214;
  assign n8216 = ~n1208 & n8215;
  assign n8217 = ~n8213 & ~n8216;
  assign n8226 = n8225 ^ n8217;
  assign n8227 = ~n5579 & n5814;
  assign n8228 = ~n1208 & n5824;
  assign n8229 = ~n1414 & n5817;
  assign n8230 = ~n8228 & ~n8229;
  assign n8231 = ~n1097 & n6295;
  assign n8232 = n8230 & ~n8231;
  assign n8233 = ~n8227 & n8232;
  assign n8234 = n8233 ^ x12;
  assign n8235 = n5748 & n8234;
  assign n8236 = ~n1319 & n8235;
  assign n8237 = n5630 & n5813;
  assign n8238 = ~n1414 & n5812;
  assign n8239 = ~n8237 & n8238;
  assign n8240 = ~n1319 & n5824;
  assign n8241 = ~n8239 & ~n8240;
  assign n8242 = n5634 & n5814;
  assign n8243 = ~n5817 & ~n8242;
  assign n8244 = ~n1208 & ~n8243;
  assign n8245 = n8241 & ~n8244;
  assign n8246 = ~n1208 & n5812;
  assign n8247 = n1319 & ~n8246;
  assign n8248 = n5823 & ~n8247;
  assign n8249 = x11 & ~n8248;
  assign n8250 = n8245 & n8249;
  assign n8251 = n8233 & n8250;
  assign n8252 = ~n8236 & ~n8251;
  assign n8253 = n8252 ^ n8225;
  assign n8254 = ~n8226 & n8253;
  assign n8255 = n8254 ^ n8252;
  assign n8256 = n8255 ^ n8207;
  assign n8257 = ~n8208 & n8256;
  assign n8258 = n8257 ^ n8255;
  assign n8259 = n8258 ^ n8196;
  assign n8260 = n8197 & ~n8259;
  assign n8261 = n8260 ^ n8258;
  assign n8262 = ~n8186 & ~n8261;
  assign n8263 = ~n5069 & n5814;
  assign n8264 = ~n734 & n5824;
  assign n8265 = ~n1638 & n6295;
  assign n8266 = ~n8264 & ~n8265;
  assign n8267 = ~n1544 & n5817;
  assign n8268 = n8266 & ~n8267;
  assign n8269 = ~n8263 & n8268;
  assign n8270 = n8269 ^ x11;
  assign n8271 = n7952 ^ n7899;
  assign n8272 = ~n8270 & n8271;
  assign n8273 = ~n8183 & ~n8185;
  assign n8274 = ~n8272 & ~n8273;
  assign n8275 = ~n8262 & n8274;
  assign n8276 = n8270 & ~n8271;
  assign n8277 = ~n8275 & ~n8276;
  assign n8278 = n7955 ^ n7882;
  assign n8279 = n8277 & ~n8278;
  assign n8280 = n7958 ^ n7865;
  assign n8281 = ~n8279 & n8280;
  assign n8282 = n5350 & n5813;
  assign n8283 = n8282 ^ n1798;
  assign n8284 = n5812 & ~n8283;
  assign n8285 = ~n1726 & n5817;
  assign n8286 = ~n1638 & n5824;
  assign n8287 = ~n8285 & ~n8286;
  assign n8288 = ~n8284 & n8287;
  assign n8289 = n8288 ^ x11;
  assign n8290 = ~n8281 & ~n8289;
  assign n8291 = ~n8277 & n8278;
  assign n8292 = ~n5703 & n5814;
  assign n8293 = ~n1726 & n6295;
  assign n8294 = ~n1638 & n5817;
  assign n8295 = ~n8293 & ~n8294;
  assign n8296 = ~n1544 & n5824;
  assign n8297 = n8295 & ~n8296;
  assign n8298 = ~n8292 & n8297;
  assign n8299 = n8298 ^ x11;
  assign n8300 = n8298 ^ n8288;
  assign n8301 = n8280 & n8300;
  assign n8302 = ~n8299 & n8301;
  assign n8303 = n8302 ^ n8299;
  assign n8304 = ~n8291 & ~n8303;
  assign n8305 = n8279 & ~n8280;
  assign n8306 = ~n8304 & ~n8305;
  assign n8307 = ~n8290 & n8306;
  assign n8308 = n8307 ^ n8174;
  assign n8309 = n8175 & ~n8308;
  assign n8310 = n8309 ^ n8307;
  assign n8311 = n8310 ^ n8164;
  assign n8312 = ~n8165 & n8311;
  assign n8313 = n8312 ^ n8310;
  assign n8322 = n8321 ^ n8313;
  assign n8323 = n7967 ^ n7812;
  assign n8324 = n8323 ^ n8321;
  assign n8325 = n8322 & n8324;
  assign n8326 = n8325 ^ n8313;
  assign n8327 = n8326 ^ n8154;
  assign n8328 = ~n8155 & n8327;
  assign n8329 = n8328 ^ n8326;
  assign n8330 = n8145 & n8329;
  assign n8331 = ~n4253 & n5814;
  assign n8332 = ~n2065 & n5824;
  assign n8333 = ~n2247 & n6295;
  assign n8334 = ~n8332 & ~n8333;
  assign n8335 = ~n2175 & n5817;
  assign n8336 = n8334 & ~n8335;
  assign n8337 = ~n8331 & n8336;
  assign n8338 = n8337 ^ x11;
  assign n8339 = n8329 & n8338;
  assign n8340 = ~n8330 & ~n8339;
  assign n8341 = n7976 ^ n7767;
  assign n8342 = ~n4323 & n5814;
  assign n8343 = ~n2357 & n6295;
  assign n8344 = ~n2247 & n5817;
  assign n8345 = ~n8343 & ~n8344;
  assign n8346 = ~n2175 & n5824;
  assign n8347 = n8345 & ~n8346;
  assign n8348 = ~n8342 & n8347;
  assign n8349 = n8341 & n8348;
  assign n8350 = n8145 & n8337;
  assign n8351 = ~n8349 & ~n8350;
  assign n8352 = n8340 & n8351;
  assign n8353 = ~n8341 & ~n8348;
  assign n8354 = ~x11 & ~n8353;
  assign n8355 = ~n8352 & n8354;
  assign n8356 = n8341 & ~n8348;
  assign n8357 = n8145 & ~n8337;
  assign n8358 = ~n8356 & ~n8357;
  assign n8359 = n8340 & n8358;
  assign n8360 = ~n8341 & n8348;
  assign n8361 = x11 & ~n8360;
  assign n8362 = ~n8359 & n8361;
  assign n8363 = ~n8355 & ~n8362;
  assign n8144 = n7979 ^ n7751;
  assign n8364 = n8363 ^ n8144;
  assign n8365 = ~n4293 & n5814;
  assign n8366 = ~n2423 & n6295;
  assign n8367 = ~n2247 & n5824;
  assign n8368 = ~n8366 & ~n8367;
  assign n8369 = ~n2357 & n5817;
  assign n8370 = n8368 & ~n8369;
  assign n8371 = ~n8365 & n8370;
  assign n8372 = n8371 ^ x11;
  assign n8373 = n8372 ^ n8144;
  assign n8374 = ~n8364 & ~n8373;
  assign n8375 = n8374 ^ n8363;
  assign n8376 = n8375 ^ n8142;
  assign n8377 = ~n8143 & ~n8376;
  assign n8378 = n8377 ^ n8375;
  assign n8379 = n8378 ^ n8132;
  assign n8380 = n8133 & n8379;
  assign n8381 = n8380 ^ n8378;
  assign n8382 = n8381 ^ n8122;
  assign n8383 = ~n8123 & ~n8382;
  assign n8384 = n8383 ^ n8381;
  assign n8385 = n8384 ^ n8112;
  assign n8386 = ~n8113 & ~n8385;
  assign n8387 = n8386 ^ n8384;
  assign n8388 = n8387 ^ n8102;
  assign n8389 = n8103 & n8388;
  assign n8390 = n8389 ^ n8387;
  assign n8391 = n8390 ^ n8092;
  assign n8392 = n8093 & n8391;
  assign n8393 = n8392 ^ n8390;
  assign n8394 = n8393 ^ n8082;
  assign n8395 = ~n8083 & ~n8394;
  assign n8396 = n8395 ^ n8393;
  assign n8397 = n8396 ^ n8072;
  assign n8398 = n8073 & n8397;
  assign n8399 = n8398 ^ n8396;
  assign n8400 = n8399 ^ n8062;
  assign n8401 = ~n8063 & ~n8400;
  assign n8402 = n8401 ^ n8399;
  assign n8403 = n8402 ^ n8052;
  assign n8404 = n8053 & n8403;
  assign n8405 = n8404 ^ n8402;
  assign n8406 = n8405 ^ n8042;
  assign n8407 = n8043 & n8406;
  assign n8408 = n8407 ^ n8405;
  assign n8419 = n8418 ^ n8408;
  assign n7513 = x5 ^ x4;
  assign n7514 = x3 ^ x2;
  assign n7515 = n7513 & n7514;
  assign n8025 = ~n3879 & n7515;
  assign n7517 = x4 ^ x3;
  assign n7518 = ~n7514 & n7517;
  assign n7519 = ~n7514 & ~n7518;
  assign n7520 = n7513 & n7519;
  assign n8026 = ~n3404 & n7520;
  assign n8027 = ~n3431 & n7518;
  assign n8028 = ~n8026 & ~n8027;
  assign n8029 = ~n7513 & n7514;
  assign n8030 = ~n3875 & n8029;
  assign n8031 = n8028 & ~n8030;
  assign n8032 = ~n8025 & n8031;
  assign n8033 = n8032 ^ x5;
  assign n8420 = n8419 ^ n8033;
  assign n8422 = n3198 & n6304;
  assign n8423 = n8422 ^ n3270;
  assign n8424 = n6305 & ~n8423;
  assign n8425 = ~n3098 & n6316;
  assign n8426 = ~n3196 & n6309;
  assign n8427 = ~n8425 & ~n8426;
  assign n8428 = ~n8424 & n8427;
  assign n8429 = n8428 ^ x8;
  assign n8421 = n8405 ^ n8043;
  assign n8430 = n8429 ^ n8421;
  assign n8439 = n8402 ^ n8053;
  assign n8431 = n3647 & n6306;
  assign n8432 = ~n2954 & n6316;
  assign n8433 = ~n3196 & n7168;
  assign n8434 = ~n8432 & ~n8433;
  assign n8435 = ~n3098 & n6309;
  assign n8436 = n8434 & ~n8435;
  assign n8437 = ~n8431 & n8436;
  assign n8438 = n8437 ^ x8;
  assign n8440 = n8439 ^ n8438;
  assign n8449 = n8399 ^ n8063;
  assign n8441 = ~n3974 & n6306;
  assign n8442 = ~n2954 & n6309;
  assign n8443 = ~n3037 & n6316;
  assign n8444 = ~n8442 & ~n8443;
  assign n8445 = ~n3098 & n7168;
  assign n8446 = n8444 & ~n8445;
  assign n8447 = ~n8441 & n8446;
  assign n8448 = n8447 ^ x8;
  assign n8450 = n8449 ^ n8448;
  assign n8834 = n8396 ^ n8073;
  assign n8459 = n8393 ^ n8083;
  assign n8451 = ~n3632 & n6306;
  assign n8452 = ~n368 & n6309;
  assign n8453 = ~n3037 & n7168;
  assign n8454 = ~n8452 & ~n8453;
  assign n8455 = ~n566 & n6316;
  assign n8456 = n8454 & ~n8455;
  assign n8457 = ~n8451 & n8456;
  assign n8458 = n8457 ^ x8;
  assign n8460 = n8459 ^ n8458;
  assign n8469 = n8390 ^ n8093;
  assign n8461 = n3749 & n6306;
  assign n8462 = ~n368 & n7168;
  assign n8463 = ~n2861 & n6316;
  assign n8464 = ~n8462 & ~n8463;
  assign n8465 = ~n566 & n6309;
  assign n8466 = n8464 & ~n8465;
  assign n8467 = ~n8461 & n8466;
  assign n8468 = n8467 ^ x8;
  assign n8470 = n8469 ^ n8468;
  assign n8479 = n8387 ^ n8103;
  assign n8471 = ~n3666 & n6306;
  assign n8472 = ~n2718 & n6316;
  assign n8473 = ~n2861 & n6309;
  assign n8474 = ~n8472 & ~n8473;
  assign n8475 = ~n566 & n7168;
  assign n8476 = n8474 & ~n8475;
  assign n8477 = ~n8471 & n8476;
  assign n8478 = n8477 ^ x8;
  assign n8480 = n8479 ^ n8478;
  assign n8489 = n8384 ^ n8113;
  assign n8481 = ~n4466 & n6306;
  assign n8482 = ~n2718 & n6309;
  assign n8483 = ~n2861 & n7168;
  assign n8484 = ~n2786 & n6316;
  assign n8485 = ~n8483 & ~n8484;
  assign n8486 = ~n8482 & n8485;
  assign n8487 = ~n8481 & n8486;
  assign n8488 = n8487 ^ x8;
  assign n8490 = n8489 ^ n8488;
  assign n8499 = n8381 ^ n8123;
  assign n8491 = ~n4495 & n6306;
  assign n8492 = ~n2718 & n7168;
  assign n8493 = ~n2786 & n6309;
  assign n8494 = ~n2669 & n6316;
  assign n8495 = ~n8493 & ~n8494;
  assign n8496 = ~n8492 & n8495;
  assign n8497 = ~n8491 & n8496;
  assign n8498 = n8497 ^ x8;
  assign n8500 = n8499 ^ n8498;
  assign n8502 = ~n4653 & n6306;
  assign n8503 = ~n2574 & n6316;
  assign n8504 = ~n2786 & n7168;
  assign n8505 = ~n2669 & n6309;
  assign n8506 = ~n8504 & ~n8505;
  assign n8507 = ~n8503 & n8506;
  assign n8508 = ~n8502 & n8507;
  assign n8509 = n8508 ^ x8;
  assign n8501 = n8378 ^ n8133;
  assign n8510 = n8509 ^ n8501;
  assign n8519 = n8375 ^ n8143;
  assign n8511 = ~n4453 & n6306;
  assign n8512 = ~n2612 & n6316;
  assign n8513 = ~n2669 & n7168;
  assign n8514 = ~n8512 & ~n8513;
  assign n8515 = ~n2574 & n6309;
  assign n8516 = n8514 & ~n8515;
  assign n8517 = ~n8511 & n8516;
  assign n8518 = n8517 ^ x8;
  assign n8520 = n8519 ^ n8518;
  assign n8529 = n8372 ^ n8364;
  assign n8521 = ~n4312 & n6306;
  assign n8522 = ~n2574 & n7168;
  assign n8523 = ~n2482 & n6316;
  assign n8524 = ~n8522 & ~n8523;
  assign n8525 = ~n2612 & n6309;
  assign n8526 = n8524 & ~n8525;
  assign n8527 = ~n8521 & n8526;
  assign n8528 = n8527 ^ x8;
  assign n8530 = n8529 ^ n8528;
  assign n8544 = n8348 ^ n8341;
  assign n8539 = n8329 ^ n8145;
  assign n8540 = n8145 ^ x11;
  assign n8541 = n8540 ^ n8337;
  assign n8542 = ~n8539 & n8541;
  assign n8543 = n8542 ^ n8337;
  assign n8545 = n8544 ^ n8543;
  assign n8531 = ~n4334 & n6306;
  assign n8532 = ~n2482 & n6309;
  assign n8533 = ~n2423 & n6316;
  assign n8534 = ~n8532 & ~n8533;
  assign n8535 = ~n2612 & n7168;
  assign n8536 = n8534 & ~n8535;
  assign n8537 = ~n8531 & n8536;
  assign n8538 = n8537 ^ x8;
  assign n8546 = n8545 ^ n8538;
  assign n8555 = n8539 ^ n8338;
  assign n8547 = ~n4434 & n6306;
  assign n8548 = ~n2423 & n6309;
  assign n8549 = ~n2482 & n7168;
  assign n8550 = ~n8548 & ~n8549;
  assign n8551 = ~n2357 & n6316;
  assign n8552 = n8550 & ~n8551;
  assign n8553 = ~n8547 & n8552;
  assign n8554 = n8553 ^ x8;
  assign n8556 = n8555 ^ n8554;
  assign n8557 = ~n4293 & n6306;
  assign n8558 = ~n2423 & n7168;
  assign n8559 = ~n2247 & n6316;
  assign n8560 = ~n8558 & ~n8559;
  assign n8561 = ~n2357 & n6309;
  assign n8562 = n8560 & ~n8561;
  assign n8563 = ~n8557 & n8562;
  assign n8564 = n8563 ^ x8;
  assign n8573 = n8323 ^ n8322;
  assign n8565 = ~n4323 & n6306;
  assign n8566 = ~n2175 & n6316;
  assign n8567 = ~n2247 & n6309;
  assign n8568 = ~n8566 & ~n8567;
  assign n8569 = ~n2357 & n7168;
  assign n8570 = n8568 & ~n8569;
  assign n8571 = ~n8565 & n8570;
  assign n8572 = n8571 ^ x8;
  assign n8574 = n8573 ^ n8572;
  assign n8583 = n8310 ^ n8165;
  assign n8575 = ~n4253 & n6306;
  assign n8576 = ~n2065 & n6316;
  assign n8577 = ~n2175 & n6309;
  assign n8578 = ~n8576 & ~n8577;
  assign n8579 = ~n2247 & n7168;
  assign n8580 = n8578 & ~n8579;
  assign n8581 = ~n8575 & n8580;
  assign n8582 = n8581 ^ x8;
  assign n8584 = n8583 ^ n8582;
  assign n8586 = ~n4507 & n6306;
  assign n8587 = ~n2175 & n7168;
  assign n8588 = ~n1974 & n6316;
  assign n8589 = ~n8587 & ~n8588;
  assign n8590 = ~n2065 & n6309;
  assign n8591 = n8589 & ~n8590;
  assign n8592 = ~n8586 & n8591;
  assign n8593 = n8592 ^ x8;
  assign n8585 = n8307 ^ n8175;
  assign n8594 = n8593 ^ n8585;
  assign n8608 = n8288 ^ n8280;
  assign n8603 = n8278 ^ n8277;
  assign n8604 = n8278 ^ x11;
  assign n8605 = n8604 ^ n8298;
  assign n8606 = n8603 & n8605;
  assign n8607 = n8606 ^ n8298;
  assign n8609 = n8608 ^ n8607;
  assign n8595 = ~n5167 & n6306;
  assign n8596 = ~n2065 & n7168;
  assign n8597 = ~n1974 & n6309;
  assign n8598 = ~n8596 & ~n8597;
  assign n8599 = ~n1878 & n6316;
  assign n8600 = n8598 & ~n8599;
  assign n8601 = ~n8595 & n8600;
  assign n8602 = n8601 ^ x8;
  assign n8610 = n8609 ^ n8602;
  assign n8619 = n8603 ^ n8299;
  assign n8611 = ~n5923 & n6306;
  assign n8612 = ~n1798 & n6316;
  assign n8613 = ~n1974 & n7168;
  assign n8614 = ~n8612 & ~n8613;
  assign n8615 = ~n1878 & n6309;
  assign n8616 = n8614 & ~n8615;
  assign n8617 = ~n8611 & n8616;
  assign n8618 = n8617 ^ x8;
  assign n8620 = n8619 ^ n8618;
  assign n8630 = n8183 ^ n7949;
  assign n8631 = ~n7945 & ~n8261;
  assign n8632 = ~n7950 & ~n8631;
  assign n8633 = n8632 ^ n7949;
  assign n8634 = ~n8630 & n8633;
  assign n8635 = n8261 ^ n7944;
  assign n8636 = ~n8184 & n8635;
  assign n8637 = n8630 & n8636;
  assign n8638 = n8637 ^ n8630;
  assign n8639 = ~n8634 & ~n8638;
  assign n8629 = n8270 ^ n7899;
  assign n8640 = n8639 ^ n8629;
  assign n8621 = ~n5371 & n6306;
  assign n8622 = ~n1798 & n6309;
  assign n8623 = ~n1726 & n6316;
  assign n8624 = ~n8622 & ~n8623;
  assign n8625 = ~n1878 & n7168;
  assign n8626 = n8624 & ~n8625;
  assign n8627 = ~n8621 & n8626;
  assign n8628 = n8627 ^ x8;
  assign n8641 = n8640 ^ n8628;
  assign n8644 = ~n5351 & n6306;
  assign n8645 = ~n1726 & n6309;
  assign n8646 = ~n1638 & n6316;
  assign n8647 = ~n8645 & ~n8646;
  assign n8648 = ~n1798 & n7168;
  assign n8649 = n8647 & ~n8648;
  assign n8650 = ~n8644 & n8649;
  assign n8651 = n8650 ^ x8;
  assign n8642 = n8185 ^ n8183;
  assign n8643 = n8642 ^ n8261;
  assign n8652 = n8651 ^ n8643;
  assign n8661 = n8258 ^ n8197;
  assign n8653 = ~n5703 & n6306;
  assign n8654 = ~n1726 & n7168;
  assign n8655 = ~n1638 & n6309;
  assign n8656 = ~n1544 & n6316;
  assign n8657 = ~n8655 & ~n8656;
  assign n8658 = ~n8654 & n8657;
  assign n8659 = ~n8653 & n8658;
  assign n8660 = n8659 ^ x8;
  assign n8662 = n8661 ^ n8660;
  assign n8671 = n8255 ^ n8208;
  assign n8663 = ~n5069 & n6306;
  assign n8664 = ~n734 & n6316;
  assign n8665 = ~n1544 & n6309;
  assign n8666 = ~n8664 & ~n8665;
  assign n8667 = ~n1638 & n7168;
  assign n8668 = n8666 & ~n8667;
  assign n8669 = ~n8663 & n8668;
  assign n8670 = n8669 ^ x8;
  assign n8672 = n8671 ^ n8670;
  assign n8681 = n8252 ^ n8226;
  assign n8673 = ~n5416 & n6306;
  assign n8674 = ~n882 & n6316;
  assign n8675 = ~n734 & n6309;
  assign n8676 = ~n1544 & n7168;
  assign n8677 = ~n8675 & ~n8676;
  assign n8678 = ~n8674 & n8677;
  assign n8679 = ~n8673 & n8678;
  assign n8680 = n8679 ^ x8;
  assign n8682 = n8681 ^ n8680;
  assign n8690 = ~n5465 & n6306;
  assign n8691 = ~n882 & n6309;
  assign n8692 = ~n734 & n7168;
  assign n8693 = ~n8691 & ~n8692;
  assign n8694 = ~n970 & n6316;
  assign n8695 = n8693 & ~n8694;
  assign n8696 = ~n8690 & n8695;
  assign n8697 = n8696 ^ x8;
  assign n8685 = ~x12 & ~n1319;
  assign n8683 = ~n1319 & n5748;
  assign n8684 = n8683 ^ x11;
  assign n8686 = n8685 ^ n8684;
  assign n8687 = ~n8250 & n8686;
  assign n8688 = n8687 ^ n8685;
  assign n8689 = n8688 ^ n8233;
  assign n8698 = n8697 ^ n8689;
  assign n8701 = ~n5481 & n6306;
  assign n8702 = ~n970 & n6309;
  assign n8703 = ~n1097 & n6316;
  assign n8704 = ~n8702 & ~n8703;
  assign n8705 = ~n882 & n7168;
  assign n8706 = n8704 & ~n8705;
  assign n8707 = ~n8701 & n8706;
  assign n8708 = n8707 ^ x8;
  assign n8699 = x11 & n8248;
  assign n8700 = n8699 ^ n8245;
  assign n8709 = n8708 ^ n8700;
  assign n8719 = ~n5564 & n6306;
  assign n8720 = ~n1097 & n6309;
  assign n8721 = ~n1414 & n6316;
  assign n8722 = ~n8720 & ~n8721;
  assign n8723 = ~n970 & n7168;
  assign n8724 = n8722 & ~n8723;
  assign n8725 = ~n8719 & n8724;
  assign n8726 = n8725 ^ x8;
  assign n8710 = ~n1208 & ~n5819;
  assign n8711 = x10 & ~n5821;
  assign n8712 = ~n8710 & n8711;
  assign n8713 = ~x10 & n5821;
  assign n8714 = ~n8712 & ~n8713;
  assign n8715 = x10 & ~n1319;
  assign n8716 = n8246 & ~n8715;
  assign n8717 = n8714 & ~n8716;
  assign n8718 = ~n8247 & ~n8717;
  assign n8727 = n8726 ^ n8718;
  assign n8728 = ~n5579 & n6306;
  assign n8729 = ~n1097 & n7168;
  assign n8730 = ~n1414 & n6309;
  assign n8731 = ~n8729 & ~n8730;
  assign n8732 = ~n1208 & n6316;
  assign n8733 = n8731 & ~n8732;
  assign n8734 = ~n8728 & n8733;
  assign n8735 = n8734 ^ x9;
  assign n8736 = n5812 & n8735;
  assign n8737 = ~n1319 & n8736;
  assign n8738 = n5630 & n6304;
  assign n8739 = ~n1414 & n6305;
  assign n8740 = ~n8738 & n8739;
  assign n8741 = ~n1319 & n6316;
  assign n8742 = ~n8740 & ~n8741;
  assign n8743 = n5634 & n6306;
  assign n8744 = ~n6309 & ~n8743;
  assign n8745 = ~n1208 & ~n8744;
  assign n8746 = n8742 & ~n8745;
  assign n8747 = ~n1208 & n6305;
  assign n8748 = ~n1319 & n6315;
  assign n8749 = ~n8747 & ~n8748;
  assign n8750 = x8 & n8749;
  assign n8751 = n8746 & n8750;
  assign n8752 = n8734 & n8751;
  assign n8753 = ~n8737 & ~n8752;
  assign n8754 = n8753 ^ n8726;
  assign n8755 = n8727 & n8754;
  assign n8756 = n8755 ^ n8753;
  assign n8757 = n8756 ^ n8708;
  assign n8758 = ~n8709 & n8757;
  assign n8759 = n8758 ^ n8756;
  assign n8760 = n8759 ^ n8697;
  assign n8761 = ~n8698 & n8760;
  assign n8762 = n8761 ^ n8759;
  assign n8763 = n8762 ^ n8681;
  assign n8764 = ~n8682 & n8763;
  assign n8765 = n8764 ^ n8762;
  assign n8766 = n8765 ^ n8671;
  assign n8767 = ~n8672 & n8766;
  assign n8768 = n8767 ^ n8765;
  assign n8769 = n8768 ^ n8661;
  assign n8770 = n8662 & ~n8769;
  assign n8771 = n8770 ^ n8768;
  assign n8772 = n8771 ^ n8651;
  assign n8773 = ~n8652 & n8772;
  assign n8774 = n8773 ^ n8771;
  assign n8775 = n8774 ^ n8640;
  assign n8776 = n8641 & ~n8775;
  assign n8777 = n8776 ^ n8774;
  assign n8778 = n8777 ^ n8619;
  assign n8779 = n8620 & ~n8778;
  assign n8780 = n8779 ^ n8777;
  assign n8781 = n8780 ^ n8609;
  assign n8782 = ~n8610 & n8781;
  assign n8783 = n8782 ^ n8780;
  assign n8784 = n8783 ^ n8593;
  assign n8785 = n8594 & n8784;
  assign n8786 = n8785 ^ n8783;
  assign n8787 = n8786 ^ n8583;
  assign n8788 = ~n8584 & n8787;
  assign n8789 = n8788 ^ n8786;
  assign n8790 = n8789 ^ n8573;
  assign n8791 = n8574 & ~n8790;
  assign n8792 = n8791 ^ n8789;
  assign n8793 = n8564 & n8792;
  assign n8794 = n8326 ^ n8155;
  assign n8795 = ~n8573 & n8789;
  assign n8796 = n8571 ^ n8563;
  assign n8797 = ~n8572 & ~n8796;
  assign n8798 = ~n8795 & n8797;
  assign n8799 = n8794 & ~n8798;
  assign n8800 = n8573 & ~n8789;
  assign n8801 = ~n8564 & n8800;
  assign n8802 = n8799 & ~n8801;
  assign n8803 = ~n8793 & ~n8802;
  assign n8804 = n8803 ^ n8555;
  assign n8805 = ~n8556 & ~n8804;
  assign n8806 = n8805 ^ n8803;
  assign n8807 = n8806 ^ n8545;
  assign n8808 = ~n8546 & ~n8807;
  assign n8809 = n8808 ^ n8806;
  assign n8810 = n8809 ^ n8529;
  assign n8811 = n8530 & n8810;
  assign n8812 = n8811 ^ n8809;
  assign n8813 = n8812 ^ n8519;
  assign n8814 = n8520 & n8813;
  assign n8815 = n8814 ^ n8812;
  assign n8816 = n8815 ^ n8509;
  assign n8817 = ~n8510 & ~n8816;
  assign n8818 = n8817 ^ n8815;
  assign n8819 = n8818 ^ n8499;
  assign n8820 = n8500 & n8819;
  assign n8821 = n8820 ^ n8818;
  assign n8822 = n8821 ^ n8489;
  assign n8823 = n8490 & n8822;
  assign n8824 = n8823 ^ n8821;
  assign n8825 = n8824 ^ n8479;
  assign n8826 = ~n8480 & ~n8825;
  assign n8827 = n8826 ^ n8824;
  assign n8828 = n8827 ^ n8469;
  assign n8829 = ~n8470 & ~n8828;
  assign n8830 = n8829 ^ n8827;
  assign n8831 = n8830 ^ n8459;
  assign n8832 = n8460 & n8831;
  assign n8833 = n8832 ^ n8830;
  assign n8835 = n8834 ^ n8833;
  assign n8836 = ~n3777 & n6306;
  assign n8837 = ~n2954 & n7168;
  assign n8838 = ~n3037 & n6309;
  assign n8839 = ~n8837 & ~n8838;
  assign n8840 = ~n368 & n6316;
  assign n8841 = n8839 & ~n8840;
  assign n8842 = ~n8836 & n8841;
  assign n8843 = n8842 ^ x8;
  assign n8844 = n8843 ^ n8834;
  assign n8845 = ~n8835 & ~n8844;
  assign n8846 = n8845 ^ n8833;
  assign n8847 = n8846 ^ n8449;
  assign n8848 = n8450 & n8847;
  assign n8849 = n8848 ^ n8846;
  assign n8850 = n8849 ^ n8439;
  assign n8851 = ~n8440 & ~n8850;
  assign n8852 = n8851 ^ n8849;
  assign n8853 = n8852 ^ n8429;
  assign n8854 = ~n8430 & ~n8853;
  assign n8855 = n8854 ^ n8852;
  assign n8856 = n8855 ^ n8419;
  assign n8857 = n8420 & n8856;
  assign n8858 = n8857 ^ n8855;
  assign n8859 = n8417 ^ n8408;
  assign n8860 = ~n8418 & ~n8859;
  assign n8861 = n8860 ^ n8408;
  assign n8862 = n8858 & n8861;
  assign n8016 = n8015 ^ n7555;
  assign n8017 = ~n7556 & n8016;
  assign n8018 = n8017 ^ n8015;
  assign n7534 = n7504 ^ n7192;
  assign n7526 = ~n5770 & n6306;
  assign n7527 = ~n3270 & n6316;
  assign n7528 = ~n3351 & n6309;
  assign n7529 = ~n3404 & n7168;
  assign n7530 = ~n7528 & ~n7529;
  assign n7531 = ~n7527 & n7530;
  assign n7532 = ~n7526 & n7531;
  assign n7533 = n7532 ^ x8;
  assign n7535 = n7534 ^ n7533;
  assign n8863 = n8018 ^ n7535;
  assign n8864 = n8862 & n8863;
  assign n8865 = n5758 & n7515;
  assign n8866 = ~n3875 & n7518;
  assign n8867 = ~n3431 & n7520;
  assign n8868 = ~n8866 & ~n8867;
  assign n8869 = ~n8865 & n8868;
  assign n8870 = n8869 ^ x5;
  assign n8871 = n8864 & ~n8870;
  assign n8019 = n8018 ^ n7534;
  assign n8020 = n7535 & ~n8019;
  assign n8021 = n8020 ^ n8018;
  assign n7524 = n7507 ^ n7182;
  assign n7516 = n6285 & n7515;
  assign n7521 = ~n3875 & n7520;
  assign n7522 = ~n7516 & ~n7521;
  assign n7523 = n7522 ^ x5;
  assign n7525 = n7524 ^ n7523;
  assign n8872 = n8021 ^ n7525;
  assign n8873 = ~n8871 & n8872;
  assign n8874 = ~n8858 & ~n8861;
  assign n8875 = ~n8863 & n8874;
  assign n8876 = ~n8870 & ~n8875;
  assign n8877 = n8861 ^ n8858;
  assign n8878 = n8863 ^ n8861;
  assign n8879 = n8877 & ~n8878;
  assign n8880 = n8879 ^ n8858;
  assign n8881 = ~n8876 & ~n8880;
  assign n8882 = ~n8873 & ~n8881;
  assign n8906 = n8855 ^ n8420;
  assign n8893 = ~n3432 & n7515;
  assign n8894 = ~n3404 & n7518;
  assign n8895 = ~n3351 & n7520;
  assign n8896 = ~n8894 & ~n8895;
  assign n8897 = ~n3431 & n8029;
  assign n8898 = n8896 & ~n8897;
  assign n8899 = ~n8893 & n8898;
  assign n8900 = n8899 ^ x5;
  assign n8883 = x0 & x1;
  assign n8884 = ~n3875 & n8883;
  assign n8885 = ~n3876 & n8884;
  assign n8886 = x1 & x2;
  assign n8887 = x2 & n3875;
  assign n8888 = ~n8886 & ~n8887;
  assign n8889 = ~n8885 & n8888;
  assign n8890 = x0 & x2;
  assign n8891 = n3876 & n8890;
  assign n8892 = n8889 & ~n8891;
  assign n8901 = n8900 ^ n8892;
  assign n8902 = n8852 ^ n8430;
  assign n8903 = n8902 ^ n8900;
  assign n8904 = ~n8901 & ~n8903;
  assign n8905 = n8904 ^ n8902;
  assign n8907 = n8906 ^ n8905;
  assign n8908 = n8849 ^ n8440;
  assign n8909 = ~n3410 & ~n3876;
  assign n8910 = n3875 & ~n8909;
  assign n8911 = ~n6285 & ~n8910;
  assign n8912 = n8890 & ~n8911;
  assign n8913 = n3877 & n8883;
  assign n8914 = ~n8886 & ~n8913;
  assign n8915 = n3875 & ~n8914;
  assign n8916 = x1 & ~n3875;
  assign n8917 = x2 & n3431;
  assign n8918 = ~n8916 & ~n8917;
  assign n33 = x2 ^ x1;
  assign n8919 = ~x0 & n33;
  assign n8920 = ~n8918 & n8919;
  assign n8921 = ~n8915 & ~n8920;
  assign n8922 = ~n8912 & n8921;
  assign n8923 = n8884 & ~n8909;
  assign n8924 = ~n8887 & ~n8923;
  assign n8925 = n3431 & ~n8924;
  assign n8926 = n8922 & ~n8925;
  assign n8927 = ~n8908 & n8926;
  assign n9448 = ~x0 & ~x1;
  assign n9877 = x2 & n3404;
  assign n9878 = n9448 & n9877;
  assign n9378 = ~x0 & x1;
  assign n9879 = n3431 ^ x2;
  assign n9880 = n9378 & ~n9879;
  assign n9881 = ~n9878 & ~n9880;
  assign n9882 = n33 & ~n3878;
  assign n9883 = n9882 ^ x1;
  assign n9884 = n9883 ^ n3875;
  assign n9885 = x0 & ~n9884;
  assign n9886 = n9881 & ~n9885;
  assign n9340 = n8843 ^ n8835;
  assign n9332 = ~n3271 & n7515;
  assign n9333 = ~n3098 & n7520;
  assign n9334 = ~n3196 & n7518;
  assign n9335 = ~n9333 & ~n9334;
  assign n9336 = ~n3270 & n8029;
  assign n9337 = n9335 & ~n9336;
  assign n9338 = ~n9332 & n9337;
  assign n9339 = n9338 ^ x5;
  assign n9341 = n9340 ^ n9339;
  assign n8947 = n8830 ^ n8460;
  assign n8939 = n3647 & n7515;
  assign n8940 = ~n3098 & n7518;
  assign n8941 = ~n3196 & n8029;
  assign n8942 = ~n8940 & ~n8941;
  assign n8943 = ~n2954 & n7520;
  assign n8944 = n8942 & ~n8943;
  assign n8945 = ~n8939 & n8944;
  assign n8946 = n8945 ^ x5;
  assign n8948 = n8947 ^ n8946;
  assign n8957 = n8827 ^ n8470;
  assign n8949 = ~n3974 & n7515;
  assign n8950 = ~n2954 & n7518;
  assign n8951 = ~n3098 & n8029;
  assign n8952 = ~n8950 & ~n8951;
  assign n8953 = ~n3037 & n7520;
  assign n8954 = n8952 & ~n8953;
  assign n8955 = ~n8949 & n8954;
  assign n8956 = n8955 ^ x5;
  assign n8958 = n8957 ^ n8956;
  assign n8967 = n8824 ^ n8480;
  assign n8959 = ~n3777 & n7515;
  assign n8960 = ~n2954 & n8029;
  assign n8961 = ~n368 & n7520;
  assign n8962 = ~n8960 & ~n8961;
  assign n8963 = ~n3037 & n7518;
  assign n8964 = n8962 & ~n8963;
  assign n8965 = ~n8959 & n8964;
  assign n8966 = n8965 ^ x5;
  assign n8968 = n8967 ^ n8966;
  assign n8977 = n8821 ^ n8490;
  assign n8969 = ~n3632 & n7515;
  assign n8970 = ~n368 & n7518;
  assign n8971 = ~n3037 & n8029;
  assign n8972 = ~n8970 & ~n8971;
  assign n8973 = ~n566 & n7520;
  assign n8974 = n8972 & ~n8973;
  assign n8975 = ~n8969 & n8974;
  assign n8976 = n8975 ^ x5;
  assign n8978 = n8977 ^ n8976;
  assign n8979 = n8818 ^ n8500;
  assign n8980 = ~n3748 & n7513;
  assign n8981 = n8980 ^ n368;
  assign n8982 = n7514 & ~n8981;
  assign n8983 = ~n566 & n7518;
  assign n8984 = ~n2861 & n7520;
  assign n8985 = ~n8983 & ~n8984;
  assign n8986 = ~n8982 & n8985;
  assign n8987 = n8986 ^ x5;
  assign n8988 = n8979 & n8987;
  assign n8989 = n8815 ^ n8510;
  assign n8998 = n8812 ^ n8520;
  assign n8990 = ~n4466 & n7515;
  assign n8991 = ~n2718 & n7518;
  assign n8992 = ~n2861 & n8029;
  assign n8993 = ~n2786 & n7520;
  assign n8994 = ~n8992 & ~n8993;
  assign n8995 = ~n8991 & n8994;
  assign n8996 = ~n8990 & n8995;
  assign n8997 = n8996 ^ x5;
  assign n8999 = n8998 ^ n8997;
  assign n9001 = ~n4495 & n7515;
  assign n9002 = ~n2718 & n8029;
  assign n9003 = ~n2669 & n7520;
  assign n9004 = ~n2786 & n7518;
  assign n9005 = ~n9003 & ~n9004;
  assign n9006 = ~n9002 & n9005;
  assign n9007 = ~n9001 & n9006;
  assign n9008 = n9007 ^ x5;
  assign n9000 = n8809 ^ n8530;
  assign n9009 = n9008 ^ n9000;
  assign n9018 = n8806 ^ n8546;
  assign n9010 = ~n4653 & n7515;
  assign n9011 = ~n2574 & n7520;
  assign n9012 = ~n2786 & n8029;
  assign n9013 = ~n2669 & n7518;
  assign n9014 = ~n9012 & ~n9013;
  assign n9015 = ~n9011 & n9014;
  assign n9016 = ~n9010 & n9015;
  assign n9017 = n9016 ^ x5;
  assign n9019 = n9018 ^ n9017;
  assign n9028 = n8803 ^ n8556;
  assign n9020 = n4452 & n7513;
  assign n9021 = n9020 ^ n2669;
  assign n9022 = n7514 & ~n9021;
  assign n9023 = ~n2612 & n7520;
  assign n9024 = ~n2574 & n7518;
  assign n9025 = ~n9023 & ~n9024;
  assign n9026 = ~n9022 & n9025;
  assign n9027 = n9026 ^ x5;
  assign n9029 = n9028 ^ n9027;
  assign n9038 = n8794 ^ n8564;
  assign n9039 = n9038 ^ n8792;
  assign n9030 = ~n4312 & n7515;
  assign n9031 = ~n2612 & n7518;
  assign n9032 = ~n2482 & n7520;
  assign n9033 = ~n9031 & ~n9032;
  assign n9034 = ~n2574 & n8029;
  assign n9035 = n9033 & ~n9034;
  assign n9036 = ~n9030 & n9035;
  assign n9037 = n9036 ^ x5;
  assign n9040 = n9039 ^ n9037;
  assign n9049 = n8789 ^ n8574;
  assign n9041 = ~n4334 & n7515;
  assign n9042 = ~n2612 & n8029;
  assign n9043 = ~n2423 & n7520;
  assign n9044 = ~n9042 & ~n9043;
  assign n9045 = ~n2482 & n7518;
  assign n9046 = n9044 & ~n9045;
  assign n9047 = ~n9041 & n9046;
  assign n9048 = n9047 ^ x5;
  assign n9050 = n9049 ^ n9048;
  assign n9059 = n8786 ^ n8584;
  assign n9051 = ~n4434 & n7515;
  assign n9052 = ~n2482 & n8029;
  assign n9053 = ~n2423 & n7518;
  assign n9054 = ~n9052 & ~n9053;
  assign n9055 = ~n2357 & n7520;
  assign n9056 = n9054 & ~n9055;
  assign n9057 = ~n9051 & n9056;
  assign n9058 = n9057 ^ x5;
  assign n9060 = n9059 ^ n9058;
  assign n9069 = n8783 ^ n8594;
  assign n9061 = ~n4293 & n7515;
  assign n9062 = ~n2423 & n8029;
  assign n9063 = ~n2247 & n7520;
  assign n9064 = ~n9062 & ~n9063;
  assign n9065 = ~n2357 & n7518;
  assign n9066 = n9064 & ~n9065;
  assign n9067 = ~n9061 & n9066;
  assign n9068 = n9067 ^ x5;
  assign n9070 = n9069 ^ n9068;
  assign n9079 = n8780 ^ n8610;
  assign n9071 = ~n4323 & n7515;
  assign n9072 = ~n2357 & n8029;
  assign n9073 = ~n2247 & n7518;
  assign n9074 = ~n9072 & ~n9073;
  assign n9075 = ~n2175 & n7520;
  assign n9076 = n9074 & ~n9075;
  assign n9077 = ~n9071 & n9076;
  assign n9078 = n9077 ^ x5;
  assign n9080 = n9079 ^ n9078;
  assign n9089 = n8777 ^ n8620;
  assign n9081 = ~n4253 & n7515;
  assign n9082 = ~n2065 & n7520;
  assign n9083 = ~n2175 & n7518;
  assign n9084 = ~n9082 & ~n9083;
  assign n9085 = ~n2247 & n8029;
  assign n9086 = n9084 & ~n9085;
  assign n9087 = ~n9081 & n9086;
  assign n9088 = n9087 ^ x5;
  assign n9090 = n9089 ^ n9088;
  assign n9099 = n8774 ^ n8641;
  assign n9091 = ~n4507 & n7515;
  assign n9092 = ~n2065 & n7518;
  assign n9093 = ~n2175 & n8029;
  assign n9094 = ~n9092 & ~n9093;
  assign n9095 = ~n1974 & n7520;
  assign n9096 = n9094 & ~n9095;
  assign n9097 = ~n9091 & n9096;
  assign n9098 = n9097 ^ x5;
  assign n9100 = n9099 ^ n9098;
  assign n9109 = n8771 ^ n8652;
  assign n9101 = ~n5167 & n7515;
  assign n9102 = ~n2065 & n8029;
  assign n9103 = ~n1974 & n7518;
  assign n9104 = ~n9102 & ~n9103;
  assign n9105 = ~n1878 & n7520;
  assign n9106 = n9104 & ~n9105;
  assign n9107 = ~n9101 & n9106;
  assign n9108 = n9107 ^ x5;
  assign n9110 = n9109 ^ n9108;
  assign n9119 = n8768 ^ n8662;
  assign n9111 = ~n5923 & n7515;
  assign n9112 = ~n1798 & n7520;
  assign n9113 = ~n1974 & n8029;
  assign n9114 = ~n9112 & ~n9113;
  assign n9115 = ~n1878 & n7518;
  assign n9116 = n9114 & ~n9115;
  assign n9117 = ~n9111 & n9116;
  assign n9118 = n9117 ^ x5;
  assign n9120 = n9119 ^ n9118;
  assign n9129 = n8765 ^ n8672;
  assign n9121 = ~n5371 & n7515;
  assign n9122 = ~n1798 & n7518;
  assign n9123 = ~n1878 & n8029;
  assign n9124 = ~n9122 & ~n9123;
  assign n9125 = ~n1726 & n7520;
  assign n9126 = n9124 & ~n9125;
  assign n9127 = ~n9121 & n9126;
  assign n9128 = n9127 ^ x5;
  assign n9130 = n9129 ^ n9128;
  assign n9139 = n8762 ^ n8682;
  assign n9131 = ~n5351 & n7515;
  assign n9132 = ~n1798 & n8029;
  assign n9133 = ~n1638 & n7520;
  assign n9134 = ~n9132 & ~n9133;
  assign n9135 = ~n1726 & n7518;
  assign n9136 = n9134 & ~n9135;
  assign n9137 = ~n9131 & n9136;
  assign n9138 = n9137 ^ x5;
  assign n9140 = n9139 ^ n9138;
  assign n9149 = n8759 ^ n8698;
  assign n9141 = ~n5703 & n7515;
  assign n9142 = ~n1726 & n8029;
  assign n9143 = ~n1638 & n7518;
  assign n9144 = ~n9142 & ~n9143;
  assign n9145 = ~n1544 & n7520;
  assign n9146 = n9144 & ~n9145;
  assign n9147 = ~n9141 & n9146;
  assign n9148 = n9147 ^ x5;
  assign n9150 = n9149 ^ n9148;
  assign n9159 = n8756 ^ n8709;
  assign n9151 = ~n5069 & n7515;
  assign n9152 = ~n734 & n7520;
  assign n9153 = ~n1638 & n8029;
  assign n9154 = ~n9152 & ~n9153;
  assign n9155 = ~n1544 & n7518;
  assign n9156 = n9154 & ~n9155;
  assign n9157 = ~n9151 & n9156;
  assign n9158 = n9157 ^ x5;
  assign n9160 = n9159 ^ n9158;
  assign n9162 = ~n5416 & n7515;
  assign n9163 = ~n882 & n7520;
  assign n9164 = ~n1544 & n8029;
  assign n9165 = ~n9163 & ~n9164;
  assign n9166 = ~n734 & n7518;
  assign n9167 = n9165 & ~n9166;
  assign n9168 = ~n9162 & n9167;
  assign n9169 = n9168 ^ x5;
  assign n9161 = n8753 ^ n8727;
  assign n9170 = n9169 ^ n9161;
  assign n9175 = ~n5465 & n7515;
  assign n9176 = ~n970 & n7520;
  assign n9177 = ~n882 & n7518;
  assign n9178 = ~n9176 & ~n9177;
  assign n9179 = ~n734 & n8029;
  assign n9180 = n9178 & ~n9179;
  assign n9181 = ~n9175 & n9180;
  assign n9182 = n9181 ^ x5;
  assign n9171 = ~n1319 & n5812;
  assign n9172 = n9171 ^ x8;
  assign n9173 = n9172 ^ n8751;
  assign n9174 = n9173 ^ n8734;
  assign n9183 = n9182 ^ n9174;
  assign n9186 = ~n5481 & n7515;
  assign n9187 = ~n882 & n8029;
  assign n9188 = ~n970 & n7518;
  assign n9189 = ~n9187 & ~n9188;
  assign n9190 = ~n1097 & n7520;
  assign n9191 = n9189 & ~n9190;
  assign n9192 = ~n9186 & n9191;
  assign n9193 = n9192 ^ x5;
  assign n9184 = x8 & ~n8749;
  assign n9185 = n9184 ^ n8746;
  assign n9194 = n9193 ^ n9185;
  assign n9204 = ~n5564 & n7515;
  assign n9205 = ~n1097 & n7518;
  assign n9206 = ~n1414 & n7520;
  assign n9207 = ~n9205 & ~n9206;
  assign n9208 = ~n970 & n8029;
  assign n9209 = n9207 & ~n9208;
  assign n9210 = ~n9204 & n9209;
  assign n9211 = n9210 ^ x5;
  assign n9195 = ~x7 & n6311;
  assign n9196 = ~n1208 & ~n6313;
  assign n9197 = x7 & ~n6311;
  assign n9198 = ~n9196 & n9197;
  assign n9199 = ~n9195 & ~n9198;
  assign n9200 = ~n1319 & ~n9199;
  assign n9201 = x7 & ~n1319;
  assign n9202 = n8747 & ~n9201;
  assign n9203 = ~n9200 & ~n9202;
  assign n9212 = n9211 ^ n9203;
  assign n9213 = ~n5579 & n7515;
  assign n9214 = ~n1097 & n8029;
  assign n9215 = ~n1414 & n7518;
  assign n9216 = ~n9214 & ~n9215;
  assign n9217 = ~n1208 & n7520;
  assign n9218 = n9216 & ~n9217;
  assign n9219 = ~n9213 & n9218;
  assign n9222 = n5630 & n7513;
  assign n9223 = ~n1414 & n7514;
  assign n9224 = ~n9222 & n9223;
  assign n9225 = ~n1319 & n7520;
  assign n9226 = ~n9224 & ~n9225;
  assign n9227 = n5634 & n7515;
  assign n9228 = ~n7518 & ~n9227;
  assign n9229 = ~n1208 & ~n9228;
  assign n9230 = n9226 & ~n9229;
  assign n9231 = ~n1208 & n7514;
  assign n9232 = n1319 & ~n9231;
  assign n9233 = ~n7519 & ~n9232;
  assign n9234 = x5 & ~n9233;
  assign n9235 = n9230 & n9234;
  assign n9236 = x5 & ~x6;
  assign n9237 = ~n1319 & n9236;
  assign n9238 = ~n9235 & ~n9237;
  assign n9220 = ~x5 & x6;
  assign n9221 = ~n1319 & n9220;
  assign n9239 = n9238 ^ n9221;
  assign n9240 = ~n9219 & ~n9239;
  assign n9241 = n9240 ^ n9238;
  assign n9242 = n9241 ^ n9203;
  assign n9243 = n9212 & ~n9242;
  assign n9244 = n9243 ^ n9211;
  assign n9245 = n9244 ^ n9193;
  assign n9246 = ~n9194 & n9245;
  assign n9247 = n9246 ^ n9244;
  assign n9248 = n9247 ^ n9182;
  assign n9249 = ~n9183 & n9248;
  assign n9250 = n9249 ^ n9247;
  assign n9251 = n9250 ^ n9169;
  assign n9252 = n9170 & n9251;
  assign n9253 = n9252 ^ n9250;
  assign n9254 = n9253 ^ n9159;
  assign n9255 = ~n9160 & n9254;
  assign n9256 = n9255 ^ n9253;
  assign n9257 = n9256 ^ n9149;
  assign n9258 = ~n9150 & n9257;
  assign n9259 = n9258 ^ n9256;
  assign n9260 = n9259 ^ n9139;
  assign n9261 = ~n9140 & n9260;
  assign n9262 = n9261 ^ n9259;
  assign n9263 = n9262 ^ n9129;
  assign n9264 = ~n9130 & n9263;
  assign n9265 = n9264 ^ n9262;
  assign n9266 = n9265 ^ n9119;
  assign n9267 = n9120 & ~n9266;
  assign n9268 = n9267 ^ n9265;
  assign n9269 = n9268 ^ n9109;
  assign n9270 = ~n9110 & n9269;
  assign n9271 = n9270 ^ n9268;
  assign n9272 = n9271 ^ n9099;
  assign n9273 = n9100 & ~n9272;
  assign n9274 = n9273 ^ n9271;
  assign n9275 = n9274 ^ n9089;
  assign n9276 = n9090 & ~n9275;
  assign n9277 = n9276 ^ n9274;
  assign n9278 = n9277 ^ n9079;
  assign n9279 = ~n9080 & n9278;
  assign n9280 = n9279 ^ n9277;
  assign n9281 = n9280 ^ n9069;
  assign n9282 = n9070 & ~n9281;
  assign n9283 = n9282 ^ n9280;
  assign n9284 = n9283 ^ n9058;
  assign n9285 = n9060 & ~n9284;
  assign n9286 = n9285 ^ n9059;
  assign n9287 = n9286 ^ n9048;
  assign n9288 = ~n9050 & ~n9287;
  assign n9289 = n9288 ^ n9049;
  assign n9290 = n9289 ^ n9037;
  assign n9291 = n9040 & n9290;
  assign n9292 = n9291 ^ n9039;
  assign n9293 = n9292 ^ n9027;
  assign n9294 = ~n9029 & ~n9293;
  assign n9295 = n9294 ^ n9028;
  assign n9296 = n9295 ^ n9017;
  assign n9297 = ~n9019 & n9296;
  assign n9298 = n9297 ^ n9018;
  assign n9299 = n9298 ^ n9008;
  assign n9300 = ~n9009 & ~n9299;
  assign n9301 = n9300 ^ n9298;
  assign n9302 = n9301 ^ n8998;
  assign n9303 = ~n8999 & ~n9302;
  assign n9304 = n9303 ^ n9301;
  assign n9305 = ~n8989 & ~n9304;
  assign n9306 = ~n8988 & ~n9305;
  assign n9307 = n8989 & n9304;
  assign n9308 = ~n3666 & n7515;
  assign n9309 = ~n2718 & n7520;
  assign n9310 = ~n2861 & n7518;
  assign n9311 = ~n9309 & ~n9310;
  assign n9312 = ~n566 & n8029;
  assign n9313 = n9311 & ~n9312;
  assign n9314 = ~n9308 & n9313;
  assign n9315 = n9314 ^ x5;
  assign n9316 = ~n9307 & n9315;
  assign n9317 = n9306 & ~n9316;
  assign n9318 = ~n8979 & ~n8987;
  assign n9319 = ~n9317 & ~n9318;
  assign n9320 = n9319 ^ n8977;
  assign n9321 = ~n8978 & n9320;
  assign n9322 = n9321 ^ n9319;
  assign n9323 = n9322 ^ n8967;
  assign n9324 = n8968 & ~n9323;
  assign n9325 = n9324 ^ n9322;
  assign n9326 = n9325 ^ n8957;
  assign n9327 = n8958 & ~n9326;
  assign n9328 = n9327 ^ n9325;
  assign n9329 = n9328 ^ n8947;
  assign n9330 = ~n8948 & n9329;
  assign n9331 = n9330 ^ n9328;
  assign n9342 = n9341 ^ n9331;
  assign n8933 = n33 & ~n3411;
  assign n8934 = n8933 ^ x1;
  assign n8935 = n8934 ^ n3431;
  assign n8929 = n3404 ^ x2;
  assign n8928 = x2 & n3351;
  assign n8930 = n8929 ^ n8928;
  assign n8931 = ~x1 & ~n8930;
  assign n8932 = n8931 ^ n8929;
  assign n8936 = n8935 ^ n8932;
  assign n8937 = ~x0 & n8936;
  assign n8938 = n8937 ^ n8935;
  assign n9343 = n9342 ^ n8938;
  assign n9355 = n9328 ^ n8948;
  assign n9349 = n33 & ~n5769;
  assign n9350 = n9349 ^ x1;
  assign n9351 = n9350 ^ n3404;
  assign n9344 = n3351 ^ x2;
  assign n9345 = x1 & ~n9344;
  assign n9346 = ~x1 & x2;
  assign n9347 = n3270 & n9346;
  assign n9348 = ~n9345 & ~n9347;
  assign n9352 = n9351 ^ n9348;
  assign n9353 = ~x0 & n9352;
  assign n9354 = n9353 ^ n9351;
  assign n9356 = n9355 ^ n9354;
  assign n9367 = n9325 ^ n8958;
  assign n9361 = n33 & ~n3988;
  assign n9362 = n9361 ^ x1;
  assign n9363 = n9362 ^ n3351;
  assign n9357 = n3270 ^ x2;
  assign n9358 = x1 & ~n9357;
  assign n9359 = n3196 & n9346;
  assign n9360 = ~n9358 & ~n9359;
  assign n9364 = n9363 ^ n9360;
  assign n9365 = ~x0 & n9364;
  assign n9366 = n9365 ^ n9363;
  assign n9368 = n9367 ^ n9366;
  assign n9370 = n9319 ^ n8978;
  assign n9372 = n3196 ^ x2;
  assign n9371 = n3196 ^ x1;
  assign n9373 = n9372 ^ n9371;
  assign n9374 = ~n3107 & n9373;
  assign n9375 = n9374 ^ n9372;
  assign n9376 = x0 & ~n9375;
  assign n9377 = n3098 ^ x2;
  assign n9379 = ~n9377 & n9378;
  assign n9380 = ~x0 & n9346;
  assign n9381 = n2954 & n9380;
  assign n9382 = ~n9379 & ~n9381;
  assign n9383 = ~n9376 & n9382;
  assign n9384 = n9370 & n9383;
  assign n9385 = n8987 ^ n8979;
  assign n9386 = n9304 ^ n8989;
  assign n9387 = ~n9315 & n9386;
  assign n9388 = n9385 & n9387;
  assign n9390 = n9385 ^ n9307;
  assign n9389 = n9315 & ~n9386;
  assign n9391 = n9390 ^ n9389;
  assign n9396 = n33 & ~n3973;
  assign n9397 = n9396 ^ x1;
  assign n9398 = n9397 ^ n3098;
  assign n9392 = n2954 ^ x2;
  assign n9393 = x1 & ~n9392;
  assign n9394 = n3037 & n9346;
  assign n9395 = ~n9393 & ~n9394;
  assign n9399 = n9398 ^ n9395;
  assign n9400 = ~x0 & n9399;
  assign n9401 = n9400 ^ n9398;
  assign n9402 = n9401 ^ n9389;
  assign n9403 = ~n9391 & ~n9402;
  assign n9404 = n9403 ^ n9390;
  assign n9405 = ~n9388 & n9404;
  assign n9406 = n9388 & n9401;
  assign n9418 = n9301 ^ n8999;
  assign n9408 = n3037 ^ x1;
  assign n9407 = n3037 ^ x2;
  assign n9409 = n9408 ^ n9407;
  assign n9410 = ~n3631 & n9409;
  assign n9411 = n9410 ^ n9408;
  assign n9412 = x0 & ~n9411;
  assign n9413 = n368 ^ x2;
  assign n9414 = n9378 & ~n9413;
  assign n9415 = n566 & n9380;
  assign n9416 = ~n9414 & ~n9415;
  assign n9417 = ~n9412 & n9416;
  assign n9419 = n9418 ^ n9417;
  assign n9813 = n9298 ^ n9009;
  assign n9797 = n9295 ^ n9019;
  assign n9437 = n9292 ^ n9029;
  assign n9427 = x2 & ~n4466;
  assign n9428 = ~x2 & n2861;
  assign n9429 = x0 & ~n9428;
  assign n9430 = ~n9427 & n9429;
  assign n9431 = ~x0 & x2;
  assign n9432 = n2786 & n9431;
  assign n9433 = ~n9430 & ~n9432;
  assign n9420 = ~x2 & n4466;
  assign n9421 = x2 & ~n2861;
  assign n9422 = x0 & ~n9421;
  assign n9423 = ~n9420 & n9422;
  assign n9424 = n2718 ^ x2;
  assign n9425 = ~x0 & ~n9424;
  assign n9426 = ~n9423 & ~n9425;
  assign n9434 = n9433 ^ n9426;
  assign n9435 = x1 & n9434;
  assign n9436 = n9435 ^ n9433;
  assign n9438 = n9437 ^ n9436;
  assign n9777 = n9289 ^ n9040;
  assign n9762 = n9286 ^ n9050;
  assign n9747 = n9283 ^ n9060;
  assign n9734 = n9280 ^ n9070;
  assign n9718 = n9277 ^ n9080;
  assign n9702 = n9274 ^ n9090;
  assign n9687 = n9271 ^ n9100;
  assign n9440 = n9265 ^ n9120;
  assign n9441 = n2247 ^ x1;
  assign n9442 = n4252 & ~n9441;
  assign n9443 = x0 & ~n9442;
  assign n9444 = n2247 ^ x2;
  assign n9445 = ~n4252 & ~n9444;
  assign n9446 = n9443 & ~n9445;
  assign n9447 = x2 & n2065;
  assign n9449 = ~n9447 & n9448;
  assign n9450 = n2175 ^ x2;
  assign n9451 = n9378 & n9450;
  assign n9452 = ~n9449 & ~n9451;
  assign n9453 = ~n9446 & n9452;
  assign n9454 = ~n9440 & ~n9453;
  assign n9455 = n9262 ^ n9130;
  assign n9456 = n2175 ^ x1;
  assign n9457 = n9456 ^ n9450;
  assign n9458 = n4506 & n9457;
  assign n9459 = n9458 ^ n9450;
  assign n9460 = x0 & n9459;
  assign n9461 = n2065 ^ x2;
  assign n9462 = n9378 & n9461;
  assign n9463 = x2 & n1974;
  assign n9464 = n9448 & ~n9463;
  assign n9465 = ~n9462 & ~n9464;
  assign n9466 = ~n9460 & n9465;
  assign n9467 = n9455 & ~n9466;
  assign n9468 = ~n9454 & ~n9467;
  assign n9469 = ~n9455 & n9466;
  assign n9655 = n9259 ^ n9140;
  assign n9640 = n9256 ^ n9150;
  assign n9471 = n9250 ^ n9170;
  assign n9472 = n33 & ~n5350;
  assign n9473 = n9472 ^ x1;
  assign n9474 = n9473 ^ n1798;
  assign n9475 = x0 & n9474;
  assign n9476 = n1726 ^ x2;
  assign n9477 = n9378 & n9476;
  assign n9478 = x2 & n1638;
  assign n9479 = n9448 & ~n9478;
  assign n9480 = ~n9477 & ~n9479;
  assign n9481 = ~n9475 & n9480;
  assign n9482 = n9471 & n9481;
  assign n9483 = n9247 ^ n9183;
  assign n9488 = n33 & ~n5702;
  assign n9489 = n9488 ^ x1;
  assign n9490 = n9489 ^ n1726;
  assign n9484 = n1638 ^ x2;
  assign n9485 = x1 & ~n9484;
  assign n9486 = n1544 & n9346;
  assign n9487 = ~n9485 & ~n9486;
  assign n9491 = n9490 ^ n9487;
  assign n9492 = ~x0 & n9491;
  assign n9493 = n9492 ^ n9490;
  assign n9494 = ~n9483 & ~n9493;
  assign n9495 = ~n9482 & ~n9494;
  assign n9496 = n9241 ^ n9212;
  assign n9504 = x2 & ~n5416;
  assign n9505 = ~x2 & n1544;
  assign n9506 = x0 & ~n9505;
  assign n9507 = ~n9504 & n9506;
  assign n9508 = n882 & n9431;
  assign n9509 = ~n9507 & ~n9508;
  assign n9497 = ~x2 & n5416;
  assign n9498 = x2 & ~n1544;
  assign n9499 = x0 & ~n9498;
  assign n9500 = ~n9497 & n9499;
  assign n9501 = n734 ^ x2;
  assign n9502 = ~x0 & ~n9501;
  assign n9503 = ~n9500 & ~n9502;
  assign n9510 = n9509 ^ n9503;
  assign n9511 = x1 & n9510;
  assign n9512 = n9511 ^ n9509;
  assign n9513 = n9496 & n9512;
  assign n9514 = x5 & n9233;
  assign n9515 = n9514 ^ n9230;
  assign n9521 = n33 & ~n5480;
  assign n9522 = n9521 ^ x1;
  assign n9523 = n9522 ^ n882;
  assign n9517 = x2 & n1097;
  assign n9516 = n970 ^ x2;
  assign n9518 = n9517 ^ n9516;
  assign n9519 = x1 & ~n9518;
  assign n9520 = n9519 ^ n9517;
  assign n9524 = n9523 ^ n9520;
  assign n9525 = ~x0 & ~n9524;
  assign n9526 = n9525 ^ n9523;
  assign n9527 = n9515 & n9526;
  assign n9539 = n33 & ~n5578;
  assign n9540 = n9539 ^ x1;
  assign n9541 = n9540 ^ n1097;
  assign n9542 = x0 & n9541;
  assign n9543 = x0 & n7514;
  assign n9544 = n1414 ^ x3;
  assign n9545 = n7514 & n9544;
  assign n9546 = x1 & n9545;
  assign n9547 = ~n9543 & ~n9546;
  assign n9548 = ~n1319 & ~n9547;
  assign n9549 = x3 & ~n1319;
  assign n9550 = n9448 & ~n9549;
  assign n9551 = ~n5634 & ~n9550;
  assign n9552 = x2 & n1208;
  assign n9553 = ~n9551 & n9552;
  assign n9554 = ~n9548 & ~n9553;
  assign n9555 = ~n9542 & ~n9554;
  assign n9528 = x2 & x3;
  assign n9529 = ~x4 & n9528;
  assign n9530 = ~x2 & ~x3;
  assign n9531 = ~n1208 & ~n9530;
  assign n9532 = x4 & ~n9528;
  assign n9533 = ~n9531 & n9532;
  assign n9534 = ~n9529 & ~n9533;
  assign n9535 = x4 & ~n1319;
  assign n9536 = n9231 & ~n9535;
  assign n9537 = n9534 & ~n9536;
  assign n9538 = ~n9232 & ~n9537;
  assign n9556 = n9555 ^ n9538;
  assign n9561 = n33 & ~n5563;
  assign n9562 = n9561 ^ x1;
  assign n9563 = n9562 ^ n970;
  assign n9557 = n1097 ^ x2;
  assign n9558 = x1 & ~n9557;
  assign n9559 = n1414 & n9346;
  assign n9560 = ~n9558 & ~n9559;
  assign n9564 = n9563 ^ n9560;
  assign n9565 = ~x0 & n9564;
  assign n9566 = n9565 ^ n9563;
  assign n9567 = n9566 ^ n9538;
  assign n9568 = n9556 & n9567;
  assign n9569 = n9568 ^ n9555;
  assign n9570 = ~n9527 & n9569;
  assign n9571 = ~n9515 & ~n9526;
  assign n9572 = x1 & ~n1419;
  assign n9573 = ~n734 & ~n9572;
  assign n9574 = n734 & n1418;
  assign n9575 = x0 & ~n9574;
  assign n9576 = x1 & n734;
  assign n9577 = n882 & n9576;
  assign n9578 = ~n2362 & ~n9577;
  assign n9579 = n9575 & n9578;
  assign n9580 = ~n9573 & n9579;
  assign n9581 = x1 & ~n882;
  assign n9582 = ~n9575 & ~n9581;
  assign n9583 = ~x2 & ~n9582;
  assign n9584 = ~n9580 & n9583;
  assign n9585 = ~x1 & n5464;
  assign n9586 = n9585 ^ n734;
  assign n9587 = n8890 & n9586;
  assign n9588 = ~x1 & ~n970;
  assign n9589 = n9431 & ~n9588;
  assign n9590 = ~n9581 & n9589;
  assign n9591 = ~n9587 & ~n9590;
  assign n9592 = ~n9584 & n9591;
  assign n9593 = ~x6 & ~n1319;
  assign n9594 = n9593 ^ n9235;
  assign n9595 = ~x5 & n1319;
  assign n9596 = ~n9594 & ~n9595;
  assign n9597 = n9596 ^ n9219;
  assign n9598 = ~n9592 & ~n9597;
  assign n9599 = ~n9571 & ~n9598;
  assign n9600 = ~n9570 & n9599;
  assign n9601 = n9592 & n9597;
  assign n9602 = ~n9600 & ~n9601;
  assign n9603 = ~n9513 & n9602;
  assign n9604 = n33 & ~n5068;
  assign n9605 = n9604 ^ x1;
  assign n9606 = n9605 ^ n1638;
  assign n9607 = x0 & n9606;
  assign n9608 = x2 & n734;
  assign n9609 = n9448 & ~n9608;
  assign n9610 = n1544 ^ x2;
  assign n9611 = n9378 & n9610;
  assign n9612 = ~n9609 & ~n9611;
  assign n9613 = ~n9607 & n9612;
  assign n9614 = n9244 ^ n9194;
  assign n9615 = n9613 & ~n9614;
  assign n9616 = ~n9496 & ~n9512;
  assign n9617 = ~n9615 & ~n9616;
  assign n9618 = ~n9603 & n9617;
  assign n9619 = n9483 & n9493;
  assign n9620 = ~n9613 & n9614;
  assign n9621 = ~n9619 & ~n9620;
  assign n9622 = ~n9618 & n9621;
  assign n9623 = n9495 & ~n9622;
  assign n9624 = ~n9471 & ~n9481;
  assign n9625 = ~n9623 & ~n9624;
  assign n9470 = n9253 ^ n9160;
  assign n9626 = n9625 ^ n9470;
  assign n9631 = n33 & ~n5023;
  assign n9632 = n9631 ^ x1;
  assign n9633 = n9632 ^ n1878;
  assign n9627 = x1 & ~n1798;
  assign n9628 = ~n1726 & n9346;
  assign n9629 = ~n9627 & ~n9628;
  assign n9630 = n9629 ^ x2;
  assign n9634 = n9633 ^ n9630;
  assign n9635 = ~x0 & n9634;
  assign n9636 = n9635 ^ n9633;
  assign n9637 = n9636 ^ n9470;
  assign n9638 = ~n9626 & ~n9637;
  assign n9639 = n9638 ^ n9625;
  assign n9641 = n9640 ^ n9639;
  assign n9646 = n33 & ~n4592;
  assign n9647 = n9646 ^ x1;
  assign n9648 = n9647 ^ n1974;
  assign n9642 = n1878 ^ x2;
  assign n9643 = x1 & ~n9642;
  assign n9644 = n1798 & n9346;
  assign n9645 = ~n9643 & ~n9644;
  assign n9649 = n9648 ^ n9645;
  assign n9650 = ~x0 & n9649;
  assign n9651 = n9650 ^ n9648;
  assign n9652 = n9651 ^ n9640;
  assign n9653 = ~n9641 & ~n9652;
  assign n9654 = n9653 ^ n9639;
  assign n9656 = n9655 ^ n9654;
  assign n9657 = x2 & n1878;
  assign n9658 = n9448 & ~n9657;
  assign n9659 = n1974 ^ x2;
  assign n9660 = n9378 & n9659;
  assign n9661 = ~n9658 & ~n9660;
  assign n9662 = n33 & ~n5166;
  assign n9663 = n9662 ^ x1;
  assign n9664 = n9663 ^ n2065;
  assign n9665 = x0 & n9664;
  assign n9666 = n9661 & ~n9665;
  assign n9667 = n9666 ^ n9655;
  assign n9668 = ~n9656 & n9667;
  assign n9669 = n9668 ^ n9654;
  assign n9670 = ~n9469 & ~n9669;
  assign n9671 = n9468 & ~n9670;
  assign n9672 = n9440 & n9453;
  assign n9673 = ~n9671 & ~n9672;
  assign n9439 = n9268 ^ n9110;
  assign n9674 = n9673 ^ n9439;
  assign n9678 = n33 & ~n4322;
  assign n9679 = n9678 ^ x1;
  assign n9680 = n9679 ^ n2357;
  assign n9675 = n2175 & n9346;
  assign n9676 = x1 & ~n9444;
  assign n9677 = ~n9675 & ~n9676;
  assign n9681 = n9680 ^ n9677;
  assign n9682 = ~x0 & n9681;
  assign n9683 = n9682 ^ n9680;
  assign n9684 = n9683 ^ n9439;
  assign n9685 = n9674 & ~n9684;
  assign n9686 = n9685 ^ n9673;
  assign n9688 = n9687 ^ n9686;
  assign n9689 = n33 & ~n4292;
  assign n9690 = n9689 ^ x1;
  assign n9691 = n9690 ^ n2423;
  assign n9692 = x0 & n9691;
  assign n9693 = n2357 ^ x2;
  assign n9694 = x1 & ~n9693;
  assign n9695 = ~x0 & ~n9694;
  assign n9696 = n2247 & n9346;
  assign n9697 = n9695 & ~n9696;
  assign n9698 = ~n9692 & ~n9697;
  assign n9699 = n9698 ^ n9687;
  assign n9700 = ~n9688 & ~n9699;
  assign n9701 = n9700 ^ n9686;
  assign n9703 = n9702 ^ n9701;
  assign n9705 = n2482 ^ x1;
  assign n9704 = n2482 ^ x2;
  assign n9706 = n9705 ^ n9704;
  assign n9707 = ~n4433 & n9706;
  assign n9708 = n9707 ^ n9705;
  assign n9709 = x0 & ~n9708;
  assign n9710 = n2423 ^ x2;
  assign n9711 = n9378 & ~n9710;
  assign n9712 = n2357 & n9380;
  assign n9713 = ~n9711 & ~n9712;
  assign n9714 = ~n9709 & n9713;
  assign n9715 = n9714 ^ n9702;
  assign n9716 = ~n9703 & n9715;
  assign n9717 = n9716 ^ n9701;
  assign n9719 = n9718 ^ n9717;
  assign n9721 = n2612 ^ x2;
  assign n9720 = n2612 ^ x1;
  assign n9722 = n9721 ^ n9720;
  assign n9723 = n4333 & n9722;
  assign n9724 = n9723 ^ n9721;
  assign n9725 = x0 & n9724;
  assign n9726 = n9378 & n9704;
  assign n9727 = x2 & n2423;
  assign n9728 = n9448 & ~n9727;
  assign n9729 = ~n9726 & ~n9728;
  assign n9730 = ~n9725 & n9729;
  assign n9731 = n9730 ^ n9718;
  assign n9732 = n9719 & n9731;
  assign n9733 = n9732 ^ n9717;
  assign n9735 = n9734 ^ n9733;
  assign n9736 = n33 & ~n4311;
  assign n9737 = n9736 ^ x1;
  assign n9738 = n9737 ^ n2574;
  assign n9739 = x0 & ~n9738;
  assign n9740 = n9378 & ~n9721;
  assign n9741 = n2482 & n9380;
  assign n9742 = ~n9740 & ~n9741;
  assign n9743 = ~n9739 & n9742;
  assign n9744 = n9743 ^ n9734;
  assign n9745 = ~n9735 & n9744;
  assign n9746 = n9745 ^ n9733;
  assign n9748 = n9747 ^ n9746;
  assign n9749 = n33 & ~n4452;
  assign n9750 = n9749 ^ x1;
  assign n9751 = n9750 ^ n2669;
  assign n9752 = x0 & ~n9751;
  assign n9753 = x1 & ~n2574;
  assign n9754 = n9753 ^ x2;
  assign n9755 = ~x1 & ~n2612;
  assign n9756 = ~x0 & ~n9755;
  assign n9757 = n9754 & n9756;
  assign n9758 = ~n9752 & ~n9757;
  assign n9759 = n9758 ^ n9747;
  assign n9760 = n9748 & ~n9759;
  assign n9761 = n9760 ^ n9746;
  assign n9763 = n9762 ^ n9761;
  assign n9768 = n33 & ~n4652;
  assign n9769 = n9768 ^ x1;
  assign n9770 = n9769 ^ n2786;
  assign n9764 = n2669 ^ x2;
  assign n9765 = x1 & ~n9764;
  assign n9766 = n2574 & n9346;
  assign n9767 = ~n9765 & ~n9766;
  assign n9771 = n9770 ^ n9767;
  assign n9772 = ~x0 & n9771;
  assign n9773 = n9772 ^ n9770;
  assign n9774 = n9773 ^ n9762;
  assign n9775 = ~n9763 & n9774;
  assign n9776 = n9775 ^ n9761;
  assign n9778 = n9777 ^ n9776;
  assign n9784 = n2718 ^ x1;
  assign n9785 = n9784 ^ n9424;
  assign n9786 = n4494 & n9785;
  assign n9787 = n9786 ^ n9424;
  assign n9780 = x2 & n2669;
  assign n9779 = n2786 ^ x2;
  assign n9781 = n9780 ^ n9779;
  assign n9782 = x1 & ~n9781;
  assign n9783 = n9782 ^ n9780;
  assign n9788 = n9787 ^ n9783;
  assign n9789 = ~x0 & ~n9788;
  assign n9790 = n9789 ^ n9787;
  assign n9791 = n9790 ^ n9777;
  assign n9792 = ~n9778 & n9791;
  assign n9793 = n9792 ^ n9776;
  assign n9794 = n9793 ^ n9436;
  assign n9795 = ~n9438 & ~n9794;
  assign n9796 = n9795 ^ n9437;
  assign n9798 = n9797 ^ n9796;
  assign n9804 = n33 & ~n3665;
  assign n9805 = n9804 ^ x1;
  assign n9806 = n9805 ^ n566;
  assign n9800 = x2 & n2718;
  assign n9799 = n2861 ^ x2;
  assign n9801 = n9800 ^ n9799;
  assign n9802 = x1 & ~n9801;
  assign n9803 = n9802 ^ n9800;
  assign n9807 = n9806 ^ n9803;
  assign n9808 = ~x0 & ~n9807;
  assign n9809 = n9808 ^ n9806;
  assign n9810 = n9809 ^ n9797;
  assign n9811 = ~n9798 & ~n9810;
  assign n9812 = n9811 ^ n9796;
  assign n9814 = n9813 ^ n9812;
  assign n9815 = n368 ^ x1;
  assign n9816 = n9815 ^ n9413;
  assign n9817 = ~n3748 & n9816;
  assign n9818 = n9817 ^ n9413;
  assign n9819 = x0 & n9818;
  assign n9820 = n566 ^ x2;
  assign n9821 = x1 & ~n9820;
  assign n9822 = n2861 & n9346;
  assign n9823 = ~x0 & ~n9822;
  assign n9824 = ~n9821 & n9823;
  assign n9825 = ~n9819 & ~n9824;
  assign n9826 = n9825 ^ n9813;
  assign n9827 = n9814 & ~n9826;
  assign n9828 = n9827 ^ n9812;
  assign n9829 = n9828 ^ n9417;
  assign n9830 = ~n9419 & n9829;
  assign n9831 = n9830 ^ n9418;
  assign n9835 = n33 & ~n3776;
  assign n9836 = n9835 ^ x1;
  assign n9837 = n9836 ^ n2954;
  assign n9832 = n368 & n9346;
  assign n9833 = x1 & ~n9407;
  assign n9834 = ~n9832 & ~n9833;
  assign n9838 = n9837 ^ n9834;
  assign n9839 = ~x0 & n9838;
  assign n9840 = n9839 ^ n9837;
  assign n9841 = n9831 & ~n9840;
  assign n9842 = ~n9406 & n9841;
  assign n9843 = ~n9405 & ~n9842;
  assign n9844 = ~n9384 & ~n9843;
  assign n9845 = ~n9831 & n9840;
  assign n9846 = n9845 ^ n9401;
  assign n9847 = ~n9387 & ~n9390;
  assign n9848 = n9847 ^ n9845;
  assign n9849 = n9846 & ~n9848;
  assign n9850 = n9849 ^ n9401;
  assign n9851 = n9844 & ~n9850;
  assign n9852 = ~n9370 & ~n9383;
  assign n9853 = ~n9851 & ~n9852;
  assign n9369 = n9322 ^ n8968;
  assign n9854 = n9853 ^ n9369;
  assign n9855 = n3270 ^ x1;
  assign n9856 = n9855 ^ n9357;
  assign n9857 = n3198 & n9856;
  assign n9858 = n9857 ^ n9357;
  assign n9859 = x0 & n9858;
  assign n9860 = x2 & n3098;
  assign n9861 = n9448 & ~n9860;
  assign n9862 = n9372 & n9378;
  assign n9863 = ~n9861 & ~n9862;
  assign n9864 = ~n9859 & n9863;
  assign n9865 = n9864 ^ n9369;
  assign n9866 = ~n9854 & ~n9865;
  assign n9867 = n9866 ^ n9853;
  assign n9868 = n9867 ^ n9367;
  assign n9869 = n9368 & ~n9868;
  assign n9870 = n9869 ^ n9867;
  assign n9871 = n9870 ^ n9355;
  assign n9872 = ~n9356 & n9871;
  assign n9873 = n9872 ^ n9870;
  assign n9874 = n9873 ^ n9342;
  assign n9875 = n9343 & ~n9874;
  assign n9876 = n9875 ^ n9873;
  assign n9887 = n9886 ^ n9876;
  assign n9892 = ~n3989 & n7515;
  assign n9893 = ~n3270 & n7518;
  assign n9894 = ~n3196 & n7520;
  assign n9895 = ~n3351 & n8029;
  assign n9896 = ~n9894 & ~n9895;
  assign n9897 = ~n9893 & n9896;
  assign n9898 = ~n9892 & n9897;
  assign n9899 = n9898 ^ x5;
  assign n9889 = n9340 ^ n9331;
  assign n9890 = n9341 & ~n9889;
  assign n9891 = n9890 ^ n9331;
  assign n9900 = n9899 ^ n9891;
  assign n9888 = n8846 ^ n8450;
  assign n9901 = n9900 ^ n9888;
  assign n9902 = n9901 ^ n9886;
  assign n9903 = n9887 & ~n9902;
  assign n9904 = n9903 ^ n9876;
  assign n9905 = ~n8927 & ~n9904;
  assign n9906 = n8902 ^ n8901;
  assign n9907 = ~n5770 & n7515;
  assign n9908 = ~n3270 & n7520;
  assign n9909 = ~n3404 & n8029;
  assign n9910 = ~n3351 & n7518;
  assign n9911 = ~n9909 & ~n9910;
  assign n9912 = ~n9908 & n9911;
  assign n9913 = ~n9907 & n9912;
  assign n9914 = n9913 ^ x5;
  assign n9915 = n9899 ^ n9888;
  assign n9916 = n9900 & ~n9915;
  assign n9917 = n9916 ^ n9891;
  assign n9918 = n9914 & n9917;
  assign n9919 = n8908 & ~n8926;
  assign n9920 = ~n9918 & ~n9919;
  assign n9921 = n9906 & n9920;
  assign n9922 = n9921 ^ n9919;
  assign n9923 = ~n9905 & ~n9922;
  assign n9924 = ~n9918 & n9919;
  assign n9925 = ~n9906 & ~n9924;
  assign n9926 = ~n9904 & ~n9925;
  assign n9927 = ~n8927 & n9906;
  assign n9928 = ~n9914 & ~n9917;
  assign n9929 = ~n9927 & ~n9928;
  assign n9930 = ~n9926 & n9929;
  assign n9931 = ~n9923 & ~n9930;
  assign n9932 = n9931 ^ n8906;
  assign n9933 = n8907 & ~n9932;
  assign n9934 = n9933 ^ n9931;
  assign n9935 = ~n8882 & ~n9934;
  assign n9936 = ~n8864 & n8870;
  assign n9937 = n8880 & ~n9936;
  assign n9938 = n8872 & ~n9937;
  assign n9939 = n8870 & n8875;
  assign n9940 = ~n9938 & ~n9939;
  assign n9941 = ~n9935 & n9940;
  assign n8022 = n8021 ^ n7524;
  assign n8023 = ~n7525 & n8022;
  assign n8024 = n8023 ^ n8021;
  assign n9942 = n9941 ^ n8024;
  assign n9943 = n7132 ^ n6851;
  assign n9944 = n9943 ^ n8024;
  assign n9945 = ~n9942 & ~n9944;
  assign n9946 = n9945 ^ n9941;
  assign n9947 = ~n7512 & n9946;
  assign n9948 = ~n8024 & n9941;
  assign n9949 = ~n9943 & n9948;
  assign n9950 = ~n7163 & ~n9949;
  assign n9951 = n8024 & ~n9941;
  assign n9952 = n9943 & n9951;
  assign n9953 = n7172 & ~n7510;
  assign n9954 = ~n9952 & ~n9953;
  assign n9955 = ~n9950 & n9954;
  assign n9956 = ~n9947 & ~n9955;
  assign n9957 = n7163 & n7511;
  assign n9958 = n9956 & ~n9957;
  assign n9959 = n9958 ^ n7138;
  assign n9960 = ~n7162 & n9959;
  assign n9961 = n9960 ^ n9958;
  assign n9962 = ~n6303 & n9961;
  assign n9963 = n7159 ^ n7142;
  assign n9964 = n7160 & ~n9963;
  assign n9965 = n9964 ^ n7145;
  assign n9966 = n7157 ^ n7148;
  assign n9967 = ~n7158 & n9966;
  assign n9968 = n9967 ^ n7148;
  assign n9969 = ~n9965 & ~n9968;
  assign n9970 = n6293 & n6302;
  assign n9971 = n9969 & ~n9970;
  assign n9972 = n6258 ^ n6016;
  assign n9973 = ~n9970 & n9972;
  assign n9974 = ~n9971 & ~n9973;
  assign n9975 = ~n9962 & ~n9974;
  assign n9976 = n9969 & n9972;
  assign n9977 = ~n9975 & ~n9976;
  assign n9978 = n9961 & ~n9973;
  assign n9979 = n9965 & n9968;
  assign n9980 = ~n6303 & ~n9972;
  assign n9981 = ~n9979 & ~n9980;
  assign n9982 = ~n9978 & n9981;
  assign n9983 = n9977 & ~n9982;
  assign n9984 = n9983 ^ n6261;
  assign n9985 = n6292 & ~n9984;
  assign n9986 = n9985 ^ n9983;
  assign n9987 = ~n5811 & ~n9986;
  assign n9991 = n6289 ^ n6281;
  assign n9992 = ~n6290 & n9991;
  assign n9993 = n9992 ^ n6284;
  assign n9988 = n6279 ^ n6264;
  assign n9989 = ~n6280 & n9988;
  assign n9990 = n9989 ^ n6264;
  assign n9994 = n9993 ^ n9990;
  assign n5736 = n5735 ^ n5298;
  assign n5737 = ~n5299 & ~n5736;
  assign n5738 = n5737 ^ n5735;
  assign n5286 = n5189 ^ n4991;
  assign n5278 = ~n3974 & n4673;
  assign n5279 = ~n3098 & n4688;
  assign n5280 = ~n2954 & n4685;
  assign n5281 = ~n5279 & ~n5280;
  assign n5282 = ~n3037 & ~n4681;
  assign n5283 = n5281 & ~n5282;
  assign n5284 = ~n5278 & n5283;
  assign n5285 = n5284 ^ x20;
  assign n5287 = n5286 ^ n5285;
  assign n5275 = n5274 ^ n5265;
  assign n5276 = n5266 & ~n5275;
  assign n5277 = n5276 ^ n5264;
  assign n5288 = n5287 ^ n5277;
  assign n5210 = ~n3989 & n4963;
  assign n5211 = ~n3270 & n4976;
  assign n5212 = ~n3351 & n4972;
  assign n5213 = ~n3196 & n4970;
  assign n5214 = ~n5212 & ~n5213;
  assign n5215 = ~n5211 & n5214;
  assign n5216 = ~n5210 & n5215;
  assign n5217 = n5216 ^ x17;
  assign n5289 = n5288 ^ n5217;
  assign n9995 = n5738 ^ n5289;
  assign n9996 = n9995 ^ n9990;
  assign n9997 = n9994 & n9996;
  assign n9998 = n9997 ^ n9993;
  assign n9999 = ~n9987 & ~n9998;
  assign n5790 = n5202 ^ n5201;
  assign n5771 = ~x17 & n4961;
  assign n5772 = ~n5770 & n5771;
  assign n5773 = ~n3270 & n4970;
  assign n5774 = ~n3351 & n4976;
  assign n5775 = ~n5773 & ~n5774;
  assign n5776 = x17 & n5775;
  assign n5777 = n3404 & n5776;
  assign n5778 = x16 & ~n5777;
  assign n5779 = ~n5772 & n5778;
  assign n5780 = n5770 & n5776;
  assign n5781 = ~n3404 & n5771;
  assign n5782 = ~x16 & ~n5781;
  assign n5783 = ~n5780 & n5782;
  assign n5784 = ~n5779 & ~n5783;
  assign n5785 = x17 & ~n4961;
  assign n5786 = n5785 ^ x17;
  assign n5787 = n5775 & ~n5786;
  assign n5788 = n5787 ^ x17;
  assign n5789 = ~n5784 & n5788;
  assign n5791 = n5790 ^ n5789;
  assign n5766 = n5286 ^ n5277;
  assign n5767 = n5287 & ~n5766;
  assign n5768 = n5767 ^ n5277;
  assign n5792 = n5791 ^ n5768;
  assign n5747 = ~n3875 & ~n5746;
  assign n5753 = ~n3431 & n5752;
  assign n5754 = ~n5747 & ~n5753;
  assign n5755 = x14 & ~n5754;
  assign n5759 = n5748 & n5758;
  assign n5760 = ~x14 & n5754;
  assign n5761 = n5760 ^ x13;
  assign n5762 = ~n5759 & ~n5761;
  assign n5763 = n5762 ^ x13;
  assign n5764 = ~n5755 & n5763;
  assign n5739 = n5738 ^ n5288;
  assign n5740 = n5289 & n5739;
  assign n5741 = n5740 ^ n5738;
  assign n5765 = n5764 ^ n5741;
  assign n10000 = n5792 ^ n5765;
  assign n10001 = ~n9999 & n10000;
  assign n10002 = n9987 & n9998;
  assign n10003 = n5811 & n9986;
  assign n10004 = n9990 & n9993;
  assign n10005 = ~n9995 & n10004;
  assign n10006 = ~n10000 & ~n10005;
  assign n10007 = ~n9990 & ~n9993;
  assign n10008 = n9995 & n10007;
  assign n10009 = ~n10006 & ~n10008;
  assign n10010 = ~n10003 & n10009;
  assign n10011 = ~n10002 & ~n10010;
  assign n10012 = ~n10001 & n10011;
  assign n5793 = n5792 ^ n5764;
  assign n5794 = n5765 & ~n5793;
  assign n5795 = n5794 ^ n5741;
  assign n10013 = n10012 ^ n5795;
  assign n10028 = n5205 ^ n4981;
  assign n10017 = ~x13 & ~n3875;
  assign n10018 = ~n3876 & ~n10017;
  assign n10019 = ~n5742 & ~n10018;
  assign n10020 = x14 & n3876;
  assign n10021 = n10019 & ~n10020;
  assign n10022 = n5744 ^ x14;
  assign n10023 = n5744 ^ x13;
  assign n10024 = ~n10022 & n10023;
  assign n10025 = ~n3875 & n10024;
  assign n10026 = n10025 ^ x14;
  assign n10027 = ~n10021 & n10026;
  assign n10029 = n10028 ^ n10027;
  assign n10014 = n5789 ^ n5768;
  assign n10015 = ~n5791 & ~n10014;
  assign n10016 = n10015 ^ n5790;
  assign n10030 = n10029 ^ n10016;
  assign n10031 = n10030 ^ n5795;
  assign n10032 = ~n10013 & n10031;
  assign n10033 = n10032 ^ n10012;
  assign n10034 = ~n5209 & ~n10033;
  assign n10035 = ~n3879 & n4963;
  assign n10036 = ~n3404 & n4970;
  assign n10037 = ~n3431 & n4976;
  assign n10038 = ~n10036 & ~n10037;
  assign n10039 = ~n3875 & n4972;
  assign n10040 = n10038 & ~n10039;
  assign n10041 = ~n10035 & n10040;
  assign n10042 = n10041 ^ x17;
  assign n10043 = n10028 ^ n10016;
  assign n10044 = n10029 & ~n10043;
  assign n10045 = n10044 ^ n10016;
  assign n10046 = n10042 & ~n10045;
  assign n10170 = n4673 & ~n5770;
  assign n10171 = ~n3270 & ~n4681;
  assign n10172 = ~n3351 & n4685;
  assign n10173 = ~n3404 & n4688;
  assign n10174 = ~n10172 & ~n10173;
  assign n10175 = ~n10171 & n10174;
  assign n10176 = ~n10170 & n10175;
  assign n10177 = n10176 ^ x20;
  assign n10167 = n4957 ^ n4864;
  assign n10168 = ~n4873 & n10167;
  assign n10169 = n10168 ^ n4957;
  assign n10178 = n10177 ^ n10169;
  assign n10148 = n4801 & n4825;
  assign n10149 = n4923 & ~n4933;
  assign n10150 = n10148 & ~n10149;
  assign n10151 = ~n4923 & n4933;
  assign n10152 = n4428 & ~n10151;
  assign n10153 = ~n10150 & n10152;
  assign n10154 = ~n4801 & ~n4825;
  assign n10155 = n10154 ^ n4933;
  assign n10156 = ~n4428 & ~n4923;
  assign n10157 = n10156 ^ n4933;
  assign n10158 = ~n10155 & n10157;
  assign n10159 = n10158 ^ n10154;
  assign n10160 = ~n10153 & ~n10159;
  assign n10137 = n41 & n4453;
  assign n10138 = n91 & n2574;
  assign n10139 = x31 & ~n10138;
  assign n10140 = ~n4931 & n10139;
  assign n10141 = ~n10137 & n10140;
  assign n10142 = n54 & ~n2574;
  assign n10143 = n41 & ~n2669;
  assign n10144 = ~n10142 & ~n10143;
  assign n10145 = ~x31 & ~n10144;
  assign n10146 = ~n10141 & ~n10145;
  assign n10104 = ~n1266 & n10103;
  assign n10105 = ~n627 & n1156;
  assign n10106 = n1874 & n4118;
  assign n10107 = n3038 & n10106;
  assign n10108 = n10105 & n10107;
  assign n10109 = n726 & n3699;
  assign n10110 = n10108 & n10109;
  assign n10111 = ~n506 & ~n540;
  assign n10112 = n2138 & n10111;
  assign n10113 = n457 & n883;
  assign n10114 = n10112 & n10113;
  assign n10115 = ~n416 & n1992;
  assign n10116 = n10114 & n10115;
  assign n10117 = n1189 & n10116;
  assign n10118 = n10110 & n10117;
  assign n10119 = n2159 & n3113;
  assign n10120 = n123 & n302;
  assign n10121 = n10119 & n10120;
  assign n10122 = n1738 & n10121;
  assign n10123 = ~n429 & ~n552;
  assign n10124 = ~n185 & ~n243;
  assign n10125 = n10123 & n10124;
  assign n10126 = ~n292 & ~n541;
  assign n10127 = ~n136 & ~n843;
  assign n10128 = n10126 & n10127;
  assign n10129 = n10125 & n10128;
  assign n10130 = n3174 & n4003;
  assign n10131 = n10129 & n10130;
  assign n10132 = n10122 & n10131;
  assign n10133 = n4378 & n10132;
  assign n10134 = n10118 & n10133;
  assign n10135 = n10104 & n10134;
  assign n10087 = n4428 ^ x14;
  assign n10088 = n4922 ^ n4428;
  assign n10089 = n10087 & ~n10088;
  assign n10090 = n10089 ^ x14;
  assign n10136 = n10135 ^ n10090;
  assign n10147 = n10146 ^ n10136;
  assign n10161 = n10160 ^ n10147;
  assign n10079 = n44 & ~n4466;
  assign n10080 = ~n2718 & n3277;
  assign n10081 = ~n2786 & n3275;
  assign n10082 = ~n2861 & n3280;
  assign n10083 = ~n10081 & ~n10082;
  assign n10084 = ~n10080 & n10083;
  assign n10085 = ~n10079 & n10084;
  assign n10086 = n10085 ^ x29;
  assign n10162 = n10161 ^ n10086;
  assign n10071 = n3285 & ~n3632;
  assign n10072 = ~n368 & n3435;
  assign n10073 = ~n3037 & n3437;
  assign n10074 = ~n10072 & ~n10073;
  assign n10075 = ~n566 & ~n3440;
  assign n10076 = n10074 & ~n10075;
  assign n10077 = ~n10071 & n10076;
  assign n10078 = n10077 ^ x26;
  assign n10163 = n10162 ^ n10078;
  assign n10068 = n4954 ^ n4935;
  assign n10069 = n4944 & n10068;
  assign n10070 = n10069 ^ n4954;
  assign n10164 = n10163 ^ n10070;
  assign n10060 = n3647 & n4478;
  assign n10061 = ~n2954 & n4480;
  assign n10062 = ~n3196 & n4487;
  assign n10063 = ~n10061 & ~n10062;
  assign n10064 = ~n3098 & n4484;
  assign n10065 = n10063 & ~n10064;
  assign n10066 = ~n10060 & n10065;
  assign n10067 = n10066 ^ x23;
  assign n10165 = n10164 ^ n10067;
  assign n10057 = n4955 ^ n4876;
  assign n10058 = ~n4956 & n10057;
  assign n10059 = n10058 ^ n4876;
  assign n10166 = n10165 ^ n10059;
  assign n10179 = n10178 ^ n10166;
  assign n10050 = n4963 & n5758;
  assign n10051 = ~n3875 & n4976;
  assign n10052 = ~n3431 & n4970;
  assign n10053 = ~n10051 & ~n10052;
  assign n10054 = ~n10050 & n10053;
  assign n10055 = n10054 ^ x17;
  assign n10047 = n4958 ^ n4852;
  assign n10048 = ~n4861 & n10047;
  assign n10049 = n10048 ^ n4958;
  assign n10056 = n10055 ^ n10049;
  assign n10180 = n10179 ^ n10056;
  assign n10181 = ~n10046 & ~n10180;
  assign n10182 = ~n4959 & ~n5208;
  assign n10183 = ~n10181 & ~n10182;
  assign n10184 = ~n10034 & n10183;
  assign n10185 = ~n10046 & n10182;
  assign n10186 = n10180 & ~n10185;
  assign n10187 = ~n10033 & ~n10186;
  assign n10188 = ~n5209 & ~n10180;
  assign n10189 = ~n10042 & n10045;
  assign n10190 = ~n10188 & ~n10189;
  assign n10191 = ~n10187 & n10190;
  assign n10192 = ~n10184 & ~n10191;
  assign n10193 = n10177 ^ n10166;
  assign n10194 = n10178 & ~n10193;
  assign n10195 = n10194 ^ n10169;
  assign n10196 = ~n10192 & n10195;
  assign n10208 = ~n189 & n1853;
  assign n10209 = ~n244 & n264;
  assign n10210 = n10208 & n10209;
  assign n10211 = n4360 & n4750;
  assign n10212 = n1072 & n2584;
  assign n10213 = n10211 & n10212;
  assign n10214 = n10210 & n10213;
  assign n10215 = n3027 & n10214;
  assign n10216 = n3299 & n10215;
  assign n10217 = ~n350 & ~n1135;
  assign n10218 = n1429 & n10217;
  assign n10219 = ~n57 & n1521;
  assign n10220 = n10218 & n10219;
  assign n10221 = ~n183 & n462;
  assign n10222 = n10220 & n10221;
  assign n10223 = n1541 & n10222;
  assign n10224 = n941 & n10223;
  assign n10225 = n3134 & n10224;
  assign n10226 = n10216 & n10225;
  assign n10227 = ~n10090 & ~n10135;
  assign n10228 = ~n10146 & n10227;
  assign n10353 = ~n10226 & n10228;
  assign n10229 = n10090 & n10135;
  assign n10230 = n10146 & n10229;
  assign n10354 = n10226 & n10230;
  assign n10355 = ~n10353 & ~n10354;
  assign n10334 = n2502 & n3136;
  assign n10335 = n1961 & n1976;
  assign n10336 = n2402 & n10335;
  assign n10337 = ~n83 & ~n296;
  assign n10338 = ~n375 & ~n541;
  assign n10339 = n10337 & n10338;
  assign n10340 = ~n216 & n1085;
  assign n10341 = n10339 & n10340;
  assign n10342 = n10336 & n10341;
  assign n10343 = n10334 & n10342;
  assign n10344 = n601 & n4208;
  assign n10345 = ~n344 & ~n627;
  assign n10346 = n2022 & n10345;
  assign n10347 = n10344 & n10346;
  assign n10348 = n5526 & n10347;
  assign n10349 = n10343 & n10348;
  assign n10350 = n5679 & n10349;
  assign n10351 = n2905 & n10350;
  assign n10352 = n10351 ^ x17;
  assign n10356 = n10355 ^ n10352;
  assign n10324 = n41 & ~n4495;
  assign n10233 = n54 & ~n2669;
  assign n10325 = n91 & ~n2786;
  assign n10326 = ~n10233 & ~n10325;
  assign n10327 = ~n10324 & n10326;
  assign n10328 = x31 & ~n10327;
  assign n10329 = ~n54 & n2718;
  assign n10330 = n54 & n2786;
  assign n10331 = n3640 & ~n10330;
  assign n10332 = ~n10329 & n10331;
  assign n10333 = ~n10328 & ~n10332;
  assign n10357 = n10356 ^ n10333;
  assign n10316 = n44 & n3749;
  assign n10317 = ~n566 & n3277;
  assign n10318 = ~n2861 & n3275;
  assign n10319 = ~n10317 & ~n10318;
  assign n10320 = ~n368 & n3280;
  assign n10321 = n10319 & ~n10320;
  assign n10322 = ~n10316 & n10321;
  assign n10323 = n10322 ^ x29;
  assign n10358 = n10357 ^ n10323;
  assign n10243 = n44 & ~n3666;
  assign n10244 = ~n2718 & n3275;
  assign n10245 = ~n2861 & n3277;
  assign n10246 = ~n10244 & ~n10245;
  assign n10247 = ~n566 & n3280;
  assign n10248 = n10246 & ~n10247;
  assign n10249 = ~n10243 & n10248;
  assign n10250 = n10249 ^ x29;
  assign n10236 = n41 & ~n4653;
  assign n10237 = n91 & ~n2669;
  assign n10238 = ~n10142 & ~n10237;
  assign n10239 = ~n10236 & n10238;
  assign n10234 = n41 & ~n2786;
  assign n10235 = ~n10233 & ~n10234;
  assign n10240 = n10239 ^ n10235;
  assign n10241 = ~x31 & n10240;
  assign n10242 = n10241 ^ n10239;
  assign n10251 = n10250 ^ n10242;
  assign n10231 = ~n10228 & ~n10230;
  assign n10232 = n10231 ^ n10226;
  assign n10313 = n10242 ^ n10232;
  assign n10314 = n10251 & n10313;
  assign n10315 = n10314 ^ n10250;
  assign n10359 = n10358 ^ n10315;
  assign n10305 = n3285 & ~n3974;
  assign n10306 = ~n2954 & n3435;
  assign n10307 = ~n3037 & ~n3440;
  assign n10308 = ~n10306 & ~n10307;
  assign n10309 = ~n3098 & n3437;
  assign n10310 = n10308 & ~n10309;
  assign n10311 = ~n10305 & n10310;
  assign n10312 = n10311 ^ x26;
  assign n10360 = n10359 ^ n10312;
  assign n10256 = n3285 & ~n3777;
  assign n10257 = ~n368 & ~n3440;
  assign n10258 = ~n3037 & n3435;
  assign n10259 = ~n10257 & ~n10258;
  assign n10260 = ~n2954 & n3437;
  assign n10261 = n10259 & ~n10260;
  assign n10262 = ~n10256 & n10261;
  assign n10263 = n10262 ^ x26;
  assign n10253 = n10147 ^ n10086;
  assign n10254 = ~n10161 & n10253;
  assign n10255 = n10254 ^ n10160;
  assign n10264 = n10263 ^ n10255;
  assign n10252 = n10251 ^ n10232;
  assign n10302 = n10263 ^ n10252;
  assign n10303 = n10264 & n10302;
  assign n10304 = n10303 ^ n10255;
  assign n10361 = n10360 ^ n10304;
  assign n10294 = ~n3989 & n4478;
  assign n10295 = ~n3270 & n4484;
  assign n10296 = ~n3351 & n4487;
  assign n10297 = ~n3196 & n4480;
  assign n10298 = ~n10296 & ~n10297;
  assign n10299 = ~n10295 & n10298;
  assign n10300 = ~n10294 & n10299;
  assign n10301 = n10300 ^ x23;
  assign n10362 = n10361 ^ n10301;
  assign n10266 = ~n3271 & n4478;
  assign n10267 = ~n3098 & n4480;
  assign n10268 = ~n3196 & n4484;
  assign n10269 = ~n10267 & ~n10268;
  assign n10270 = ~n3270 & n4487;
  assign n10271 = n10269 & ~n10270;
  assign n10272 = ~n10266 & n10271;
  assign n10273 = n10272 ^ x23;
  assign n10265 = n10264 ^ n10252;
  assign n10274 = n10273 ^ n10265;
  assign n10205 = n10162 ^ n10070;
  assign n10206 = n10163 & n10205;
  assign n10207 = n10206 ^ n10070;
  assign n10291 = n10273 ^ n10207;
  assign n10292 = n10274 & ~n10291;
  assign n10293 = n10292 ^ n10207;
  assign n10363 = n10362 ^ n10293;
  assign n10283 = ~n3879 & n4673;
  assign n10284 = ~n3404 & ~n4681;
  assign n10285 = ~n3431 & n4685;
  assign n10286 = ~n10284 & ~n10285;
  assign n10287 = ~n3875 & n4688;
  assign n10288 = n10286 & ~n10287;
  assign n10289 = ~n10283 & n10288;
  assign n10290 = n10289 ^ x20;
  assign n10364 = n10363 ^ n10290;
  assign n10275 = n10274 ^ n10207;
  assign n10197 = ~n3432 & n4673;
  assign n10198 = ~n3404 & n4685;
  assign n10199 = ~n3431 & n4688;
  assign n10200 = ~n10198 & ~n10199;
  assign n10201 = ~n3351 & ~n4681;
  assign n10202 = n10200 & ~n10201;
  assign n10203 = ~n10197 & n10202;
  assign n10204 = n10203 ^ x20;
  assign n10276 = n10275 ^ n10204;
  assign n10277 = n10164 ^ n10059;
  assign n10278 = ~n10165 & n10277;
  assign n10279 = n10278 ^ n10059;
  assign n10280 = n10279 ^ n10275;
  assign n10281 = ~n10276 & n10280;
  assign n10282 = n10281 ^ n10279;
  assign n10365 = n10364 ^ n10282;
  assign n10366 = ~n10196 & n10365;
  assign n10367 = n4963 & n6285;
  assign n10368 = ~n3875 & n4970;
  assign n10369 = ~n10367 & ~n10368;
  assign n10370 = n10369 ^ x17;
  assign n10371 = n10179 ^ n10049;
  assign n10372 = ~n10056 & n10371;
  assign n10373 = n10372 ^ n10179;
  assign n10374 = ~n10370 & ~n10373;
  assign n10375 = n10279 ^ n10276;
  assign n10376 = ~n10374 & n10375;
  assign n10377 = n10370 & n10373;
  assign n10378 = ~n10376 & ~n10377;
  assign n10379 = ~n10366 & ~n10378;
  assign n10380 = n10192 & ~n10195;
  assign n10381 = n10373 ^ n10365;
  assign n10382 = n10375 ^ n10370;
  assign n10383 = n10373 ^ n10370;
  assign n10384 = ~n10382 & ~n10383;
  assign n10385 = ~n10381 & n10384;
  assign n10386 = n10385 ^ n10365;
  assign n10387 = ~n10380 & ~n10386;
  assign n10388 = n10196 & ~n10365;
  assign n10389 = ~n10387 & ~n10388;
  assign n10390 = ~n10379 & n10389;
  assign n10391 = n4673 & n5758;
  assign n10392 = ~n3875 & n4685;
  assign n10393 = ~n3431 & ~n4681;
  assign n10394 = ~n10392 & ~n10393;
  assign n10395 = ~n10391 & n10394;
  assign n10396 = n10395 ^ x20;
  assign n10397 = n10390 & ~n10396;
  assign n10444 = ~n10333 & ~n10354;
  assign n10445 = ~n10353 & ~n10444;
  assign n10446 = ~n10352 & ~n10445;
  assign n10447 = n10226 & n10352;
  assign n10448 = ~n10228 & ~n10447;
  assign n10449 = ~n10333 & ~n10448;
  assign n10450 = ~n10230 & n10447;
  assign n10451 = ~n10449 & ~n10450;
  assign n10452 = ~n10446 & n10451;
  assign n10433 = n41 & n4466;
  assign n10434 = n91 & n2718;
  assign n10435 = x31 & ~n10330;
  assign n10436 = ~n10434 & n10435;
  assign n10437 = ~n10433 & n10436;
  assign n10438 = ~n2718 & n3671;
  assign n10439 = ~n2861 & n3676;
  assign n10440 = ~n10438 & ~n10439;
  assign n10441 = ~n10437 & n10440;
  assign n10428 = n10226 ^ x17;
  assign n10429 = n10351 ^ n10226;
  assign n10430 = n10428 & ~n10429;
  assign n10431 = n10430 ^ x17;
  assign n3457 = n1406 & n1492;
  assign n3459 = n1101 & n3458;
  assign n3460 = n3457 & n3459;
  assign n3461 = ~n458 & ~n790;
  assign n3462 = ~n359 & n3461;
  assign n3463 = n3460 & n3462;
  assign n3464 = n2817 & n2827;
  assign n3465 = n430 & n842;
  assign n3466 = n3464 & n3465;
  assign n3467 = n3463 & n3466;
  assign n3468 = n1897 & n3467;
  assign n3469 = n3456 & n3468;
  assign n3470 = ~n432 & n3361;
  assign n3474 = n3472 & n3473;
  assign n3475 = n3471 & n3474;
  assign n3476 = n3470 & n3475;
  assign n3477 = n2523 & n3476;
  assign n3478 = ~n263 & ~n358;
  assign n3479 = n673 & n3478;
  assign n3480 = ~n231 & n3130;
  assign n3481 = n3479 & n3480;
  assign n3483 = n1275 & n3482;
  assign n3484 = n3481 & n3483;
  assign n3485 = n3477 & n3484;
  assign n3486 = n3469 & n3485;
  assign n3487 = ~n319 & n3375;
  assign n3488 = n1121 & n3487;
  assign n3489 = n1305 & n1941;
  assign n3490 = n1665 & n1678;
  assign n3491 = n3489 & n3490;
  assign n3492 = n3488 & n3491;
  assign n3493 = ~n504 & ~n627;
  assign n3494 = ~n218 & ~n791;
  assign n3495 = n3493 & n3494;
  assign n3496 = n1528 & n3495;
  assign n3497 = n3492 & n3496;
  assign n3498 = n636 & n3235;
  assign n3501 = n3499 & n3500;
  assign n3502 = n3498 & n3501;
  assign n3503 = n3497 & n3502;
  assign n3504 = n2259 & n3503;
  assign n3505 = n3486 & n3504;
  assign n10432 = n10431 ^ n3505;
  assign n10442 = n10441 ^ n10432;
  assign n10420 = n44 & ~n3632;
  assign n10421 = ~n368 & n3277;
  assign n10422 = ~n3037 & n3280;
  assign n10423 = ~n10421 & ~n10422;
  assign n10424 = ~n566 & n3275;
  assign n10425 = n10423 & ~n10424;
  assign n10426 = ~n10420 & n10425;
  assign n10427 = n10426 ^ x29;
  assign n10443 = n10442 ^ n10427;
  assign n10453 = n10452 ^ n10443;
  assign n10412 = n3285 & n3647;
  assign n10413 = ~n2954 & ~n3440;
  assign n10414 = ~n3196 & n3437;
  assign n10415 = ~n10413 & ~n10414;
  assign n10416 = ~n3098 & n3435;
  assign n10417 = n10415 & ~n10416;
  assign n10418 = ~n10412 & n10417;
  assign n10419 = n10418 ^ x26;
  assign n10454 = n10453 ^ n10419;
  assign n10409 = n10357 ^ n10315;
  assign n10410 = ~n10358 & n10409;
  assign n10411 = n10410 ^ n10315;
  assign n10455 = n10454 ^ n10411;
  assign n10401 = n4478 & ~n5770;
  assign n10402 = ~n3270 & n4480;
  assign n10403 = ~n3351 & n4484;
  assign n10404 = ~n3404 & n4487;
  assign n10405 = ~n10403 & ~n10404;
  assign n10406 = ~n10402 & n10405;
  assign n10407 = ~n10401 & n10406;
  assign n10408 = n10407 ^ x23;
  assign n10456 = n10455 ^ n10408;
  assign n10398 = n10359 ^ n10304;
  assign n10399 = ~n10360 & n10398;
  assign n10400 = n10399 ^ n10304;
  assign n10457 = n10456 ^ n10400;
  assign n10458 = n10363 ^ n10282;
  assign n10459 = n10364 & ~n10458;
  assign n10460 = n10459 ^ n10282;
  assign n10461 = n10457 & ~n10460;
  assign n10462 = n10361 ^ n10293;
  assign n10463 = ~n10362 & ~n10462;
  assign n10464 = n10463 ^ n10293;
  assign n10465 = n10461 & n10464;
  assign n10466 = ~n10397 & ~n10465;
  assign n10506 = ~n10431 & ~n10441;
  assign n10507 = n10427 & n10452;
  assign n10508 = ~n10427 & ~n10452;
  assign n10509 = ~n3505 & ~n10508;
  assign n10510 = ~n10507 & ~n10509;
  assign n10511 = n10506 & n10510;
  assign n10512 = ~n3505 & ~n10506;
  assign n10513 = n10507 & n10512;
  assign n10514 = n10431 & n10441;
  assign n10515 = n10507 & n10514;
  assign n10516 = ~n10513 & ~n10515;
  assign n10517 = n10514 ^ n10508;
  assign n10518 = n10514 ^ n3505;
  assign n10519 = n10517 & n10518;
  assign n10520 = n10516 & n10519;
  assign n10521 = n10520 ^ n10516;
  assign n10522 = ~n10511 & n10521;
  assign n3680 = n520 & n2067;
  assign n3681 = ~n57 & n3680;
  assign n3682 = ~n136 & n1554;
  assign n3683 = n2964 & n3682;
  assign n3684 = n3681 & n3683;
  assign n3686 = ~n370 & ~n800;
  assign n3687 = n3685 & n3686;
  assign n3688 = ~n343 & ~n750;
  assign n3689 = n3687 & n3688;
  assign n3690 = ~n237 & ~n320;
  assign n3691 = ~n218 & n3690;
  assign n3692 = n3689 & n3691;
  assign n3693 = n3684 & n3692;
  assign n3694 = ~n272 & n2402;
  assign n3695 = n2163 & n3694;
  assign n3696 = ~n500 & n1238;
  assign n3697 = ~n327 & n3696;
  assign n3698 = n3695 & n3697;
  assign n3701 = n1085 & n1438;
  assign n3702 = n2170 & n3156;
  assign n3703 = n3701 & n3702;
  assign n3704 = n3700 & n3703;
  assign n3705 = n3698 & n3704;
  assign n3706 = n3693 & n3705;
  assign n3731 = n448 & n1453;
  assign n3732 = n1043 & n2544;
  assign n3733 = n2773 & n3732;
  assign n3734 = ~n375 & ~n1227;
  assign n3735 = n419 & n3734;
  assign n3736 = n3733 & n3735;
  assign n3532 = ~n243 & ~n314;
  assign n3739 = n3532 & n3738;
  assign n3740 = n3737 & n3739;
  assign n3741 = n1802 & n3740;
  assign n3742 = n3736 & n3741;
  assign n3743 = n3731 & n3742;
  assign n3744 = n3730 & n3743;
  assign n3745 = n3706 & n3744;
  assign n10504 = n3745 ^ n3505;
  assign n3668 = ~n3666 & n3667;
  assign n3670 = ~n2718 & n3669;
  assign n3674 = ~n2861 & ~n3673;
  assign n3675 = ~n3670 & ~n3674;
  assign n3677 = ~n566 & n3676;
  assign n3678 = n3675 & ~n3677;
  assign n3679 = ~n3668 & n3678;
  assign n10505 = n10504 ^ n3679;
  assign n10523 = n10522 ^ n10505;
  assign n10495 = ~n3271 & n3285;
  assign n10496 = ~n3098 & ~n3440;
  assign n10497 = ~n3196 & n3435;
  assign n10498 = ~n10496 & ~n10497;
  assign n10499 = ~n3270 & n3437;
  assign n10500 = n10498 & ~n10499;
  assign n10501 = ~n10495 & n10500;
  assign n10502 = n10501 ^ x26;
  assign n10487 = n44 & ~n3777;
  assign n10488 = ~n368 & n3275;
  assign n10489 = ~n3037 & n3277;
  assign n10490 = ~n10488 & ~n10489;
  assign n10491 = ~n2954 & n3280;
  assign n10492 = n10490 & ~n10491;
  assign n10493 = ~n10487 & n10492;
  assign n10494 = n10493 ^ x29;
  assign n10503 = n10502 ^ n10494;
  assign n10524 = n10523 ^ n10503;
  assign n10478 = ~n3432 & n4478;
  assign n10479 = ~n3404 & n4484;
  assign n10480 = ~n3351 & n4480;
  assign n10481 = ~n10479 & ~n10480;
  assign n10482 = ~n3431 & n4487;
  assign n10483 = n10481 & ~n10482;
  assign n10484 = ~n10478 & n10483;
  assign n10485 = n10484 ^ x23;
  assign n10475 = n10453 ^ n10411;
  assign n10476 = n10454 & ~n10475;
  assign n10477 = n10476 ^ n10411;
  assign n10486 = n10485 ^ n10477;
  assign n10525 = n10524 ^ n10486;
  assign n10470 = n4673 & n6285;
  assign n10471 = ~n3875 & ~n4681;
  assign n10472 = ~n10470 & ~n10471;
  assign n10473 = n10472 ^ x20;
  assign n10467 = n10455 ^ n10400;
  assign n10468 = n10456 & ~n10467;
  assign n10469 = n10468 ^ n10400;
  assign n10474 = n10473 ^ n10469;
  assign n10526 = n10525 ^ n10474;
  assign n10527 = n10460 ^ n10457;
  assign n10528 = n10464 ^ n10457;
  assign n10529 = ~n10527 & ~n10528;
  assign n10530 = n10529 ^ n10460;
  assign n10531 = ~n10526 & n10530;
  assign n10532 = ~n10466 & ~n10531;
  assign n10533 = ~n10457 & n10460;
  assign n10534 = ~n10464 & n10533;
  assign n10535 = n10526 & ~n10534;
  assign n10536 = ~n10532 & ~n10535;
  assign n10537 = ~n10390 & n10396;
  assign n10538 = n10526 & ~n10530;
  assign n10539 = n10537 & ~n10538;
  assign n10540 = ~n10536 & ~n10539;
  assign n10541 = n10525 ^ n10469;
  assign n10542 = ~n10474 & ~n10541;
  assign n10543 = n10542 ^ n10525;
  assign n10544 = ~n10540 & ~n10543;
  assign n10592 = n3285 & ~n5770;
  assign n10593 = ~n3270 & ~n3440;
  assign n10594 = ~n3351 & n3435;
  assign n10595 = ~n3404 & n3437;
  assign n10596 = ~n10594 & ~n10595;
  assign n10597 = ~n10593 & n10596;
  assign n10598 = ~n10592 & n10597;
  assign n10599 = n10598 ^ x26;
  assign n3746 = ~n3505 & ~n3745;
  assign n3747 = ~n3679 & n3746;
  assign n3750 = n3667 & n3749;
  assign n3751 = ~n566 & ~n3673;
  assign n3752 = ~n2861 & n3669;
  assign n3753 = ~n3751 & ~n3752;
  assign n3754 = ~n368 & n3676;
  assign n3755 = n3753 & ~n3754;
  assign n3756 = ~n3750 & n3755;
  assign n3757 = ~n3747 & n3756;
  assign n3758 = n3505 & n3745;
  assign n3759 = n3679 & n3758;
  assign n3507 = ~n98 & ~n504;
  assign n3508 = ~n1482 & n3507;
  assign n3509 = n965 & n3508;
  assign n3510 = ~n270 & ~n439;
  assign n3511 = n149 & n3510;
  assign n3512 = n1836 & n3511;
  assign n3513 = n3509 & n3512;
  assign n3514 = n3193 & n3513;
  assign n3515 = ~n110 & ~n592;
  assign n3516 = n2040 & n3515;
  assign n3517 = ~n263 & ~n284;
  assign n3518 = ~n87 & ~n346;
  assign n3519 = n3517 & n3518;
  assign n3520 = n3516 & n3519;
  assign n3522 = ~n327 & ~n841;
  assign n3523 = ~n751 & ~n1166;
  assign n3524 = n3522 & n3523;
  assign n3525 = n3521 & n3524;
  assign n3526 = n3520 & n3525;
  assign n3527 = n3514 & n3526;
  assign n3528 = ~n262 & n712;
  assign n3530 = n118 & n3529;
  assign n3531 = n3528 & n3530;
  assign n3533 = n1874 & n3532;
  assign n3534 = n1834 & n3533;
  assign n3535 = n3531 & n3534;
  assign n3536 = n3527 & n3535;
  assign n3559 = n1043 & n1567;
  assign n3561 = n1554 & n3560;
  assign n3562 = n3559 & n3561;
  assign n3563 = n618 & n2608;
  assign n3564 = n1153 & n2024;
  assign n3565 = n3563 & n3564;
  assign n3566 = n3562 & n3565;
  assign n3567 = ~n373 & ~n567;
  assign n3568 = ~n503 & n3567;
  assign n3569 = n802 & n2780;
  assign n3570 = n3568 & n3569;
  assign n3571 = n3566 & n3570;
  assign n3572 = n105 & n1021;
  assign n3573 = ~n234 & ~n272;
  assign n3574 = ~n403 & n3573;
  assign n3575 = n3572 & n3574;
  assign n3578 = n1058 & n2942;
  assign n3579 = n3577 & n3578;
  assign n3580 = n3575 & n3579;
  assign n3581 = n3571 & n3580;
  assign n3582 = n3558 & n3581;
  assign n3583 = n3536 & n3582;
  assign n3760 = n3583 ^ x20;
  assign n3761 = ~n3759 & ~n3760;
  assign n3762 = ~n3757 & n3761;
  assign n3763 = n3745 ^ n3679;
  assign n3764 = n3756 ^ n3745;
  assign n3765 = n3505 & n3760;
  assign n3766 = n3765 ^ n3756;
  assign n3767 = ~n3764 & ~n3766;
  assign n3768 = ~n3763 & n3767;
  assign n3769 = n3768 ^ n3765;
  assign n3770 = ~n3762 & ~n3769;
  assign n3648 = n44 & n3647;
  assign n3649 = ~n2954 & n3275;
  assign n3650 = ~n3196 & n3280;
  assign n3651 = ~n3649 & ~n3650;
  assign n3652 = ~n3098 & n3277;
  assign n3653 = n3651 & ~n3652;
  assign n3654 = ~n3648 & n3653;
  assign n3655 = n3654 ^ x29;
  assign n3633 = n41 & n3632;
  assign n3634 = n91 & n368;
  assign n3635 = x31 & ~n3634;
  assign n3636 = n54 & n566;
  assign n3637 = n3635 & ~n3636;
  assign n3638 = ~n3633 & n3637;
  assign n3639 = n54 & n368;
  assign n3641 = ~n54 & n3037;
  assign n3642 = n3640 & ~n3641;
  assign n3643 = ~n3639 & n3642;
  assign n3644 = ~n3638 & ~n3643;
  assign n3587 = ~n327 & ~n449;
  assign n3588 = ~n800 & n3587;
  assign n3589 = n1992 & n2170;
  assign n3590 = n3588 & n3589;
  assign n3591 = n235 & n453;
  assign n3592 = n3262 & n3591;
  assign n3593 = n3590 & n3592;
  assign n3594 = ~n710 & ~n791;
  assign n3595 = n1611 & n3594;
  assign n3597 = n570 & n3596;
  assign n3598 = n3595 & n3597;
  assign n3599 = n3593 & n3598;
  assign n3600 = ~n134 & ~n189;
  assign n3601 = n2123 & n3600;
  assign n3602 = ~n254 & n2404;
  assign n3603 = n3601 & n3602;
  assign n3604 = n1223 & n3603;
  assign n3605 = n3599 & n3604;
  assign n3607 = ~n155 & n3606;
  assign n3608 = n2560 & n3607;
  assign n3610 = ~n221 & ~n540;
  assign n3611 = n3609 & n3610;
  assign n3612 = ~n396 & n1209;
  assign n3613 = n3611 & n3612;
  assign n3614 = n3608 & n3613;
  assign n3615 = ~n403 & ~n628;
  assign n3616 = ~n249 & n3615;
  assign n3617 = n1398 & n3616;
  assign n3618 = ~n136 & n1043;
  assign n3619 = n3617 & n3618;
  assign n3620 = n3614 & n3619;
  assign n3621 = n1941 & n2488;
  assign n3622 = n992 & n2827;
  assign n3623 = n3621 & n3622;
  assign n3624 = ~n919 & n3623;
  assign n3625 = n3620 & n3624;
  assign n3626 = n3605 & n3625;
  assign n3627 = n2759 & n3626;
  assign n3628 = n696 & n1153;
  assign n3629 = n3627 & n3628;
  assign n3645 = n3644 ^ n3629;
  assign n3506 = n3505 ^ x20;
  assign n3584 = n3583 ^ n3505;
  assign n3585 = n3506 & ~n3584;
  assign n3586 = n3585 ^ x20;
  assign n3646 = n3645 ^ n3586;
  assign n3656 = n3655 ^ n3646;
  assign n10591 = n3770 ^ n3656;
  assign n10600 = n10599 ^ n10591;
  assign n10556 = n44 & ~n3974;
  assign n10557 = ~n2954 & n3277;
  assign n10558 = ~n3037 & n3275;
  assign n10559 = ~n10557 & ~n10558;
  assign n10560 = ~n3098 & n3280;
  assign n10561 = n10559 & ~n10560;
  assign n10562 = ~n10556 & n10561;
  assign n10563 = n10562 ^ x29;
  assign n10554 = ~n3747 & ~n3759;
  assign n10553 = n3760 ^ n3756;
  assign n10555 = n10554 ^ n10553;
  assign n10564 = n10563 ^ n10555;
  assign n10565 = n10505 & ~n10514;
  assign n10566 = ~n10510 & ~n10565;
  assign n10567 = n3505 & n10508;
  assign n10568 = ~n10505 & ~n10506;
  assign n10569 = ~n10567 & n10568;
  assign n10570 = ~n10505 & n10514;
  assign n10571 = ~n10513 & ~n10570;
  assign n10572 = ~n10569 & n10571;
  assign n10573 = ~n10566 & n10572;
  assign n10588 = n10573 ^ n10563;
  assign n10589 = ~n10564 & ~n10588;
  assign n10590 = n10589 ^ n10573;
  assign n10601 = n10600 ^ n10590;
  assign n10582 = n4478 & n5758;
  assign n10583 = ~n3875 & n4484;
  assign n10584 = ~n3431 & n4480;
  assign n10585 = ~n10583 & ~n10584;
  assign n10586 = ~n10582 & n10585;
  assign n10587 = n10586 ^ x23;
  assign n10602 = n10601 ^ n10587;
  assign n10574 = n10573 ^ n10564;
  assign n10545 = n3285 & ~n3989;
  assign n10546 = ~n3270 & n3435;
  assign n10547 = ~n3351 & n3437;
  assign n10548 = ~n3196 & ~n3440;
  assign n10549 = ~n10547 & ~n10548;
  assign n10550 = ~n10546 & n10549;
  assign n10551 = ~n10545 & n10550;
  assign n10552 = n10551 ^ x26;
  assign n10575 = n10574 ^ n10552;
  assign n10576 = n10523 ^ n10502;
  assign n10577 = ~n10503 & ~n10576;
  assign n10578 = n10577 ^ n10523;
  assign n10579 = n10578 ^ n10574;
  assign n10580 = n10575 & n10579;
  assign n10581 = n10580 ^ n10578;
  assign n10603 = n10602 ^ n10581;
  assign n10604 = ~n3879 & n4478;
  assign n10605 = ~n3404 & n4480;
  assign n10606 = ~n3875 & n4487;
  assign n10607 = ~n10605 & ~n10606;
  assign n10608 = ~n3431 & n4484;
  assign n10609 = n10607 & ~n10608;
  assign n10610 = ~n10604 & n10609;
  assign n10611 = n10610 ^ x23;
  assign n10612 = n10524 ^ n10485;
  assign n10613 = ~n10486 & ~n10612;
  assign n10614 = n10613 ^ n10524;
  assign n10615 = ~n10611 & n10614;
  assign n10616 = n10578 ^ n10575;
  assign n10617 = n10615 & ~n10616;
  assign n10618 = ~n10603 & ~n10617;
  assign n10619 = n10611 & ~n10614;
  assign n10620 = n10616 & n10619;
  assign n10621 = ~n10618 & ~n10620;
  assign n10622 = ~n10544 & n10621;
  assign n10623 = n10616 ^ n10611;
  assign n10624 = n10614 ^ n10611;
  assign n10625 = ~n10623 & ~n10624;
  assign n10626 = n10625 ^ n10614;
  assign n10627 = n10603 & n10626;
  assign n10628 = ~n10622 & ~n10627;
  assign n10629 = n10540 & n10543;
  assign n10630 = ~n10603 & ~n10626;
  assign n10631 = n10629 & ~n10630;
  assign n10632 = n10628 & ~n10631;
  assign n3845 = ~n3586 & ~n3629;
  assign n3846 = ~n3644 & n3845;
  assign n3847 = n3586 & n3629;
  assign n3848 = n3644 & n3847;
  assign n3849 = ~n3846 & ~n3848;
  assign n3797 = ~n166 & ~n312;
  assign n3798 = ~n109 & n3797;
  assign n3799 = n1046 & n3798;
  assign n3800 = ~n740 & ~n800;
  assign n3801 = ~n382 & n3800;
  assign n3802 = n464 & n3801;
  assign n3803 = n3799 & n3802;
  assign n3804 = n1392 & n3803;
  assign n3811 = n251 & n3019;
  assign n3814 = n3812 & n3813;
  assign n3815 = n3811 & n3814;
  assign n3816 = ~n87 & ~n691;
  assign n3817 = ~n156 & n3816;
  assign n3818 = n3815 & n3817;
  assign n3819 = n3810 & n3818;
  assign n3820 = n3804 & n3819;
  assign n3821 = n3796 & n3820;
  assign n3822 = ~n256 & n902;
  assign n3823 = n187 & n3822;
  assign n3825 = n1817 & n3824;
  assign n3826 = n2307 & n3825;
  assign n3827 = n3823 & n3826;
  assign n3829 = n1006 & n3828;
  assign n3830 = ~n330 & ~n361;
  assign n3831 = ~n518 & n3830;
  assign n3832 = n834 & n934;
  assign n3833 = n3831 & n3832;
  assign n3834 = n3829 & n3833;
  assign n3835 = n3827 & n3834;
  assign n3837 = ~n535 & ~n627;
  assign n3838 = ~n506 & n3837;
  assign n3839 = n3836 & n3838;
  assign n3840 = ~n197 & n1847;
  assign n3841 = n3839 & n3840;
  assign n3842 = n1963 & n3841;
  assign n3843 = n3835 & n3842;
  assign n3844 = n3821 & n3843;
  assign n3850 = n3849 ^ n3844;
  assign n3778 = n41 & n3777;
  assign n3779 = n91 & n3037;
  assign n3780 = x31 & ~n3779;
  assign n3781 = ~n3639 & n3780;
  assign n3782 = ~n3778 & n3781;
  assign n3783 = ~n54 & n2954;
  assign n3784 = n54 & n3037;
  assign n3785 = n3640 & ~n3784;
  assign n3786 = ~n3783 & n3785;
  assign n3787 = ~n3782 & ~n3786;
  assign n3851 = n3850 ^ n3787;
  assign n3771 = n3770 ^ n3655;
  assign n3772 = n3656 & n3771;
  assign n3773 = n3772 ^ n3770;
  assign n3852 = n3851 ^ n3773;
  assign n3433 = n3285 & ~n3432;
  assign n3436 = ~n3404 & n3435;
  assign n3438 = ~n3431 & n3437;
  assign n3439 = ~n3436 & ~n3438;
  assign n3441 = ~n3351 & ~n3440;
  assign n3442 = n3439 & ~n3441;
  assign n3443 = ~n3433 & n3442;
  assign n3444 = n3443 ^ x26;
  assign n3272 = n44 & ~n3271;
  assign n3276 = ~n3098 & n3275;
  assign n3278 = ~n3196 & n3277;
  assign n3279 = ~n3276 & ~n3278;
  assign n3281 = ~n3270 & n3280;
  assign n3282 = n3279 & ~n3281;
  assign n3283 = ~n3272 & n3282;
  assign n3284 = n3283 ^ x29;
  assign n3445 = n3444 ^ n3284;
  assign n10633 = n3852 ^ n3445;
  assign n3990 = n44 & ~n3989;
  assign n3991 = ~n3270 & n3277;
  assign n3992 = ~n3196 & n3275;
  assign n3993 = n3280 & ~n3351;
  assign n3994 = ~n3992 & ~n3993;
  assign n3995 = ~n3991 & n3994;
  assign n3996 = ~n3990 & n3995;
  assign n3997 = n3996 ^ x29;
  assign n3984 = n3844 & ~n3848;
  assign n3985 = ~n3846 & ~n3984;
  assign n3975 = n41 & n3974;
  assign n3976 = n91 & n2954;
  assign n3977 = x31 & ~n3784;
  assign n3978 = ~n3976 & n3977;
  assign n3979 = ~n3975 & n3978;
  assign n3980 = ~n3098 & n3676;
  assign n3981 = ~n2954 & n3671;
  assign n3982 = ~n3980 & ~n3981;
  assign n3983 = ~n3979 & n3982;
  assign n3986 = n3985 ^ n3983;
  assign n3915 = n168 & n1212;
  assign n3916 = n3022 & n3915;
  assign n3917 = n3914 & n3916;
  assign n3918 = ~n266 & n1091;
  assign n3919 = n3000 & n3918;
  assign n3920 = n3917 & n3919;
  assign n3921 = ~n322 & ~n369;
  assign n3922 = ~n337 & n3921;
  assign n3923 = n2544 & n3922;
  assign n3924 = n454 & n3923;
  assign n3926 = ~n514 & ~n640;
  assign n3927 = ~n689 & n3926;
  assign n3928 = n1274 & n2623;
  assign n3929 = n3927 & n3928;
  assign n3930 = n3925 & n3929;
  assign n3931 = n3924 & n3930;
  assign n3932 = n3920 & n3931;
  assign n3933 = n3911 & n3932;
  assign n3934 = n2282 & n3933;
  assign n3936 = ~n208 & ~n800;
  assign n3937 = n3935 & n3936;
  assign n3938 = ~n111 & ~n412;
  assign n3939 = n3937 & n3938;
  assign n3940 = ~n128 & n271;
  assign n3941 = n2344 & n2694;
  assign n3942 = n3940 & n3941;
  assign n3943 = n3939 & n3942;
  assign n3944 = n2517 & n3943;
  assign n3945 = ~n231 & ~n1005;
  assign n3946 = n1530 & n3945;
  assign n3947 = ~n221 & ~n627;
  assign n3948 = n3946 & n3947;
  assign n3949 = ~n553 & ~n659;
  assign n3950 = n3552 & n3949;
  assign n3951 = n3948 & n3950;
  assign n3952 = n771 & n982;
  assign n3953 = ~n560 & n3576;
  assign n3954 = n3952 & n3953;
  assign n3955 = n3951 & n3954;
  assign n3956 = n3944 & n3955;
  assign n3957 = ~n109 & ~n428;
  assign n3958 = ~n152 & n3957;
  assign n3959 = ~n353 & ~n1345;
  assign n3960 = n485 & n3959;
  assign n3961 = n3958 & n3960;
  assign n3962 = ~n331 & n1360;
  assign n3963 = ~n245 & ~n358;
  assign n3964 = n1314 & n3963;
  assign n3965 = n3962 & n3964;
  assign n3966 = n3961 & n3965;
  assign n3967 = n2335 & n3966;
  assign n3968 = n3956 & n3967;
  assign n3969 = n3934 & n3968;
  assign n3891 = n3844 ^ x23;
  assign n3970 = n3969 ^ n3891;
  assign n3987 = n3986 ^ n3970;
  assign n3998 = n3997 ^ n3987;
  assign n3888 = n3850 ^ n3773;
  assign n3889 = n3851 & ~n3888;
  assign n3890 = n3889 ^ n3773;
  assign n3999 = n3998 ^ n3890;
  assign n3880 = n3285 & ~n3879;
  assign n3881 = ~n3404 & ~n3440;
  assign n3882 = ~n3431 & n3435;
  assign n3883 = ~n3881 & ~n3882;
  assign n3884 = n3437 & ~n3875;
  assign n3885 = n3883 & ~n3884;
  assign n3886 = ~n3880 & n3885;
  assign n3887 = n3886 ^ x26;
  assign n4000 = n3999 ^ n3887;
  assign n3853 = n3852 ^ n3284;
  assign n3854 = n3445 & n3853;
  assign n3855 = n3854 ^ n3444;
  assign n4001 = n4000 ^ n3855;
  assign n10637 = n4478 & n6285;
  assign n10638 = ~n3875 & n4480;
  assign n10639 = ~n10637 & ~n10638;
  assign n10640 = n10639 ^ x23;
  assign n10634 = n10599 ^ n10590;
  assign n10635 = n10600 & ~n10634;
  assign n10636 = n10635 ^ n10590;
  assign n10641 = n10640 ^ n10636;
  assign n10642 = n10601 ^ n10581;
  assign n10643 = ~n10602 & ~n10642;
  assign n10644 = n10643 ^ n10581;
  assign n10645 = n10644 ^ n10636;
  assign n10646 = n10641 & n10645;
  assign n10647 = n10646 ^ n10644;
  assign n10946 = ~n4001 & n10647;
  assign n10947 = ~n10633 & ~n10946;
  assign n10649 = ~n10636 & n10640;
  assign n10650 = ~n10644 & n10649;
  assign n10653 = n10636 & ~n10640;
  assign n10654 = n10644 & n10653;
  assign n10948 = n4001 & ~n10654;
  assign n10949 = ~n10650 & ~n10948;
  assign n10950 = ~n10947 & n10949;
  assign n10951 = n10632 & ~n10950;
  assign n10952 = ~n10633 & ~n10949;
  assign n10953 = n4001 & ~n10647;
  assign n10954 = ~n10952 & ~n10953;
  assign n10955 = ~n10951 & n10954;
  assign n10884 = n3997 ^ n3890;
  assign n10885 = ~n3998 & n10884;
  assign n10886 = n10885 ^ n3890;
  assign n10937 = n3285 & n5758;
  assign n10938 = n3435 & ~n3875;
  assign n10939 = ~n3431 & ~n3440;
  assign n10940 = ~n10938 & ~n10939;
  assign n10941 = ~n10937 & n10940;
  assign n10942 = n10941 ^ x26;
  assign n11200 = n10886 & n10942;
  assign n11422 = n10955 & ~n11200;
  assign n10881 = n3999 ^ n3855;
  assign n10882 = ~n4000 & n10881;
  assign n10883 = n10882 ^ n3855;
  assign n10932 = n3983 ^ n3970;
  assign n10933 = n3986 & ~n10932;
  assign n10934 = n10933 ^ n3985;
  assign n10929 = n3969 ^ n3844;
  assign n10930 = n3891 & ~n10929;
  assign n10931 = n10930 ^ x23;
  assign n10935 = n10934 ^ n10931;
  assign n10920 = n44 & ~n5770;
  assign n10921 = ~n3270 & n3275;
  assign n10922 = n3277 & ~n3351;
  assign n10923 = n3280 & ~n3404;
  assign n10924 = ~n10922 & ~n10923;
  assign n10925 = ~n10921 & n10924;
  assign n10926 = ~n10920 & n10925;
  assign n10927 = n10926 ^ x29;
  assign n10909 = n41 & ~n3647;
  assign n10910 = n91 & n3098;
  assign n10911 = x31 & ~n10910;
  assign n10912 = n54 & n2954;
  assign n10913 = n10911 & ~n10912;
  assign n10914 = ~n10909 & n10913;
  assign n10915 = ~n3098 & n3671;
  assign n10916 = ~n3196 & n3676;
  assign n10917 = ~n10915 & ~n10916;
  assign n10918 = ~n10914 & n10917;
  assign n10919 = n10918 ^ n10908;
  assign n10928 = n10927 ^ n10919;
  assign n10936 = n10935 ^ n10928;
  assign n11197 = n10883 & ~n10936;
  assign n11198 = ~n10886 & ~n10942;
  assign n11204 = n11197 & ~n11198;
  assign n11180 = ~n10931 & ~n10934;
  assign n11181 = n10927 & ~n11180;
  assign n11182 = n10931 & n10934;
  assign n11183 = ~n11181 & ~n11182;
  assign n11185 = n10908 & ~n10918;
  assign n11184 = ~n10908 & n10918;
  assign n11186 = n11185 ^ n11184;
  assign n11187 = n11183 & n11186;
  assign n11188 = n11187 ^ n11185;
  assign n11189 = n10931 ^ n10927;
  assign n11190 = n10934 ^ n10927;
  assign n11191 = ~n11189 & ~n11190;
  assign n11192 = ~n10919 & n11191;
  assign n11193 = n11192 ^ n10919;
  assign n11194 = ~n11188 & n11193;
  assign n11178 = n11177 ^ n10908;
  assign n11179 = n11178 ^ n11130;
  assign n11195 = n11194 ^ n11179;
  assign n11097 = n44 & ~n3432;
  assign n11098 = n3275 & ~n3351;
  assign n11099 = n3280 ^ n3277;
  assign n11100 = n3404 & n11099;
  assign n11101 = n11100 ^ n3277;
  assign n11102 = ~n11098 & ~n11101;
  assign n11103 = ~n11097 & n11102;
  assign n11104 = n11103 ^ x29;
  assign n11093 = n3285 & n6285;
  assign n11094 = ~n3440 & ~n3875;
  assign n11095 = ~n11093 & ~n11094;
  assign n11096 = n11095 ^ x26;
  assign n11105 = n11104 ^ n11096;
  assign n11196 = n11195 ^ n11105;
  assign n11423 = ~n11196 & ~n11198;
  assign n11424 = ~n11204 & ~n11423;
  assign n11425 = ~n11422 & ~n11424;
  assign n11426 = ~n11196 & n11197;
  assign n11427 = ~n11425 & ~n11426;
  assign n11428 = n10955 & ~n11423;
  assign n11201 = ~n10883 & n10936;
  assign n11429 = n11196 & ~n11200;
  assign n11430 = ~n11201 & ~n11429;
  assign n11431 = ~n11428 & n11430;
  assign n11432 = n11427 & ~n11431;
  assign n11433 = n10927 ^ n10918;
  assign n11434 = n11179 ^ n10908;
  assign n11435 = n10919 & ~n11434;
  assign n11436 = ~n11433 & n11435;
  assign n11437 = n11436 ^ n11179;
  assign n11438 = ~n11180 & n11437;
  assign n11439 = n11182 ^ n11179;
  assign n11440 = n10919 & n11433;
  assign n11441 = n11440 ^ n10927;
  assign n11442 = n11441 ^ n11179;
  assign n11443 = n11439 & ~n11442;
  assign n11444 = n11443 ^ n11182;
  assign n11445 = ~n11438 & ~n11444;
  assign n11449 = n11353 ^ n11352;
  assign n11446 = n11130 ^ n10908;
  assign n11447 = n11177 ^ n11130;
  assign n11448 = n11446 & n11447;
  assign n11450 = n11449 ^ n11448;
  assign n11451 = n11445 & ~n11450;
  assign n11452 = ~n11432 & ~n11451;
  assign n11453 = ~n11445 & n11450;
  assign n11454 = n44 & ~n3879;
  assign n11455 = n3404 & ~n3875;
  assign n11456 = ~n3277 & ~n11455;
  assign n11457 = n3431 & ~n3875;
  assign n11458 = ~n3275 & ~n11457;
  assign n11459 = n11458 ^ n3431;
  assign n11460 = n11456 & n11459;
  assign n11461 = n11460 ^ n3431;
  assign n11462 = ~n11454 & n11461;
  assign n11463 = n11462 ^ x29;
  assign n11464 = n11195 ^ n11104;
  assign n11465 = ~n11105 & ~n11464;
  assign n11466 = n11465 ^ n11195;
  assign n11467 = ~n11463 & n11466;
  assign n11468 = n11365 ^ n11342;
  assign n11469 = ~n11467 & ~n11468;
  assign n11470 = ~n11453 & ~n11469;
  assign n11471 = ~n11452 & n11470;
  assign n11472 = n11453 & ~n11467;
  assign n11473 = n11468 & ~n11472;
  assign n11474 = ~n11432 & ~n11473;
  assign n11475 = n11463 & ~n11466;
  assign n11476 = ~n11451 & ~n11468;
  assign n11477 = ~n11475 & ~n11476;
  assign n11478 = ~n11474 & n11477;
  assign n11479 = ~n11471 & ~n11478;
  assign n11735 = n11479 ^ n11420;
  assign n11736 = n11421 & ~n11735;
  assign n11737 = n11736 ^ n11479;
  assign n11762 = n41 & ~n3879;
  assign n11763 = n54 & ~n3404;
  assign n11764 = n91 & ~n3431;
  assign n11765 = ~n11763 & ~n11764;
  assign n11766 = ~n11762 & n11765;
  assign n11767 = x31 & ~n11766;
  assign n11860 = n11737 & ~n11767;
  assign n11889 = ~n11855 & ~n11860;
  assign n11890 = n11761 & ~n11889;
  assign n11738 = n11419 ^ n11377;
  assign n11739 = ~n11378 & ~n11738;
  assign n11740 = n11739 ^ n11419;
  assign n11769 = n11413 & ~n11415;
  assign n11770 = ~n11417 & ~n11769;
  assign n11859 = ~n11740 & n11770;
  assign n11857 = ~n11737 & n11767;
  assign n11891 = n11855 & ~n11857;
  assign n11892 = ~n11859 & ~n11891;
  assign n11893 = ~n11890 & n11892;
  assign n11856 = n11740 & ~n11770;
  assign n11894 = n11856 ^ n11855;
  assign n11768 = n11767 ^ n11761;
  assign n11895 = n11767 ^ n11737;
  assign n11896 = n11768 & ~n11895;
  assign n11897 = n11896 ^ n11737;
  assign n11898 = n11897 ^ n11855;
  assign n11899 = ~n11894 & ~n11898;
  assign n11900 = n11899 ^ n11856;
  assign n11901 = ~n11893 & ~n11900;
  assign n12015 = ~n11880 & n11901;
  assign n12016 = ~n11922 & ~n12015;
  assign n12017 = x26 & ~n817;
  assign n12018 = n121 & ~n12017;
  assign n12019 = ~n12016 & n12018;
  assign n13725 = x14 & n12019;
  assign n18806 = x16 & ~x17;
  assign n18807 = n13725 & n18806;
  assign n18808 = ~x14 & x17;
  assign n18809 = ~n18807 & ~n18808;
  assign n18810 = x15 & ~n18809;
  assign n18811 = x17 & n12019;
  assign n18812 = n4966 & ~n18811;
  assign n11674 = x17 & ~n4968;
  assign n18813 = ~x14 & ~x16;
  assign n18814 = n11674 & ~n18813;
  assign n18815 = ~n18812 & ~n18814;
  assign n18816 = ~n18810 & n18815;
  assign n11908 = n11839 & ~n11854;
  assign n11909 = n11901 & n11908;
  assign n11881 = ~n819 & ~n1507;
  assign n11882 = ~n2506 & n11881;
  assign n11883 = ~n3868 & n11882;
  assign n11884 = n11753 & n11883;
  assign n11885 = n3324 & n11884;
  assign n11886 = n3422 & n11885;
  assign n11910 = ~n11839 & n11854;
  assign n11911 = n11886 & ~n11910;
  assign n11912 = ~n11909 & n11911;
  assign n11913 = n11880 & ~n11901;
  assign n11914 = ~n11912 & ~n11913;
  assign n11923 = ~n11914 & ~n11922;
  assign n11933 = n121 & n11839;
  assign n11934 = ~n11850 & ~n11922;
  assign n11935 = ~n11933 & ~n11934;
  assign n11936 = ~n11854 & ~n11935;
  assign n11924 = ~n11850 & n11922;
  assign n11925 = ~n11839 & n11924;
  assign n11926 = n11850 & ~n11886;
  assign n11927 = ~n11925 & ~n11926;
  assign n11928 = n11854 & ~n11927;
  assign n11929 = ~n11839 & n11850;
  assign n11930 = ~n11924 & ~n11929;
  assign n11931 = ~n11886 & ~n11930;
  assign n11932 = ~n11928 & ~n11931;
  assign n11937 = n11936 ^ n11932;
  assign n11938 = ~n11901 & ~n11937;
  assign n11939 = n11938 ^ n11936;
  assign n11940 = ~n11923 & ~n11939;
  assign n11858 = n11856 & n11857;
  assign n11861 = n11859 & n11860;
  assign n11862 = ~n11858 & ~n11861;
  assign n11863 = n11770 ^ n11767;
  assign n11864 = n11770 ^ n11740;
  assign n11865 = n11863 & ~n11864;
  assign n11866 = n11865 ^ n11740;
  assign n11868 = n11737 & ~n11866;
  assign n11869 = ~n11767 & n11859;
  assign n11870 = ~n11868 & ~n11869;
  assign n11867 = ~n11737 & n11866;
  assign n11871 = n11870 ^ n11867;
  assign n11872 = ~n11761 & ~n11871;
  assign n11873 = n11872 ^ n11870;
  assign n11874 = n11862 & n11873;
  assign n11875 = n11874 ^ n11855;
  assign n11771 = n11770 ^ n11768;
  assign n11772 = n11771 ^ n11740;
  assign n11773 = n11772 ^ n11737;
  assign n11480 = n11479 ^ n11421;
  assign n11488 = ~n11472 & ~n11475;
  assign n11489 = n11452 & ~n11488;
  assign n11490 = n11451 & ~n11475;
  assign n11491 = ~n11453 & n11467;
  assign n11492 = ~n11490 & ~n11491;
  assign n11493 = n11432 & ~n11492;
  assign n11494 = n11466 ^ n11445;
  assign n11483 = n11463 ^ n11450;
  assign n11495 = n11450 ^ n11445;
  assign n11496 = ~n11483 & n11495;
  assign n11497 = ~n11494 & n11496;
  assign n11498 = ~n11493 & ~n11497;
  assign n11499 = ~n11489 & n11498;
  assign n11500 = n11499 ^ n11468;
  assign n11484 = n11483 ^ n11445;
  assign n11485 = n11484 ^ n11466;
  assign n11486 = n11485 ^ n11432;
  assign n11205 = ~n11200 & ~n11204;
  assign n11206 = ~n11201 & ~n11205;
  assign n11199 = ~n11197 & n11198;
  assign n11202 = ~n11200 & n11201;
  assign n11203 = ~n11199 & ~n11202;
  assign n11207 = n11206 ^ n11203;
  assign n11208 = n10955 & ~n11207;
  assign n11209 = n11208 ^ n11206;
  assign n11210 = n10886 ^ n10883;
  assign n10943 = n10942 ^ n10936;
  assign n11211 = n10942 ^ n10886;
  assign n11212 = n10943 & ~n11211;
  assign n11213 = ~n11210 & n11212;
  assign n11214 = ~n11209 & ~n11213;
  assign n11215 = n11214 ^ n11196;
  assign n10944 = n10943 ^ n10886;
  assign n10945 = n10944 ^ n10883;
  assign n10956 = n10955 ^ n10945;
  assign n10648 = ~n10633 & ~n10647;
  assign n10651 = ~n10648 & ~n10650;
  assign n10652 = n10632 & ~n10651;
  assign n10655 = ~n10650 & ~n10654;
  assign n10656 = n10644 ^ n10633;
  assign n10657 = ~n10655 & ~n10656;
  assign n10658 = ~n10652 & ~n10657;
  assign n10659 = ~n10633 & ~n10654;
  assign n10660 = n10647 & ~n10659;
  assign n10661 = ~n10632 & n10660;
  assign n10662 = n10658 & ~n10661;
  assign n10663 = n10662 ^ n4001;
  assign n10666 = n10615 & n10629;
  assign n10667 = n10544 & n10619;
  assign n10668 = ~n10666 & ~n10667;
  assign n10669 = n10620 ^ n10617;
  assign n10670 = ~n10543 & n10669;
  assign n10671 = n10670 ^ n10617;
  assign n10672 = ~n10543 & ~n10615;
  assign n10673 = ~n10619 & ~n10672;
  assign n10674 = n10673 ^ n10616;
  assign n10675 = n10673 ^ n10540;
  assign n10676 = n10674 & ~n10675;
  assign n10677 = ~n10671 & n10676;
  assign n10678 = n10677 ^ n10671;
  assign n10679 = n10668 & ~n10678;
  assign n10680 = n10679 ^ n10603;
  assign n11216 = n10663 & ~n10680;
  assign n10664 = n10656 ^ n10641;
  assign n10665 = n10664 ^ n10632;
  assign n11217 = ~n10665 & n10956;
  assign n11218 = ~n11216 & ~n11217;
  assign n10681 = n10623 ^ n10614;
  assign n10682 = n10681 ^ n10543;
  assign n10683 = n10682 ^ n10540;
  assign n10684 = n10397 & ~n10533;
  assign n10685 = n10461 & ~n10537;
  assign n10686 = ~n10684 & ~n10685;
  assign n10687 = n10464 & ~n10686;
  assign n10688 = n10530 & n10537;
  assign n10689 = n10534 ^ n10461;
  assign n10690 = ~n10397 & n10689;
  assign n10691 = n10690 ^ n10461;
  assign n10692 = ~n10688 & ~n10691;
  assign n10693 = ~n10687 & n10692;
  assign n10694 = n10693 ^ n10526;
  assign n10695 = n10464 ^ n10396;
  assign n10696 = n10695 ^ n10457;
  assign n10697 = n10696 ^ n10460;
  assign n10698 = n10697 ^ n10390;
  assign n10699 = ~n10370 & ~n10375;
  assign n10700 = ~n10196 & n10699;
  assign n10701 = n10370 & n10375;
  assign n10702 = n10380 & ~n10701;
  assign n10703 = ~n10700 & ~n10702;
  assign n10704 = ~n10373 & ~n10703;
  assign n10705 = n10195 ^ n10192;
  assign n10706 = n10375 ^ n10195;
  assign n10707 = ~n10705 & ~n10706;
  assign n10708 = n10707 ^ n10192;
  assign n10709 = n10377 & ~n10708;
  assign n10710 = n10196 & n10376;
  assign n10711 = n10380 & n10699;
  assign n10712 = ~n10710 & ~n10711;
  assign n10713 = ~n10709 & n10712;
  assign n10714 = ~n10704 & n10713;
  assign n10715 = n10714 ^ n10365;
  assign n10716 = n10382 ^ n10195;
  assign n10717 = n10716 ^ n10373;
  assign n10718 = n10717 ^ n10192;
  assign n10719 = n5208 & n10046;
  assign n10720 = ~n4959 & ~n10719;
  assign n10721 = n10045 ^ n10042;
  assign n10722 = n10045 ^ n5208;
  assign n10723 = n10721 & ~n10722;
  assign n10724 = n10723 ^ n5208;
  assign n10725 = ~n10720 & n10724;
  assign n10726 = n10033 & n10725;
  assign n10727 = ~n5208 & n10189;
  assign n10728 = ~n10719 & ~n10727;
  assign n10729 = n5208 ^ n4959;
  assign n10730 = ~n10728 & ~n10729;
  assign n10731 = ~n10726 & ~n10730;
  assign n10732 = n4959 & ~n10727;
  assign n10733 = ~n10724 & ~n10732;
  assign n10734 = ~n10033 & n10733;
  assign n10735 = n10731 & ~n10734;
  assign n10736 = n10735 ^ n10180;
  assign n10737 = n10729 ^ n10721;
  assign n10738 = n10737 ^ n10033;
  assign n10739 = n10030 ^ n10012;
  assign n10740 = n10739 ^ n5795;
  assign n10741 = ~n5811 & ~n10008;
  assign n10742 = ~n9998 & ~n10741;
  assign n10743 = n10742 ^ n10005;
  assign n10744 = n9986 & n10743;
  assign n10745 = n10744 ^ n10005;
  assign n10746 = ~n10002 & ~n10745;
  assign n10747 = n10008 ^ n10005;
  assign n10748 = n5811 & n10747;
  assign n10749 = n10748 ^ n10005;
  assign n10750 = n10746 & ~n10749;
  assign n10751 = n10750 ^ n10000;
  assign n10752 = n10740 & n10751;
  assign n10753 = n9995 ^ n5811;
  assign n10754 = n10753 ^ n9990;
  assign n10755 = n10754 ^ n9993;
  assign n10756 = n10755 ^ n9986;
  assign n10757 = n9983 ^ n6292;
  assign n10758 = n9961 & n9965;
  assign n10763 = n6303 & ~n9968;
  assign n10759 = n6302 ^ n6293;
  assign n10760 = n9968 ^ n6302;
  assign n10761 = n10759 & ~n10760;
  assign n10762 = n10761 ^ n6293;
  assign n10764 = n10763 ^ n10762;
  assign n10765 = ~n10758 & n10764;
  assign n10766 = n10765 ^ n10762;
  assign n10767 = ~n9961 & ~n9965;
  assign n10768 = n9968 & n9970;
  assign n10769 = n10768 ^ n10762;
  assign n10770 = ~n10767 & ~n10769;
  assign n10771 = n10770 ^ n10762;
  assign n10772 = ~n10766 & n10771;
  assign n10773 = n10772 ^ n9972;
  assign n10774 = n10759 ^ n9968;
  assign n10775 = n10774 ^ n9965;
  assign n10776 = n10775 ^ n9961;
  assign n10777 = n9958 ^ n7162;
  assign n10778 = n9949 ^ n9946;
  assign n10779 = ~n9953 & ~n10778;
  assign n10780 = n10779 ^ n9946;
  assign n10781 = n9952 ^ n9946;
  assign n10782 = ~n7511 & n10781;
  assign n10783 = n10782 ^ n9946;
  assign n10784 = n10780 & ~n10783;
  assign n10785 = n10784 ^ n7163;
  assign n10786 = n7510 ^ n7172;
  assign n10787 = n10786 ^ n9943;
  assign n10788 = n10787 ^ n8024;
  assign n10789 = n10788 ^ n9941;
  assign n10790 = n9934 & n9937;
  assign n10791 = ~n8871 & ~n10790;
  assign n10792 = n8881 & ~n9934;
  assign n10793 = ~n9939 & ~n10792;
  assign n10794 = n10791 & n10793;
  assign n10795 = n10794 ^ n8872;
  assign n10796 = n8870 ^ n8863;
  assign n10797 = n10796 ^ n8861;
  assign n10798 = n10797 ^ n8858;
  assign n10799 = n10798 ^ n9934;
  assign n10800 = n9931 ^ n8907;
  assign n10801 = n8927 & ~n9928;
  assign n10802 = n9918 & ~n9919;
  assign n10803 = ~n10801 & ~n10802;
  assign n10804 = n9904 & ~n10803;
  assign n10805 = n8926 ^ n8908;
  assign n10806 = n9917 ^ n8926;
  assign n10807 = n9917 ^ n9914;
  assign n10808 = ~n10806 & ~n10807;
  assign n10809 = n10805 & n10808;
  assign n10810 = ~n10804 & ~n10809;
  assign n10811 = ~n8927 & n9928;
  assign n10812 = ~n9924 & ~n10811;
  assign n10813 = ~n9904 & ~n10812;
  assign n10814 = n10810 & ~n10813;
  assign n10815 = n10814 ^ n9906;
  assign n10816 = n9914 ^ n8926;
  assign n10817 = n10816 ^ n8908;
  assign n10818 = n10817 ^ n9917;
  assign n10819 = n10818 ^ n9904;
  assign n10820 = n9901 ^ n9887;
  assign n10821 = n9873 ^ n9343;
  assign n10822 = n9870 ^ n9356;
  assign n10823 = ~n9354 & ~n9355;
  assign n10824 = n10823 ^ n9343;
  assign n10825 = n9867 ^ n9368;
  assign n10826 = n10824 & ~n10825;
  assign n10827 = ~n10822 & ~n10826;
  assign n10828 = ~n10821 & ~n10827;
  assign n10829 = ~n10820 & ~n10828;
  assign n10830 = ~n10819 & ~n10829;
  assign n10831 = n10815 & ~n10830;
  assign n10832 = n10800 & ~n10831;
  assign n10833 = ~n10799 & ~n10832;
  assign n10834 = n10795 & ~n10833;
  assign n10835 = ~n10789 & ~n10834;
  assign n10836 = ~n10785 & ~n10835;
  assign n10837 = ~n10777 & ~n10836;
  assign n10838 = n10776 & ~n10837;
  assign n10839 = n10773 & ~n10838;
  assign n10840 = ~n10757 & ~n10839;
  assign n10841 = ~n10756 & ~n10840;
  assign n10842 = n10740 & n10841;
  assign n10843 = ~n10752 & ~n10842;
  assign n10844 = ~n10738 & n10843;
  assign n10845 = ~n10736 & ~n10844;
  assign n10846 = ~n10718 & ~n10845;
  assign n10847 = n10715 & ~n10846;
  assign n10848 = ~n10698 & ~n10847;
  assign n10849 = n10694 & ~n10848;
  assign n10850 = ~n10683 & ~n10849;
  assign n10853 = n10821 & ~n10822;
  assign n10854 = n10820 & ~n10853;
  assign n10855 = n10819 & ~n10854;
  assign n10856 = ~n10815 & ~n10855;
  assign n10857 = ~n10800 & ~n10856;
  assign n10858 = n10799 & ~n10857;
  assign n10859 = ~n10795 & ~n10858;
  assign n10860 = n10789 & ~n10859;
  assign n10861 = n10785 & ~n10860;
  assign n10862 = n10777 & ~n10861;
  assign n10863 = ~n10776 & ~n10862;
  assign n10864 = ~n10773 & ~n10863;
  assign n10865 = n10757 & ~n10864;
  assign n10866 = n10756 & ~n10865;
  assign n10867 = n10751 & ~n10866;
  assign n10868 = ~n10740 & ~n10867;
  assign n10869 = n10738 & ~n10868;
  assign n10870 = n10736 & ~n10869;
  assign n10871 = n10718 & ~n10870;
  assign n10872 = ~n10715 & ~n10871;
  assign n10873 = n10698 & ~n10872;
  assign n10874 = ~n10694 & ~n10873;
  assign n10875 = n10683 & ~n10874;
  assign n10876 = ~n10680 & ~n10875;
  assign n11219 = ~n10850 & ~n10876;
  assign n11220 = ~n11218 & ~n11219;
  assign n11221 = n10665 & ~n10956;
  assign n11222 = n10663 & ~n11221;
  assign n11223 = ~n10665 & ~n10680;
  assign n11224 = n10956 & n11223;
  assign n11225 = ~n11222 & ~n11224;
  assign n11226 = ~n11220 & n11225;
  assign n11502 = n10956 & ~n11226;
  assign n11503 = n11215 & ~n11502;
  assign n11504 = ~n11486 & ~n11503;
  assign n11505 = n11500 & ~n11504;
  assign n11774 = ~n11480 & ~n11505;
  assign n11876 = ~n11773 & ~n11774;
  assign n11877 = n11875 & ~n11876;
  assign n11887 = n11886 ^ n11850;
  assign n11888 = n11887 ^ n11880;
  assign n11902 = n11901 ^ n11888;
  assign n11903 = ~n11877 & n11902;
  assign n11481 = ~n10956 & n11226;
  assign n11482 = ~n11215 & ~n11481;
  assign n11487 = ~n11482 & n11486;
  assign n11501 = ~n11487 & ~n11500;
  assign n11775 = n11480 & ~n11501;
  assign n11904 = n11773 & ~n11775;
  assign n11905 = ~n11875 & ~n11904;
  assign n11906 = ~n11902 & ~n11905;
  assign n11907 = ~n11903 & ~n11906;
  assign n11941 = n11940 ^ n11907;
  assign n12668 = n4673 & ~n11941;
  assign n12669 = n4688 & ~n11940;
  assign n12670 = n4685 & n11902;
  assign n12671 = ~n4681 & ~n11875;
  assign n12672 = ~n12670 & ~n12671;
  assign n12673 = ~n12669 & n12672;
  assign n12674 = ~n12668 & n12673;
  assign n12675 = n12674 ^ x20;
  assign n11776 = ~n11774 & ~n11775;
  assign n11777 = n11776 ^ n11773;
  assign n12658 = n4478 & ~n11777;
  assign n12659 = n4487 & ~n11773;
  assign n12660 = n4480 & n11500;
  assign n12661 = n4484 & n11480;
  assign n12662 = ~n12660 & ~n12661;
  assign n12663 = ~n12659 & n12662;
  assign n12664 = ~n12658 & n12663;
  assign n12665 = n12664 ^ x23;
  assign n11703 = ~n11482 & ~n11503;
  assign n11704 = n11703 ^ n11486;
  assign n12383 = n3285 & n11704;
  assign n12384 = n3437 & n11486;
  assign n12385 = n3435 & n11215;
  assign n12386 = ~n3440 & ~n10956;
  assign n12387 = ~n12385 & ~n12386;
  assign n12388 = ~n12384 & n12387;
  assign n12389 = ~n12383 & n12388;
  assign n12390 = n12389 ^ x26;
  assign n10851 = n10680 & ~n10850;
  assign n10852 = ~n10665 & ~n10851;
  assign n10877 = n10665 & ~n10876;
  assign n11693 = ~n10852 & ~n10877;
  assign n11694 = n11693 ^ n10663;
  assign n12372 = n44 & ~n11694;
  assign n12373 = n3280 & ~n10663;
  assign n12374 = n3275 & n10680;
  assign n12375 = n3277 & n10665;
  assign n12376 = ~n12374 & ~n12375;
  assign n12377 = ~n12373 & n12376;
  assign n12378 = ~n12372 & n12377;
  assign n12379 = n12378 ^ x29;
  assign n12033 = ~n10847 & ~n10872;
  assign n12034 = n12033 ^ n10698;
  assign n12035 = n41 & ~n12034;
  assign n12036 = n91 & ~n10715;
  assign n12037 = n54 & ~n10718;
  assign n12038 = ~n12036 & ~n12037;
  assign n12039 = ~n12035 & n12038;
  assign n12030 = n54 & n10715;
  assign n12031 = n41 & n10698;
  assign n12032 = ~n12030 & ~n12031;
  assign n12040 = n12039 ^ n12032;
  assign n12041 = ~x31 & ~n12040;
  assign n12042 = n12041 ^ n12039;
  assign n12043 = ~n582 & ~n640;
  assign n12044 = ~n93 & ~n901;
  assign n12045 = n12043 & n12044;
  assign n12046 = n1821 & n12045;
  assign n12047 = n3577 & n12046;
  assign n12048 = ~n432 & ~n1135;
  assign n12049 = n828 & n1205;
  assign n12050 = n12048 & n12049;
  assign n12051 = n12047 & n12050;
  assign n12052 = ~n257 & n4750;
  assign n12053 = ~n296 & n602;
  assign n12054 = n658 & n12053;
  assign n12055 = n12052 & n12054;
  assign n12056 = n870 & n2854;
  assign n12057 = ~n209 & ~n314;
  assign n12058 = n1598 & n12057;
  assign n12059 = ~n557 & ~n740;
  assign n12060 = n2817 & n12059;
  assign n12061 = n12058 & n12060;
  assign n12062 = n12056 & n12061;
  assign n12063 = n12055 & n12062;
  assign n12064 = n3841 & n12063;
  assign n12065 = n12051 & n12064;
  assign n12066 = n2151 & n2570;
  assign n12067 = n3473 & n12066;
  assign n12068 = n2774 & n12067;
  assign n12069 = n144 & n2577;
  assign n12070 = ~n975 & n4058;
  assign n12071 = ~n51 & ~n309;
  assign n12072 = n12070 & n12071;
  assign n12073 = n12069 & n12072;
  assign n12074 = n12068 & n12073;
  assign n12075 = ~n812 & n856;
  assign n12076 = n338 & n355;
  assign n12077 = n1091 & n2935;
  assign n12078 = n12076 & n12077;
  assign n12079 = n12075 & n12078;
  assign n12080 = n12074 & n12079;
  assign n12081 = n1685 & n12080;
  assign n12082 = n12065 & n12081;
  assign n12359 = ~n12042 & n12082;
  assign n11575 = ~x13 & n5744;
  assign n11576 = x13 & n5742;
  assign n11577 = x14 & ~n11576;
  assign n11578 = ~n11575 & ~n11577;
  assign n11555 = ~n209 & ~n750;
  assign n11556 = ~n148 & ~n244;
  assign n11557 = n1153 & n11556;
  assign n11558 = n11555 & n11557;
  assign n11559 = n3607 & n3918;
  assign n11560 = n11558 & n11559;
  assign n11561 = n563 & n4389;
  assign n11562 = n11560 & n11561;
  assign n11563 = ~n308 & ~n656;
  assign n11564 = n532 & n11563;
  assign n11565 = n2385 & n4554;
  assign n11566 = n11564 & n11565;
  assign n11567 = n1085 & n2298;
  assign n11568 = n2433 & n4417;
  assign n11569 = n11567 & n11568;
  assign n11570 = n11566 & n11569;
  assign n11571 = n11562 & n11570;
  assign n11572 = n2054 & n11571;
  assign n11573 = n2030 & n5412;
  assign n11574 = n11572 & n11573;
  assign n11579 = n11578 ^ n11574;
  assign n12086 = ~n10848 & ~n10873;
  assign n12087 = n12086 ^ n10694;
  assign n12088 = n41 & n12087;
  assign n12089 = n91 & n10698;
  assign n12090 = x31 & ~n12089;
  assign n12091 = ~n12030 & n12090;
  assign n12092 = ~n12088 & n12091;
  assign n12093 = n41 & n10694;
  assign n11601 = n54 & n10698;
  assign n12094 = ~x31 & ~n11601;
  assign n12095 = ~n12093 & n12094;
  assign n12096 = ~n12092 & ~n12095;
  assign n12360 = n11579 & n12096;
  assign n12361 = n12359 & ~n12360;
  assign n11580 = ~n1060 & n2982;
  assign n11581 = n4033 & n11580;
  assign n11582 = n1660 & n4566;
  assign n11583 = ~n146 & ~n683;
  assign n11584 = n11582 & n11583;
  assign n11585 = n2493 & n3127;
  assign n11586 = n2791 & n11585;
  assign n11587 = n11584 & n11586;
  assign n11588 = ~n714 & n4277;
  assign n11589 = n11587 & n11588;
  assign n11590 = n2549 & n11589;
  assign n11591 = n1138 & n11590;
  assign n11592 = n11581 & n11591;
  assign n11593 = n2931 & n11592;
  assign n12362 = ~n11579 & ~n12096;
  assign n12363 = n11593 & ~n12362;
  assign n12364 = ~n12361 & n12363;
  assign n12365 = n12042 & ~n12082;
  assign n12366 = n12365 ^ n12096;
  assign n12367 = ~n11579 & ~n11593;
  assign n12368 = n12367 ^ n12096;
  assign n12369 = n12366 & ~n12368;
  assign n12370 = n12369 ^ n12365;
  assign n12371 = ~n12364 & ~n12370;
  assign n12380 = n12379 ^ n12371;
  assign n11598 = ~n10849 & ~n10874;
  assign n11599 = n11598 ^ n10683;
  assign n11600 = ~n54 & n11599;
  assign n11234 = x31 & ~n91;
  assign n11602 = n11234 & ~n11601;
  assign n11603 = ~n11600 & n11602;
  assign n11604 = n54 & n10694;
  assign n11605 = ~x31 & ~n11604;
  assign n11606 = n41 & n10683;
  assign n11607 = n11605 & ~n11606;
  assign n11608 = n3672 & ~n10694;
  assign n11609 = ~n11607 & ~n11608;
  assign n11610 = ~n11603 & n11609;
  assign n11594 = n11593 ^ n11578;
  assign n11595 = ~n11579 & n11594;
  assign n11596 = n11595 ^ n11593;
  assign n11517 = ~n567 & ~n710;
  assign n11518 = n2385 & n11517;
  assign n11519 = ~n167 & ~n244;
  assign n11520 = ~n428 & ~n550;
  assign n11521 = n11519 & n11520;
  assign n11522 = n11518 & n11521;
  assign n11523 = ~n298 & ~n975;
  assign n11524 = n3560 & n11523;
  assign n11525 = n483 & n11524;
  assign n11526 = n11522 & n11525;
  assign n11527 = ~n683 & ~n841;
  assign n11528 = n3310 & n11527;
  assign n11529 = ~n183 & ~n630;
  assign n11530 = n11528 & n11529;
  assign n11531 = n5087 & n11530;
  assign n11532 = n11526 & n11531;
  assign n11533 = n4427 & n11532;
  assign n11534 = ~n344 & n1180;
  assign n11535 = n11533 & n11534;
  assign n11536 = n2843 & n3059;
  assign n11537 = n4373 & n11536;
  assign n11538 = n1212 & n1944;
  assign n11539 = n990 & n1116;
  assign n11540 = n11538 & n11539;
  assign n11541 = n11537 & n11540;
  assign n11542 = n2104 & n5381;
  assign n11543 = n536 & n3904;
  assign n11544 = n11542 & n11543;
  assign n11545 = n892 & n2227;
  assign n11546 = n1451 & n11545;
  assign n11547 = n11544 & n11546;
  assign n11548 = n4157 & n10127;
  assign n11549 = n2711 & n11548;
  assign n11550 = n4532 & n11549;
  assign n11551 = n11547 & n11550;
  assign n11552 = n11541 & n11551;
  assign n11553 = n1279 & n11552;
  assign n11554 = n11535 & n11553;
  assign n11597 = n11596 ^ n11554;
  assign n12358 = n11610 ^ n11597;
  assign n12381 = n12380 ^ n12358;
  assign n12099 = ~n10851 & ~n10876;
  assign n12100 = n12099 ^ n10665;
  assign n12101 = n44 & n12100;
  assign n12102 = n3277 & n10680;
  assign n12103 = n3275 & n10683;
  assign n12104 = ~n12102 & ~n12103;
  assign n12105 = n3280 & n10665;
  assign n12106 = n12104 & ~n12105;
  assign n12107 = ~n12101 & n12106;
  assign n12108 = n12107 ^ x29;
  assign n12097 = n12096 ^ n11579;
  assign n12083 = n12082 ^ n12042;
  assign n12084 = n12042 ^ n11593;
  assign n12085 = n12083 & n12084;
  assign n12098 = n12097 ^ n12085;
  assign n12109 = n12108 ^ n12098;
  assign n12110 = ~n10846 & ~n10871;
  assign n12111 = n12110 ^ n10715;
  assign n12112 = n41 & ~n12111;
  assign n12113 = n54 & n10736;
  assign n12114 = n91 & ~n10718;
  assign n12115 = x31 & ~n12114;
  assign n12116 = ~n12113 & n12115;
  assign n12117 = ~n12112 & n12116;
  assign n12118 = n3676 & n10715;
  assign n12119 = n3671 & n10718;
  assign n12120 = ~n12118 & ~n12119;
  assign n12121 = ~n12117 & n12120;
  assign n12124 = n289 & n2538;
  assign n12125 = n4626 & n12124;
  assign n10977 = ~n167 & n4397;
  assign n12126 = n1232 & n10977;
  assign n12127 = n2733 & n2929;
  assign n12128 = n12126 & n12127;
  assign n12129 = ~n330 & ~n344;
  assign n12130 = ~n336 & n12129;
  assign n12131 = ~n199 & ~n440;
  assign n12132 = n12130 & n12131;
  assign n12133 = n2503 & n12132;
  assign n12134 = n305 & n413;
  assign n11970 = ~n146 & ~n850;
  assign n12135 = n1567 & n11970;
  assign n12136 = n12134 & n12135;
  assign n12137 = n12133 & n12136;
  assign n12138 = n12128 & n12137;
  assign n12139 = n3134 & n12138;
  assign n12140 = n12125 & n12139;
  assign n12122 = ~x11 & n5823;
  assign n12123 = n12122 ^ n5822;
  assign n12141 = n12140 ^ n12123;
  assign n12142 = ~n163 & ~n442;
  assign n12143 = ~n405 & ~n531;
  assign n12144 = n12142 & n12143;
  assign n12145 = ~n64 & ~n409;
  assign n12146 = n12144 & n12145;
  assign n12147 = n1716 & n2392;
  assign n12148 = n398 & n12147;
  assign n12149 = n12146 & n12148;
  assign n12150 = ~n151 & n1286;
  assign n12151 = n12149 & n12150;
  assign n12152 = ~n202 & ~n369;
  assign n12153 = n4019 & n12152;
  assign n12154 = n2325 & n12153;
  assign n12155 = n2225 & n3499;
  assign n12156 = n393 & n1197;
  assign n12157 = n2795 & n4066;
  assign n12158 = n12156 & n12157;
  assign n12159 = n12155 & n12158;
  assign n12160 = n12154 & n12159;
  assign n12161 = n856 & n994;
  assign n12162 = ~n111 & ~n218;
  assign n12163 = ~n375 & ~n525;
  assign n12164 = n12162 & n12163;
  assign n12165 = n12161 & n12164;
  assign n12166 = n1014 & n1755;
  assign n12167 = ~n206 & n1567;
  assign n12168 = n12166 & n12167;
  assign n12169 = n12165 & n12168;
  assign n12170 = n12160 & n12169;
  assign n12171 = n5065 & n12170;
  assign n12172 = n1249 & n12171;
  assign n12173 = n12151 & n12172;
  assign n12174 = n12173 ^ n12123;
  assign n12175 = ~n12141 & n12174;
  assign n12176 = n12175 ^ n12173;
  assign n12177 = ~n12121 & ~n12176;
  assign n12329 = n12176 ^ n11593;
  assign n12330 = n12329 ^ n12121;
  assign n12179 = ~n10845 & ~n10870;
  assign n12180 = n12179 ^ n10718;
  assign n12181 = n41 & ~n12180;
  assign n12182 = n91 & n10736;
  assign n12183 = x31 & ~n54;
  assign n12184 = x31 & n10738;
  assign n12185 = ~n12183 & ~n12184;
  assign n12186 = ~n12182 & ~n12185;
  assign n12187 = ~n12181 & n12186;
  assign n12188 = n3640 & ~n12113;
  assign n12189 = ~n54 & ~n10718;
  assign n12190 = n12188 & ~n12189;
  assign n12191 = ~n12187 & ~n12190;
  assign n12178 = n12173 ^ n12141;
  assign n12192 = n12191 ^ n12178;
  assign n12193 = n10843 & ~n10868;
  assign n12194 = n12193 ^ n10738;
  assign n12195 = n41 & ~n12194;
  assign n12196 = n91 & ~n10740;
  assign n12197 = ~n12195 & ~n12196;
  assign n12198 = x31 & ~n12197;
  assign n12199 = n41 & n10738;
  assign n12200 = n54 & n10740;
  assign n12201 = ~x31 & ~n12200;
  assign n12202 = ~n12199 & n12201;
  assign n12203 = n3669 & ~n10751;
  assign n12204 = ~n12202 & ~n12203;
  assign n12205 = ~n12198 & n12204;
  assign n12208 = ~n429 & n2085;
  assign n12209 = n1021 & n2214;
  assign n12210 = n12208 & n12209;
  assign n12211 = n483 & n1286;
  assign n12212 = ~n492 & n12211;
  assign n12213 = n12210 & n12212;
  assign n12214 = n1733 & n12213;
  assign n12215 = n135 & n2076;
  assign n12216 = ~n424 & ~n442;
  assign n12217 = n12215 & n12216;
  assign n12218 = ~n270 & ~n710;
  assign n12219 = ~n303 & ~n540;
  assign n12220 = n12218 & n12219;
  assign n12221 = n577 & n12220;
  assign n12222 = n12217 & n12221;
  assign n12223 = n5101 & n12222;
  assign n12224 = n1460 & n2704;
  assign n12225 = ~n359 & ~n375;
  assign n12226 = ~n217 & ~n330;
  assign n12227 = n12225 & n12226;
  assign n12228 = n12224 & n12227;
  assign n12229 = ~n93 & ~n221;
  assign n12230 = n2521 & n12229;
  assign n12231 = ~n616 & n3004;
  assign n12232 = n12230 & n12231;
  assign n12233 = n12228 & n12232;
  assign n12234 = n12223 & n12233;
  assign n12235 = n12214 & n12234;
  assign n12236 = n2568 & n11279;
  assign n12237 = n12235 & n12236;
  assign n12206 = ~x8 & n6315;
  assign n12207 = n12206 ^ n6312;
  assign n12238 = n12237 ^ n12207;
  assign n12239 = ~n278 & ~n506;
  assign n12240 = n1958 & n12239;
  assign n12241 = ~n185 & ~n550;
  assign n12242 = n10895 & n12241;
  assign n12243 = n12240 & n12242;
  assign n12244 = n5676 & n12243;
  assign n12245 = n282 & n1521;
  assign n12246 = n430 & n498;
  assign n12247 = n12245 & n12246;
  assign n12248 = n12244 & n12247;
  assign n12249 = n1817 & n11251;
  assign n12250 = n519 & ~n623;
  assign n12251 = n12249 & n12250;
  assign n12252 = n611 & n1785;
  assign n12253 = n1859 & n12252;
  assign n12254 = n12251 & n12253;
  assign n12255 = n144 & n2896;
  assign n12256 = n1328 & n10126;
  assign n12257 = n12255 & n12256;
  assign n12258 = n3496 & n12257;
  assign n12259 = n12254 & n12258;
  assign n12260 = n12248 & n12259;
  assign n12261 = n813 & n2683;
  assign n12262 = ~n146 & ~n322;
  assign n12263 = ~n98 & n12262;
  assign n12264 = n2976 & n12263;
  assign n12265 = n12261 & n12264;
  assign n12266 = n12260 & n12265;
  assign n12267 = ~n93 & ~n492;
  assign n12268 = ~n99 & n12267;
  assign n12269 = n1560 & n3417;
  assign n12270 = n12268 & n12269;
  assign n12271 = n2993 & n12270;
  assign n12272 = n1792 & n4916;
  assign n12273 = n105 & n2293;
  assign n12274 = n12272 & n12273;
  assign n12275 = n12271 & n12274;
  assign n12276 = ~n256 & n12275;
  assign n12277 = n12266 & n12276;
  assign n12278 = n3628 & n12277;
  assign n12279 = n12278 ^ n12207;
  assign n12280 = ~n12238 & n12279;
  assign n12281 = n12280 ^ n12278;
  assign n12282 = ~n12205 & n12281;
  assign n12283 = n12173 & ~n12282;
  assign n12284 = n12205 & ~n12281;
  assign n12285 = ~n12173 & ~n12284;
  assign n12286 = ~n202 & ~n616;
  assign n12287 = n11970 & n12286;
  assign n12288 = n4527 & n12287;
  assign n12289 = n2432 & n11400;
  assign n12290 = n834 & n12289;
  assign n12291 = n12288 & n12290;
  assign n12292 = ~n544 & ~n799;
  assign n12293 = ~n417 & n12292;
  assign n12294 = n450 & n12293;
  assign n12295 = n329 & n12294;
  assign n12296 = n12291 & n12295;
  assign n12297 = n219 & ~n647;
  assign n12298 = ~n238 & ~n1166;
  assign n12299 = n2593 & n12298;
  assign n12300 = n12297 & n12299;
  assign n12301 = n860 & n1225;
  assign n12302 = ~n375 & n2392;
  assign n12303 = n12301 & n12302;
  assign n12304 = n12300 & n12303;
  assign n12305 = n12296 & n12304;
  assign n12306 = n1813 & n12305;
  assign n12307 = n537 & n12069;
  assign n11040 = ~n222 & ~n1060;
  assign n12308 = n2848 & n11040;
  assign n12309 = n2240 & n2308;
  assign n12310 = n12308 & n12309;
  assign n12311 = n12307 & n12310;
  assign n12312 = n2207 & n3075;
  assign n12313 = n2723 & n12312;
  assign n12314 = n12311 & n12313;
  assign n12315 = ~n361 & ~n710;
  assign n12316 = ~n819 & n12315;
  assign n12317 = n1221 & n2384;
  assign n12318 = n12316 & n12317;
  assign n12319 = n933 & n12318;
  assign n12320 = n688 & n12319;
  assign n12321 = n12314 & n12320;
  assign n12322 = n10132 & n12321;
  assign n12323 = n12306 & n12322;
  assign n12324 = ~n12285 & ~n12323;
  assign n12325 = ~n12283 & ~n12324;
  assign n12326 = n12325 ^ n12191;
  assign n12327 = ~n12192 & n12326;
  assign n12328 = n12327 ^ n12325;
  assign n12331 = n12330 ^ n12328;
  assign n12332 = n44 & n11599;
  assign n12333 = n3277 & n10694;
  assign n12334 = n3275 & n10698;
  assign n12335 = ~n12333 & ~n12334;
  assign n12336 = n3280 & n10683;
  assign n12337 = n12335 & ~n12336;
  assign n12338 = ~n12332 & n12337;
  assign n12339 = n12338 ^ x29;
  assign n12340 = n12339 ^ n12330;
  assign n12341 = n12331 & ~n12340;
  assign n12342 = n12341 ^ n12339;
  assign n12343 = n12083 & n12342;
  assign n12344 = n12177 & ~n12343;
  assign n12345 = ~n12083 & ~n12342;
  assign n12346 = ~n11593 & ~n12345;
  assign n12347 = ~n12344 & n12346;
  assign n12348 = n12121 & n12176;
  assign n12349 = n12348 ^ n12342;
  assign n12350 = n11593 & ~n12083;
  assign n12351 = n12350 ^ n12348;
  assign n12352 = n12349 & ~n12351;
  assign n12353 = n12352 ^ n12342;
  assign n12354 = ~n12347 & ~n12353;
  assign n12355 = n12354 ^ n12108;
  assign n12356 = ~n12109 & ~n12355;
  assign n12357 = n12356 ^ n12354;
  assign n12382 = n12381 ^ n12357;
  assign n12656 = n12390 ^ n12382;
  assign n11227 = n11226 ^ n11215;
  assign n12460 = n11227 ^ n10956;
  assign n12558 = n3285 & ~n12460;
  assign n12559 = n3437 & n11215;
  assign n12560 = ~n3440 & ~n10663;
  assign n12561 = n3435 & ~n10956;
  assign n12562 = ~n12560 & ~n12561;
  assign n12563 = ~n12559 & n12562;
  assign n12564 = ~n12558 & n12563;
  assign n12565 = n12564 ^ x26;
  assign n12557 = n12354 ^ n12109;
  assign n12566 = n12565 ^ n12557;
  assign n12533 = n12176 ^ n12121;
  assign n12534 = ~n12329 & ~n12533;
  assign n12535 = n12534 ^ n12083;
  assign n12536 = n12535 ^ n12342;
  assign n11616 = ~n10850 & ~n10875;
  assign n12524 = n11616 ^ n10680;
  assign n12525 = n44 & n12524;
  assign n12526 = n3280 & n10680;
  assign n12527 = n3277 & n10683;
  assign n12528 = n3275 & n10694;
  assign n12529 = ~n12527 & ~n12528;
  assign n12530 = ~n12526 & n12529;
  assign n12531 = ~n12525 & n12530;
  assign n12532 = n12531 ^ x29;
  assign n12537 = n12536 ^ n12532;
  assign n10878 = n10877 ^ n10852;
  assign n10879 = ~n10663 & n10878;
  assign n10880 = n10879 ^ n10877;
  assign n10957 = n10956 ^ n10880;
  assign n12417 = ~x26 & n735;
  assign n12538 = ~n10957 & n12417;
  assign n12539 = n3435 & ~n10663;
  assign n12540 = ~n3440 & n10665;
  assign n12541 = ~n12539 & ~n12540;
  assign n12542 = x26 & n12541;
  assign n12543 = n10956 & n12542;
  assign n12544 = ~n12538 & ~n12543;
  assign n12545 = x25 & n12544;
  assign n12546 = n10957 & n12542;
  assign n12547 = ~n10956 & n12417;
  assign n12548 = ~x25 & ~n12547;
  assign n12549 = ~n12546 & n12548;
  assign n12550 = ~n12545 & ~n12549;
  assign n12431 = x26 & ~n735;
  assign n12432 = n12431 ^ x26;
  assign n12551 = ~n12432 & n12541;
  assign n12552 = n12551 ^ x26;
  assign n12553 = ~n12550 & n12552;
  assign n12554 = n12553 ^ n12536;
  assign n12555 = n12537 & ~n12554;
  assign n12556 = n12555 ^ n12553;
  assign n12653 = n12565 ^ n12556;
  assign n12654 = n12566 & n12653;
  assign n12655 = n12654 ^ n12556;
  assign n12657 = n12656 ^ n12655;
  assign n12666 = n12665 ^ n12657;
  assign n11506 = ~n11501 & ~n11505;
  assign n11507 = n11506 ^ n11480;
  assign n12568 = n4478 & n11507;
  assign n12569 = n4487 & n11480;
  assign n12570 = n4484 & n11500;
  assign n12571 = ~n12569 & ~n12570;
  assign n12572 = n4480 & n11486;
  assign n12573 = n12571 & ~n12572;
  assign n12574 = ~n12568 & n12573;
  assign n12575 = n12574 ^ x23;
  assign n12567 = n12566 ^ n12556;
  assign n12576 = n12575 ^ n12567;
  assign n12637 = n12553 ^ n12537;
  assign n12624 = n3285 & ~n11694;
  assign n12625 = n3437 & ~n10663;
  assign n12626 = ~n3440 & n10680;
  assign n12627 = n3435 & n10665;
  assign n12628 = ~n12626 & ~n12627;
  assign n12629 = ~n12625 & n12628;
  assign n12630 = ~n12624 & n12629;
  assign n12631 = n12630 ^ x26;
  assign n12578 = n44 & n12087;
  assign n12579 = n3280 & n10694;
  assign n12580 = n3275 & n10715;
  assign n12581 = n3277 & n10698;
  assign n12582 = ~n12580 & ~n12581;
  assign n12583 = ~n12579 & n12582;
  assign n12584 = ~n12578 & n12583;
  assign n12585 = n12584 ^ x29;
  assign n12577 = n12325 ^ n12192;
  assign n12586 = n12585 ^ n12577;
  assign n12466 = ~x29 & n42;
  assign n12599 = n12034 & n12466;
  assign n12600 = n3277 & n10715;
  assign n12601 = n3275 & n10718;
  assign n12602 = ~n12600 & ~n12601;
  assign n12603 = x29 & n12602;
  assign n12604 = ~n10698 & n12603;
  assign n12605 = ~n12599 & ~n12604;
  assign n12606 = x28 & n12605;
  assign n12607 = ~n12034 & n12603;
  assign n12608 = n10698 & n12466;
  assign n12609 = ~x28 & ~n12608;
  assign n12610 = ~n12607 & n12609;
  assign n12611 = ~n12606 & ~n12610;
  assign n12475 = x29 & ~n42;
  assign n12476 = n12475 ^ x29;
  assign n12612 = ~n12476 & n12602;
  assign n12613 = n12612 ^ x29;
  assign n12614 = ~n12611 & n12613;
  assign n12587 = ~x31 & ~n10736;
  assign n12588 = n41 & ~n12587;
  assign n12589 = ~n5354 & ~n10738;
  assign n12590 = n3669 & ~n10740;
  assign n12591 = ~x31 & n91;
  assign n12592 = ~n12590 & ~n12591;
  assign n12593 = ~n12589 & n12592;
  assign n12594 = ~n12588 & n12593;
  assign n12595 = ~n10844 & ~n10869;
  assign n12596 = n12595 ^ n10736;
  assign n12597 = n3667 & ~n12596;
  assign n12598 = ~n12594 & ~n12597;
  assign n12615 = n12614 ^ n12598;
  assign n12616 = ~n12283 & ~n12285;
  assign n12617 = n12616 ^ n12323;
  assign n12618 = n12617 ^ n12598;
  assign n12619 = n12615 & ~n12618;
  assign n12620 = n12619 ^ n12614;
  assign n12621 = n12620 ^ n12585;
  assign n12622 = ~n12586 & n12621;
  assign n12623 = n12622 ^ n12620;
  assign n12632 = n12631 ^ n12623;
  assign n12633 = n12339 ^ n12331;
  assign n12634 = n12633 ^ n12623;
  assign n12635 = n12632 & n12634;
  assign n12636 = n12635 ^ n12631;
  assign n12638 = n12637 ^ n12636;
  assign n11956 = ~n11487 & ~n11504;
  assign n11957 = n11956 ^ n11500;
  assign n12639 = n4478 & n11957;
  assign n12640 = n4487 & n11500;
  assign n12641 = n4484 & n11486;
  assign n12642 = n4480 & n11215;
  assign n12643 = ~n12641 & ~n12642;
  assign n12644 = ~n12640 & n12643;
  assign n12645 = ~n12639 & n12644;
  assign n12646 = n12645 ^ x23;
  assign n12647 = n12646 ^ n12637;
  assign n12648 = n12638 & ~n12647;
  assign n12649 = n12648 ^ n12646;
  assign n12650 = n12649 ^ n12575;
  assign n12651 = n12576 & n12650;
  assign n12652 = n12651 ^ n12649;
  assign n12667 = n12666 ^ n12652;
  assign n18805 = n12675 ^ n12667;
  assign n18828 = n18816 ^ n18805;
  assign n17382 = ~n11903 & n11940;
  assign n17383 = ~n12019 & ~n17382;
  assign n18775 = n4963 & n17383;
  assign n18776 = n4970 & ~n11940;
  assign n18777 = n4976 & ~n12019;
  assign n18778 = ~n4972 & ~n18777;
  assign n18779 = ~n18776 & n18778;
  assign n18780 = ~n18775 & n18779;
  assign n18781 = n18780 ^ x17;
  assign n12503 = ~n11877 & ~n11905;
  assign n12504 = n12503 ^ n11902;
  assign n18765 = n4673 & n12504;
  assign n18766 = n4688 & n11902;
  assign n18767 = n4685 & ~n11875;
  assign n18768 = ~n4681 & ~n11773;
  assign n18769 = ~n18767 & ~n18768;
  assign n18770 = ~n18766 & n18769;
  assign n18771 = ~n18765 & n18770;
  assign n18772 = n18771 ^ x20;
  assign n18764 = n12649 ^ n12576;
  assign n18773 = n18772 ^ n18764;
  assign n13067 = n12646 ^ n12638;
  assign n13041 = n12633 ^ n12632;
  assign n13025 = n3285 & n12100;
  assign n13026 = n3437 & n10665;
  assign n13027 = n3435 & n10680;
  assign n13028 = ~n13026 & ~n13027;
  assign n13029 = ~n3440 & n10683;
  assign n13030 = n13028 & ~n13029;
  assign n13031 = ~n13025 & n13030;
  assign n13032 = n13031 ^ x26;
  assign n13024 = n12620 ^ n12586;
  assign n13033 = n13032 ^ n13024;
  assign n12989 = n12617 ^ n12615;
  assign n12962 = n12281 ^ n12173;
  assign n12963 = n12962 ^ n12205;
  assign n12702 = ~n10840 & ~n10865;
  assign n12703 = n12702 ^ n10756;
  assign n12704 = n41 & ~n12703;
  assign n12705 = n54 & n10773;
  assign n12706 = n91 & n10757;
  assign n12707 = ~n12705 & ~n12706;
  assign n12708 = ~n12704 & n12707;
  assign n12709 = x31 & ~n12708;
  assign n12710 = n3676 & ~n10756;
  assign n12711 = n3671 & n10757;
  assign n12712 = ~n12710 & ~n12711;
  assign n12713 = ~n12709 & n12712;
  assign n12714 = n485 & n1172;
  assign n12715 = n542 & ~n919;
  assign n12716 = n12714 & n12715;
  assign n12717 = n360 & n4534;
  assign n12718 = n12716 & n12717;
  assign n11084 = ~n269 & ~n920;
  assign n12719 = n2384 & n4407;
  assign n12720 = n11084 & n12719;
  assign n12721 = n3070 & n12720;
  assign n12722 = n12718 & n12721;
  assign n12723 = n10115 & n11567;
  assign n12724 = n11169 & n12723;
  assign n12725 = n1364 & n12724;
  assign n12726 = n12722 & n12725;
  assign n12727 = ~n208 & n12299;
  assign n12728 = ~n265 & n1225;
  assign n12729 = n12727 & n12728;
  assign n12730 = ~n127 & n3543;
  assign n12731 = n995 & n12730;
  assign n10986 = ~n74 & ~n120;
  assign n12732 = n10986 & n11304;
  assign n12733 = n191 & n12732;
  assign n12734 = n12731 & n12733;
  assign n12735 = n12729 & n12734;
  assign n12736 = n12726 & n12735;
  assign n12737 = n255 & n3738;
  assign n12738 = n3538 & n12737;
  assign n12739 = n5546 & n12738;
  assign n12740 = n3951 & n12739;
  assign n12741 = ~n117 & ~n687;
  assign n12742 = n157 & n12741;
  assign n12743 = ~n138 & ~n452;
  assign n12744 = n2310 & n12743;
  assign n12745 = n12742 & n12744;
  assign n12746 = n5040 & n12745;
  assign n12747 = n12740 & n12746;
  assign n12748 = n12151 & n12747;
  assign n12749 = n12736 & n12748;
  assign n12750 = ~x2 & ~n9448;
  assign n12751 = x3 & x4;
  assign n12752 = x5 & ~n12751;
  assign n12753 = x2 & ~n12752;
  assign n12754 = ~x3 & ~x4;
  assign n12755 = ~x5 & ~n12754;
  assign n12756 = ~n12753 & ~n12755;
  assign n12757 = ~n12750 & n12756;
  assign n12758 = n12749 & ~n12757;
  assign n12759 = n12750 & n12755;
  assign n12760 = ~n12758 & ~n12759;
  assign n12761 = n12713 & ~n12760;
  assign n12762 = n12278 & ~n12761;
  assign n12763 = ~n12713 & n12760;
  assign n12764 = ~n12278 & ~n12763;
  assign n12765 = n1567 & ~n2506;
  assign n12766 = n999 & n1614;
  assign n12767 = n12765 & n12766;
  assign n12768 = n3696 & n12767;
  assign n12769 = n365 & n12768;
  assign n12770 = n2308 & n12143;
  assign n12771 = ~n1215 & n12770;
  assign n12772 = n274 & n2570;
  assign n12773 = n3610 & n11517;
  assign n12774 = n12772 & n12773;
  assign n12775 = n12771 & n12774;
  assign n12776 = n3053 & n12775;
  assign n12777 = n12769 & n12776;
  assign n12778 = n2062 & n12777;
  assign n12779 = n1829 & n12778;
  assign n12780 = ~n12764 & ~n12779;
  assign n12781 = ~n12762 & ~n12780;
  assign n12701 = n12278 ^ n12238;
  assign n12782 = n12781 ^ n12701;
  assign n12783 = ~n54 & n10842;
  assign n12784 = ~n10841 & ~n10865;
  assign n12785 = ~n54 & n12784;
  assign n12786 = ~n10756 & ~n12785;
  assign n12787 = ~n10740 & ~n12786;
  assign n12788 = ~n91 & ~n12787;
  assign n12789 = ~n12783 & n12788;
  assign n12790 = ~n10751 & ~n12789;
  assign n12791 = n41 & n10867;
  assign n12792 = ~n10740 & n12791;
  assign n12793 = ~n12790 & ~n12792;
  assign n12794 = x31 & ~n10756;
  assign n12795 = ~n91 & n12784;
  assign n12796 = n10752 & n12795;
  assign n12797 = n12183 & ~n12796;
  assign n12798 = ~n12794 & ~n12797;
  assign n12799 = n12793 & ~n12798;
  assign n12800 = n3676 & n10740;
  assign n12801 = n3671 & n10751;
  assign n12802 = ~n12800 & ~n12801;
  assign n12803 = ~n12799 & n12802;
  assign n12959 = n12803 ^ n12781;
  assign n12960 = ~n12782 & n12959;
  assign n12961 = n12960 ^ n12803;
  assign n12964 = n12963 ^ n12961;
  assign n12965 = n44 & n12111;
  assign n12966 = n3280 & n10715;
  assign n12967 = n3275 & ~n10736;
  assign n12968 = n3277 & n10718;
  assign n12969 = ~n12967 & ~n12968;
  assign n12970 = ~n12966 & n12969;
  assign n12971 = ~n12965 & n12970;
  assign n12972 = n12971 ^ x29;
  assign n12986 = n12972 ^ n12963;
  assign n12987 = ~n12964 & n12986;
  assign n12988 = n12987 ^ n12972;
  assign n12990 = n12989 ^ n12988;
  assign n12991 = n3285 & n12524;
  assign n12992 = n3437 & n10680;
  assign n12993 = n3435 & n10683;
  assign n12994 = ~n3440 & n10694;
  assign n12995 = ~n12993 & ~n12994;
  assign n12996 = ~n12992 & n12995;
  assign n12997 = ~n12991 & n12996;
  assign n12998 = n12997 ^ x26;
  assign n13021 = n12998 ^ n12989;
  assign n13022 = ~n12990 & n13021;
  assign n13023 = n13022 ^ n12998;
  assign n13038 = n13024 ^ n13023;
  assign n13039 = n13033 & ~n13038;
  assign n13040 = n13039 ^ n13032;
  assign n13042 = n13041 ^ n13040;
  assign n13043 = n4478 & n11704;
  assign n13044 = n4487 & n11486;
  assign n13045 = n4484 & n11215;
  assign n13046 = n4480 & ~n10956;
  assign n13047 = ~n13045 & ~n13046;
  assign n13048 = ~n13044 & n13047;
  assign n13049 = ~n13043 & n13048;
  assign n13050 = n13049 ^ x23;
  assign n13064 = n13050 ^ n13041;
  assign n13065 = n13042 & ~n13064;
  assign n13066 = n13065 ^ n13050;
  assign n13068 = n13067 ^ n13066;
  assign n11999 = ~n11876 & ~n11904;
  assign n12000 = n11999 ^ n11875;
  assign n13069 = n4673 & ~n12000;
  assign n13070 = n4688 & ~n11875;
  assign n13071 = n4685 & ~n11773;
  assign n13072 = ~n4681 & n11480;
  assign n13073 = ~n13071 & ~n13072;
  assign n13074 = ~n13070 & n13073;
  assign n13075 = ~n13069 & n13074;
  assign n13076 = n13075 ^ x20;
  assign n18761 = n13076 ^ n13066;
  assign n18762 = n13068 & n18761;
  assign n18763 = n18762 ^ n13076;
  assign n18774 = n18773 ^ n18763;
  assign n18782 = n18781 ^ n18774;
  assign n13077 = n13076 ^ n13068;
  assign n13051 = n13050 ^ n13042;
  assign n13012 = n4478 & ~n12460;
  assign n13013 = n4487 & n11215;
  assign n13014 = n4480 & ~n10663;
  assign n13015 = n4484 & ~n10956;
  assign n13016 = ~n13014 & ~n13015;
  assign n13017 = ~n13013 & n13016;
  assign n13018 = ~n13012 & n13017;
  assign n13019 = n13018 ^ x23;
  assign n12999 = n12998 ^ n12990;
  assign n12973 = n12972 ^ n12964;
  assign n12805 = n44 & n12180;
  assign n12806 = n3277 & ~n10736;
  assign n12807 = n3275 & n10738;
  assign n12808 = ~n12806 & ~n12807;
  assign n12809 = n3280 & n10718;
  assign n12810 = n12808 & ~n12809;
  assign n12811 = ~n12805 & n12810;
  assign n12812 = n12811 ^ x29;
  assign n12804 = n12803 ^ n12782;
  assign n12813 = n12812 ^ n12804;
  assign n12939 = ~n10841 & ~n10866;
  assign n12940 = n12939 ^ n10751;
  assign n12941 = n41 & ~n12940;
  assign n12942 = ~n11234 & ~n12794;
  assign n12943 = n54 & ~n10757;
  assign n12944 = ~n12942 & ~n12943;
  assign n12945 = ~n12941 & n12944;
  assign n12946 = n3676 & n10751;
  assign n12947 = n3671 & ~n10756;
  assign n12948 = ~n12946 & ~n12947;
  assign n12949 = ~n12945 & n12948;
  assign n12925 = n12760 ^ n12278;
  assign n12926 = n12925 ^ n12713;
  assign n12817 = ~n10839 & ~n10864;
  assign n12818 = n12817 ^ n10757;
  assign n12819 = n41 & n12818;
  assign n12820 = n91 & n10773;
  assign n12821 = n54 & ~n10776;
  assign n12822 = x31 & ~n12821;
  assign n12823 = ~n12820 & n12822;
  assign n12824 = ~n12819 & n12823;
  assign n12825 = n41 & n10757;
  assign n12826 = ~n12705 & ~n12825;
  assign n12827 = ~x31 & n12826;
  assign n12828 = ~n12824 & ~n12827;
  assign n12814 = n12755 ^ n12750;
  assign n12815 = ~n12753 & ~n12814;
  assign n12816 = n12815 ^ n12749;
  assign n12829 = n12828 ^ n12816;
  assign n12830 = n54 & ~n10789;
  assign n12831 = ~n10836 & ~n10861;
  assign n12832 = n12831 ^ n10777;
  assign n12833 = n41 & ~n12832;
  assign n12834 = ~n12830 & ~n12833;
  assign n12835 = x31 & ~n12834;
  assign n12836 = ~n3673 & n10785;
  assign n12837 = n3676 & ~n10777;
  assign n12838 = ~n12836 & ~n12837;
  assign n12839 = ~n12835 & n12838;
  assign n12840 = n857 & n4381;
  assign n12841 = ~n171 & ~n541;
  assign n12842 = n3128 & n12841;
  assign n12843 = n12840 & n12842;
  assign n12844 = n635 & ~n797;
  assign n12845 = n4056 & n12844;
  assign n12846 = n12843 & n12845;
  assign n12847 = ~n627 & ~n683;
  assign n12848 = n2404 & n12847;
  assign n12849 = n311 & n12848;
  assign n12850 = n12846 & n12849;
  assign n12851 = ~n418 & n900;
  assign n12852 = n1538 & n1805;
  assign n12853 = n4208 & n12852;
  assign n12854 = n12851 & n12853;
  assign n12855 = n2164 & n12854;
  assign n12856 = n12850 & n12855;
  assign n12857 = ~n344 & ~n452;
  assign n12858 = n2255 & n12857;
  assign n12859 = n5666 & n12858;
  assign n12860 = n12856 & n12859;
  assign n11023 = n473 & n3176;
  assign n11024 = ~n292 & n1492;
  assign n11025 = n1906 & n11024;
  assign n11026 = n11023 & n11025;
  assign n11027 = n1180 & n2104;
  assign n11028 = ~n640 & ~n850;
  assign n11029 = n11027 & n11028;
  assign n11030 = ~n390 & ~n929;
  assign n11031 = ~n750 & n11030;
  assign n11032 = n1141 & n2207;
  assign n11033 = n11031 & n11032;
  assign n11034 = n11029 & n11033;
  assign n11035 = n11026 & n11034;
  assign n11036 = n1852 & n11035;
  assign n12861 = ~n396 & n1273;
  assign n12862 = n2155 & n12861;
  assign n12863 = n12299 & n12862;
  assign n12864 = ~n254 & ~n666;
  assign n12865 = n5659 & n12864;
  assign n12866 = n2344 & n5520;
  assign n12867 = n3127 & n12866;
  assign n12868 = n12865 & n12867;
  assign n12869 = n1717 & n1911;
  assign n12870 = n493 & n2662;
  assign n12871 = n12869 & n12870;
  assign n12872 = ~n174 & ~n293;
  assign n12873 = n2300 & n12872;
  assign n12874 = n12871 & n12873;
  assign n12875 = n12868 & n12874;
  assign n12876 = n12863 & n12875;
  assign n12877 = n11036 & n12876;
  assign n12878 = n12860 & n12877;
  assign n12879 = n12839 & n12878;
  assign n12880 = n12750 & ~n12879;
  assign n12881 = ~n12839 & ~n12878;
  assign n12882 = ~n12750 & ~n12881;
  assign n12883 = n1263 & n11523;
  assign n12884 = n11139 & n12883;
  assign n12885 = n435 & n12884;
  assign n12886 = ~n227 & n1072;
  assign n12887 = n5394 & n12886;
  assign n12888 = n2698 & n12887;
  assign n12889 = n12885 & n12888;
  assign n11800 = ~n115 & ~n361;
  assign n11801 = ~n443 & n11800;
  assign n11802 = n279 & n11801;
  assign n12890 = n2923 & n4750;
  assign n12891 = n934 & n3113;
  assign n12892 = n12890 & n12891;
  assign n12893 = ~n517 & ~n567;
  assign n12894 = n4077 & n12893;
  assign n12895 = n235 & ~n320;
  assign n12896 = n12894 & n12895;
  assign n12897 = n12892 & n12896;
  assign n12898 = n11802 & n12897;
  assign n12899 = n12889 & n12898;
  assign n12900 = n12736 & n12899;
  assign n12901 = ~n12882 & ~n12900;
  assign n12902 = ~n12880 & ~n12901;
  assign n12903 = n12902 ^ n12750;
  assign n12904 = n1306 & n4417;
  assign n12905 = n602 & n12904;
  assign n12906 = n1255 & n12905;
  assign n12907 = n618 & n12142;
  assign n12908 = ~n475 & ~n652;
  assign n12909 = n279 & n12908;
  assign n12910 = n12907 & n12909;
  assign n11066 = n1328 & n1887;
  assign n12911 = ~n527 & ~n751;
  assign n12912 = ~n304 & n12911;
  assign n12913 = n11066 & n12912;
  assign n12914 = n12910 & n12913;
  assign n12915 = n12906 & n12914;
  assign n12916 = n4542 & n12915;
  assign n12917 = n3224 & n12916;
  assign n12918 = n3821 & n12917;
  assign n12919 = n12918 ^ n12902;
  assign n12920 = ~n12903 & ~n12919;
  assign n12921 = n12920 ^ n12750;
  assign n12922 = n12921 ^ n12828;
  assign n12923 = ~n12829 & n12922;
  assign n12924 = n12923 ^ n12921;
  assign n12927 = n12926 ^ n12924;
  assign n12928 = n44 & n12194;
  assign n12929 = n3280 & n10738;
  assign n12930 = n3277 & n10740;
  assign n12931 = n3275 & n10751;
  assign n12932 = ~n12930 & ~n12931;
  assign n12933 = ~n12929 & n12932;
  assign n12934 = ~n12928 & n12933;
  assign n12935 = n12934 ^ x29;
  assign n12936 = n12935 ^ n12924;
  assign n12937 = n12927 & ~n12936;
  assign n12938 = n12937 ^ n12935;
  assign n12950 = n12949 ^ n12938;
  assign n12951 = ~n12762 & ~n12764;
  assign n12952 = n12951 ^ n12779;
  assign n12953 = n12952 ^ n12949;
  assign n12954 = n12950 & ~n12953;
  assign n12955 = n12954 ^ n12938;
  assign n12956 = n12955 ^ n12812;
  assign n12957 = ~n12813 & n12956;
  assign n12958 = n12957 ^ n12955;
  assign n12974 = n12973 ^ n12958;
  assign n12975 = n3285 & n11599;
  assign n12976 = n3435 & n10694;
  assign n12977 = ~n3440 & n10698;
  assign n12978 = ~n12976 & ~n12977;
  assign n12979 = n3437 & n10683;
  assign n12980 = n12978 & ~n12979;
  assign n12981 = ~n12975 & n12980;
  assign n12982 = n12981 ^ x26;
  assign n12983 = n12982 ^ n12973;
  assign n12984 = ~n12974 & n12983;
  assign n12985 = n12984 ^ n12982;
  assign n13000 = n12999 ^ n12985;
  assign n13001 = n4478 & ~n10957;
  assign n13002 = n4484 & ~n10663;
  assign n13003 = n4487 & ~n10956;
  assign n13004 = n4480 & n10665;
  assign n13005 = ~n13003 & ~n13004;
  assign n13006 = ~n13002 & n13005;
  assign n13007 = ~n13001 & n13006;
  assign n13008 = n13007 ^ x23;
  assign n13009 = n13008 ^ n12999;
  assign n13010 = ~n13000 & n13009;
  assign n13011 = n13010 ^ n13008;
  assign n13020 = n13019 ^ n13011;
  assign n13034 = n13033 ^ n13023;
  assign n13035 = n13034 ^ n13011;
  assign n13036 = n13020 & ~n13035;
  assign n13037 = n13036 ^ n13019;
  assign n13052 = n13051 ^ n13037;
  assign n13053 = n4673 & ~n11777;
  assign n13054 = n4688 & ~n11773;
  assign n13055 = ~n4681 & n11500;
  assign n13056 = n4685 & n11480;
  assign n13057 = ~n13055 & ~n13056;
  assign n13058 = ~n13054 & n13057;
  assign n13059 = ~n13053 & n13058;
  assign n13060 = n13059 ^ x20;
  assign n13061 = n13060 ^ n13051;
  assign n13062 = n13052 & ~n13061;
  assign n13063 = n13062 ^ n13060;
  assign n13078 = n13077 ^ n13063;
  assign n12011 = n11906 ^ n11903;
  assign n12012 = ~n11940 & n12011;
  assign n12013 = n12012 ^ n11903;
  assign n13079 = n4962 & n12013;
  assign n13080 = n4961 & ~n12019;
  assign n13081 = ~n13079 & n13080;
  assign n13082 = n4976 & ~n11940;
  assign n13083 = n4970 & n11902;
  assign n13084 = ~n13082 & ~n13083;
  assign n13085 = ~n13081 & n13084;
  assign n13086 = n13085 ^ x17;
  assign n18758 = n13086 ^ n13077;
  assign n18759 = n13078 & ~n18758;
  assign n18760 = n18759 ^ n13086;
  assign n18818 = n18781 ^ n18760;
  assign n18819 = n18782 & n18818;
  assign n18820 = n18819 ^ n18760;
  assign n18829 = n18820 ^ n18805;
  assign n18830 = ~n18828 & ~n18829;
  assign n18831 = n18830 ^ n18820;
  assign n13087 = n13086 ^ n13078;
  assign n13719 = x13 & ~x14;
  assign n13720 = x11 & n12019;
  assign n13721 = n13719 & n13720;
  assign n13722 = ~x11 & x14;
  assign n13723 = ~n13721 & ~n13722;
  assign n13724 = x12 & ~n13723;
  assign n13726 = n11575 & ~n13725;
  assign n13727 = ~x11 & ~x13;
  assign n13728 = n11577 & ~n13727;
  assign n13729 = ~n13726 & ~n13728;
  assign n13730 = ~n13724 & n13729;
  assign n13689 = n4673 & n11507;
  assign n13690 = n4688 & n11480;
  assign n13691 = n4685 & n11500;
  assign n13692 = ~n13690 & ~n13691;
  assign n13693 = ~n4681 & n11486;
  assign n13694 = n13692 & ~n13693;
  assign n13695 = ~n13689 & n13694;
  assign n13696 = n13695 ^ x20;
  assign n13688 = n13034 ^ n13020;
  assign n13697 = n13696 ^ n13688;
  assign n13651 = n13008 ^ n13000;
  assign n13625 = n12982 ^ n12974;
  assign n13118 = n3285 & n12087;
  assign n13119 = n3437 & n10694;
  assign n13120 = ~n3440 & n10715;
  assign n13121 = n3435 & n10698;
  assign n13122 = ~n13120 & ~n13121;
  assign n13123 = ~n13119 & n13122;
  assign n13124 = ~n13118 & n13123;
  assign n13125 = n13124 ^ x26;
  assign n13117 = n12955 ^ n12813;
  assign n13126 = n13125 ^ n13117;
  assign n13096 = n12952 ^ n12950;
  assign n13088 = n44 & ~n12596;
  assign n13089 = n3280 & ~n10736;
  assign n13090 = n3277 & n10738;
  assign n13091 = n3275 & n10740;
  assign n13092 = ~n13090 & ~n13091;
  assign n13093 = ~n13089 & n13092;
  assign n13094 = ~n13088 & n13093;
  assign n13095 = n13094 ^ x29;
  assign n13097 = n13096 ^ n13095;
  assign n13098 = n12034 & n12417;
  assign n13099 = n3435 & n10715;
  assign n13100 = ~n3440 & n10718;
  assign n13101 = ~n13099 & ~n13100;
  assign n13102 = x26 & n13101;
  assign n13103 = ~n10698 & n13102;
  assign n13104 = ~n13098 & ~n13103;
  assign n13105 = x25 & n13104;
  assign n13106 = ~n12034 & n13102;
  assign n13107 = n10698 & n12417;
  assign n13108 = ~x25 & ~n13107;
  assign n13109 = ~n13106 & n13108;
  assign n13110 = ~n13105 & ~n13109;
  assign n13111 = ~n12432 & n13101;
  assign n13112 = n13111 ^ x26;
  assign n13113 = ~n13110 & n13112;
  assign n13114 = n13113 ^ n13096;
  assign n13115 = ~n13097 & n13114;
  assign n13116 = n13115 ^ n13113;
  assign n13622 = n13125 ^ n13116;
  assign n13623 = ~n13126 & n13622;
  assign n13624 = n13623 ^ n13116;
  assign n13626 = n13625 ^ n13624;
  assign n13627 = n4478 & ~n11694;
  assign n13628 = n4487 & ~n10663;
  assign n13629 = n4480 & n10680;
  assign n13630 = n4484 & n10665;
  assign n13631 = ~n13629 & ~n13630;
  assign n13632 = ~n13628 & n13631;
  assign n13633 = ~n13627 & n13632;
  assign n13634 = n13633 ^ x23;
  assign n13648 = n13634 ^ n13624;
  assign n13649 = ~n13626 & n13648;
  assign n13650 = n13649 ^ n13634;
  assign n13652 = n13651 ^ n13650;
  assign n13653 = ~x20 & n4671;
  assign n13654 = n11957 & n13653;
  assign n13655 = n4685 & n11486;
  assign n13656 = ~n4681 & n11215;
  assign n13657 = ~n13655 & ~n13656;
  assign n13658 = x20 & n13657;
  assign n13659 = ~n11500 & n13658;
  assign n13660 = x19 & ~n13659;
  assign n13661 = ~n13654 & n13660;
  assign n13662 = ~n11957 & n13658;
  assign n13663 = n11500 & n13653;
  assign n13664 = ~x19 & ~n13663;
  assign n13665 = ~n13662 & n13664;
  assign n13666 = ~n13661 & ~n13665;
  assign n13667 = x20 & ~n4671;
  assign n13668 = n13667 ^ x20;
  assign n13669 = n13657 & ~n13668;
  assign n13670 = n13669 ^ x20;
  assign n13671 = ~n13666 & n13670;
  assign n13685 = n13671 ^ n13651;
  assign n13686 = ~n13652 & n13685;
  assign n13687 = n13686 ^ n13671;
  assign n13698 = n13697 ^ n13687;
  assign n13672 = n13671 ^ n13652;
  assign n13635 = n13634 ^ n13626;
  assign n13128 = n4478 & n12100;
  assign n13129 = n4484 & n10680;
  assign n13130 = n4480 & n10683;
  assign n13131 = ~n13129 & ~n13130;
  assign n13132 = n4487 & n10665;
  assign n13133 = n13131 & ~n13132;
  assign n13134 = ~n13128 & n13133;
  assign n13135 = n13134 ^ x23;
  assign n13127 = n13126 ^ n13116;
  assign n13136 = n13135 ^ n13127;
  assign n13606 = n13113 ^ n13097;
  assign n13593 = n12935 ^ n12927;
  assign n13138 = n10866 ^ n10841;
  assign n13139 = ~n10751 & n13138;
  assign n13140 = n13139 ^ n10866;
  assign n13141 = n13140 ^ n10740;
  assign n13142 = n44 & n13141;
  assign n13143 = n3280 & n10740;
  assign n13144 = n3277 & n10751;
  assign n13145 = n3275 & ~n10756;
  assign n13146 = ~n13144 & ~n13145;
  assign n13147 = ~n13143 & n13146;
  assign n13148 = ~n13142 & n13147;
  assign n13149 = n13148 ^ x29;
  assign n13137 = n12921 ^ n12829;
  assign n13150 = n13149 ^ n13137;
  assign n13163 = n12918 ^ n12750;
  assign n13164 = n13163 ^ n12902;
  assign n13151 = n41 & n10773;
  assign n13152 = ~n12821 & ~n13151;
  assign n13153 = ~x31 & ~n13152;
  assign n13154 = ~n10838 & ~n10863;
  assign n13155 = n13154 ^ n10773;
  assign n13156 = n41 & ~n13155;
  assign n13157 = n91 & n10776;
  assign n13158 = n54 & n10777;
  assign n13159 = x31 & ~n13158;
  assign n13160 = ~n13157 & n13159;
  assign n13161 = ~n13156 & n13160;
  assign n13162 = ~n13153 & ~n13161;
  assign n13165 = n13164 ^ n13162;
  assign n13175 = ~n12880 & ~n12882;
  assign n13176 = n13175 ^ n12900;
  assign n13166 = ~n10837 & ~n10862;
  assign n13167 = n13166 ^ n10776;
  assign n13168 = n3667 & ~n13167;
  assign n13169 = n3676 & ~n10776;
  assign n13170 = n3669 & n10785;
  assign n13171 = ~n3673 & ~n10777;
  assign n13172 = ~n13170 & ~n13171;
  assign n13173 = ~n13169 & n13172;
  assign n13174 = ~n13168 & n13173;
  assign n13177 = n13176 ^ n13174;
  assign n13570 = n12878 ^ n12750;
  assign n13571 = n13570 ^ n12839;
  assign n13196 = ~n10835 & ~n10860;
  assign n13197 = n13196 ^ n10785;
  assign n13198 = n41 & n13197;
  assign n13199 = n54 & ~n10795;
  assign n13200 = x31 & ~n13199;
  assign n13201 = n91 & ~n10789;
  assign n13202 = n13200 & ~n13201;
  assign n13203 = ~n13198 & n13202;
  assign n13204 = n41 & n10785;
  assign n13205 = ~x31 & ~n12830;
  assign n13206 = ~n13204 & n13205;
  assign n13207 = ~n13203 & ~n13206;
  assign n13178 = n142 & n574;
  assign n13179 = n123 & ~n13178;
  assign n13180 = n3578 & n13179;
  assign n13181 = n184 & n379;
  assign n13182 = ~n582 & n13181;
  assign n13183 = n13180 & n13182;
  assign n13184 = ~n312 & n673;
  assign n13185 = n10902 & n13184;
  assign n13186 = n1276 & n13185;
  assign n13187 = n13183 & n13186;
  assign n13188 = n2271 & n11148;
  assign n13189 = n1569 & n12241;
  assign n13190 = n13188 & n13189;
  assign n13191 = n12154 & n13190;
  assign n13192 = n1494 & n13191;
  assign n13193 = n13187 & n13192;
  assign n13194 = n2859 & n13193;
  assign n13195 = n4749 & n13194;
  assign n13208 = n13207 ^ n13195;
  assign n13223 = ~n10834 & ~n10859;
  assign n13224 = n13223 ^ n10789;
  assign n13225 = n41 & ~n13224;
  assign n13226 = n91 & ~n10795;
  assign n13227 = n54 & ~n10799;
  assign n13228 = x31 & ~n13227;
  assign n13229 = ~n13226 & n13228;
  assign n13230 = ~n13225 & n13229;
  assign n13231 = n41 & ~n10789;
  assign n13232 = ~n13199 & ~n13231;
  assign n13233 = ~x31 & n13232;
  assign n13234 = ~n13230 & ~n13233;
  assign n13209 = ~n560 & ~n928;
  assign n13210 = ~n2506 & n13209;
  assign n13211 = n519 & n2022;
  assign n13212 = n13210 & n13211;
  assign n10968 = n267 & ~n301;
  assign n13213 = n2094 & n10968;
  assign n13214 = n13212 & n13213;
  assign n13215 = n1134 & n1306;
  assign n13216 = n3936 & n13215;
  assign n13217 = n753 & n13216;
  assign n13218 = n13214 & n13217;
  assign n13219 = n5096 & n11307;
  assign n13220 = n13218 & n13219;
  assign n13221 = n490 & n13220;
  assign n13222 = n1939 & n13221;
  assign n13235 = n13234 ^ n13222;
  assign n13248 = ~n656 & n1866;
  assign n13249 = n4358 & n10896;
  assign n13250 = n13248 & n13249;
  assign n13251 = n2182 & n11040;
  assign n13252 = n591 & n1976;
  assign n13253 = n13251 & n13252;
  assign n13254 = n13250 & n13253;
  assign n13255 = n2096 & n4397;
  assign n13256 = n1811 & n13255;
  assign n13257 = n13254 & n13256;
  assign n13258 = n1012 & n13257;
  assign n13259 = n2142 & n13258;
  assign n13260 = n12860 & n13259;
  assign n13238 = ~n10833 & ~n10858;
  assign n13239 = n13238 ^ n10795;
  assign n13240 = n41 & n13239;
  assign n13241 = n91 & n10799;
  assign n13242 = n54 & n10800;
  assign n13243 = ~n13241 & ~n13242;
  assign n13244 = ~n13240 & n13243;
  assign n13236 = n41 & ~n10795;
  assign n13237 = ~n13227 & ~n13236;
  assign n13245 = n13244 ^ n13237;
  assign n13246 = ~x31 & ~n13245;
  assign n13247 = n13246 ^ n13244;
  assign n13261 = n13260 ^ n13247;
  assign n13277 = ~n10832 & ~n10857;
  assign n13278 = n13277 ^ n10799;
  assign n13279 = x31 & n13278;
  assign n13280 = ~x31 & n10799;
  assign n13281 = n41 & ~n13280;
  assign n13282 = ~n13279 & n13281;
  assign n13283 = n54 & n10815;
  assign n13284 = x31 & n13283;
  assign n13285 = ~n3673 & ~n10800;
  assign n13286 = ~n13284 & ~n13285;
  assign n13287 = ~n13282 & n13286;
  assign n13262 = ~n216 & ~n2506;
  assign n13263 = n2813 & n13262;
  assign n13264 = n2096 & n2855;
  assign n13265 = n13263 & n13264;
  assign n13266 = n1782 & n2923;
  assign n13267 = n1342 & n13266;
  assign n13268 = n11291 & n13267;
  assign n13269 = n13265 & n13268;
  assign n13270 = ~n164 & n4226;
  assign n13271 = ~n104 & n1854;
  assign n13272 = n13270 & n13271;
  assign n13273 = n3526 & n13272;
  assign n13274 = n13269 & n13273;
  assign n13275 = n3150 & n13274;
  assign n13276 = n3934 & n13275;
  assign n13288 = n13287 ^ n13276;
  assign n13340 = ~n10831 & ~n10856;
  assign n13341 = n13340 ^ n10800;
  assign n13342 = n41 & ~n13341;
  assign n13343 = n91 & n10815;
  assign n13344 = n54 & n10819;
  assign n13345 = x31 & ~n13344;
  assign n13346 = ~n13343 & n13345;
  assign n13347 = ~n13342 & n13346;
  assign n13348 = n41 & ~n10800;
  assign n13349 = ~x31 & ~n13348;
  assign n13350 = ~n13283 & n13349;
  assign n13351 = ~n13347 & ~n13350;
  assign n13289 = n889 & n3472;
  assign n13290 = n393 & n13289;
  assign n13291 = n3570 & n13290;
  assign n13292 = n5511 & n13291;
  assign n13293 = n3518 & n12847;
  assign n13294 = ~n250 & ~n458;
  assign n13295 = ~n128 & ~n605;
  assign n13296 = n13294 & n13295;
  assign n13297 = n13293 & n13296;
  assign n13298 = n2419 & n12052;
  assign n13299 = n13297 & n13298;
  assign n13300 = n13292 & n13299;
  assign n13301 = n679 & n13300;
  assign n13302 = ~n652 & ~n948;
  assign n13303 = n11843 & n13302;
  assign n13304 = n2160 & n2550;
  assign n13305 = n13303 & n13304;
  assign n13306 = n5392 & n13305;
  assign n13307 = ~n308 & ~n428;
  assign n13308 = n934 & n13307;
  assign n13309 = n13306 & n13308;
  assign n13310 = ~n166 & ~n689;
  assign n13311 = n10888 & n13310;
  assign n13312 = n2465 & n13311;
  assign n13313 = n3618 & n13312;
  assign n13314 = n1113 & n13313;
  assign n13315 = n12051 & n13314;
  assign n13316 = n13309 & n13315;
  assign n13317 = n5618 & n11141;
  assign n13318 = n519 & n1406;
  assign n13319 = n321 & n1520;
  assign n13320 = n13318 & n13319;
  assign n13321 = n13317 & n13320;
  assign n13322 = n363 & n2529;
  assign n13323 = n602 & n2975;
  assign n13324 = n13322 & n13323;
  assign n13325 = n4115 & n5121;
  assign n13326 = n598 & n13325;
  assign n13327 = n13324 & n13326;
  assign n13328 = n13321 & n13327;
  assign n13329 = n108 & n1467;
  assign n13330 = ~x24 & ~n818;
  assign n13331 = n116 & n13330;
  assign n13332 = ~n13329 & ~n13331;
  assign n13333 = x26 & ~n13332;
  assign n13334 = ~n761 & ~n5451;
  assign n13335 = n108 & ~n13334;
  assign n13336 = ~n13333 & ~n13335;
  assign n13337 = n13328 & n13336;
  assign n13338 = n13316 & n13337;
  assign n13339 = n13301 & n13338;
  assign n13352 = n13351 ^ n13339;
  assign n13386 = ~n10830 & ~n10855;
  assign n13387 = n13386 ^ n10815;
  assign n13388 = n41 & ~n13387;
  assign n13389 = n91 & ~n10819;
  assign n13390 = n54 & n10820;
  assign n13391 = x31 & ~n13390;
  assign n13392 = ~n13389 & n13391;
  assign n13393 = ~n13388 & n13392;
  assign n13394 = n41 & n10815;
  assign n13395 = ~n13344 & ~n13394;
  assign n13396 = ~x31 & ~n13395;
  assign n13397 = ~n13393 & ~n13396;
  assign n13353 = ~n141 & ~n148;
  assign n13354 = ~n369 & ~n843;
  assign n13355 = n13353 & n13354;
  assign n13356 = n2832 & n13355;
  assign n13357 = n964 & n11016;
  assign n13358 = n1072 & n1554;
  assign n13359 = n13357 & n13358;
  assign n13360 = n13356 & n13359;
  assign n13361 = n255 & n1961;
  assign n13362 = n1992 & n3068;
  assign n13363 = n13361 & n13362;
  assign n13364 = n13360 & n13363;
  assign n13365 = n2480 & n12214;
  assign n13366 = n13364 & n13365;
  assign n13367 = ~n190 & ~n529;
  assign n13368 = ~n359 & n13367;
  assign n13369 = n1728 & n13368;
  assign n13370 = n3004 & n10346;
  assign n13371 = n13369 & n13370;
  assign n13372 = n3471 & n3893;
  assign n13373 = n3936 & n13372;
  assign n13374 = n2051 & n2654;
  assign n13375 = n1014 & n1787;
  assign n13376 = n13374 & n13375;
  assign n13377 = n13373 & n13376;
  assign n13378 = n13371 & n13377;
  assign n13379 = n11274 & n12075;
  assign n13380 = ~n362 & ~n385;
  assign n13381 = n13379 & n13380;
  assign n13382 = n2021 & n13381;
  assign n13383 = n13378 & n13382;
  assign n13384 = n11164 & n13383;
  assign n13385 = n13366 & n13384;
  assign n13398 = n13397 ^ n13385;
  assign n13428 = ~n10829 & ~n10854;
  assign n13429 = n13428 ^ n10819;
  assign n13430 = n41 & n13429;
  assign n13431 = n54 & n10821;
  assign n13432 = n91 & ~n10820;
  assign n13433 = ~n13431 & ~n13432;
  assign n13434 = ~n13430 & n13433;
  assign n13435 = x31 & ~n13434;
  assign n13436 = ~n54 & ~n10819;
  assign n13437 = n3640 & ~n13390;
  assign n13438 = ~n13436 & n13437;
  assign n13439 = ~n13435 & ~n13438;
  assign n13399 = ~n901 & n2401;
  assign n13400 = n5121 & n13399;
  assign n13401 = n522 & n13400;
  assign n13402 = n4775 & n10219;
  assign n13403 = n13401 & n13402;
  assign n13404 = n651 & n12208;
  assign n13405 = ~n155 & n1212;
  assign n13406 = n13404 & n13405;
  assign n13407 = n13403 & n13406;
  assign n13408 = n638 & n13407;
  assign n13409 = n2323 & n13408;
  assign n13410 = n2326 & n11555;
  assign n13411 = n3019 & n13410;
  assign n13412 = n2074 & n3111;
  assign n13413 = n3560 & n12048;
  assign n13414 = n13412 & n13413;
  assign n13415 = n13411 & n13414;
  assign n13416 = ~n74 & ~n347;
  assign n13417 = ~n138 & n13416;
  assign n13418 = n1041 & n13417;
  assign n13419 = n13415 & n13418;
  assign n13420 = ~n269 & ~n666;
  assign n13421 = ~n171 & ~n300;
  assign n13422 = n13420 & n13421;
  assign n13423 = n3413 & n13422;
  assign n13424 = n813 & n13423;
  assign n13425 = n12319 & n13424;
  assign n13426 = n13419 & n13425;
  assign n13427 = n13409 & n13426;
  assign n13440 = n13439 ^ n13427;
  assign n13454 = n10827 ^ n10820;
  assign n13455 = ~n91 & ~n13454;
  assign n13456 = ~n54 & ~n10821;
  assign n13457 = ~n13455 & n13456;
  assign n13458 = n10821 & ~n13454;
  assign n13459 = n41 & n13458;
  assign n13460 = ~n13457 & ~n13459;
  assign n13461 = x31 & ~n13460;
  assign n13462 = n41 & ~n10820;
  assign n13463 = ~x31 & ~n13431;
  assign n13464 = ~n13462 & n13463;
  assign n13465 = n3669 & n10822;
  assign n13466 = ~n13464 & ~n13465;
  assign n13467 = ~n13461 & n13466;
  assign n13441 = ~n3302 & n5427;
  assign n13442 = n1376 & n13441;
  assign n13443 = ~n313 & ~n416;
  assign n13444 = n990 & n13443;
  assign n13445 = n955 & n3004;
  assign n13446 = n13444 & n13445;
  assign n13447 = n1586 & n3962;
  assign n13448 = n13446 & n13447;
  assign n13449 = n4211 & n13448;
  assign n13450 = n13442 & n13449;
  assign n13451 = n11321 & n11408;
  assign n13452 = n13450 & n13451;
  assign n13453 = n3558 & n13452;
  assign n13468 = n13467 ^ n13453;
  assign n13495 = n41 & ~n10822;
  assign n13496 = n5636 & n10825;
  assign n13497 = ~n13495 & ~n13496;
  assign n13498 = ~n10822 & n10825;
  assign n13499 = n3667 & n13498;
  assign n13500 = ~n13497 & ~n13499;
  assign n13501 = ~n166 & ~n245;
  assign n13502 = ~n656 & n13501;
  assign n13503 = n1352 & n13502;
  assign n13504 = n1144 & n13503;
  assign n13505 = n13272 & n13504;
  assign n13506 = n194 & ~n841;
  assign n13507 = ~n334 & ~n354;
  assign n13508 = n13506 & n13507;
  assign n13509 = n1857 & n4387;
  assign n13510 = n13508 & n13509;
  assign n13511 = n13505 & n13510;
  assign n13512 = n3309 & n3470;
  assign n13513 = n11250 & n12297;
  assign n13514 = n13512 & n13513;
  assign n13515 = n13511 & n13514;
  assign n13516 = ~n560 & ~n666;
  assign n13517 = n999 & n13516;
  assign n13518 = n12844 & n13517;
  assign n13519 = n4015 & n11318;
  assign n13520 = n13518 & n13519;
  assign n13521 = n1667 & n1707;
  assign n13522 = n13520 & n13521;
  assign n13523 = n5560 & n13522;
  assign n13524 = n774 & n13523;
  assign n13525 = n13515 & n13524;
  assign n13473 = ~n189 & ~n549;
  assign n13526 = n2212 & n4109;
  assign n13527 = n13473 & n13526;
  assign n13528 = n3227 & n13527;
  assign n13529 = n13525 & n13528;
  assign n13530 = n13500 & ~n13529;
  assign n13469 = n1855 & n11155;
  assign n13470 = n2377 & n2993;
  assign n13471 = n13469 & n13470;
  assign n13472 = n2270 & n4077;
  assign n13474 = n3020 & n13473;
  assign n13475 = n13472 & n13474;
  assign n13476 = ~n518 & ~n680;
  assign n13477 = ~n273 & ~n442;
  assign n13478 = n13476 & n13477;
  assign n13479 = n4056 & n13478;
  assign n13480 = n13475 & n13479;
  assign n13481 = n13471 & n13480;
  assign n13482 = n12868 & n13481;
  assign n13483 = ~n190 & ~n557;
  assign n13484 = ~n797 & n13483;
  assign n13485 = n1853 & n2461;
  assign n13486 = n13484 & n13485;
  assign n13487 = n1031 & n13486;
  assign n11001 = ~n57 & ~n293;
  assign n13488 = ~n617 & ~n791;
  assign n13489 = n2055 & n13488;
  assign n13490 = n11001 & n13489;
  assign n13491 = n1790 & n13490;
  assign n13492 = n13487 & n13491;
  assign n13493 = n13482 & n13492;
  assign n13494 = n12306 & n13493;
  assign n13531 = n13530 ^ n13494;
  assign n13532 = ~n10822 & ~n10825;
  assign n13533 = ~n10821 & n13532;
  assign n13534 = ~n10822 & ~n11234;
  assign n13535 = ~n13533 & ~n13534;
  assign n13536 = n5636 & ~n13535;
  assign n13537 = x31 & n13532;
  assign n13538 = n10821 & ~n13537;
  assign n13539 = n41 & n13538;
  assign n13540 = n3669 & n10825;
  assign n13541 = ~n13539 & ~n13540;
  assign n13542 = ~n13536 & n13541;
  assign n13543 = n13542 ^ n13530;
  assign n13544 = n13531 & ~n13543;
  assign n13545 = n13544 ^ n13542;
  assign n13546 = n13545 ^ n13453;
  assign n13547 = ~n13468 & ~n13546;
  assign n13548 = n13547 ^ n13467;
  assign n13549 = n13548 ^ n13439;
  assign n13550 = ~n13440 & ~n13549;
  assign n13551 = n13550 ^ n13548;
  assign n13552 = n13551 ^ n13397;
  assign n13553 = ~n13398 & ~n13552;
  assign n13554 = n13553 ^ n13551;
  assign n13555 = n13554 ^ n13351;
  assign n13556 = n13352 & n13555;
  assign n13557 = n13556 ^ n13554;
  assign n13558 = n13557 ^ n13287;
  assign n13559 = ~n13288 & ~n13558;
  assign n13560 = n13559 ^ n13557;
  assign n13561 = n13560 ^ n13247;
  assign n13562 = n13261 & n13561;
  assign n13563 = n13562 ^ n13560;
  assign n13564 = n13563 ^ n13234;
  assign n13565 = n13235 & n13564;
  assign n13566 = n13565 ^ n13563;
  assign n13567 = n13566 ^ n13207;
  assign n13568 = n13208 & n13567;
  assign n13569 = n13568 ^ n13566;
  assign n13572 = n13571 ^ n13569;
  assign n13573 = n44 & n12818;
  assign n13574 = n3280 & n10757;
  assign n13575 = n3275 & ~n10776;
  assign n13576 = ~n13574 & ~n13575;
  assign n13577 = n3277 & n10773;
  assign n13578 = n13576 & ~n13577;
  assign n13579 = ~n13573 & n13578;
  assign n13580 = n13579 ^ x29;
  assign n13581 = n13580 ^ n13569;
  assign n13582 = ~n13572 & ~n13581;
  assign n13583 = n13582 ^ n13580;
  assign n13584 = n13583 ^ n13176;
  assign n13585 = ~n13177 & n13584;
  assign n13586 = n13585 ^ n13583;
  assign n13587 = n13586 ^ n13164;
  assign n13588 = n13165 & ~n13587;
  assign n13589 = n13588 ^ n13586;
  assign n13590 = n13589 ^ n13149;
  assign n13591 = n13150 & n13590;
  assign n13592 = n13591 ^ n13589;
  assign n13594 = n13593 ^ n13592;
  assign n13595 = n3285 & n12111;
  assign n13596 = n3437 & n10715;
  assign n13597 = ~n3440 & ~n10736;
  assign n13598 = n3435 & n10718;
  assign n13599 = ~n13597 & ~n13598;
  assign n13600 = ~n13596 & n13599;
  assign n13601 = ~n13595 & n13600;
  assign n13602 = n13601 ^ x26;
  assign n13603 = n13602 ^ n13592;
  assign n13604 = n13594 & n13603;
  assign n13605 = n13604 ^ n13602;
  assign n13607 = n13606 ^ n13605;
  assign n13608 = n4478 & n12524;
  assign n13609 = n4487 & n10680;
  assign n13610 = n4484 & n10683;
  assign n13611 = n4480 & n10694;
  assign n13612 = ~n13610 & ~n13611;
  assign n13613 = ~n13609 & n13612;
  assign n13614 = ~n13608 & n13613;
  assign n13615 = n13614 ^ x23;
  assign n13616 = n13615 ^ n13606;
  assign n13617 = ~n13607 & n13616;
  assign n13618 = n13617 ^ n13615;
  assign n13619 = n13618 ^ n13127;
  assign n13620 = n13136 & ~n13619;
  assign n13621 = n13620 ^ n13135;
  assign n13636 = n13635 ^ n13621;
  assign n13637 = n4673 & n11704;
  assign n13638 = n4688 & n11486;
  assign n13639 = n4685 & n11215;
  assign n13640 = ~n4681 & ~n10956;
  assign n13641 = ~n13639 & ~n13640;
  assign n13642 = ~n13638 & n13641;
  assign n13643 = ~n13637 & n13642;
  assign n13644 = n13643 ^ x20;
  assign n13645 = n13644 ^ n13621;
  assign n13646 = ~n13636 & n13645;
  assign n13647 = n13646 ^ n13644;
  assign n13673 = n13672 ^ n13647;
  assign n13674 = n4963 & ~n12000;
  assign n13675 = n4972 & ~n11875;
  assign n13676 = n4976 & ~n11773;
  assign n13677 = n4970 & n11480;
  assign n13678 = ~n13676 & ~n13677;
  assign n13679 = ~n13675 & n13678;
  assign n13680 = ~n13674 & n13679;
  assign n13681 = n13680 ^ x17;
  assign n13682 = n13681 ^ n13672;
  assign n13683 = ~n13673 & n13682;
  assign n13684 = n13683 ^ n13681;
  assign n13699 = n13698 ^ n13684;
  assign n13700 = n5771 & n12504;
  assign n13701 = n4976 & ~n11875;
  assign n13702 = n4970 & ~n11773;
  assign n13703 = ~n13701 & ~n13702;
  assign n13704 = x17 & n13703;
  assign n13705 = ~n11902 & n13704;
  assign n13706 = ~n13700 & ~n13705;
  assign n13707 = x16 & n13706;
  assign n13708 = ~n12504 & n13704;
  assign n13709 = n5771 & n11902;
  assign n13710 = ~x16 & ~n13709;
  assign n13711 = ~n13708 & n13710;
  assign n13712 = ~n13707 & ~n13711;
  assign n13713 = ~n5786 & n13703;
  assign n13714 = n13713 ^ x17;
  assign n13715 = ~n13712 & n13714;
  assign n13716 = n13715 ^ n13684;
  assign n13717 = ~n13699 & n13716;
  assign n13718 = n13717 ^ n13715;
  assign n13731 = n13730 ^ n13718;
  assign n13737 = n5771 & ~n11941;
  assign n13738 = n4976 & n11902;
  assign n13739 = n4970 & ~n11875;
  assign n13740 = ~n13738 & ~n13739;
  assign n13741 = x17 & n13740;
  assign n13742 = n11940 & n13741;
  assign n13743 = x16 & ~n13742;
  assign n13744 = ~n13737 & n13743;
  assign n13745 = n11941 & n13741;
  assign n13746 = n5771 & ~n11940;
  assign n13747 = ~x16 & ~n13746;
  assign n13748 = ~n13745 & n13747;
  assign n13749 = ~n13744 & ~n13748;
  assign n13750 = ~n5786 & n13740;
  assign n13751 = n13750 ^ x17;
  assign n13752 = ~n13749 & n13751;
  assign n13735 = n13060 ^ n13052;
  assign n13732 = n13696 ^ n13687;
  assign n13733 = ~n13697 & n13732;
  assign n13734 = n13733 ^ n13687;
  assign n13736 = n13735 ^ n13734;
  assign n13753 = n13752 ^ n13736;
  assign n13754 = n13753 ^ n13718;
  assign n13755 = n13731 & ~n13754;
  assign n13756 = n13755 ^ n13753;
  assign n13757 = n13087 & n13756;
  assign n13758 = n13753 ^ n13731;
  assign n13863 = ~n12013 & ~n12019;
  assign n13864 = n7860 & n13863;
  assign n13865 = ~n5746 & ~n11940;
  assign n13866 = n5752 & n11902;
  assign n13867 = ~n13865 & ~n13866;
  assign n13868 = n5748 & ~n12019;
  assign n13869 = ~x14 & ~n13868;
  assign n13870 = n13867 & n13869;
  assign n13871 = ~n13864 & ~n13870;
  assign n13872 = x13 & n13868;
  assign n13873 = n12013 & n13872;
  assign n13874 = x14 & ~n13867;
  assign n13875 = ~n13873 & ~n13874;
  assign n13876 = n13871 & n13875;
  assign n13861 = n13681 ^ n13673;
  assign n13848 = n13644 ^ n13636;
  assign n13835 = n4673 & ~n12460;
  assign n13836 = n4688 & n11215;
  assign n13837 = ~n4681 & ~n10663;
  assign n13838 = n4685 & ~n10956;
  assign n13839 = ~n13837 & ~n13838;
  assign n13840 = ~n13836 & n13839;
  assign n13841 = ~n13835 & n13840;
  assign n13842 = n13841 ^ x20;
  assign n13822 = n13615 ^ n13607;
  assign n13809 = n13602 ^ n13594;
  assign n13788 = n12180 & n12417;
  assign n13789 = n3435 & ~n10736;
  assign n13790 = ~n3440 & n10738;
  assign n13791 = ~n13789 & ~n13790;
  assign n13792 = x26 & n13791;
  assign n13793 = ~n10718 & n13792;
  assign n13794 = ~n13788 & ~n13793;
  assign n13795 = x25 & n13794;
  assign n13796 = ~n12180 & n13792;
  assign n13797 = n10718 & n12417;
  assign n13798 = ~x25 & ~n13797;
  assign n13799 = ~n13796 & n13798;
  assign n13800 = ~n13795 & ~n13799;
  assign n13801 = ~n12432 & n13791;
  assign n13802 = n13801 ^ x26;
  assign n13803 = ~n13800 & n13802;
  assign n13767 = n13586 ^ n13165;
  assign n13759 = n44 & n12940;
  assign n13760 = n3280 & n10751;
  assign n13761 = n3277 & ~n10756;
  assign n13762 = n3275 & n10757;
  assign n13763 = ~n13761 & ~n13762;
  assign n13764 = ~n13760 & n13763;
  assign n13765 = ~n13759 & n13764;
  assign n13766 = n13765 ^ x29;
  assign n13768 = n13767 ^ n13766;
  assign n13769 = n12417 & ~n12596;
  assign n13770 = n3435 & n10738;
  assign n13771 = ~n3440 & n10740;
  assign n13772 = ~n13770 & ~n13771;
  assign n13773 = x26 & n13772;
  assign n13774 = n10736 & n13773;
  assign n13775 = x25 & ~n13774;
  assign n13776 = ~n13769 & n13775;
  assign n13777 = n12596 & n13773;
  assign n13778 = ~n10736 & n12417;
  assign n13779 = ~x25 & ~n13778;
  assign n13780 = ~n13777 & n13779;
  assign n13781 = ~n13776 & ~n13780;
  assign n13782 = ~n12432 & n13772;
  assign n13783 = n13782 ^ x26;
  assign n13784 = ~n13781 & n13783;
  assign n13785 = n13784 ^ n13767;
  assign n13786 = n13768 & ~n13785;
  assign n13787 = n13786 ^ n13784;
  assign n13804 = n13803 ^ n13787;
  assign n13805 = n13589 ^ n13150;
  assign n13806 = n13805 ^ n13787;
  assign n13807 = n13804 & n13806;
  assign n13808 = n13807 ^ n13803;
  assign n13810 = n13809 ^ n13808;
  assign n13811 = n4478 & n11599;
  assign n13812 = n4484 & n10694;
  assign n13813 = n4480 & n10698;
  assign n13814 = ~n13812 & ~n13813;
  assign n13815 = n4487 & n10683;
  assign n13816 = n13814 & ~n13815;
  assign n13817 = ~n13811 & n13816;
  assign n13818 = n13817 ^ x23;
  assign n13819 = n13818 ^ n13808;
  assign n13820 = n13810 & n13819;
  assign n13821 = n13820 ^ n13818;
  assign n13823 = n13822 ^ n13821;
  assign n13824 = n4673 & ~n10957;
  assign n13825 = n4685 & ~n10663;
  assign n13826 = n4688 & ~n10956;
  assign n13827 = ~n4681 & n10665;
  assign n13828 = ~n13826 & ~n13827;
  assign n13829 = ~n13825 & n13828;
  assign n13830 = ~n13824 & n13829;
  assign n13831 = n13830 ^ x20;
  assign n13832 = n13831 ^ n13822;
  assign n13833 = ~n13823 & n13832;
  assign n13834 = n13833 ^ n13831;
  assign n13843 = n13842 ^ n13834;
  assign n13844 = n13618 ^ n13136;
  assign n13845 = n13844 ^ n13842;
  assign n13846 = n13843 & ~n13845;
  assign n13847 = n13846 ^ n13834;
  assign n13849 = n13848 ^ n13847;
  assign n13850 = n4963 & ~n11777;
  assign n13851 = n4972 & ~n11773;
  assign n13852 = n4970 & n11500;
  assign n13853 = n4976 & n11480;
  assign n13854 = ~n13852 & ~n13853;
  assign n13855 = ~n13851 & n13854;
  assign n13856 = ~n13850 & n13855;
  assign n13857 = n13856 ^ x17;
  assign n13858 = n13857 ^ n13848;
  assign n13859 = ~n13849 & n13858;
  assign n13860 = n13859 ^ n13857;
  assign n13862 = n13861 ^ n13860;
  assign n13877 = n13876 ^ n13862;
  assign n13878 = n13877 ^ n12123;
  assign n13981 = n13857 ^ n13849;
  assign n13880 = n5771 & n11507;
  assign n13881 = n4976 & n11500;
  assign n13882 = n4970 & n11486;
  assign n13883 = ~n13881 & ~n13882;
  assign n13884 = x17 & n13883;
  assign n13885 = ~n11480 & n13884;
  assign n13886 = x16 & ~n13885;
  assign n13887 = ~n13880 & n13886;
  assign n13888 = ~n11507 & n13884;
  assign n13889 = n5771 & n11480;
  assign n13890 = ~x16 & ~n13889;
  assign n13891 = ~n13888 & n13890;
  assign n13892 = ~n13887 & ~n13891;
  assign n13893 = ~n5786 & n13883;
  assign n13894 = n13893 ^ x17;
  assign n13895 = ~n13892 & n13894;
  assign n13879 = n13844 ^ n13843;
  assign n13896 = n13895 ^ n13879;
  assign n13965 = n13831 ^ n13823;
  assign n13952 = n13818 ^ n13810;
  assign n13931 = n13805 ^ n13804;
  assign n13918 = n13784 ^ n13768;
  assign n13905 = n13583 ^ n13177;
  assign n13897 = n44 & ~n12703;
  assign n13898 = n3280 & ~n10756;
  assign n13899 = n3277 & n10757;
  assign n13900 = n3275 & n10773;
  assign n13901 = ~n13899 & ~n13900;
  assign n13902 = ~n13898 & n13901;
  assign n13903 = ~n13897 & n13902;
  assign n13904 = n13903 ^ x29;
  assign n13906 = n13905 ^ n13904;
  assign n13907 = n3285 & n12194;
  assign n13908 = n3437 & n10738;
  assign n13909 = n3435 & n10740;
  assign n13910 = ~n3440 & n10751;
  assign n13911 = ~n13909 & ~n13910;
  assign n13912 = ~n13908 & n13911;
  assign n13913 = ~n13907 & n13912;
  assign n13914 = n13913 ^ x26;
  assign n13915 = n13914 ^ n13905;
  assign n13916 = ~n13906 & n13915;
  assign n13917 = n13916 ^ n13914;
  assign n13919 = n13918 ^ n13917;
  assign n13920 = n4478 & n12034;
  assign n13921 = n4484 & n10715;
  assign n13922 = n4487 & n10698;
  assign n13923 = n4480 & n10718;
  assign n13924 = ~n13922 & ~n13923;
  assign n13925 = ~n13921 & n13924;
  assign n13926 = ~n13920 & n13925;
  assign n13927 = n13926 ^ x23;
  assign n13928 = n13927 ^ n13918;
  assign n13929 = n13919 & ~n13928;
  assign n13930 = n13929 ^ n13927;
  assign n13932 = n13931 ^ n13930;
  assign n12502 = ~x23 & n4476;
  assign n13933 = n12087 & n12502;
  assign n13934 = n4480 & n10715;
  assign n13935 = n4484 & n10698;
  assign n13936 = ~n13934 & ~n13935;
  assign n13937 = x23 & n13936;
  assign n13938 = ~n10694 & n13937;
  assign n13939 = x22 & ~n13938;
  assign n13940 = ~n13933 & n13939;
  assign n13941 = ~n12087 & n13937;
  assign n13942 = n10694 & n12502;
  assign n13943 = ~x22 & ~n13942;
  assign n13944 = ~n13941 & n13943;
  assign n13945 = ~n13940 & ~n13944;
  assign n12518 = x23 & ~n4476;
  assign n12519 = n12518 ^ x23;
  assign n13946 = ~n12519 & n13936;
  assign n13947 = n13946 ^ x23;
  assign n13948 = ~n13945 & n13947;
  assign n13949 = n13948 ^ n13930;
  assign n13950 = n13932 & n13949;
  assign n13951 = n13950 ^ n13948;
  assign n13953 = n13952 ^ n13951;
  assign n13954 = n4673 & ~n11694;
  assign n13955 = n4688 & ~n10663;
  assign n13956 = ~n4681 & n10680;
  assign n13957 = n4685 & n10665;
  assign n13958 = ~n13956 & ~n13957;
  assign n13959 = ~n13955 & n13958;
  assign n13960 = ~n13954 & n13959;
  assign n13961 = n13960 ^ x20;
  assign n13962 = n13961 ^ n13951;
  assign n13963 = n13953 & n13962;
  assign n13964 = n13963 ^ n13961;
  assign n13966 = n13965 ^ n13964;
  assign n13967 = n4963 & n11957;
  assign n13968 = n4972 & n11500;
  assign n13969 = n4976 & n11486;
  assign n13970 = n4970 & n11215;
  assign n13971 = ~n13969 & ~n13970;
  assign n13972 = ~n13968 & n13971;
  assign n13973 = ~n13967 & n13972;
  assign n13974 = n13973 ^ x17;
  assign n13975 = n13974 ^ n13965;
  assign n13976 = ~n13966 & n13975;
  assign n13977 = n13976 ^ n13974;
  assign n13978 = n13977 ^ n13879;
  assign n13979 = n13896 & ~n13978;
  assign n13980 = n13979 ^ n13895;
  assign n13982 = n13981 ^ n13980;
  assign n13995 = n5749 & ~n11907;
  assign n13996 = n13995 ^ x13;
  assign n13997 = n13996 ^ n11940;
  assign n13983 = ~x13 & n11902;
  assign n13984 = x12 & ~n13983;
  assign n13985 = x13 & ~n11875;
  assign n13986 = ~x14 & n13985;
  assign n13987 = n13984 & ~n13986;
  assign n13988 = x13 & n11902;
  assign n13989 = ~x13 & x14;
  assign n13990 = ~n11875 & n13989;
  assign n13991 = ~x12 & ~n13990;
  assign n13992 = ~n13988 & n13991;
  assign n13993 = ~n13987 & ~n13992;
  assign n13994 = n13993 ^ x14;
  assign n13998 = n13997 ^ n13994;
  assign n13999 = ~n5748 & ~n13998;
  assign n14000 = n13999 ^ n13997;
  assign n14001 = n14000 ^ n13980;
  assign n14002 = ~n13982 & n14001;
  assign n14003 = n14002 ^ n14000;
  assign n14004 = n14003 ^ n13877;
  assign n14005 = n13878 & n14004;
  assign n14006 = n14005 ^ n12123;
  assign n14007 = n13876 ^ n13861;
  assign n14008 = ~n13862 & ~n14007;
  assign n14009 = n14008 ^ n13876;
  assign n14010 = n14006 & n14009;
  assign n14011 = n13758 & ~n14010;
  assign n14302 = n14003 ^ n12123;
  assign n14303 = n14302 ^ n13877;
  assign n14019 = n14000 ^ n13982;
  assign n14012 = n5820 & n13720;
  assign n14013 = ~n12123 & ~n14012;
  assign n14014 = x8 & n12019;
  assign n14015 = x10 & ~x11;
  assign n14016 = n14014 & n14015;
  assign n14017 = x9 & n14016;
  assign n14018 = ~n14013 & ~n14017;
  assign n14020 = n14019 ^ n14018;
  assign n14280 = ~x13 & n12504;
  assign n14281 = x14 & ~n13988;
  assign n14282 = ~n14280 & n14281;
  assign n14283 = ~n5746 & ~n11875;
  assign n14284 = n5752 & ~n11773;
  assign n14285 = ~n14283 & ~n14284;
  assign n14286 = ~n7559 & n14285;
  assign n14287 = ~n14282 & n14286;
  assign n14288 = x14 & ~n14285;
  assign n14289 = ~n14287 & ~n14288;
  assign n14290 = x13 & n12503;
  assign n14291 = n14290 ^ n11902;
  assign n14292 = n6033 & n14291;
  assign n14293 = ~n14289 & ~n14292;
  assign n14251 = n13974 ^ n13966;
  assign n14238 = n13961 ^ n13953;
  assign n14022 = n4673 & n12100;
  assign n14023 = n4685 & n10680;
  assign n14024 = ~n4681 & n10683;
  assign n14025 = ~n14023 & ~n14024;
  assign n14026 = n4688 & n10665;
  assign n14027 = n14025 & ~n14026;
  assign n14028 = ~n14022 & n14027;
  assign n14029 = n14028 ^ x20;
  assign n14021 = n13948 ^ n13932;
  assign n14030 = n14029 ^ n14021;
  assign n14222 = n13927 ^ n13919;
  assign n14209 = n13914 ^ n13906;
  assign n14039 = n13563 ^ n13235;
  assign n14040 = n44 & ~n13167;
  assign n14041 = n3280 & ~n10776;
  assign n14042 = n3277 & ~n10777;
  assign n14043 = n3275 & n10785;
  assign n14044 = ~n14042 & ~n14043;
  assign n14045 = ~n14041 & n14044;
  assign n14046 = ~n14040 & n14045;
  assign n14047 = n14046 ^ x29;
  assign n14048 = ~n14039 & ~n14047;
  assign n14050 = n44 & ~n12832;
  assign n14051 = n3280 & ~n10777;
  assign n14052 = n3275 & ~n10789;
  assign n14053 = ~n14051 & ~n14052;
  assign n14054 = n3277 & n10785;
  assign n14055 = n14053 & ~n14054;
  assign n14056 = ~n14050 & n14055;
  assign n14057 = n14056 ^ x29;
  assign n14049 = n13560 ^ n13261;
  assign n14058 = n14057 ^ n14049;
  assign n14060 = n44 & n13197;
  assign n14061 = n3280 & n10785;
  assign n14062 = n3277 & ~n10789;
  assign n14063 = n3275 & ~n10795;
  assign n14064 = ~n14062 & ~n14063;
  assign n14065 = ~n14061 & n14064;
  assign n14066 = ~n14060 & n14065;
  assign n14067 = n14066 ^ x29;
  assign n14059 = n13557 ^ n13288;
  assign n14068 = n14067 ^ n14059;
  assign n14077 = n13554 ^ n13352;
  assign n14069 = n44 & ~n13224;
  assign n14070 = n3280 & ~n10789;
  assign n14071 = n3275 & ~n10799;
  assign n14072 = ~n14070 & ~n14071;
  assign n14073 = n3277 & ~n10795;
  assign n14074 = n14072 & ~n14073;
  assign n14075 = ~n14069 & n14074;
  assign n14076 = n14075 ^ x29;
  assign n14078 = n14077 ^ n14076;
  assign n14080 = n44 & ~n13239;
  assign n14081 = n3280 & ~n10795;
  assign n14082 = n3277 & ~n10799;
  assign n14083 = n3275 & ~n10800;
  assign n14084 = ~n14082 & ~n14083;
  assign n14085 = ~n14081 & n14084;
  assign n14086 = ~n14080 & n14085;
  assign n14087 = n14086 ^ x29;
  assign n14079 = n13551 ^ n13398;
  assign n14088 = n14087 ^ n14079;
  assign n14090 = n44 & ~n13278;
  assign n14091 = n3280 & ~n10799;
  assign n14092 = n3277 & ~n10800;
  assign n14093 = n3275 & n10815;
  assign n14094 = ~n14092 & ~n14093;
  assign n14095 = ~n14091 & n14094;
  assign n14096 = ~n14090 & n14095;
  assign n14097 = n14096 ^ x29;
  assign n14089 = n13548 ^ n13440;
  assign n14098 = n14097 ^ n14089;
  assign n14100 = n44 & ~n13341;
  assign n14101 = n3280 & ~n10800;
  assign n14102 = n3275 & n10819;
  assign n14103 = ~n14101 & ~n14102;
  assign n14104 = n3277 & n10815;
  assign n14105 = n14103 & ~n14104;
  assign n14106 = ~n14100 & n14105;
  assign n14107 = n14106 ^ x29;
  assign n14099 = n13545 ^ n13468;
  assign n14108 = n14107 ^ n14099;
  assign n14149 = n13542 ^ n13531;
  assign n14110 = n10827 ^ n10821;
  assign n14111 = n14110 ^ n10820;
  assign n14112 = n44 & ~n14111;
  assign n14113 = n3280 & ~n10820;
  assign n14114 = n3277 & n10821;
  assign n14115 = n3275 & ~n10822;
  assign n14116 = ~n14114 & ~n14115;
  assign n14117 = ~n14113 & n14116;
  assign n14118 = ~n14112 & n14117;
  assign n14119 = n14118 ^ x29;
  assign n14120 = n13532 ^ n10821;
  assign n14121 = n44 & n14120;
  assign n14122 = n3280 & n10821;
  assign n14123 = n3277 & ~n10822;
  assign n14124 = n3275 & n10825;
  assign n14125 = ~n14123 & ~n14124;
  assign n14126 = ~n14122 & n14125;
  assign n14127 = ~n14121 & n14126;
  assign n14128 = n10822 & ~n10825;
  assign n14129 = n3277 & n10825;
  assign n14130 = ~n42 & ~n14129;
  assign n14131 = ~n14128 & ~n14130;
  assign n14132 = x29 & ~n14131;
  assign n14133 = n14127 & n14132;
  assign n14134 = n41 & n10825;
  assign n14135 = ~n14133 & ~n14134;
  assign n14136 = ~n14119 & ~n14135;
  assign n14109 = n13529 ^ n13500;
  assign n14137 = n14136 ^ n14109;
  assign n14138 = n44 & n13429;
  assign n14139 = n3280 & n10819;
  assign n14140 = n3277 & ~n10820;
  assign n14141 = n3275 & n10821;
  assign n14142 = ~n14140 & ~n14141;
  assign n14143 = ~n14139 & n14142;
  assign n14144 = ~n14138 & n14143;
  assign n14145 = n14144 ^ x29;
  assign n14146 = n14145 ^ n14136;
  assign n14147 = n14137 & ~n14146;
  assign n14148 = n14147 ^ n14145;
  assign n14150 = n14149 ^ n14148;
  assign n14151 = n44 & n13387;
  assign n14152 = n3280 & n10815;
  assign n14153 = n3277 & n10819;
  assign n14154 = n3275 & ~n10820;
  assign n14155 = ~n14153 & ~n14154;
  assign n14156 = ~n14152 & n14155;
  assign n14157 = ~n14151 & n14156;
  assign n14158 = n14157 ^ x29;
  assign n14159 = n14158 ^ n14149;
  assign n14160 = ~n14150 & n14159;
  assign n14161 = n14160 ^ n14148;
  assign n14162 = n14161 ^ n14107;
  assign n14163 = n14108 & n14162;
  assign n14164 = n14163 ^ n14161;
  assign n14165 = n14164 ^ n14097;
  assign n14166 = n14098 & n14165;
  assign n14167 = n14166 ^ n14164;
  assign n14168 = n14167 ^ n14087;
  assign n14169 = n14088 & n14168;
  assign n14170 = n14169 ^ n14167;
  assign n14171 = n14170 ^ n14077;
  assign n14172 = ~n14078 & n14171;
  assign n14173 = n14172 ^ n14170;
  assign n14174 = n14173 ^ n14067;
  assign n14175 = n14068 & n14174;
  assign n14176 = n14175 ^ n14173;
  assign n14177 = n14176 ^ n14057;
  assign n14178 = ~n14058 & n14177;
  assign n14179 = n14178 ^ n14176;
  assign n14180 = ~n14048 & n14179;
  assign n14181 = n13566 ^ n13208;
  assign n14182 = n44 & n13155;
  assign n14183 = n3280 & n10773;
  assign n14184 = n3277 & ~n10776;
  assign n14185 = n3275 & ~n10777;
  assign n14186 = ~n14184 & ~n14185;
  assign n14187 = ~n14183 & n14186;
  assign n14188 = ~n14182 & n14187;
  assign n14189 = n14181 & ~n14188;
  assign n14190 = n14039 & ~n14046;
  assign n14191 = ~n14189 & ~n14190;
  assign n14192 = ~n14180 & n14191;
  assign n14193 = ~n14181 & n14188;
  assign n14194 = x29 & ~n14193;
  assign n14195 = ~n14192 & n14194;
  assign n14196 = n14181 & n14188;
  assign n14197 = n14039 & n14046;
  assign n14198 = ~n14196 & ~n14197;
  assign n14199 = ~n14180 & n14198;
  assign n14200 = ~n14181 & ~n14188;
  assign n14201 = ~x29 & ~n14200;
  assign n14202 = ~n14199 & n14201;
  assign n14203 = ~n14195 & ~n14202;
  assign n14031 = n3285 & n13141;
  assign n14032 = n3437 & n10740;
  assign n14033 = n3435 & n10751;
  assign n14034 = ~n3440 & ~n10756;
  assign n14035 = ~n14033 & ~n14034;
  assign n14036 = ~n14032 & n14035;
  assign n14037 = ~n14031 & n14036;
  assign n14038 = n14037 ^ x26;
  assign n14204 = n14203 ^ n14038;
  assign n14205 = n13580 ^ n13572;
  assign n14206 = n14205 ^ n14038;
  assign n14207 = ~n14204 & ~n14206;
  assign n14208 = n14207 ^ n14203;
  assign n14210 = n14209 ^ n14208;
  assign n14211 = n4478 & n12111;
  assign n14212 = n4487 & n10715;
  assign n14213 = n4480 & ~n10736;
  assign n14214 = n4484 & n10718;
  assign n14215 = ~n14213 & ~n14214;
  assign n14216 = ~n14212 & n14215;
  assign n14217 = ~n14211 & n14216;
  assign n14218 = n14217 ^ x23;
  assign n14219 = n14218 ^ n14209;
  assign n14220 = n14210 & n14219;
  assign n14221 = n14220 ^ n14218;
  assign n14223 = n14222 ^ n14221;
  assign n14224 = n4673 & n12524;
  assign n14225 = n4688 & n10680;
  assign n14226 = n4685 & n10683;
  assign n14227 = ~n4681 & n10694;
  assign n14228 = ~n14226 & ~n14227;
  assign n14229 = ~n14225 & n14228;
  assign n14230 = ~n14224 & n14229;
  assign n14231 = n14230 ^ x20;
  assign n14232 = n14231 ^ n14222;
  assign n14233 = n14223 & ~n14232;
  assign n14234 = n14233 ^ n14231;
  assign n14235 = n14234 ^ n14021;
  assign n14236 = ~n14030 & n14235;
  assign n14237 = n14236 ^ n14029;
  assign n14239 = n14238 ^ n14237;
  assign n14240 = n4963 & n11704;
  assign n14241 = n4972 & n11486;
  assign n14242 = n4976 & n11215;
  assign n14243 = n4970 & ~n10956;
  assign n14244 = ~n14242 & ~n14243;
  assign n14245 = ~n14241 & n14244;
  assign n14246 = ~n14240 & n14245;
  assign n14247 = n14246 ^ x17;
  assign n14248 = n14247 ^ n14237;
  assign n14249 = n14239 & n14248;
  assign n14250 = n14249 ^ n14247;
  assign n14252 = n14251 ^ n14250;
  assign n14253 = ~x13 & ~n12000;
  assign n14254 = ~x14 & ~n11999;
  assign n14255 = n5748 & ~n14254;
  assign n14256 = ~n14253 & n14255;
  assign n14257 = ~n13985 & n14256;
  assign n14258 = ~x11 & ~n11773;
  assign n14259 = x11 & ~x14;
  assign n14260 = n11480 & n14259;
  assign n14261 = ~n14258 & ~n14260;
  assign n14262 = x13 & ~n14261;
  assign n14263 = n5742 & n11773;
  assign n14264 = n11480 & n13989;
  assign n14265 = n5744 & ~n14264;
  assign n14266 = ~n14263 & ~n14265;
  assign n14267 = ~n11576 & n14266;
  assign n14268 = ~n14262 & ~n14267;
  assign n14269 = n14268 ^ x14;
  assign n14270 = x13 & n11999;
  assign n14271 = n14270 ^ n11875;
  assign n14272 = n5748 & n14271;
  assign n14273 = ~n14268 & n14272;
  assign n14274 = ~n14269 & n14273;
  assign n14275 = n14274 ^ n14269;
  assign n14276 = ~n14257 & n14275;
  assign n14277 = n14276 ^ n14250;
  assign n14278 = ~n14252 & n14277;
  assign n14279 = n14278 ^ n14276;
  assign n14294 = n14293 ^ n14279;
  assign n14295 = n13977 ^ n13896;
  assign n14296 = n14295 ^ n14293;
  assign n14297 = n14294 & ~n14296;
  assign n14298 = n14297 ^ n14279;
  assign n14299 = n14298 ^ n14019;
  assign n14300 = n14020 & n14299;
  assign n14301 = n14300 ^ n14298;
  assign n14304 = n14303 ^ n14301;
  assign n14305 = n14295 ^ n14294;
  assign n14627 = n5813 & n12013;
  assign n14628 = n5812 & ~n12019;
  assign n14629 = ~n14627 & n14628;
  assign n14630 = n5817 & ~n11940;
  assign n14631 = n5824 & n11902;
  assign n14632 = ~n14630 & ~n14631;
  assign n14633 = ~n14629 & n14632;
  assign n14634 = n14633 ^ x11;
  assign n14625 = n14276 ^ n14252;
  assign n14604 = n14247 ^ n14239;
  assign n14583 = n14234 ^ n14030;
  assign n14570 = n14231 ^ n14223;
  assign n14557 = n14218 ^ n14210;
  assign n14307 = n4478 & n12180;
  assign n14308 = n4487 & n10718;
  assign n14309 = n4480 & n10738;
  assign n14310 = ~n14308 & ~n14309;
  assign n14311 = n4484 & ~n10736;
  assign n14312 = n14310 & ~n14311;
  assign n14313 = ~n14307 & n14312;
  assign n14314 = n14313 ^ x23;
  assign n14306 = n14205 ^ n14204;
  assign n14315 = n14314 ^ n14306;
  assign n14329 = n14188 ^ n14181;
  assign n14324 = n14179 ^ n14039;
  assign n14325 = n14039 ^ x29;
  assign n14326 = n14325 ^ n14046;
  assign n14327 = ~n14324 & n14326;
  assign n14328 = n14327 ^ n14046;
  assign n14330 = n14329 ^ n14328;
  assign n14316 = n3285 & n12940;
  assign n14317 = n3437 & n10751;
  assign n14318 = n3435 & ~n10756;
  assign n14319 = ~n3440 & n10757;
  assign n14320 = ~n14318 & ~n14319;
  assign n14321 = ~n14317 & n14320;
  assign n14322 = ~n14316 & n14321;
  assign n14323 = n14322 ^ x26;
  assign n14331 = n14330 ^ n14323;
  assign n14340 = n14324 ^ n14047;
  assign n14332 = n3285 & ~n12703;
  assign n14333 = n3437 & ~n10756;
  assign n14334 = n3435 & n10757;
  assign n14335 = ~n3440 & n10773;
  assign n14336 = ~n14334 & ~n14335;
  assign n14337 = ~n14333 & n14336;
  assign n14338 = ~n14332 & n14337;
  assign n14339 = n14338 ^ x26;
  assign n14341 = n14340 ^ n14339;
  assign n14350 = n14176 ^ n14058;
  assign n14342 = n3285 & n12818;
  assign n14343 = n3437 & n10757;
  assign n14344 = ~n3440 & ~n10776;
  assign n14345 = ~n14343 & ~n14344;
  assign n14346 = n3435 & n10773;
  assign n14347 = n14345 & ~n14346;
  assign n14348 = ~n14342 & n14347;
  assign n14349 = n14348 ^ x26;
  assign n14351 = n14350 ^ n14349;
  assign n14353 = n3285 & n13155;
  assign n14354 = n3437 & n10773;
  assign n14355 = n3435 & ~n10776;
  assign n14356 = ~n3440 & ~n10777;
  assign n14357 = ~n14355 & ~n14356;
  assign n14358 = ~n14354 & n14357;
  assign n14359 = ~n14353 & n14358;
  assign n14360 = n14359 ^ x26;
  assign n14352 = n14173 ^ n14068;
  assign n14361 = n14360 ^ n14352;
  assign n14363 = n3285 & ~n13167;
  assign n14364 = n3437 & ~n10776;
  assign n14365 = n3435 & ~n10777;
  assign n14366 = ~n3440 & n10785;
  assign n14367 = ~n14365 & ~n14366;
  assign n14368 = ~n14364 & n14367;
  assign n14369 = ~n14363 & n14368;
  assign n14370 = n14369 ^ x26;
  assign n14362 = n14170 ^ n14078;
  assign n14371 = n14370 ^ n14362;
  assign n14373 = n3285 & ~n12832;
  assign n14374 = n3437 & ~n10777;
  assign n14375 = ~n3440 & ~n10789;
  assign n14376 = ~n14374 & ~n14375;
  assign n14377 = n3435 & n10785;
  assign n14378 = n14376 & ~n14377;
  assign n14379 = ~n14373 & n14378;
  assign n14380 = n14379 ^ x26;
  assign n14372 = n14167 ^ n14088;
  assign n14381 = n14380 ^ n14372;
  assign n14515 = n12417 & n13197;
  assign n14516 = ~n3440 & ~n10795;
  assign n14517 = n3435 & ~n10789;
  assign n14518 = ~n14516 & ~n14517;
  assign n14519 = x26 & n14518;
  assign n14520 = ~n10785 & n14519;
  assign n14521 = x25 & ~n14520;
  assign n14522 = ~n14515 & n14521;
  assign n14523 = ~n13197 & n14519;
  assign n14524 = n10785 & n12417;
  assign n14525 = ~x25 & ~n14524;
  assign n14526 = ~n14523 & n14525;
  assign n14527 = ~n14522 & ~n14526;
  assign n14528 = ~n12432 & n14518;
  assign n14529 = n14528 ^ x26;
  assign n14530 = ~n14527 & n14529;
  assign n14383 = n12417 & ~n13224;
  assign n14384 = n3435 & ~n10795;
  assign n14385 = ~n3440 & ~n10799;
  assign n14386 = ~n14384 & ~n14385;
  assign n14387 = x26 & n14386;
  assign n14388 = n10789 & n14387;
  assign n14389 = ~n14383 & ~n14388;
  assign n14390 = x25 & n14389;
  assign n14391 = n13224 & n14387;
  assign n14392 = ~n10789 & n12417;
  assign n14393 = ~x25 & ~n14392;
  assign n14394 = ~n14391 & n14393;
  assign n14395 = ~n14390 & ~n14394;
  assign n14396 = ~n12432 & n14386;
  assign n14397 = n14396 ^ x26;
  assign n14398 = ~n14395 & n14397;
  assign n14382 = n14161 ^ n14108;
  assign n14399 = n14398 ^ n14382;
  assign n14401 = n3285 & ~n13239;
  assign n14402 = n3437 & ~n10795;
  assign n14403 = n3435 & ~n10799;
  assign n14404 = ~n3440 & ~n10800;
  assign n14405 = ~n14403 & ~n14404;
  assign n14406 = ~n14402 & n14405;
  assign n14407 = ~n14401 & n14406;
  assign n14408 = n14407 ^ x26;
  assign n14400 = n14158 ^ n14150;
  assign n14409 = n14408 ^ n14400;
  assign n14488 = n12417 & ~n13278;
  assign n14489 = ~n3440 & n10815;
  assign n14490 = n3435 & ~n10800;
  assign n14491 = ~n14489 & ~n14490;
  assign n14492 = x26 & n14491;
  assign n14493 = n10799 & n14492;
  assign n14494 = x25 & ~n14493;
  assign n14495 = ~n14488 & n14494;
  assign n14496 = n13278 & n14492;
  assign n14497 = ~n10799 & n12417;
  assign n14498 = ~x25 & ~n14497;
  assign n14499 = ~n14496 & n14498;
  assign n14500 = ~n14495 & ~n14499;
  assign n14501 = ~n12432 & n14491;
  assign n14502 = n14501 ^ x26;
  assign n14503 = ~n14500 & n14502;
  assign n14418 = n3285 & ~n13341;
  assign n14419 = n3437 & ~n10800;
  assign n14420 = ~n3440 & n10819;
  assign n14421 = ~n14419 & ~n14420;
  assign n14422 = n3435 & n10815;
  assign n14423 = n14421 & ~n14422;
  assign n14424 = ~n14418 & n14423;
  assign n14425 = n14424 ^ x26;
  assign n14410 = ~n14119 & ~n14133;
  assign n14411 = n91 & n14410;
  assign n14412 = n14133 ^ n14119;
  assign n14413 = ~n54 & n10825;
  assign n14414 = ~n14412 & n14413;
  assign n14415 = ~n14411 & n14414;
  assign n14416 = ~n14134 & n14412;
  assign n14417 = ~n14415 & ~n14416;
  assign n14426 = n14425 ^ n14417;
  assign n14471 = x29 & n14131;
  assign n14472 = n14471 ^ n14127;
  assign n14437 = n3285 & n13429;
  assign n14438 = n3437 & n10819;
  assign n14439 = n3435 & ~n10820;
  assign n14440 = ~n3440 & n10821;
  assign n14441 = ~n14439 & ~n14440;
  assign n14442 = ~n14438 & n14441;
  assign n14443 = ~n14437 & n14442;
  assign n14444 = n14443 ^ x26;
  assign n14427 = x26 & n77;
  assign n14428 = ~n6177 & ~n14427;
  assign n14429 = ~n10822 & n14428;
  assign n14430 = n6476 & n10825;
  assign n14431 = ~n14429 & n14430;
  assign n14432 = n42 & n10825;
  assign n14433 = x28 & n14432;
  assign n14434 = n14433 ^ n42;
  assign n14435 = ~n10822 & n14434;
  assign n14436 = ~n14431 & ~n14435;
  assign n14445 = n14444 ^ n14436;
  assign n14446 = n3285 & ~n14111;
  assign n14447 = n3437 & ~n10820;
  assign n14448 = n3435 & n10821;
  assign n14449 = ~n3440 & ~n10822;
  assign n14450 = ~n14448 & ~n14449;
  assign n14451 = ~n14447 & n14450;
  assign n14452 = ~n14446 & n14451;
  assign n14453 = n14452 ^ x26;
  assign n14454 = n3285 & n14120;
  assign n14455 = n3437 & n10821;
  assign n14456 = n3435 & ~n10822;
  assign n14457 = ~n3440 & n10825;
  assign n14458 = ~n14456 & ~n14457;
  assign n14459 = ~n14455 & n14458;
  assign n14460 = ~n14454 & n14459;
  assign n14461 = n735 & ~n10822;
  assign n14462 = ~n6509 & n10825;
  assign n14463 = ~n14461 & ~n14462;
  assign n14464 = x26 & n14463;
  assign n14465 = n14460 & n14464;
  assign n14466 = ~n14432 & ~n14465;
  assign n14467 = ~n14453 & ~n14466;
  assign n14468 = n14467 ^ n14436;
  assign n14469 = n14445 & n14468;
  assign n14470 = n14469 ^ n14444;
  assign n14473 = n14472 ^ n14470;
  assign n14474 = n3285 & n13387;
  assign n14475 = n3437 & n10815;
  assign n14476 = n3435 & n10819;
  assign n14477 = ~n3440 & ~n10820;
  assign n14478 = ~n14476 & ~n14477;
  assign n14479 = ~n14475 & n14478;
  assign n14480 = ~n14474 & n14479;
  assign n14481 = n14480 ^ x26;
  assign n14482 = n14481 ^ n14472;
  assign n14483 = n14473 & ~n14482;
  assign n14484 = n14483 ^ n14470;
  assign n14485 = n14484 ^ n14425;
  assign n14486 = n14426 & n14485;
  assign n14487 = n14486 ^ n14484;
  assign n14504 = n14503 ^ n14487;
  assign n14505 = n14145 ^ n14137;
  assign n14506 = n14505 ^ n14503;
  assign n14507 = n14504 & n14506;
  assign n14508 = n14507 ^ n14487;
  assign n14509 = n14508 ^ n14408;
  assign n14510 = n14409 & n14509;
  assign n14511 = n14510 ^ n14508;
  assign n14512 = n14511 ^ n14398;
  assign n14513 = n14399 & n14512;
  assign n14514 = n14513 ^ n14511;
  assign n14531 = n14530 ^ n14514;
  assign n14532 = n14164 ^ n14098;
  assign n14533 = n14532 ^ n14514;
  assign n14534 = n14531 & n14533;
  assign n14535 = n14534 ^ n14530;
  assign n14536 = n14535 ^ n14380;
  assign n14537 = n14381 & n14536;
  assign n14538 = n14537 ^ n14535;
  assign n14539 = n14538 ^ n14370;
  assign n14540 = ~n14371 & n14539;
  assign n14541 = n14540 ^ n14538;
  assign n14542 = n14541 ^ n14360;
  assign n14543 = n14361 & n14542;
  assign n14544 = n14543 ^ n14541;
  assign n14545 = n14544 ^ n14350;
  assign n14546 = ~n14351 & n14545;
  assign n14547 = n14546 ^ n14544;
  assign n14548 = n14547 ^ n14340;
  assign n14549 = ~n14341 & n14548;
  assign n14550 = n14549 ^ n14547;
  assign n14551 = n14550 ^ n14330;
  assign n14552 = ~n14331 & n14551;
  assign n14553 = n14552 ^ n14550;
  assign n14554 = n14553 ^ n14306;
  assign n14555 = ~n14315 & n14554;
  assign n14556 = n14555 ^ n14314;
  assign n14558 = n14557 ^ n14556;
  assign n14559 = n4673 & n11599;
  assign n14560 = n4685 & n10694;
  assign n14561 = ~n4681 & n10698;
  assign n14562 = ~n14560 & ~n14561;
  assign n14563 = n4688 & n10683;
  assign n14564 = n14562 & ~n14563;
  assign n14565 = ~n14559 & n14564;
  assign n14566 = n14565 ^ x20;
  assign n14567 = n14566 ^ n14557;
  assign n14568 = n14558 & ~n14567;
  assign n14569 = n14568 ^ n14566;
  assign n14571 = n14570 ^ n14569;
  assign n14572 = n4963 & ~n10957;
  assign n14573 = n4976 & ~n10663;
  assign n14574 = n4972 & ~n10956;
  assign n14575 = n4970 & n10665;
  assign n14576 = ~n14574 & ~n14575;
  assign n14577 = ~n14573 & n14576;
  assign n14578 = ~n14572 & n14577;
  assign n14579 = n14578 ^ x17;
  assign n14580 = n14579 ^ n14570;
  assign n14581 = n14571 & ~n14580;
  assign n14582 = n14581 ^ n14579;
  assign n14584 = n14583 ^ n14582;
  assign n14592 = n5771 & ~n12460;
  assign n14585 = n4970 & ~n10663;
  assign n14586 = n4976 & ~n10956;
  assign n14587 = ~n14585 & ~n14586;
  assign n14588 = x17 & n14587;
  assign n14593 = ~n11215 & n14588;
  assign n14594 = ~n14592 & ~n14593;
  assign n14589 = n12460 & n14588;
  assign n14590 = n5771 & n11215;
  assign n14591 = ~n14589 & ~n14590;
  assign n14595 = n14594 ^ n14591;
  assign n14596 = ~x16 & n14595;
  assign n14597 = n14596 ^ n14594;
  assign n14598 = ~n5786 & n14587;
  assign n14599 = n14598 ^ x17;
  assign n14600 = n14597 & n14599;
  assign n14601 = n14600 ^ n14582;
  assign n14602 = n14584 & n14601;
  assign n14603 = n14602 ^ n14600;
  assign n14605 = n14604 ^ n14603;
  assign n14606 = n6033 & ~n11777;
  assign n14607 = ~n5746 & n11480;
  assign n14608 = n5752 & n11500;
  assign n14609 = ~n14607 & ~n14608;
  assign n14610 = x14 & n14609;
  assign n14611 = n11773 & n14610;
  assign n14612 = x13 & ~n14611;
  assign n14613 = ~n14606 & n14612;
  assign n14614 = n11777 & n14610;
  assign n14615 = n6033 & ~n11773;
  assign n14616 = ~x13 & ~n14615;
  assign n14617 = ~n14614 & n14616;
  assign n14618 = ~n14613 & ~n14617;
  assign n14619 = ~n7589 & n14609;
  assign n14620 = n14619 ^ x14;
  assign n14621 = ~n14618 & n14620;
  assign n14622 = n14621 ^ n14603;
  assign n14623 = n14605 & n14622;
  assign n14624 = n14623 ^ n14621;
  assign n14626 = n14625 ^ n14624;
  assign n14635 = n14634 ^ n14626;
  assign n14636 = n14635 ^ n12207;
  assign n14970 = n14621 ^ n14605;
  assign n14949 = n5749 & ~n11506;
  assign n14950 = n14949 ^ x13;
  assign n14951 = n14950 ^ n11480;
  assign n14952 = n5748 & ~n14951;
  assign n14953 = n11500 & n13989;
  assign n14954 = ~n11486 & n13719;
  assign n14955 = ~n14953 & ~n14954;
  assign n14956 = n5742 & ~n14955;
  assign n14941 = x12 & x13;
  assign n14942 = n6048 & ~n14941;
  assign n14939 = ~x12 & ~x13;
  assign n14957 = n11500 & ~n14939;
  assign n14958 = n14942 & ~n14957;
  assign n14959 = ~n14956 & ~n14958;
  assign n14933 = ~x13 & n11486;
  assign n14928 = x13 & x14;
  assign n14960 = n11500 & n14928;
  assign n14961 = ~n14933 & ~n14960;
  assign n14962 = n5744 & ~n14961;
  assign n14963 = n14959 & ~n14962;
  assign n14964 = ~n14952 & n14963;
  assign n14921 = n14579 ^ n14571;
  assign n14908 = n14566 ^ n14558;
  assign n14638 = n4673 & n12087;
  assign n14639 = n4688 & n10694;
  assign n14640 = ~n4681 & n10715;
  assign n14641 = n4685 & n10698;
  assign n14642 = ~n14640 & ~n14641;
  assign n14643 = ~n14639 & n14642;
  assign n14644 = ~n14638 & n14643;
  assign n14645 = n14644 ^ x20;
  assign n14637 = n14553 ^ n14315;
  assign n14646 = n14645 ^ n14637;
  assign n14648 = n4478 & ~n12596;
  assign n14649 = n4487 & ~n10736;
  assign n14650 = n4484 & n10738;
  assign n14651 = n4480 & n10740;
  assign n14652 = ~n14650 & ~n14651;
  assign n14653 = ~n14649 & n14652;
  assign n14654 = ~n14648 & n14653;
  assign n14655 = n14654 ^ x23;
  assign n14647 = n14550 ^ n14331;
  assign n14656 = n14655 ^ n14647;
  assign n14658 = n4478 & n12194;
  assign n14659 = n4487 & n10738;
  assign n14660 = n4484 & n10740;
  assign n14661 = n4480 & n10751;
  assign n14662 = ~n14660 & ~n14661;
  assign n14663 = ~n14659 & n14662;
  assign n14664 = ~n14658 & n14663;
  assign n14665 = n14664 ^ x23;
  assign n14657 = n14547 ^ n14341;
  assign n14666 = n14665 ^ n14657;
  assign n14668 = n4478 & n13141;
  assign n14669 = n4487 & n10740;
  assign n14670 = n4484 & n10751;
  assign n14671 = n4480 & ~n10756;
  assign n14672 = ~n14670 & ~n14671;
  assign n14673 = ~n14669 & n14672;
  assign n14674 = ~n14668 & n14673;
  assign n14675 = n14674 ^ x23;
  assign n14667 = n14544 ^ n14351;
  assign n14676 = n14675 ^ n14667;
  assign n14678 = n4478 & n12940;
  assign n14679 = n4487 & n10751;
  assign n14680 = n4484 & ~n10756;
  assign n14681 = n4480 & n10757;
  assign n14682 = ~n14680 & ~n14681;
  assign n14683 = ~n14679 & n14682;
  assign n14684 = ~n14678 & n14683;
  assign n14685 = n14684 ^ x23;
  assign n14677 = n14541 ^ n14361;
  assign n14686 = n14685 ^ n14677;
  assign n14688 = n4478 & ~n12703;
  assign n14689 = n4487 & ~n10756;
  assign n14690 = n4484 & n10757;
  assign n14691 = n4480 & n10773;
  assign n14692 = ~n14690 & ~n14691;
  assign n14693 = ~n14689 & n14692;
  assign n14694 = ~n14688 & n14693;
  assign n14695 = n14694 ^ x23;
  assign n14687 = n14538 ^ n14371;
  assign n14696 = n14695 ^ n14687;
  assign n14698 = n4478 & n12818;
  assign n14699 = n4487 & n10757;
  assign n14700 = n4480 & ~n10776;
  assign n14701 = ~n14699 & ~n14700;
  assign n14702 = n4484 & n10773;
  assign n14703 = n14701 & ~n14702;
  assign n14704 = ~n14698 & n14703;
  assign n14705 = n14704 ^ x23;
  assign n14697 = n14535 ^ n14381;
  assign n14706 = n14705 ^ n14697;
  assign n14708 = n4478 & n13155;
  assign n14709 = n4487 & n10773;
  assign n14710 = n4484 & ~n10776;
  assign n14711 = n4480 & ~n10777;
  assign n14712 = ~n14710 & ~n14711;
  assign n14713 = ~n14709 & n14712;
  assign n14714 = ~n14708 & n14713;
  assign n14715 = n14714 ^ x23;
  assign n14707 = n14532 ^ n14531;
  assign n14716 = n14715 ^ n14707;
  assign n14718 = n4478 & ~n13167;
  assign n14719 = n4487 & ~n10776;
  assign n14720 = n4484 & ~n10777;
  assign n14721 = n4480 & n10785;
  assign n14722 = ~n14720 & ~n14721;
  assign n14723 = ~n14719 & n14722;
  assign n14724 = ~n14718 & n14723;
  assign n14725 = n14724 ^ x23;
  assign n14717 = n14511 ^ n14399;
  assign n14726 = n14725 ^ n14717;
  assign n14727 = n14505 ^ n14504;
  assign n14729 = ~x22 & ~n13224;
  assign n14730 = x22 & ~n10789;
  assign n14731 = x23 & ~n14730;
  assign n14732 = ~n14729 & n14731;
  assign n14733 = ~n12518 & ~n14732;
  assign n14734 = n4484 & ~n10795;
  assign n14735 = n4480 & ~n10799;
  assign n14736 = ~n14734 & ~n14735;
  assign n14737 = ~n14733 & n14736;
  assign n14738 = x22 & n4476;
  assign n14739 = ~n13224 & n14738;
  assign n14740 = ~x22 & n4476;
  assign n14741 = ~n10789 & n14740;
  assign n14742 = n14736 & ~n14741;
  assign n14743 = ~n14739 & n14742;
  assign n14744 = ~x23 & ~n14743;
  assign n14745 = ~n14737 & ~n14744;
  assign n14728 = n14484 ^ n14426;
  assign n14746 = n14745 ^ n14728;
  assign n14828 = n12502 & ~n13239;
  assign n14829 = n4484 & ~n10799;
  assign n14830 = n4480 & ~n10800;
  assign n14831 = ~n14829 & ~n14830;
  assign n14832 = x23 & n14831;
  assign n14833 = n10795 & n14832;
  assign n14834 = x22 & ~n14833;
  assign n14835 = ~n14828 & n14834;
  assign n14836 = n13239 & n14832;
  assign n14837 = ~n10795 & n12502;
  assign n14838 = ~x22 & ~n14837;
  assign n14839 = ~n14836 & n14838;
  assign n14840 = ~n14835 & ~n14839;
  assign n14841 = ~n12519 & n14831;
  assign n14842 = n14841 ^ x23;
  assign n14843 = ~n14840 & n14842;
  assign n14748 = n4478 & ~n13278;
  assign n14749 = n4487 & ~n10799;
  assign n14750 = n4484 & ~n10800;
  assign n14751 = n4480 & n10815;
  assign n14752 = ~n14750 & ~n14751;
  assign n14753 = ~n14749 & n14752;
  assign n14754 = ~n14748 & n14753;
  assign n14755 = n14754 ^ x23;
  assign n14747 = n14467 ^ n14445;
  assign n14756 = n14755 ^ n14747;
  assign n14759 = n4478 & ~n13341;
  assign n14760 = n4487 & ~n10800;
  assign n14761 = n4480 & n10819;
  assign n14762 = ~n14760 & ~n14761;
  assign n14763 = n4484 & n10815;
  assign n14764 = n14762 & ~n14763;
  assign n14765 = ~n14759 & n14764;
  assign n14766 = n14765 ^ x23;
  assign n14757 = n14465 ^ n14432;
  assign n14758 = n14757 ^ n14453;
  assign n14767 = n14766 ^ n14758;
  assign n14808 = x26 & ~n14463;
  assign n14809 = n14808 ^ n14460;
  assign n14773 = n4478 & ~n14111;
  assign n14774 = n4487 & ~n10820;
  assign n14775 = n4484 & n10821;
  assign n14776 = n4480 & ~n10822;
  assign n14777 = ~n14775 & ~n14776;
  assign n14778 = ~n14774 & n14777;
  assign n14779 = ~n14773 & n14778;
  assign n14780 = n14779 ^ x23;
  assign n14781 = n4478 & n14120;
  assign n14782 = n4487 & n10821;
  assign n14783 = n4484 & ~n10822;
  assign n14784 = n4480 & n10825;
  assign n14785 = ~n14783 & ~n14784;
  assign n14786 = ~n14782 & n14785;
  assign n14787 = ~n14781 & n14786;
  assign n14788 = n4476 & ~n10822;
  assign n14789 = n38 & n10825;
  assign n14790 = ~n14788 & ~n14789;
  assign n14791 = x23 & n14790;
  assign n14792 = n14787 & n14791;
  assign n14793 = n735 & n10825;
  assign n14794 = ~n14792 & ~n14793;
  assign n14795 = ~n14780 & ~n14794;
  assign n14769 = n6715 & n10825;
  assign n14768 = x25 & n10825;
  assign n14770 = n14769 ^ n14768;
  assign n14771 = n14461 & ~n14770;
  assign n14772 = n14771 ^ n14769;
  assign n14796 = n14795 ^ n14772;
  assign n14797 = n4478 & n13429;
  assign n14798 = n4487 & n10819;
  assign n14799 = n4484 & ~n10820;
  assign n14800 = n4480 & n10821;
  assign n14801 = ~n14799 & ~n14800;
  assign n14802 = ~n14798 & n14801;
  assign n14803 = ~n14797 & n14802;
  assign n14804 = n14803 ^ x23;
  assign n14805 = n14804 ^ n14795;
  assign n14806 = ~n14796 & ~n14805;
  assign n14807 = n14806 ^ n14804;
  assign n14810 = n14809 ^ n14807;
  assign n14811 = n4478 & n13387;
  assign n14812 = n4487 & n10815;
  assign n14813 = n4484 & n10819;
  assign n14814 = n4480 & ~n10820;
  assign n14815 = ~n14813 & ~n14814;
  assign n14816 = ~n14812 & n14815;
  assign n14817 = ~n14811 & n14816;
  assign n14818 = n14817 ^ x23;
  assign n14819 = n14818 ^ n14807;
  assign n14820 = ~n14810 & n14819;
  assign n14821 = n14820 ^ n14818;
  assign n14822 = n14821 ^ n14758;
  assign n14823 = n14767 & ~n14822;
  assign n14824 = n14823 ^ n14766;
  assign n14825 = n14824 ^ n14755;
  assign n14826 = n14756 & n14825;
  assign n14827 = n14826 ^ n14824;
  assign n14844 = n14843 ^ n14827;
  assign n14845 = n14481 ^ n14473;
  assign n14846 = n14845 ^ n14843;
  assign n14847 = n14844 & ~n14846;
  assign n14848 = n14847 ^ n14827;
  assign n14849 = n14848 ^ n14745;
  assign n14850 = n14746 & n14849;
  assign n14851 = n14850 ^ n14848;
  assign n14852 = ~n14727 & n14851;
  assign n14853 = n4478 & n13197;
  assign n14854 = n4487 & n10785;
  assign n14855 = n4484 & ~n10789;
  assign n14856 = n4480 & ~n10795;
  assign n14857 = ~n14855 & ~n14856;
  assign n14858 = ~n14854 & n14857;
  assign n14859 = ~n14853 & n14858;
  assign n14860 = n14859 ^ x23;
  assign n14861 = n14508 ^ n14409;
  assign n14862 = n4478 & ~n12832;
  assign n14863 = n4487 & ~n10777;
  assign n14864 = n4480 & ~n10789;
  assign n14865 = ~n14863 & ~n14864;
  assign n14866 = n4484 & n10785;
  assign n14867 = n14865 & ~n14866;
  assign n14868 = ~n14862 & n14867;
  assign n14869 = n14868 ^ n14859;
  assign n14870 = ~n14861 & n14869;
  assign n14871 = ~n14860 & n14870;
  assign n14872 = n14871 ^ n14860;
  assign n14873 = ~n14852 & ~n14872;
  assign n14874 = n14727 & ~n14851;
  assign n14875 = n14874 ^ n14861;
  assign n14876 = n14868 ^ x23;
  assign n14877 = n14876 ^ n14861;
  assign n14878 = n14875 & n14877;
  assign n14879 = n14878 ^ n14874;
  assign n14880 = ~n14873 & ~n14879;
  assign n14881 = n14880 ^ n14725;
  assign n14882 = n14726 & n14881;
  assign n14883 = n14882 ^ n14880;
  assign n14884 = n14883 ^ n14715;
  assign n14885 = n14716 & n14884;
  assign n14886 = n14885 ^ n14883;
  assign n14887 = n14886 ^ n14705;
  assign n14888 = n14706 & n14887;
  assign n14889 = n14888 ^ n14886;
  assign n14890 = n14889 ^ n14695;
  assign n14891 = ~n14696 & n14890;
  assign n14892 = n14891 ^ n14889;
  assign n14893 = n14892 ^ n14685;
  assign n14894 = n14686 & n14893;
  assign n14895 = n14894 ^ n14892;
  assign n14896 = n14895 ^ n14675;
  assign n14897 = ~n14676 & n14896;
  assign n14898 = n14897 ^ n14895;
  assign n14899 = n14898 ^ n14665;
  assign n14900 = ~n14666 & n14899;
  assign n14901 = n14900 ^ n14898;
  assign n14902 = n14901 ^ n14655;
  assign n14903 = ~n14656 & n14902;
  assign n14904 = n14903 ^ n14901;
  assign n14905 = n14904 ^ n14645;
  assign n14906 = n14646 & n14905;
  assign n14907 = n14906 ^ n14904;
  assign n14909 = n14908 ^ n14907;
  assign n14910 = n4963 & ~n11694;
  assign n14911 = n4972 & ~n10663;
  assign n14912 = n4970 & n10680;
  assign n14913 = n4976 & n10665;
  assign n14914 = ~n14912 & ~n14913;
  assign n14915 = ~n14911 & n14914;
  assign n14916 = ~n14910 & n14915;
  assign n14917 = n14916 ^ x17;
  assign n14918 = n14917 ^ n14907;
  assign n14919 = n14909 & n14918;
  assign n14920 = n14919 ^ n14917;
  assign n14922 = n14921 ^ n14920;
  assign n14923 = n5749 & ~n11956;
  assign n14924 = n14923 ^ x13;
  assign n14925 = n14924 ^ n11500;
  assign n14926 = n5748 & ~n14925;
  assign n14927 = ~x13 & n11215;
  assign n14929 = n11486 & n14928;
  assign n14930 = ~n14927 & ~n14929;
  assign n14931 = ~x12 & ~n14930;
  assign n14932 = x13 & ~n11215;
  assign n14934 = ~n14932 & ~n14933;
  assign n14935 = x12 & n5749;
  assign n14936 = ~n14934 & n14935;
  assign n14937 = ~n14931 & ~n14936;
  assign n14938 = ~n5748 & ~n14937;
  assign n14940 = n11486 & ~n14939;
  assign n14943 = ~n14940 & n14942;
  assign n14944 = ~n14938 & ~n14943;
  assign n14945 = ~n14926 & n14944;
  assign n14946 = n14945 ^ n14921;
  assign n14947 = n14922 & n14946;
  assign n14948 = n14947 ^ n14945;
  assign n14965 = n14964 ^ n14948;
  assign n14966 = n14600 ^ n14584;
  assign n14967 = n14966 ^ n14964;
  assign n14968 = n14965 & ~n14967;
  assign n14969 = n14968 ^ n14948;
  assign n14971 = n14970 ^ n14969;
  assign n14972 = n7536 & ~n11941;
  assign n14973 = n5817 & n11902;
  assign n14974 = n5824 & ~n11875;
  assign n14975 = ~n14973 & ~n14974;
  assign n14976 = x11 & n14975;
  assign n14977 = n11940 & n14976;
  assign n14978 = x10 & ~n14977;
  assign n14979 = ~n14972 & n14978;
  assign n14980 = n11941 & n14976;
  assign n14981 = n7536 & ~n11940;
  assign n14982 = ~x10 & ~n14981;
  assign n14983 = ~n14980 & n14982;
  assign n14984 = ~n14979 & ~n14983;
  assign n14985 = ~n7551 & n14975;
  assign n14986 = n14985 ^ x11;
  assign n14987 = ~n14984 & n14986;
  assign n14988 = n14987 ^ n14969;
  assign n14989 = ~n14971 & ~n14988;
  assign n14990 = n14989 ^ n14987;
  assign n14991 = n14990 ^ n12207;
  assign n14992 = ~n14636 & n14991;
  assign n14993 = n14992 ^ n14635;
  assign n14994 = ~n14305 & ~n14993;
  assign n15371 = n14990 ^ n14636;
  assign n15360 = n6314 & ~n14014;
  assign n15361 = n6311 & n6316;
  assign n15362 = n12019 & n15361;
  assign n15363 = x8 & n6315;
  assign n15364 = ~n15362 & ~n15363;
  assign n15365 = ~n15360 & n15364;
  assign n15347 = n5814 & n12504;
  assign n15348 = n6295 & n11902;
  assign n15349 = n5817 & ~n11875;
  assign n15350 = n5824 & ~n11773;
  assign n15351 = ~n15349 & ~n15350;
  assign n15352 = ~n15348 & n15351;
  assign n15353 = ~n15347 & n15352;
  assign n15354 = n15353 ^ x11;
  assign n15334 = n14945 ^ n14922;
  assign n15315 = n14917 ^ n14909;
  assign n14996 = n4963 & n12100;
  assign n14997 = n4976 & n10680;
  assign n14998 = n4970 & n10683;
  assign n14999 = ~n14997 & ~n14998;
  assign n15000 = n4972 & n10665;
  assign n15001 = n14999 & ~n15000;
  assign n15002 = ~n14996 & n15001;
  assign n15003 = n15002 ^ x17;
  assign n14995 = n14904 ^ n14646;
  assign n15004 = n15003 ^ n14995;
  assign n15013 = n14901 ^ n14656;
  assign n15005 = n4673 & n12034;
  assign n15006 = n4685 & n10715;
  assign n15007 = n4688 & n10698;
  assign n15008 = ~n4681 & n10718;
  assign n15009 = ~n15007 & ~n15008;
  assign n15010 = ~n15006 & n15009;
  assign n15011 = ~n15005 & n15010;
  assign n15012 = n15011 ^ x20;
  assign n15014 = n15013 ^ n15012;
  assign n15016 = n4673 & n12111;
  assign n15017 = n4688 & n10715;
  assign n15018 = ~n4681 & ~n10736;
  assign n15019 = n4685 & n10718;
  assign n15020 = ~n15018 & ~n15019;
  assign n15021 = ~n15017 & n15020;
  assign n15022 = ~n15016 & n15021;
  assign n15023 = n15022 ^ x20;
  assign n15015 = n14898 ^ n14666;
  assign n15024 = n15023 ^ n15015;
  assign n15026 = n4673 & n12180;
  assign n15027 = n4685 & ~n10736;
  assign n15028 = n4688 & n10718;
  assign n15029 = ~n15027 & ~n15028;
  assign n15030 = ~n4681 & n10738;
  assign n15031 = n15029 & ~n15030;
  assign n15032 = ~n15026 & n15031;
  assign n15033 = n15032 ^ x20;
  assign n15025 = n14895 ^ n14676;
  assign n15034 = n15033 ^ n15025;
  assign n15043 = n14892 ^ n14686;
  assign n15035 = n4673 & ~n12596;
  assign n15036 = n4688 & ~n10736;
  assign n15037 = n4685 & n10738;
  assign n15038 = ~n4681 & n10740;
  assign n15039 = ~n15037 & ~n15038;
  assign n15040 = ~n15036 & n15039;
  assign n15041 = ~n15035 & n15040;
  assign n15042 = n15041 ^ x20;
  assign n15044 = n15043 ^ n15042;
  assign n15046 = n4673 & n12194;
  assign n15047 = n4688 & n10738;
  assign n15048 = n4685 & n10740;
  assign n15049 = ~n4681 & n10751;
  assign n15050 = ~n15048 & ~n15049;
  assign n15051 = ~n15047 & n15050;
  assign n15052 = ~n15046 & n15051;
  assign n15053 = n15052 ^ x20;
  assign n15045 = n14889 ^ n14696;
  assign n15054 = n15053 ^ n15045;
  assign n15055 = n4673 & n13141;
  assign n15056 = n4688 & n10740;
  assign n15057 = n4685 & n10751;
  assign n15058 = ~n4681 & ~n10756;
  assign n15059 = ~n15057 & ~n15058;
  assign n15060 = ~n15056 & n15059;
  assign n15061 = ~n15055 & n15060;
  assign n15062 = n14886 ^ n14706;
  assign n15063 = ~n15061 & n15062;
  assign n15271 = n4673 & n12940;
  assign n15272 = n4688 & n10751;
  assign n15273 = n4685 & ~n10756;
  assign n15274 = ~n4681 & n10757;
  assign n15275 = ~n15273 & ~n15274;
  assign n15276 = ~n15272 & n15275;
  assign n15277 = ~n15271 & n15276;
  assign n15065 = n4673 & ~n12703;
  assign n15066 = n4688 & ~n10756;
  assign n15067 = n4685 & n10757;
  assign n15068 = ~n4681 & n10773;
  assign n15069 = ~n15067 & ~n15068;
  assign n15070 = ~n15066 & n15069;
  assign n15071 = ~n15065 & n15070;
  assign n15072 = n15071 ^ x20;
  assign n15064 = n14880 ^ n14726;
  assign n15073 = n15072 ^ n15064;
  assign n15081 = n4673 & n12818;
  assign n15082 = n4688 & n10757;
  assign n15083 = ~n4681 & ~n10776;
  assign n15084 = ~n15082 & ~n15083;
  assign n15085 = n4685 & n10773;
  assign n15086 = n15084 & ~n15085;
  assign n15087 = ~n15081 & n15086;
  assign n15088 = n15087 ^ x20;
  assign n15079 = n14868 ^ n14861;
  assign n15074 = n14851 ^ n14727;
  assign n15075 = n14727 ^ x23;
  assign n15076 = n15075 ^ n14859;
  assign n15077 = n15074 & ~n15076;
  assign n15078 = n15077 ^ n14859;
  assign n15080 = n15079 ^ n15078;
  assign n15089 = n15088 ^ n15080;
  assign n15091 = n4673 & n13155;
  assign n15092 = n4688 & n10773;
  assign n15093 = n4685 & ~n10776;
  assign n15094 = ~n4681 & ~n10777;
  assign n15095 = ~n15093 & ~n15094;
  assign n15096 = ~n15092 & n15095;
  assign n15097 = ~n15091 & n15096;
  assign n15098 = n15097 ^ x20;
  assign n15090 = n15074 ^ n14860;
  assign n15099 = n15098 ^ n15090;
  assign n15101 = n4673 & ~n13167;
  assign n15102 = n4688 & ~n10776;
  assign n15103 = n4685 & ~n10777;
  assign n15104 = ~n4681 & n10785;
  assign n15105 = ~n15103 & ~n15104;
  assign n15106 = ~n15102 & n15105;
  assign n15107 = ~n15101 & n15106;
  assign n15108 = n15107 ^ x20;
  assign n15100 = n14848 ^ n14746;
  assign n15109 = n15108 ^ n15100;
  assign n15111 = n4673 & ~n12832;
  assign n15112 = n4688 & ~n10777;
  assign n15113 = ~n4681 & ~n10789;
  assign n15114 = ~n15112 & ~n15113;
  assign n15115 = n4685 & n10785;
  assign n15116 = n15114 & ~n15115;
  assign n15117 = ~n15111 & n15116;
  assign n15118 = n15117 ^ x20;
  assign n15110 = n14845 ^ n14844;
  assign n15119 = n15118 ^ n15110;
  assign n15121 = n13197 & n13653;
  assign n15122 = ~n4681 & ~n10795;
  assign n15123 = n4685 & ~n10789;
  assign n15124 = ~n15122 & ~n15123;
  assign n15125 = x20 & n15124;
  assign n15126 = ~n10785 & n15125;
  assign n15127 = x19 & ~n15126;
  assign n15128 = ~n15121 & n15127;
  assign n15129 = ~n13197 & n15125;
  assign n15130 = n10785 & n13653;
  assign n15131 = ~x19 & ~n15130;
  assign n15132 = ~n15129 & n15131;
  assign n15133 = ~n15128 & ~n15132;
  assign n15134 = ~n13668 & n15124;
  assign n15135 = n15134 ^ x20;
  assign n15136 = ~n15133 & n15135;
  assign n15120 = n14824 ^ n14756;
  assign n15137 = n15136 ^ n15120;
  assign n15139 = n4673 & ~n13224;
  assign n15140 = n4688 & ~n10789;
  assign n15141 = ~n4681 & ~n10799;
  assign n15142 = ~n15140 & ~n15141;
  assign n15143 = n4685 & ~n10795;
  assign n15144 = n15142 & ~n15143;
  assign n15145 = ~n15139 & n15144;
  assign n15146 = n15145 ^ x20;
  assign n15138 = n14821 ^ n14767;
  assign n15147 = n15146 ^ n15138;
  assign n15149 = n4673 & ~n13239;
  assign n15150 = n4688 & ~n10795;
  assign n15151 = n4685 & ~n10799;
  assign n15152 = ~n4681 & ~n10800;
  assign n15153 = ~n15151 & ~n15152;
  assign n15154 = ~n15150 & n15153;
  assign n15155 = ~n15149 & n15154;
  assign n15156 = n15155 ^ x20;
  assign n15148 = n14818 ^ n14810;
  assign n15157 = n15156 ^ n15148;
  assign n15159 = n4673 & ~n13278;
  assign n15160 = n4688 & ~n10799;
  assign n15161 = n4685 & ~n10800;
  assign n15162 = ~n4681 & n10815;
  assign n15163 = ~n15161 & ~n15162;
  assign n15164 = ~n15160 & n15163;
  assign n15165 = ~n15159 & n15164;
  assign n15166 = n15165 ^ x20;
  assign n15158 = n14804 ^ n14796;
  assign n15167 = n15166 ^ n15158;
  assign n15170 = n4673 & ~n13341;
  assign n15171 = n4688 & ~n10800;
  assign n15172 = ~n4681 & n10819;
  assign n15173 = ~n15171 & ~n15172;
  assign n15174 = n4685 & n10815;
  assign n15175 = n15173 & ~n15174;
  assign n15176 = ~n15170 & n15175;
  assign n15177 = n15176 ^ x20;
  assign n15168 = n14793 ^ n14792;
  assign n15169 = n15168 ^ n14780;
  assign n15178 = n15177 ^ n15169;
  assign n15219 = x23 & ~n14790;
  assign n15220 = n15219 ^ n14787;
  assign n15184 = n4673 & ~n14111;
  assign n15185 = n4688 & ~n10820;
  assign n15186 = n4685 & n10821;
  assign n15187 = ~n4681 & ~n10822;
  assign n15188 = ~n15186 & ~n15187;
  assign n15189 = ~n15185 & n15188;
  assign n15190 = ~n15184 & n15189;
  assign n15191 = n15190 ^ x20;
  assign n15192 = n4673 & n14120;
  assign n15193 = n4688 & n10821;
  assign n15194 = n4685 & ~n10822;
  assign n15195 = ~n4681 & n10825;
  assign n15196 = ~n15194 & ~n15195;
  assign n15197 = ~n15193 & n15196;
  assign n15198 = ~n15192 & n15197;
  assign n15199 = n4671 & ~n10822;
  assign n15200 = ~n7059 & n10825;
  assign n15201 = ~n15199 & ~n15200;
  assign n15202 = x20 & n15201;
  assign n15203 = n15198 & n15202;
  assign n15204 = n4476 & n10825;
  assign n15205 = ~n15203 & ~n15204;
  assign n15206 = ~n15191 & ~n15205;
  assign n15180 = x22 & n10825;
  assign n15179 = n7030 & n10825;
  assign n15181 = n15180 ^ n15179;
  assign n15182 = ~n14788 & ~n15181;
  assign n15183 = n15182 ^ n15180;
  assign n15207 = n15206 ^ n15183;
  assign n15208 = n4673 & n13429;
  assign n15209 = n4688 & n10819;
  assign n15210 = n4685 & ~n10820;
  assign n15211 = ~n4681 & n10821;
  assign n15212 = ~n15210 & ~n15211;
  assign n15213 = ~n15209 & n15212;
  assign n15214 = ~n15208 & n15213;
  assign n15215 = n15214 ^ x20;
  assign n15216 = n15215 ^ n15206;
  assign n15217 = n15207 & ~n15216;
  assign n15218 = n15217 ^ n15215;
  assign n15221 = n15220 ^ n15218;
  assign n15222 = ~x19 & ~n13387;
  assign n15223 = x19 & ~n10815;
  assign n15224 = n4671 & ~n15223;
  assign n15225 = ~n15222 & n15224;
  assign n15226 = n4685 & n10819;
  assign n15227 = ~n4681 & ~n10820;
  assign n15228 = ~n15226 & ~n15227;
  assign n15229 = x20 & n15228;
  assign n15230 = ~n15225 & n15229;
  assign n15231 = x19 & ~n13387;
  assign n15232 = ~x19 & ~n10815;
  assign n15233 = n13653 & ~n15232;
  assign n15234 = ~n15231 & n15233;
  assign n15235 = ~x20 & ~n15228;
  assign n15236 = ~n15234 & ~n15235;
  assign n15237 = ~n15230 & n15236;
  assign n15238 = n15237 ^ n15218;
  assign n15239 = n15221 & ~n15238;
  assign n15240 = n15239 ^ n15220;
  assign n15241 = n15240 ^ n15177;
  assign n15242 = ~n15178 & n15241;
  assign n15243 = n15242 ^ n15240;
  assign n15244 = n15243 ^ n15166;
  assign n15245 = ~n15167 & n15244;
  assign n15246 = n15245 ^ n15243;
  assign n15247 = n15246 ^ n15156;
  assign n15248 = ~n15157 & n15247;
  assign n15249 = n15248 ^ n15246;
  assign n15250 = n15249 ^ n15146;
  assign n15251 = ~n15147 & n15250;
  assign n15252 = n15251 ^ n15249;
  assign n15253 = n15252 ^ n15136;
  assign n15254 = n15137 & n15253;
  assign n15255 = n15254 ^ n15252;
  assign n15256 = n15255 ^ n15118;
  assign n15257 = ~n15119 & n15256;
  assign n15258 = n15257 ^ n15255;
  assign n15259 = n15258 ^ n15108;
  assign n15260 = n15109 & n15259;
  assign n15261 = n15260 ^ n15258;
  assign n15262 = n15261 ^ n15098;
  assign n15263 = n15099 & n15262;
  assign n15264 = n15263 ^ n15261;
  assign n15265 = n15264 ^ n15088;
  assign n15266 = n15089 & n15265;
  assign n15267 = n15266 ^ n15264;
  assign n15268 = n15267 ^ n15072;
  assign n15269 = n15073 & n15268;
  assign n15270 = n15269 ^ n15267;
  assign n15278 = n15277 ^ n15270;
  assign n15279 = n14883 ^ n14716;
  assign n15280 = n15279 ^ n15277;
  assign n15281 = n15278 & n15280;
  assign n15282 = n15281 ^ n15270;
  assign n15283 = ~n15063 & n15282;
  assign n15284 = n15061 & ~n15062;
  assign n15285 = ~x20 & ~n15284;
  assign n15286 = ~n15283 & n15285;
  assign n15287 = n15277 & n15279;
  assign n15288 = n15270 & ~n15287;
  assign n15289 = ~n15277 & ~n15279;
  assign n15290 = ~n15288 & ~n15289;
  assign n15291 = n15061 & n15062;
  assign n15292 = ~n15290 & ~n15291;
  assign n15293 = ~n15061 & ~n15062;
  assign n15294 = x20 & ~n15293;
  assign n15295 = ~n15292 & n15294;
  assign n15296 = ~n15286 & ~n15295;
  assign n15297 = n15296 ^ n15053;
  assign n15298 = ~n15054 & n15297;
  assign n15299 = n15298 ^ n15296;
  assign n15300 = n15299 ^ n15043;
  assign n15301 = n15044 & ~n15300;
  assign n15302 = n15301 ^ n15299;
  assign n15303 = n15302 ^ n15033;
  assign n15304 = ~n15034 & n15303;
  assign n15305 = n15304 ^ n15302;
  assign n15306 = n15305 ^ n15023;
  assign n15307 = ~n15024 & n15306;
  assign n15308 = n15307 ^ n15305;
  assign n15309 = n15308 ^ n15013;
  assign n15310 = ~n15014 & n15309;
  assign n15311 = n15310 ^ n15308;
  assign n15312 = n15311 ^ n15003;
  assign n15313 = n15004 & n15312;
  assign n15314 = n15313 ^ n15311;
  assign n15316 = n15315 ^ n15314;
  assign n15317 = x13 & n11703;
  assign n15318 = n15317 ^ n11486;
  assign n15319 = n6033 & n15318;
  assign n15320 = ~n11704 & n13989;
  assign n15321 = ~n5746 & n11215;
  assign n15322 = n5752 & ~n10956;
  assign n15323 = ~n15321 & ~n15322;
  assign n15324 = ~n7559 & n15323;
  assign n15325 = ~n11486 & n14928;
  assign n15326 = n15324 & ~n15325;
  assign n15327 = ~n15320 & n15326;
  assign n15328 = x14 & ~n15323;
  assign n15329 = ~n15327 & ~n15328;
  assign n15330 = ~n15319 & ~n15329;
  assign n15331 = n15330 ^ n15314;
  assign n15332 = n15316 & n15331;
  assign n15333 = n15332 ^ n15330;
  assign n15335 = n15334 ^ n15333;
  assign n15336 = n5814 & ~n12000;
  assign n15337 = n6295 & ~n11875;
  assign n15338 = n5817 & ~n11773;
  assign n15339 = n5824 & n11480;
  assign n15340 = ~n15338 & ~n15339;
  assign n15341 = ~n15337 & n15340;
  assign n15342 = ~n15336 & n15341;
  assign n15343 = n15342 ^ x11;
  assign n15344 = n15343 ^ n15334;
  assign n15345 = ~n15335 & n15344;
  assign n15346 = n15345 ^ n15343;
  assign n15355 = n15354 ^ n15346;
  assign n15356 = n14966 ^ n14965;
  assign n15357 = n15356 ^ n15354;
  assign n15358 = n15355 & n15357;
  assign n15359 = n15358 ^ n15346;
  assign n15366 = n15365 ^ n15359;
  assign n15367 = n14987 ^ n14971;
  assign n15368 = n15367 ^ n15359;
  assign n15369 = n15366 & n15368;
  assign n15370 = n15369 ^ n15367;
  assign n15372 = n15371 ^ n15370;
  assign n17384 = n7515 & n17383;
  assign n17385 = n7520 & ~n11940;
  assign n17386 = n7518 & ~n12019;
  assign n17387 = ~n8029 & ~n17386;
  assign n17388 = ~n17385 & n17387;
  assign n17389 = ~n17384 & n17388;
  assign n17390 = n17389 ^ x5;
  assign n16805 = ~x8 & n6305;
  assign n17364 = n12504 & n16805;
  assign n17365 = n6309 & ~n11875;
  assign n17366 = n6316 & ~n11773;
  assign n17367 = ~n17365 & ~n17366;
  assign n17368 = x8 & n17367;
  assign n17369 = ~n11902 & n17368;
  assign n17370 = ~n17364 & ~n17369;
  assign n17371 = x7 & n17370;
  assign n17372 = ~n12504 & n17368;
  assign n17373 = n11902 & n16805;
  assign n17374 = ~x7 & ~n17373;
  assign n17375 = ~n17372 & n17374;
  assign n17376 = ~n17371 & ~n17375;
  assign n16819 = x8 & ~n6305;
  assign n16820 = n16819 ^ x8;
  assign n17377 = ~n16820 & n17367;
  assign n17378 = n17377 ^ x8;
  assign n17379 = ~n17376 & n17378;
  assign n17346 = n7536 & n11507;
  assign n17347 = n5817 & n11500;
  assign n17348 = n5824 & n11486;
  assign n17349 = ~n17347 & ~n17348;
  assign n17350 = x11 & n17349;
  assign n17351 = ~n11480 & n17350;
  assign n17352 = x10 & ~n17351;
  assign n17353 = ~n17346 & n17352;
  assign n17354 = ~n11507 & n17350;
  assign n17355 = n7536 & n11480;
  assign n17356 = ~x10 & ~n17355;
  assign n17357 = ~n17354 & n17356;
  assign n17358 = ~n17353 & ~n17357;
  assign n17359 = ~n7551 & n17349;
  assign n17360 = n17359 ^ x11;
  assign n17361 = ~n17358 & n17360;
  assign n17332 = n12460 ^ n11215;
  assign n17333 = x13 & ~n17332;
  assign n17334 = n17333 ^ n11215;
  assign n17335 = n6033 & n17334;
  assign n17336 = ~x13 & n12460;
  assign n17337 = n7860 & ~n14932;
  assign n17338 = ~n17336 & n17337;
  assign n17339 = n5752 & ~n10663;
  assign n17340 = ~n5746 & ~n10956;
  assign n17341 = ~n17339 & ~n17340;
  assign n17342 = n17341 ^ x14;
  assign n17343 = ~n17338 & ~n17342;
  assign n17344 = ~n17335 & ~n17343;
  assign n17330 = n15311 ^ n15004;
  assign n16760 = n15308 ^ n15014;
  assign n16752 = n4963 & n12524;
  assign n16753 = n4972 & n10680;
  assign n16754 = n4976 & n10683;
  assign n16755 = n4970 & n10694;
  assign n16756 = ~n16754 & ~n16755;
  assign n16757 = ~n16753 & n16756;
  assign n16758 = ~n16752 & n16757;
  assign n16759 = n16758 ^ x17;
  assign n16761 = n16760 ^ n16759;
  assign n16284 = n15305 ^ n15024;
  assign n16276 = n4963 & n11599;
  assign n16277 = n4976 & n10694;
  assign n16278 = n4970 & n10698;
  assign n16279 = ~n16277 & ~n16278;
  assign n16280 = n4972 & n10683;
  assign n16281 = n16279 & ~n16280;
  assign n16282 = ~n16276 & n16281;
  assign n16283 = n16282 ^ x17;
  assign n16285 = n16284 ^ n16283;
  assign n15719 = n15302 ^ n15034;
  assign n15711 = n4963 & n12087;
  assign n15712 = n4972 & n10694;
  assign n15713 = n4970 & n10715;
  assign n15714 = n4976 & n10698;
  assign n15715 = ~n15713 & ~n15714;
  assign n15716 = ~n15712 & n15715;
  assign n15717 = ~n15711 & n15716;
  assign n15718 = n15717 ^ x17;
  assign n15720 = n15719 ^ n15718;
  assign n15390 = n5771 & n12034;
  assign n15391 = n4976 & n10715;
  assign n15392 = n4970 & n10718;
  assign n15393 = ~n15391 & ~n15392;
  assign n15394 = x17 & n15393;
  assign n15395 = ~n10698 & n15394;
  assign n15396 = ~n15390 & ~n15395;
  assign n15397 = x16 & n15396;
  assign n15398 = ~n12034 & n15394;
  assign n15399 = n5771 & n10698;
  assign n15400 = ~x16 & ~n15399;
  assign n15401 = ~n15398 & n15400;
  assign n15402 = ~n15397 & ~n15401;
  assign n15403 = ~n5786 & n15393;
  assign n15404 = n15403 ^ x17;
  assign n15405 = ~n15402 & n15404;
  assign n15389 = n15299 ^ n15044;
  assign n15406 = n15405 ^ n15389;
  assign n15408 = n4963 & n12111;
  assign n15409 = n4972 & n10715;
  assign n15410 = n4970 & ~n10736;
  assign n15411 = n4976 & n10718;
  assign n15412 = ~n15410 & ~n15411;
  assign n15413 = ~n15409 & n15412;
  assign n15414 = ~n15408 & n15413;
  assign n15415 = n15414 ^ x17;
  assign n15407 = n15296 ^ n15054;
  assign n15416 = n15415 ^ n15407;
  assign n15424 = n4963 & n12180;
  assign n15425 = n4976 & ~n10736;
  assign n15426 = n4972 & n10718;
  assign n15427 = ~n15425 & ~n15426;
  assign n15428 = n4970 & n10738;
  assign n15429 = n15427 & ~n15428;
  assign n15430 = ~n15424 & n15429;
  assign n15431 = n15430 ^ x17;
  assign n15422 = n15062 ^ n15061;
  assign n15417 = n15277 ^ x20;
  assign n15418 = n15417 ^ n15279;
  assign n15419 = n15279 ^ n15270;
  assign n15420 = ~n15418 & n15419;
  assign n15421 = n15420 ^ n15277;
  assign n15423 = n15422 ^ n15421;
  assign n15432 = n15431 ^ n15423;
  assign n15436 = n4963 & ~n12596;
  assign n15437 = n4972 & ~n10736;
  assign n15438 = n4976 & n10738;
  assign n15439 = n4970 & n10740;
  assign n15440 = ~n15438 & ~n15439;
  assign n15441 = ~n15437 & n15440;
  assign n15442 = ~n15436 & n15441;
  assign n15443 = n15442 ^ x17;
  assign n15433 = n15279 ^ x20;
  assign n15434 = n15433 ^ n15277;
  assign n15435 = n15434 ^ n15270;
  assign n15444 = n15443 ^ n15435;
  assign n15446 = n4963 & n12194;
  assign n15447 = n4972 & n10738;
  assign n15448 = n4976 & n10740;
  assign n15449 = n4970 & n10751;
  assign n15450 = ~n15448 & ~n15449;
  assign n15451 = ~n15447 & n15450;
  assign n15452 = ~n15446 & n15451;
  assign n15453 = n15452 ^ x17;
  assign n15445 = n15267 ^ n15073;
  assign n15454 = n15453 ^ n15445;
  assign n15456 = n4963 & n13141;
  assign n15457 = n4972 & n10740;
  assign n15458 = n4976 & n10751;
  assign n15459 = n4970 & ~n10756;
  assign n15460 = ~n15458 & ~n15459;
  assign n15461 = ~n15457 & n15460;
  assign n15462 = ~n15456 & n15461;
  assign n15463 = n15462 ^ x17;
  assign n15455 = n15264 ^ n15089;
  assign n15464 = n15463 ^ n15455;
  assign n15466 = n4963 & n12940;
  assign n15467 = n4972 & n10751;
  assign n15468 = n4976 & ~n10756;
  assign n15469 = n4970 & n10757;
  assign n15470 = ~n15468 & ~n15469;
  assign n15471 = ~n15467 & n15470;
  assign n15472 = ~n15466 & n15471;
  assign n15473 = n15472 ^ x17;
  assign n15465 = n15261 ^ n15099;
  assign n15474 = n15473 ^ n15465;
  assign n15476 = n4963 & ~n12703;
  assign n15477 = n4972 & ~n10756;
  assign n15478 = n4976 & n10757;
  assign n15479 = n4970 & n10773;
  assign n15480 = ~n15478 & ~n15479;
  assign n15481 = ~n15477 & n15480;
  assign n15482 = ~n15476 & n15481;
  assign n15483 = n15482 ^ x17;
  assign n15475 = n15258 ^ n15109;
  assign n15484 = n15483 ^ n15475;
  assign n15486 = n4963 & n12818;
  assign n15487 = n4972 & n10757;
  assign n15488 = n4970 & ~n10776;
  assign n15489 = ~n15487 & ~n15488;
  assign n15490 = n4976 & n10773;
  assign n15491 = n15489 & ~n15490;
  assign n15492 = ~n15486 & n15491;
  assign n15493 = n15492 ^ x17;
  assign n15485 = n15255 ^ n15119;
  assign n15494 = n15493 ^ n15485;
  assign n15496 = ~x16 & n13155;
  assign n15497 = x16 & n10773;
  assign n15498 = x17 & ~n15497;
  assign n15499 = ~n15496 & n15498;
  assign n15500 = ~n5785 & ~n15499;
  assign n15501 = n4976 & ~n10776;
  assign n15502 = n4970 & ~n10777;
  assign n15503 = ~n15501 & ~n15502;
  assign n15504 = ~n15500 & n15503;
  assign n15505 = x16 & ~n13155;
  assign n15506 = ~x16 & ~n10773;
  assign n15507 = n5771 & ~n15506;
  assign n15508 = ~n15505 & n15507;
  assign n15509 = ~x17 & ~n15503;
  assign n15510 = ~n15508 & ~n15509;
  assign n15511 = ~n15504 & n15510;
  assign n15495 = n15252 ^ n15137;
  assign n15512 = n15511 ^ n15495;
  assign n15661 = n15249 ^ n15147;
  assign n15514 = n4963 & ~n12832;
  assign n15515 = n4972 & ~n10777;
  assign n15516 = n4970 & ~n10789;
  assign n15517 = ~n15515 & ~n15516;
  assign n15518 = n4976 & n10785;
  assign n15519 = n15517 & ~n15518;
  assign n15520 = ~n15514 & n15519;
  assign n15521 = n15520 ^ x17;
  assign n15513 = n15246 ^ n15157;
  assign n15522 = n15521 ^ n15513;
  assign n15524 = n4963 & n13197;
  assign n15525 = n4972 & n10785;
  assign n15526 = n4976 & ~n10789;
  assign n15527 = n4970 & ~n10795;
  assign n15528 = ~n15526 & ~n15527;
  assign n15529 = ~n15525 & n15528;
  assign n15530 = ~n15524 & n15529;
  assign n15531 = n15530 ^ x17;
  assign n15523 = n15243 ^ n15167;
  assign n15532 = n15531 ^ n15523;
  assign n15534 = n4963 & ~n13224;
  assign n15535 = n4972 & ~n10789;
  assign n15536 = n4970 & ~n10799;
  assign n15537 = ~n15535 & ~n15536;
  assign n15538 = n4976 & ~n10795;
  assign n15539 = n15537 & ~n15538;
  assign n15540 = ~n15534 & n15539;
  assign n15541 = n15540 ^ x17;
  assign n15533 = n15240 ^ n15178;
  assign n15542 = n15541 ^ n15533;
  assign n15550 = n5771 & ~n13239;
  assign n15551 = n4976 & ~n10799;
  assign n15552 = n4970 & ~n10800;
  assign n15553 = ~n15551 & ~n15552;
  assign n15554 = x17 & n15553;
  assign n15555 = n10795 & n15554;
  assign n15556 = x16 & ~n15555;
  assign n15557 = ~n15550 & n15556;
  assign n15558 = n13239 & n15554;
  assign n15559 = n5771 & ~n10795;
  assign n15560 = ~x16 & ~n15559;
  assign n15561 = ~n15558 & n15560;
  assign n15562 = ~n15557 & ~n15561;
  assign n15563 = ~n5786 & n15553;
  assign n15564 = n15563 ^ x17;
  assign n15565 = ~n15562 & n15564;
  assign n15544 = n4673 & n13387;
  assign n15545 = n4688 & n10815;
  assign n15546 = n15228 & ~n15545;
  assign n15547 = ~n15544 & n15546;
  assign n15543 = n15220 ^ x20;
  assign n15548 = n15547 ^ n15543;
  assign n15549 = n15548 ^ n15218;
  assign n15566 = n15565 ^ n15549;
  assign n15568 = n4963 & ~n13278;
  assign n15569 = n4972 & ~n10799;
  assign n15570 = n4976 & ~n10800;
  assign n15571 = n4970 & n10815;
  assign n15572 = ~n15570 & ~n15571;
  assign n15573 = ~n15569 & n15572;
  assign n15574 = ~n15568 & n15573;
  assign n15575 = n15574 ^ x17;
  assign n15567 = n15215 ^ n15207;
  assign n15576 = n15575 ^ n15567;
  assign n15579 = n4963 & ~n13341;
  assign n15580 = n4972 & ~n10800;
  assign n15581 = n4970 & n10819;
  assign n15582 = ~n15580 & ~n15581;
  assign n15583 = n4976 & n10815;
  assign n15584 = n15582 & ~n15583;
  assign n15585 = ~n15579 & n15584;
  assign n15586 = n15585 ^ x17;
  assign n15577 = n15204 ^ n15203;
  assign n15578 = n15577 ^ n15191;
  assign n15587 = n15586 ^ n15578;
  assign n15590 = n4963 & n13387;
  assign n15591 = n4972 & n10815;
  assign n15592 = n4976 & n10819;
  assign n15593 = n4970 & ~n10820;
  assign n15594 = ~n15592 & ~n15593;
  assign n15595 = ~n15591 & n15594;
  assign n15596 = ~n15590 & n15595;
  assign n15597 = n15596 ^ x17;
  assign n15588 = x20 & ~n15201;
  assign n15589 = n15588 ^ n15198;
  assign n15598 = n15597 ^ n15589;
  assign n15622 = x19 & n4671;
  assign n15623 = n13498 & n15622;
  assign n15624 = n4678 ^ x19;
  assign n15625 = n10825 & n15624;
  assign n15626 = ~n15199 & ~n15625;
  assign n15627 = ~n15623 & ~n15626;
  assign n15599 = n4963 & ~n14111;
  assign n15600 = n4972 & ~n10820;
  assign n15601 = n4976 & n10821;
  assign n15602 = n4970 & ~n10822;
  assign n15603 = ~n15601 & ~n15602;
  assign n15604 = ~n15600 & n15603;
  assign n15605 = ~n15599 & n15604;
  assign n15608 = n4963 & n14120;
  assign n15609 = n4972 & n10821;
  assign n15610 = n4970 & n10825;
  assign n15611 = ~n15609 & ~n15610;
  assign n15612 = ~n15608 & n15611;
  assign n15613 = x17 & n15612;
  assign n15614 = n4969 & ~n14128;
  assign n15615 = n15613 & ~n15614;
  assign n15616 = ~x18 & n10825;
  assign n15617 = x17 & n15616;
  assign n15618 = ~n15615 & ~n15617;
  assign n15606 = ~x17 & x18;
  assign n15607 = n10825 & n15606;
  assign n15619 = n15618 ^ n15607;
  assign n15620 = ~n15605 & ~n15619;
  assign n15621 = n15620 ^ n15618;
  assign n15628 = n15627 ^ n15621;
  assign n15629 = n4963 & n13429;
  assign n15630 = n4972 & n10819;
  assign n15631 = n4976 & ~n10820;
  assign n15632 = n4970 & n10821;
  assign n15633 = ~n15631 & ~n15632;
  assign n15634 = ~n15630 & n15633;
  assign n15635 = ~n15629 & n15634;
  assign n15636 = n15635 ^ x17;
  assign n15637 = n15636 ^ n15621;
  assign n15638 = n15628 & n15637;
  assign n15639 = n15638 ^ n15636;
  assign n15640 = n15639 ^ n15589;
  assign n15641 = n15598 & ~n15640;
  assign n15642 = n15641 ^ n15597;
  assign n15643 = n15642 ^ n15586;
  assign n15644 = ~n15587 & n15643;
  assign n15645 = n15644 ^ n15642;
  assign n15646 = n15645 ^ n15575;
  assign n15647 = n15576 & n15646;
  assign n15648 = n15647 ^ n15645;
  assign n15649 = n15648 ^ n15565;
  assign n15650 = ~n15566 & n15649;
  assign n15651 = n15650 ^ n15648;
  assign n15652 = n15651 ^ n15541;
  assign n15653 = ~n15542 & n15652;
  assign n15654 = n15653 ^ n15651;
  assign n15655 = n15654 ^ n15531;
  assign n15656 = ~n15532 & n15655;
  assign n15657 = n15656 ^ n15654;
  assign n15658 = n15657 ^ n15521;
  assign n15659 = ~n15522 & n15658;
  assign n15660 = n15659 ^ n15657;
  assign n15662 = n15661 ^ n15660;
  assign n15663 = n4970 & n10785;
  assign n15664 = n4976 & ~n10777;
  assign n15665 = ~n15663 & ~n15664;
  assign n15667 = ~n5771 & ~n10776;
  assign n15668 = ~n13166 & ~n15667;
  assign n15669 = ~x17 & n10776;
  assign n15670 = n15668 & ~n15669;
  assign n15671 = n10776 ^ x16;
  assign n15672 = n13166 & ~n15671;
  assign n15673 = ~n15670 & ~n15672;
  assign n15666 = n15665 ^ x17;
  assign n15674 = n15673 ^ n15666;
  assign n15675 = n15665 & n15674;
  assign n15676 = n4961 & n15675;
  assign n15677 = n15676 ^ n15666;
  assign n15678 = n15677 ^ n15661;
  assign n15679 = n15662 & ~n15678;
  assign n15680 = n15679 ^ n15660;
  assign n15681 = n15680 ^ n15495;
  assign n15682 = ~n15512 & n15681;
  assign n15683 = n15682 ^ n15511;
  assign n15684 = n15683 ^ n15493;
  assign n15685 = ~n15494 & n15684;
  assign n15686 = n15685 ^ n15683;
  assign n15687 = n15686 ^ n15483;
  assign n15688 = n15484 & n15687;
  assign n15689 = n15688 ^ n15686;
  assign n15690 = n15689 ^ n15473;
  assign n15691 = n15474 & n15690;
  assign n15692 = n15691 ^ n15689;
  assign n15693 = n15692 ^ n15463;
  assign n15694 = n15464 & n15693;
  assign n15695 = n15694 ^ n15692;
  assign n15696 = n15695 ^ n15453;
  assign n15697 = n15454 & n15696;
  assign n15698 = n15697 ^ n15695;
  assign n15699 = n15698 ^ n15443;
  assign n15700 = n15444 & n15699;
  assign n15701 = n15700 ^ n15698;
  assign n15702 = n15701 ^ n15431;
  assign n15703 = n15432 & n15702;
  assign n15704 = n15703 ^ n15701;
  assign n15705 = n15704 ^ n15415;
  assign n15706 = ~n15416 & n15705;
  assign n15707 = n15706 ^ n15704;
  assign n15708 = n15707 ^ n15405;
  assign n15709 = n15406 & n15708;
  assign n15710 = n15709 ^ n15707;
  assign n16273 = n15719 ^ n15710;
  assign n16274 = ~n15720 & n16273;
  assign n16275 = n16274 ^ n15710;
  assign n16749 = n16284 ^ n16275;
  assign n16750 = ~n16285 & n16749;
  assign n16751 = n16750 ^ n16275;
  assign n17327 = n16760 ^ n16751;
  assign n17328 = ~n16761 & n17327;
  assign n17329 = n17328 ^ n16751;
  assign n17331 = n17330 ^ n17329;
  assign n17345 = n17344 ^ n17331;
  assign n17362 = n17361 ^ n17345;
  assign n16763 = n6033 & ~n10957;
  assign n16764 = ~n5746 & ~n10663;
  assign n16765 = n5752 & n10665;
  assign n16766 = ~n16764 & ~n16765;
  assign n16767 = x14 & n16766;
  assign n16768 = n10956 & n16767;
  assign n16769 = ~n16763 & ~n16768;
  assign n16770 = x13 & n16769;
  assign n16771 = n10957 & n16767;
  assign n16772 = n6033 & ~n10956;
  assign n16773 = ~x13 & ~n16772;
  assign n16774 = ~n16771 & n16773;
  assign n16775 = ~n16770 & ~n16774;
  assign n16776 = ~n7589 & n16766;
  assign n16777 = n16776 ^ x14;
  assign n16778 = ~n16775 & n16777;
  assign n16762 = n16761 ^ n16751;
  assign n16779 = n16778 ^ n16762;
  assign n16287 = n6033 & ~n11694;
  assign n16288 = ~n5746 & n10665;
  assign n16289 = n5752 & n10680;
  assign n16290 = ~n16288 & ~n16289;
  assign n16291 = x14 & n16290;
  assign n16292 = n10663 & n16291;
  assign n16293 = x13 & ~n16292;
  assign n16294 = ~n16287 & n16293;
  assign n16295 = n11694 & n16291;
  assign n16296 = n6033 & ~n10663;
  assign n16297 = ~x13 & ~n16296;
  assign n16298 = ~n16295 & n16297;
  assign n16299 = ~n16294 & ~n16298;
  assign n16300 = ~n7589 & n16290;
  assign n16301 = n16300 ^ x14;
  assign n16302 = ~n16299 & n16301;
  assign n16286 = n16285 ^ n16275;
  assign n16303 = n16302 ^ n16286;
  assign n15722 = ~n10665 & ~n12099;
  assign n15723 = n6033 & ~n15722;
  assign n15724 = ~n5746 & n10680;
  assign n15725 = n5752 & n10683;
  assign n15726 = ~n15724 & ~n15725;
  assign n15727 = x14 & n15726;
  assign n15728 = ~n15723 & ~n15727;
  assign n15729 = ~x13 & n12099;
  assign n15730 = n15729 ^ n10665;
  assign n15731 = n6033 & ~n12099;
  assign n15732 = ~n15729 & n15731;
  assign n15733 = n15730 & n15732;
  assign n15734 = n15733 ^ n15730;
  assign n15735 = ~n15728 & ~n15734;
  assign n15736 = ~n7589 & n15726;
  assign n15737 = n15736 ^ x14;
  assign n15738 = ~n15735 & n15737;
  assign n15721 = n15720 ^ n15710;
  assign n15739 = n15738 ^ n15721;
  assign n15741 = n5752 & n10694;
  assign n15742 = ~n5746 & n10683;
  assign n15743 = ~n15741 & ~n15742;
  assign n15744 = x14 & n15743;
  assign n15745 = n15744 ^ x13;
  assign n15746 = ~n11616 & n15745;
  assign n15747 = n15746 ^ x13;
  assign n15748 = ~n10680 & n15747;
  assign n15749 = n5748 & ~n15748;
  assign n15750 = x13 & n11616;
  assign n11626 = n10680 & ~n11616;
  assign n15751 = ~n6033 & n11626;
  assign n15752 = n15751 ^ n10680;
  assign n15753 = ~n15750 & n15752;
  assign n15754 = n15749 & ~n15753;
  assign n15755 = ~n6048 & n15743;
  assign n15756 = ~n15754 & n15755;
  assign n15757 = ~x14 & ~n15743;
  assign n15758 = ~n15756 & ~n15757;
  assign n15740 = n15707 ^ n15406;
  assign n15759 = n15758 ^ n15740;
  assign n15761 = n6033 & n11599;
  assign n15762 = ~n5746 & n10694;
  assign n15763 = n5752 & n10698;
  assign n15764 = ~n15762 & ~n15763;
  assign n15765 = x14 & n15764;
  assign n15766 = ~n10683 & n15765;
  assign n15767 = ~n15761 & ~n15766;
  assign n15768 = x13 & n15767;
  assign n15769 = ~n11599 & n15765;
  assign n15770 = n6033 & n10683;
  assign n15771 = ~x13 & ~n15770;
  assign n15772 = ~n15769 & n15771;
  assign n15773 = ~n15768 & ~n15772;
  assign n15774 = ~n7589 & n15764;
  assign n15775 = n15774 ^ x14;
  assign n15776 = ~n15773 & n15775;
  assign n15760 = n15704 ^ n15416;
  assign n15777 = n15776 ^ n15760;
  assign n15779 = n6033 & n12087;
  assign n15780 = n5752 & n10715;
  assign n15781 = ~n5746 & n10698;
  assign n15782 = ~n15780 & ~n15781;
  assign n15783 = x14 & n15782;
  assign n15784 = ~n10694 & n15783;
  assign n15785 = x13 & ~n15784;
  assign n15786 = ~n15779 & n15785;
  assign n15787 = ~n12087 & n15783;
  assign n15788 = n6033 & n10694;
  assign n15789 = ~x13 & ~n15788;
  assign n15790 = ~n15787 & n15789;
  assign n15791 = ~n15786 & ~n15790;
  assign n15792 = ~n7589 & n15782;
  assign n15793 = n15792 ^ x14;
  assign n15794 = ~n15791 & n15793;
  assign n15778 = n15701 ^ n15432;
  assign n15795 = n15794 ^ n15778;
  assign n15797 = n6033 & n12034;
  assign n15798 = ~n5746 & n10715;
  assign n15799 = n5752 & n10718;
  assign n15800 = ~n15798 & ~n15799;
  assign n15801 = x14 & n15800;
  assign n15802 = ~n10698 & n15801;
  assign n15803 = ~n15797 & ~n15802;
  assign n15804 = x13 & n15803;
  assign n15805 = ~n12034 & n15801;
  assign n15806 = n6033 & n10698;
  assign n15807 = ~x13 & ~n15806;
  assign n15808 = ~n15805 & n15807;
  assign n15809 = ~n15804 & ~n15808;
  assign n15810 = ~n7589 & n15800;
  assign n15811 = n15810 ^ x14;
  assign n15812 = ~n15809 & n15811;
  assign n15796 = n15698 ^ n15444;
  assign n15813 = n15812 ^ n15796;
  assign n15815 = n6033 & n12111;
  assign n15816 = n5752 & ~n10736;
  assign n15817 = ~n5746 & n10718;
  assign n15818 = ~n15816 & ~n15817;
  assign n15819 = x14 & n15818;
  assign n15820 = ~n10715 & n15819;
  assign n15821 = x13 & ~n15820;
  assign n15822 = ~n15815 & n15821;
  assign n15823 = ~n12111 & n15819;
  assign n15824 = n6033 & n10715;
  assign n15825 = ~x13 & ~n15824;
  assign n15826 = ~n15823 & n15825;
  assign n15827 = ~n15822 & ~n15826;
  assign n15828 = ~n7589 & n15818;
  assign n15829 = n15828 ^ x14;
  assign n15830 = ~n15827 & n15829;
  assign n15814 = n15695 ^ n15454;
  assign n15831 = n15830 ^ n15814;
  assign n15833 = n6033 & n12180;
  assign n15834 = ~n5746 & ~n10736;
  assign n15835 = n5752 & n10738;
  assign n15836 = ~n15834 & ~n15835;
  assign n15837 = x14 & n15836;
  assign n15838 = ~n10718 & n15837;
  assign n15839 = ~n15833 & ~n15838;
  assign n15840 = x13 & n15839;
  assign n15841 = ~n12180 & n15837;
  assign n15842 = n6033 & n10718;
  assign n15843 = ~x13 & ~n15842;
  assign n15844 = ~n15841 & n15843;
  assign n15845 = ~n15840 & ~n15844;
  assign n15846 = ~n7589 & n15836;
  assign n15847 = n15846 ^ x14;
  assign n15848 = ~n15845 & n15847;
  assign n15832 = n15692 ^ n15464;
  assign n15849 = n15848 ^ n15832;
  assign n15851 = n6033 & ~n12596;
  assign n15852 = ~n5746 & n10738;
  assign n15853 = n5752 & n10740;
  assign n15854 = ~n15852 & ~n15853;
  assign n15855 = x14 & n15854;
  assign n15856 = n10736 & n15855;
  assign n15857 = x13 & ~n15856;
  assign n15858 = ~n15851 & n15857;
  assign n15859 = n12596 & n15855;
  assign n15860 = n6033 & ~n10736;
  assign n15861 = ~x13 & ~n15860;
  assign n15862 = ~n15859 & n15861;
  assign n15863 = ~n15858 & ~n15862;
  assign n15864 = ~n7589 & n15854;
  assign n15865 = n15864 ^ x14;
  assign n15866 = ~n15863 & n15865;
  assign n15850 = n15689 ^ n15474;
  assign n15867 = n15866 ^ n15850;
  assign n15869 = n6033 & n12194;
  assign n15870 = ~n5746 & n10740;
  assign n15871 = n5752 & n10751;
  assign n15872 = ~n15870 & ~n15871;
  assign n15873 = x14 & n15872;
  assign n15874 = ~n10738 & n15873;
  assign n15875 = x13 & ~n15874;
  assign n15876 = ~n15869 & n15875;
  assign n15877 = ~n12194 & n15873;
  assign n15878 = n6033 & n10738;
  assign n15879 = ~x13 & ~n15878;
  assign n15880 = ~n15877 & n15879;
  assign n15881 = ~n15876 & ~n15880;
  assign n15882 = ~n7589 & n15872;
  assign n15883 = n15882 ^ x14;
  assign n15884 = ~n15881 & n15883;
  assign n15868 = n15686 ^ n15484;
  assign n15885 = n15884 ^ n15868;
  assign n15888 = ~n5746 & n10751;
  assign n15889 = n5752 & ~n10756;
  assign n15890 = ~n15888 & ~n15889;
  assign n15891 = x14 & n15890;
  assign n15895 = ~n6033 & ~n15891;
  assign n15896 = ~n6034 & ~n13140;
  assign n15897 = n15896 ^ x13;
  assign n15898 = ~n15895 & ~n15897;
  assign n15887 = ~x13 & n13140;
  assign n15892 = n6033 & n13140;
  assign n15893 = ~n15891 & ~n15892;
  assign n15894 = ~n15887 & ~n15893;
  assign n15899 = n15898 ^ n15894;
  assign n15900 = ~n10740 & n15899;
  assign n15901 = n15900 ^ n15898;
  assign n15902 = ~n7589 & n15890;
  assign n15903 = n15902 ^ x14;
  assign n15904 = ~n15901 & n15903;
  assign n15886 = n15683 ^ n15494;
  assign n15905 = n15904 ^ n15886;
  assign n15907 = n6033 & n12940;
  assign n15908 = ~n5746 & ~n10756;
  assign n15909 = n5752 & n10757;
  assign n15910 = ~n15908 & ~n15909;
  assign n15911 = x14 & n15910;
  assign n15912 = ~n10751 & n15911;
  assign n15913 = x13 & ~n15912;
  assign n15914 = ~n15907 & n15913;
  assign n15915 = ~n12940 & n15911;
  assign n15916 = n6033 & n10751;
  assign n15917 = ~x13 & ~n15916;
  assign n15918 = ~n15915 & n15917;
  assign n15919 = ~n15914 & ~n15918;
  assign n15920 = ~n7589 & n15910;
  assign n15921 = n15920 ^ x14;
  assign n15922 = ~n15919 & n15921;
  assign n15906 = n15680 ^ n15512;
  assign n15923 = n15922 ^ n15906;
  assign n15925 = n6033 & ~n12703;
  assign n15926 = n5752 & n10773;
  assign n15927 = ~n5746 & n10757;
  assign n15928 = ~n15926 & ~n15927;
  assign n15929 = x14 & n15928;
  assign n15930 = n10756 & n15929;
  assign n15931 = x13 & ~n15930;
  assign n15932 = ~n15925 & n15931;
  assign n15933 = n12703 & n15929;
  assign n15934 = n6033 & ~n10756;
  assign n15935 = ~x13 & ~n15934;
  assign n15936 = ~n15933 & n15935;
  assign n15937 = ~n15932 & ~n15936;
  assign n15938 = ~n7589 & n15928;
  assign n15939 = n15938 ^ x14;
  assign n15940 = ~n15937 & n15939;
  assign n15924 = n15677 ^ n15662;
  assign n15941 = n15940 ^ n15924;
  assign n15943 = ~n10757 & ~n12817;
  assign n15944 = x13 & ~n10757;
  assign n15945 = ~n15943 & ~n15944;
  assign n15946 = n6033 & ~n12817;
  assign n15947 = n15945 & ~n15946;
  assign n15948 = n10757 & n12817;
  assign n15949 = ~x13 & n15948;
  assign n15950 = n15947 & ~n15949;
  assign n15951 = n5748 & ~n15943;
  assign n15952 = ~x14 & ~n15951;
  assign n15953 = ~n15950 & ~n15952;
  assign n15954 = ~n5746 & n10773;
  assign n15955 = n5752 & ~n10776;
  assign n15956 = ~n15954 & ~n15955;
  assign n15957 = ~n7559 & n15956;
  assign n15958 = ~n15953 & n15957;
  assign n15959 = x14 & ~n15956;
  assign n15960 = ~n15958 & ~n15959;
  assign n15942 = n15657 ^ n15522;
  assign n15961 = n15960 ^ n15942;
  assign n15963 = ~n13155 & n13989;
  assign n15964 = ~n10773 & n14928;
  assign n15965 = ~n7559 & ~n15964;
  assign n15966 = ~n15963 & n15965;
  assign n15967 = ~n5746 & ~n10776;
  assign n15968 = n5752 & ~n10777;
  assign n15969 = ~n15967 & ~n15968;
  assign n15970 = ~n15966 & n15969;
  assign n15971 = x13 & ~n13155;
  assign n15972 = ~x13 & ~n10773;
  assign n15973 = n6033 & ~n15972;
  assign n15974 = ~n15971 & n15973;
  assign n15975 = ~x14 & ~n15969;
  assign n15976 = ~n15974 & ~n15975;
  assign n15977 = ~n15970 & n15976;
  assign n15962 = n15654 ^ n15532;
  assign n15978 = n15977 ^ n15962;
  assign n15980 = x14 & ~n13166;
  assign n15981 = n5752 & n10785;
  assign n15982 = ~n5746 & ~n10777;
  assign n15983 = ~n15981 & ~n15982;
  assign n15984 = n15980 & n15983;
  assign n15985 = x13 & n13166;
  assign n15986 = ~n15984 & ~n15985;
  assign n15987 = n10776 & ~n15986;
  assign n15988 = ~n10776 & ~n15985;
  assign n15989 = ~n15980 & n15988;
  assign n15990 = n5748 & ~n15989;
  assign n15991 = ~n15987 & n15990;
  assign n15992 = ~n6048 & n15983;
  assign n15993 = ~n15991 & n15992;
  assign n15994 = ~x14 & ~n15983;
  assign n15995 = ~n15993 & ~n15994;
  assign n15979 = n15651 ^ n15542;
  assign n15996 = n15995 ^ n15979;
  assign n15998 = n6033 & ~n12832;
  assign n15999 = ~n5746 & n10785;
  assign n16000 = n5752 & ~n10789;
  assign n16001 = ~n15999 & ~n16000;
  assign n16002 = x14 & n16001;
  assign n16003 = n10777 & n16002;
  assign n16004 = ~n15998 & ~n16003;
  assign n16005 = x13 & n16004;
  assign n16006 = n12832 & n16002;
  assign n16007 = n6033 & ~n10777;
  assign n16008 = ~x13 & ~n16007;
  assign n16009 = ~n16006 & n16008;
  assign n16010 = ~n16005 & ~n16009;
  assign n16011 = ~n7589 & n16001;
  assign n16012 = n16011 ^ x14;
  assign n16013 = ~n16010 & n16012;
  assign n15997 = n15648 ^ n15566;
  assign n16014 = n16013 ^ n15997;
  assign n16204 = n6033 & n13197;
  assign n16205 = n5752 & ~n10795;
  assign n16206 = ~n5746 & ~n10789;
  assign n16207 = ~n16205 & ~n16206;
  assign n16208 = x14 & n16207;
  assign n16209 = ~n10785 & n16208;
  assign n16210 = x13 & ~n16209;
  assign n16211 = ~n16204 & n16210;
  assign n16212 = ~n13197 & n16208;
  assign n16213 = n6033 & n10785;
  assign n16214 = ~x13 & ~n16213;
  assign n16215 = ~n16212 & n16214;
  assign n16216 = ~n16211 & ~n16215;
  assign n16217 = ~n7589 & n16207;
  assign n16218 = n16217 ^ x14;
  assign n16219 = ~n16216 & n16218;
  assign n16016 = n6033 & ~n13224;
  assign n16017 = ~n5746 & ~n10795;
  assign n16018 = n5752 & ~n10799;
  assign n16019 = ~n16017 & ~n16018;
  assign n16020 = x14 & n16019;
  assign n16021 = n10789 & n16020;
  assign n16022 = ~n16016 & ~n16021;
  assign n16023 = x13 & n16022;
  assign n16024 = n13224 & n16020;
  assign n16025 = n6033 & ~n10789;
  assign n16026 = ~x13 & ~n16025;
  assign n16027 = ~n16024 & n16026;
  assign n16028 = ~n16023 & ~n16027;
  assign n16029 = ~n7589 & n16019;
  assign n16030 = n16029 ^ x14;
  assign n16031 = ~n16028 & n16030;
  assign n16015 = n15642 ^ n15587;
  assign n16032 = n16031 ^ n16015;
  assign n16034 = n6033 & ~n13239;
  assign n16035 = ~n5746 & ~n10799;
  assign n16036 = n5752 & ~n10800;
  assign n16037 = ~n16035 & ~n16036;
  assign n16038 = x14 & n16037;
  assign n16039 = n10795 & n16038;
  assign n16040 = x13 & ~n16039;
  assign n16041 = ~n16034 & n16040;
  assign n16042 = n13239 & n16038;
  assign n16043 = n6033 & ~n10795;
  assign n16044 = ~x13 & ~n16043;
  assign n16045 = ~n16042 & n16044;
  assign n16046 = ~n16041 & ~n16045;
  assign n16047 = ~n7589 & n16037;
  assign n16048 = n16047 ^ x14;
  assign n16049 = ~n16046 & n16048;
  assign n16033 = n15639 ^ n15598;
  assign n16050 = n16049 ^ n16033;
  assign n16052 = n6033 & ~n13278;
  assign n16053 = n5752 & n10815;
  assign n16054 = ~n5746 & ~n10800;
  assign n16055 = ~n16053 & ~n16054;
  assign n16056 = x14 & n16055;
  assign n16057 = n10799 & n16056;
  assign n16058 = x13 & ~n16057;
  assign n16059 = ~n16052 & n16058;
  assign n16060 = n13278 & n16056;
  assign n16061 = n6033 & ~n10799;
  assign n16062 = ~x13 & ~n16061;
  assign n16063 = ~n16060 & n16062;
  assign n16064 = ~n16059 & ~n16063;
  assign n16065 = ~n7589 & n16055;
  assign n16066 = n16065 ^ x14;
  assign n16067 = ~n16064 & n16066;
  assign n16051 = n15636 ^ n15628;
  assign n16068 = n16067 ^ n16051;
  assign n16073 = n10800 & ~n13340;
  assign n16074 = n6033 & ~n16073;
  assign n16075 = ~n5746 & n10815;
  assign n16076 = n5752 & n10819;
  assign n16077 = ~n16075 & ~n16076;
  assign n16078 = x14 & n16077;
  assign n16079 = ~n16074 & ~n16078;
  assign n16080 = ~x13 & n13340;
  assign n16081 = n16080 ^ n10800;
  assign n16082 = n6033 & ~n13340;
  assign n16083 = ~n16080 & n16082;
  assign n16084 = ~n16081 & n16083;
  assign n16085 = n16084 ^ n16081;
  assign n16086 = ~n16079 & n16085;
  assign n16087 = ~n7589 & n16077;
  assign n16088 = n16087 ^ x14;
  assign n16089 = ~n16086 & n16088;
  assign n16069 = n4671 & n10825;
  assign n16070 = n16069 ^ x17;
  assign n16071 = n16070 ^ n15615;
  assign n16072 = n16071 ^ n15605;
  assign n16090 = n16089 ^ n16072;
  assign n16157 = n6033 & n13387;
  assign n16158 = ~n5746 & n10819;
  assign n16159 = n5752 & ~n10820;
  assign n16160 = ~n16158 & ~n16159;
  assign n16161 = x14 & n16160;
  assign n16162 = ~n10815 & n16161;
  assign n16163 = x13 & ~n16162;
  assign n16164 = ~n16157 & n16163;
  assign n16165 = ~n13387 & n16161;
  assign n16166 = n6033 & n10815;
  assign n16167 = ~x13 & ~n16166;
  assign n16168 = ~n16165 & n16167;
  assign n16169 = ~n16164 & ~n16168;
  assign n16170 = ~n7589 & n16160;
  assign n16171 = n16170 ^ x14;
  assign n16172 = ~n16169 & n16171;
  assign n16098 = n6033 & n13429;
  assign n16099 = ~n5746 & ~n10820;
  assign n16100 = n5752 & n10821;
  assign n16101 = ~n16099 & ~n16100;
  assign n16102 = x14 & n16101;
  assign n16103 = ~n10819 & n16102;
  assign n16104 = ~n16098 & ~n16103;
  assign n16105 = x13 & n16104;
  assign n16106 = ~n13429 & n16102;
  assign n16107 = n6033 & n10819;
  assign n16108 = ~x13 & ~n16107;
  assign n16109 = ~n16106 & n16108;
  assign n16110 = ~n16105 & ~n16109;
  assign n16111 = ~n7589 & n16101;
  assign n16112 = n16111 ^ x14;
  assign n16113 = ~n16110 & n16112;
  assign n16091 = n4961 & ~n10822;
  assign n16094 = x16 & n10825;
  assign n16092 = n4967 ^ x16;
  assign n16093 = n10825 & n16092;
  assign n16095 = n16094 ^ n16093;
  assign n16096 = ~n16091 & ~n16095;
  assign n16097 = n16096 ^ n16094;
  assign n16114 = n16113 ^ n16097;
  assign n16115 = ~n6034 & ~n14110;
  assign n16116 = n16115 ^ x13;
  assign n16117 = ~n10820 & ~n16116;
  assign n16118 = n5748 & ~n16117;
  assign n16119 = x13 & n14110;
  assign n16120 = x14 & ~n14110;
  assign n16121 = ~n16119 & ~n16120;
  assign n16122 = n10820 & ~n16121;
  assign n16123 = n16118 & ~n16122;
  assign n16124 = ~n5746 & n10821;
  assign n16125 = n5752 & ~n10822;
  assign n16126 = ~n16124 & ~n16125;
  assign n16127 = ~n6048 & n16126;
  assign n16128 = ~n16123 & n16127;
  assign n16129 = ~x14 & ~n16126;
  assign n16130 = ~n16128 & ~n16129;
  assign n16131 = ~n10821 & ~n13532;
  assign n16132 = n6033 & ~n16131;
  assign n16133 = n10821 & ~n13532;
  assign n16134 = ~n5746 & ~n10822;
  assign n16135 = n5752 & n10825;
  assign n16136 = ~n16134 & ~n16135;
  assign n16137 = x14 & n16136;
  assign n16138 = ~n16133 & n16137;
  assign n16139 = ~n16132 & ~n16138;
  assign n16140 = n10821 ^ x13;
  assign n16141 = n13532 & ~n16140;
  assign n16142 = ~n16139 & ~n16141;
  assign n16143 = ~n7589 & n16136;
  assign n16144 = n16143 ^ x14;
  assign n16145 = ~n16142 & n16144;
  assign n16146 = ~n5746 & n10825;
  assign n16147 = ~n5748 & ~n16146;
  assign n16148 = ~n14128 & ~n16147;
  assign n16149 = x14 & ~n16148;
  assign n16150 = ~n16145 & n16149;
  assign n16151 = n4961 & n10825;
  assign n16152 = ~n16150 & ~n16151;
  assign n16153 = ~n16130 & ~n16152;
  assign n16154 = n16153 ^ n16097;
  assign n16155 = n16114 & n16154;
  assign n16156 = n16155 ^ n16113;
  assign n16173 = n16172 ^ n16156;
  assign n16174 = n10822 & n10825;
  assign n16175 = n15613 & n16174;
  assign n16176 = n4976 & ~n13532;
  assign n16177 = ~n16175 & n16176;
  assign n16178 = x17 & ~n14128;
  assign n16179 = n4961 & n16178;
  assign n16180 = n15612 & n16179;
  assign n16181 = ~n4976 & ~n15610;
  assign n16182 = ~n16180 & n16181;
  assign n16183 = ~n16177 & ~n16182;
  assign n16184 = ~n15612 & ~n16178;
  assign n16185 = ~x17 & n4976;
  assign n16186 = ~n10822 & n16185;
  assign n16187 = ~n16184 & ~n16186;
  assign n16188 = ~n16183 & n16187;
  assign n16189 = n16188 ^ n16172;
  assign n16190 = n16173 & ~n16189;
  assign n16191 = n16190 ^ n16156;
  assign n16192 = n16191 ^ n16072;
  assign n16193 = n16090 & ~n16192;
  assign n16194 = n16193 ^ n16089;
  assign n16195 = n16194 ^ n16067;
  assign n16196 = n16068 & n16195;
  assign n16197 = n16196 ^ n16194;
  assign n16198 = n16197 ^ n16049;
  assign n16199 = ~n16050 & n16198;
  assign n16200 = n16199 ^ n16197;
  assign n16201 = n16200 ^ n16031;
  assign n16202 = ~n16032 & n16201;
  assign n16203 = n16202 ^ n16200;
  assign n16220 = n16219 ^ n16203;
  assign n16221 = n15645 ^ n15576;
  assign n16222 = n16221 ^ n16219;
  assign n16223 = n16220 & n16222;
  assign n16224 = n16223 ^ n16203;
  assign n16225 = n16224 ^ n16013;
  assign n16226 = ~n16014 & n16225;
  assign n16227 = n16226 ^ n16224;
  assign n16228 = n16227 ^ n15995;
  assign n16229 = ~n15996 & n16228;
  assign n16230 = n16229 ^ n16227;
  assign n16231 = n16230 ^ n15977;
  assign n16232 = ~n15978 & n16231;
  assign n16233 = n16232 ^ n16230;
  assign n16234 = n16233 ^ n15942;
  assign n16235 = ~n15961 & ~n16234;
  assign n16236 = n16235 ^ n15960;
  assign n16237 = n16236 ^ n15940;
  assign n16238 = ~n15941 & ~n16237;
  assign n16239 = n16238 ^ n16236;
  assign n16240 = n16239 ^ n15922;
  assign n16241 = n15923 & ~n16240;
  assign n16242 = n16241 ^ n16239;
  assign n16243 = n16242 ^ n15904;
  assign n16244 = ~n15905 & ~n16243;
  assign n16245 = n16244 ^ n16242;
  assign n16246 = n16245 ^ n15884;
  assign n16247 = n15885 & ~n16246;
  assign n16248 = n16247 ^ n16245;
  assign n16249 = n16248 ^ n15866;
  assign n16250 = n15867 & ~n16249;
  assign n16251 = n16250 ^ n16248;
  assign n16252 = n16251 ^ n15848;
  assign n16253 = n15849 & ~n16252;
  assign n16254 = n16253 ^ n16251;
  assign n16255 = n16254 ^ n15830;
  assign n16256 = n15831 & ~n16255;
  assign n16257 = n16256 ^ n16254;
  assign n16258 = n16257 ^ n15812;
  assign n16259 = n15813 & ~n16258;
  assign n16260 = n16259 ^ n16257;
  assign n16261 = n16260 ^ n15794;
  assign n16262 = n15795 & ~n16261;
  assign n16263 = n16262 ^ n16260;
  assign n16264 = n16263 ^ n15776;
  assign n16265 = ~n15777 & ~n16264;
  assign n16266 = n16265 ^ n16263;
  assign n16267 = n16266 ^ n15758;
  assign n16268 = n15759 & ~n16267;
  assign n16269 = n16268 ^ n16266;
  assign n16270 = n16269 ^ n15738;
  assign n16271 = ~n15739 & ~n16270;
  assign n16272 = n16271 ^ n16269;
  assign n16746 = n16302 ^ n16272;
  assign n16747 = ~n16303 & ~n16746;
  assign n16748 = n16747 ^ n16272;
  assign n17324 = n16778 ^ n16748;
  assign n17325 = ~n16779 & ~n17324;
  assign n17326 = n17325 ^ n16748;
  assign n17363 = n17362 ^ n17326;
  assign n17380 = n17379 ^ n17363;
  assign n16780 = n16779 ^ n16748;
  assign n16738 = n5814 & n11957;
  assign n16739 = n6295 & n11500;
  assign n16740 = n5817 & n11486;
  assign n16741 = n5824 & n11215;
  assign n16742 = ~n16740 & ~n16741;
  assign n16743 = ~n16739 & n16742;
  assign n16744 = ~n16738 & n16743;
  assign n16745 = n16744 ^ x11;
  assign n16781 = n16780 ^ n16745;
  assign n16304 = n16303 ^ n16272;
  assign n15381 = n5814 & n11704;
  assign n15382 = n6295 & n11486;
  assign n15383 = n5817 & n11215;
  assign n15384 = n5824 & ~n10956;
  assign n15385 = ~n15383 & ~n15384;
  assign n15386 = ~n15382 & n15385;
  assign n15387 = ~n15381 & n15386;
  assign n15388 = n15387 ^ x11;
  assign n16305 = n16304 ^ n15388;
  assign n16314 = n16269 ^ n15739;
  assign n16306 = n5814 & ~n12460;
  assign n16307 = n6295 & n11215;
  assign n16308 = n5824 & ~n10663;
  assign n16309 = n5817 & ~n10956;
  assign n16310 = ~n16308 & ~n16309;
  assign n16311 = ~n16307 & n16310;
  assign n16312 = ~n16306 & n16311;
  assign n16313 = n16312 ^ x11;
  assign n16315 = n16314 ^ n16313;
  assign n16317 = n7536 & ~n10957;
  assign n16318 = n5817 & ~n10663;
  assign n16319 = n5824 & n10665;
  assign n16320 = ~n16318 & ~n16319;
  assign n16321 = x11 & n16320;
  assign n16322 = n10956 & n16321;
  assign n16323 = ~n16317 & ~n16322;
  assign n16324 = x10 & n16323;
  assign n16325 = n10957 & n16321;
  assign n16326 = n7536 & ~n10956;
  assign n16327 = ~x10 & ~n16326;
  assign n16328 = ~n16325 & n16327;
  assign n16329 = ~n16324 & ~n16328;
  assign n16330 = ~n7551 & n16320;
  assign n16331 = n16330 ^ x11;
  assign n16332 = ~n16329 & n16331;
  assign n16316 = n16266 ^ n15759;
  assign n16333 = n16332 ^ n16316;
  assign n16342 = n16263 ^ n15777;
  assign n16334 = n5814 & ~n11694;
  assign n16335 = n6295 & ~n10663;
  assign n16336 = n5824 & n10680;
  assign n16337 = n5817 & n10665;
  assign n16338 = ~n16336 & ~n16337;
  assign n16339 = ~n16335 & n16338;
  assign n16340 = ~n16334 & n16339;
  assign n16341 = n16340 ^ x11;
  assign n16343 = n16342 ^ n16341;
  assign n16352 = n16260 ^ n15795;
  assign n16344 = n5814 & n12100;
  assign n16345 = n5817 & n10680;
  assign n16346 = n5824 & n10683;
  assign n16347 = ~n16345 & ~n16346;
  assign n16348 = n6295 & n10665;
  assign n16349 = n16347 & ~n16348;
  assign n16350 = ~n16344 & n16349;
  assign n16351 = n16350 ^ x11;
  assign n16353 = n16352 ^ n16351;
  assign n16355 = n5814 & n12524;
  assign n16356 = n6295 & n10680;
  assign n16357 = n5817 & n10683;
  assign n16358 = n5824 & n10694;
  assign n16359 = ~n16357 & ~n16358;
  assign n16360 = ~n16356 & n16359;
  assign n16361 = ~n16355 & n16360;
  assign n16362 = n16361 ^ x11;
  assign n16354 = n16257 ^ n15813;
  assign n16363 = n16362 ^ n16354;
  assign n16372 = n16254 ^ n15831;
  assign n16364 = n5814 & n11599;
  assign n16365 = n5817 & n10694;
  assign n16366 = n5824 & n10698;
  assign n16367 = ~n16365 & ~n16366;
  assign n16368 = n6295 & n10683;
  assign n16369 = n16367 & ~n16368;
  assign n16370 = ~n16364 & n16369;
  assign n16371 = n16370 ^ x11;
  assign n16373 = n16372 ^ n16371;
  assign n16375 = n5814 & n12087;
  assign n16376 = n6295 & n10694;
  assign n16377 = n5824 & n10715;
  assign n16378 = n5817 & n10698;
  assign n16379 = ~n16377 & ~n16378;
  assign n16380 = ~n16376 & n16379;
  assign n16381 = ~n16375 & n16380;
  assign n16382 = n16381 ^ x11;
  assign n16374 = n16251 ^ n15849;
  assign n16383 = n16382 ^ n16374;
  assign n16385 = n5814 & n12034;
  assign n16386 = n5817 & n10715;
  assign n16387 = n6295 & n10698;
  assign n16388 = n5824 & n10718;
  assign n16389 = ~n16387 & ~n16388;
  assign n16390 = ~n16386 & n16389;
  assign n16391 = ~n16385 & n16390;
  assign n16392 = n16391 ^ x11;
  assign n16384 = n16248 ^ n15867;
  assign n16393 = n16392 ^ n16384;
  assign n16395 = n5814 & n12111;
  assign n16396 = n6295 & n10715;
  assign n16397 = n5824 & ~n10736;
  assign n16398 = n5817 & n10718;
  assign n16399 = ~n16397 & ~n16398;
  assign n16400 = ~n16396 & n16399;
  assign n16401 = ~n16395 & n16400;
  assign n16402 = n16401 ^ x11;
  assign n16394 = n16245 ^ n15885;
  assign n16403 = n16402 ^ n16394;
  assign n16412 = n16242 ^ n15905;
  assign n16404 = n5814 & n12180;
  assign n16405 = n5817 & ~n10736;
  assign n16406 = n5824 & n10738;
  assign n16407 = ~n16405 & ~n16406;
  assign n16408 = n6295 & n10718;
  assign n16409 = n16407 & ~n16408;
  assign n16410 = ~n16404 & n16409;
  assign n16411 = n16410 ^ x11;
  assign n16413 = n16412 ^ n16411;
  assign n16415 = n5814 & ~n12596;
  assign n16416 = n6295 & ~n10736;
  assign n16417 = n5817 & n10738;
  assign n16418 = n5824 & n10740;
  assign n16419 = ~n16417 & ~n16418;
  assign n16420 = ~n16416 & n16419;
  assign n16421 = ~n16415 & n16420;
  assign n16422 = n16421 ^ x11;
  assign n16414 = n16239 ^ n15923;
  assign n16423 = n16422 ^ n16414;
  assign n16425 = n5814 & n12194;
  assign n16426 = n6295 & n10738;
  assign n16427 = n5817 & n10740;
  assign n16428 = n5824 & n10751;
  assign n16429 = ~n16427 & ~n16428;
  assign n16430 = ~n16426 & n16429;
  assign n16431 = ~n16425 & n16430;
  assign n16432 = n16431 ^ x11;
  assign n16424 = n16236 ^ n15941;
  assign n16433 = n16432 ^ n16424;
  assign n16435 = n5814 & n13141;
  assign n16436 = n6295 & n10740;
  assign n16437 = n5817 & n10751;
  assign n16438 = n5824 & ~n10756;
  assign n16439 = ~n16437 & ~n16438;
  assign n16440 = ~n16436 & n16439;
  assign n16441 = ~n16435 & n16440;
  assign n16442 = n16441 ^ x11;
  assign n16434 = n16233 ^ n15961;
  assign n16443 = n16442 ^ n16434;
  assign n16445 = n5814 & n12940;
  assign n16446 = n6295 & n10751;
  assign n16447 = n5817 & ~n10756;
  assign n16448 = n5824 & n10757;
  assign n16449 = ~n16447 & ~n16448;
  assign n16450 = ~n16446 & n16449;
  assign n16451 = ~n16445 & n16450;
  assign n16452 = n16451 ^ x11;
  assign n16444 = n16230 ^ n15978;
  assign n16453 = n16452 ^ n16444;
  assign n16455 = n5814 & ~n12703;
  assign n16456 = n6295 & ~n10756;
  assign n16457 = n5817 & n10757;
  assign n16458 = n5824 & n10773;
  assign n16459 = ~n16457 & ~n16458;
  assign n16460 = ~n16456 & n16459;
  assign n16461 = ~n16455 & n16460;
  assign n16462 = n16461 ^ x11;
  assign n16454 = n16227 ^ n15996;
  assign n16463 = n16462 ^ n16454;
  assign n16465 = n5814 & n12818;
  assign n16466 = n6295 & n10757;
  assign n16467 = n5824 & ~n10776;
  assign n16468 = ~n16466 & ~n16467;
  assign n16469 = n5817 & n10773;
  assign n16470 = n16468 & ~n16469;
  assign n16471 = ~n16465 & n16470;
  assign n16472 = n16471 ^ x11;
  assign n16464 = n16224 ^ n16014;
  assign n16473 = n16472 ^ n16464;
  assign n16475 = ~x10 & n13155;
  assign n16476 = x10 & n10773;
  assign n16477 = x11 & ~n16476;
  assign n16478 = ~n16475 & n16477;
  assign n16479 = ~n7550 & ~n16478;
  assign n16480 = n5817 & ~n10776;
  assign n16481 = n5824 & ~n10777;
  assign n16482 = ~n16480 & ~n16481;
  assign n16483 = ~n16479 & n16482;
  assign n16484 = x10 & ~n13155;
  assign n16485 = ~x10 & ~n10773;
  assign n16486 = n7536 & ~n16485;
  assign n16487 = ~n16484 & n16486;
  assign n16488 = ~x11 & ~n16482;
  assign n16489 = ~n16487 & ~n16488;
  assign n16490 = ~n16483 & n16489;
  assign n16474 = n16221 ^ n16220;
  assign n16491 = n16490 ^ n16474;
  assign n16507 = n16200 ^ n16032;
  assign n16492 = n5824 & n10785;
  assign n16493 = n5817 & ~n10777;
  assign n16494 = ~n16492 & ~n16493;
  assign n16496 = ~x11 & n10776;
  assign n16497 = ~n13166 & ~n16496;
  assign n16498 = ~n7536 & ~n10776;
  assign n16499 = n16497 & ~n16498;
  assign n16500 = n10776 ^ x10;
  assign n16501 = n13166 & ~n16500;
  assign n16502 = ~n16499 & ~n16501;
  assign n16495 = n16494 ^ x11;
  assign n16503 = n16502 ^ n16495;
  assign n16504 = n16494 & n16503;
  assign n16505 = n5812 & n16504;
  assign n16506 = n16505 ^ n16495;
  assign n16508 = n16507 ^ n16506;
  assign n16510 = n7536 & ~n12832;
  assign n16511 = n5817 & n10785;
  assign n16512 = n5824 & ~n10789;
  assign n16513 = ~n16511 & ~n16512;
  assign n16514 = x11 & n16513;
  assign n16515 = n10777 & n16514;
  assign n16516 = ~n16510 & ~n16515;
  assign n16517 = x10 & n16516;
  assign n16518 = n12832 & n16514;
  assign n16519 = n7536 & ~n10777;
  assign n16520 = ~x10 & ~n16519;
  assign n16521 = ~n16518 & n16520;
  assign n16522 = ~n16517 & ~n16521;
  assign n16523 = ~n7551 & n16513;
  assign n16524 = n16523 ^ x11;
  assign n16525 = ~n16522 & n16524;
  assign n16509 = n16197 ^ n16050;
  assign n16526 = n16525 ^ n16509;
  assign n16657 = n16194 ^ n16068;
  assign n16528 = n7536 & ~n13224;
  assign n16529 = n5817 & ~n10795;
  assign n16530 = n5824 & ~n10799;
  assign n16531 = ~n16529 & ~n16530;
  assign n16532 = x11 & n16531;
  assign n16533 = n10789 & n16532;
  assign n16534 = ~n16528 & ~n16533;
  assign n16535 = x10 & n16534;
  assign n16536 = n13224 & n16532;
  assign n16537 = n7536 & ~n10789;
  assign n16538 = ~x10 & ~n16537;
  assign n16539 = ~n16536 & n16538;
  assign n16540 = ~n16535 & ~n16539;
  assign n16541 = ~n7551 & n16531;
  assign n16542 = n16541 ^ x11;
  assign n16543 = ~n16540 & n16542;
  assign n16527 = n16191 ^ n16090;
  assign n16544 = n16543 ^ n16527;
  assign n16561 = n16151 ^ n16150;
  assign n16562 = n16561 ^ n16130;
  assign n16564 = n5814 & n13387;
  assign n16565 = n6295 & n10815;
  assign n16566 = n5817 & n10819;
  assign n16567 = n5824 & ~n10820;
  assign n16568 = ~n16566 & ~n16567;
  assign n16569 = ~n16565 & n16568;
  assign n16570 = ~n16564 & n16569;
  assign n16571 = n16570 ^ x11;
  assign n16563 = n16149 ^ n16145;
  assign n16572 = n16571 ^ n16563;
  assign n16581 = ~n5744 & ~n10822;
  assign n16582 = n8210 & ~n16581;
  assign n16583 = ~n5743 & ~n16582;
  assign n16584 = n10825 & ~n16583;
  assign n16585 = n5748 & n10825;
  assign n16586 = x13 & n16585;
  assign n16587 = n16586 ^ n5748;
  assign n16588 = ~n10822 & n16587;
  assign n16589 = ~n16584 & ~n16588;
  assign n16573 = n5814 & n13429;
  assign n16574 = n6295 & n10819;
  assign n16575 = n5817 & ~n10820;
  assign n16576 = n5824 & n10821;
  assign n16577 = ~n16575 & ~n16576;
  assign n16578 = ~n16574 & n16577;
  assign n16579 = ~n16573 & n16578;
  assign n16580 = n16579 ^ x11;
  assign n16590 = n16589 ^ n16580;
  assign n16591 = n5814 & n10821;
  assign n16592 = ~n5824 & ~n16591;
  assign n16593 = n10825 & ~n16592;
  assign n16594 = n6295 & n10821;
  assign n16595 = ~n16593 & ~n16594;
  assign n16596 = ~n10853 & ~n16131;
  assign n16597 = n5814 & n16596;
  assign n16598 = n16595 & ~n16597;
  assign n16599 = x11 & n16598;
  assign n16600 = n5823 & ~n14128;
  assign n16601 = n16599 & ~n16600;
  assign n16602 = ~n16585 & ~n16601;
  assign n16603 = n5814 & ~n14111;
  assign n16604 = n6295 & ~n10820;
  assign n16605 = n5817 & n10821;
  assign n16606 = n5824 & ~n10822;
  assign n16607 = ~n16605 & ~n16606;
  assign n16608 = ~n16604 & n16607;
  assign n16609 = ~n16603 & n16608;
  assign n16610 = n16609 ^ x11;
  assign n16611 = ~n16602 & ~n16610;
  assign n16612 = n16611 ^ n16589;
  assign n16613 = ~n16590 & ~n16612;
  assign n16614 = n16613 ^ n16611;
  assign n16615 = n16614 ^ n16563;
  assign n16616 = n16572 & n16615;
  assign n16617 = n16616 ^ n16571;
  assign n16618 = ~n16562 & ~n16617;
  assign n16619 = n5814 & ~n13341;
  assign n16620 = n6295 & ~n10800;
  assign n16621 = n5824 & n10819;
  assign n16622 = ~n16620 & ~n16621;
  assign n16623 = n5817 & n10815;
  assign n16624 = n16622 & ~n16623;
  assign n16625 = ~n16619 & n16624;
  assign n16626 = n16625 ^ x11;
  assign n16627 = n16153 ^ n16113;
  assign n16628 = n16627 ^ n16097;
  assign n16629 = n5814 & ~n13278;
  assign n16630 = n6295 & ~n10799;
  assign n16631 = n5817 & ~n10800;
  assign n16632 = n5824 & n10815;
  assign n16633 = ~n16631 & ~n16632;
  assign n16634 = ~n16630 & n16633;
  assign n16635 = ~n16629 & n16634;
  assign n16636 = n16635 ^ n16625;
  assign n16637 = n16628 & n16636;
  assign n16638 = n16626 & n16637;
  assign n16639 = n16638 ^ n16626;
  assign n16640 = ~n16618 & n16639;
  assign n16641 = n16635 ^ x11;
  assign n16642 = n16641 ^ n16628;
  assign n16643 = n16562 & n16617;
  assign n16644 = n16643 ^ n16641;
  assign n16645 = ~n16642 & ~n16644;
  assign n16646 = n16645 ^ n16628;
  assign n16647 = ~n16640 & n16646;
  assign n16545 = n7536 & ~n13239;
  assign n16546 = n5817 & ~n10799;
  assign n16547 = n5824 & ~n10800;
  assign n16548 = ~n16546 & ~n16547;
  assign n16549 = x11 & n16548;
  assign n16550 = n10795 & n16549;
  assign n16551 = x10 & ~n16550;
  assign n16552 = ~n16545 & n16551;
  assign n16553 = n13239 & n16549;
  assign n16554 = n7536 & ~n10795;
  assign n16555 = ~x10 & ~n16554;
  assign n16556 = ~n16553 & n16555;
  assign n16557 = ~n16552 & ~n16556;
  assign n16558 = ~n7551 & n16548;
  assign n16559 = n16558 ^ x11;
  assign n16560 = ~n16557 & n16559;
  assign n16648 = n16647 ^ n16560;
  assign n16649 = n16188 ^ n16156;
  assign n16650 = n16649 ^ n16172;
  assign n16651 = n16650 ^ n16560;
  assign n16652 = ~n16648 & ~n16651;
  assign n16653 = n16652 ^ n16647;
  assign n16654 = n16653 ^ n16527;
  assign n16655 = n16544 & n16654;
  assign n16656 = n16655 ^ n16543;
  assign n16658 = n16657 ^ n16656;
  assign n16659 = n7536 & n13197;
  assign n16660 = n5824 & ~n10795;
  assign n16661 = n5817 & ~n10789;
  assign n16662 = ~n16660 & ~n16661;
  assign n16663 = x11 & n16662;
  assign n16664 = ~n10785 & n16663;
  assign n16665 = x10 & ~n16664;
  assign n16666 = ~n16659 & n16665;
  assign n16667 = ~n13197 & n16663;
  assign n16668 = n7536 & n10785;
  assign n16669 = ~x10 & ~n16668;
  assign n16670 = ~n16667 & n16669;
  assign n16671 = ~n16666 & ~n16670;
  assign n16672 = ~n7551 & n16662;
  assign n16673 = n16672 ^ x11;
  assign n16674 = ~n16671 & n16673;
  assign n16675 = n16674 ^ n16657;
  assign n16676 = ~n16658 & n16675;
  assign n16677 = n16676 ^ n16656;
  assign n16678 = n16677 ^ n16509;
  assign n16679 = n16526 & ~n16678;
  assign n16680 = n16679 ^ n16525;
  assign n16681 = n16680 ^ n16506;
  assign n16682 = ~n16508 & n16681;
  assign n16683 = n16682 ^ n16680;
  assign n16684 = n16683 ^ n16490;
  assign n16685 = n16491 & n16684;
  assign n16686 = n16685 ^ n16683;
  assign n16687 = n16686 ^ n16472;
  assign n16688 = ~n16473 & n16687;
  assign n16689 = n16688 ^ n16686;
  assign n16690 = n16689 ^ n16462;
  assign n16691 = ~n16463 & n16690;
  assign n16692 = n16691 ^ n16689;
  assign n16693 = n16692 ^ n16452;
  assign n16694 = ~n16453 & n16693;
  assign n16695 = n16694 ^ n16692;
  assign n16696 = n16695 ^ n16442;
  assign n16697 = n16443 & n16696;
  assign n16698 = n16697 ^ n16695;
  assign n16699 = n16698 ^ n16432;
  assign n16700 = n16433 & n16699;
  assign n16701 = n16700 ^ n16698;
  assign n16702 = n16701 ^ n16422;
  assign n16703 = ~n16423 & n16702;
  assign n16704 = n16703 ^ n16701;
  assign n16705 = n16704 ^ n16412;
  assign n16706 = n16413 & ~n16705;
  assign n16707 = n16706 ^ n16704;
  assign n16708 = n16707 ^ n16402;
  assign n16709 = ~n16403 & n16708;
  assign n16710 = n16709 ^ n16707;
  assign n16711 = n16710 ^ n16392;
  assign n16712 = ~n16393 & n16711;
  assign n16713 = n16712 ^ n16710;
  assign n16714 = n16713 ^ n16382;
  assign n16715 = ~n16383 & n16714;
  assign n16716 = n16715 ^ n16713;
  assign n16717 = n16716 ^ n16372;
  assign n16718 = ~n16373 & n16717;
  assign n16719 = n16718 ^ n16716;
  assign n16720 = n16719 ^ n16362;
  assign n16721 = ~n16363 & n16720;
  assign n16722 = n16721 ^ n16719;
  assign n16723 = n16722 ^ n16352;
  assign n16724 = ~n16353 & n16723;
  assign n16725 = n16724 ^ n16722;
  assign n16726 = n16725 ^ n16342;
  assign n16727 = n16343 & ~n16726;
  assign n16728 = n16727 ^ n16725;
  assign n16729 = n16728 ^ n16332;
  assign n16730 = ~n16333 & n16729;
  assign n16731 = n16730 ^ n16728;
  assign n16732 = n16731 ^ n16314;
  assign n16733 = n16315 & ~n16732;
  assign n16734 = n16733 ^ n16731;
  assign n16735 = n16734 ^ n16304;
  assign n16736 = n16305 & ~n16735;
  assign n16737 = n16736 ^ n16734;
  assign n17321 = n16780 ^ n16737;
  assign n17322 = n16781 & ~n17321;
  assign n17323 = n17322 ^ n16737;
  assign n17381 = n17380 ^ n17323;
  assign n17391 = n17390 ^ n17381;
  assign n16782 = n16781 ^ n16737;
  assign n15373 = n6306 & ~n12000;
  assign n15374 = n7168 & ~n11875;
  assign n15375 = n6309 & ~n11773;
  assign n15376 = n6316 & n11480;
  assign n15377 = ~n15375 & ~n15376;
  assign n15378 = ~n15374 & n15377;
  assign n15379 = ~n15373 & n15378;
  assign n15380 = n15379 ^ x8;
  assign n16783 = n16782 ^ n15380;
  assign n16792 = n16734 ^ n16305;
  assign n16784 = n6306 & ~n11777;
  assign n16785 = n7168 & ~n11773;
  assign n16786 = n6316 & n11500;
  assign n16787 = n6309 & n11480;
  assign n16788 = ~n16786 & ~n16787;
  assign n16789 = ~n16785 & n16788;
  assign n16790 = ~n16784 & n16789;
  assign n16791 = n16790 ^ x8;
  assign n16793 = n16792 ^ n16791;
  assign n16802 = n16731 ^ n16315;
  assign n16794 = n6306 & n11507;
  assign n16795 = n7168 & n11480;
  assign n16796 = n6309 & n11500;
  assign n16797 = ~n16795 & ~n16796;
  assign n16798 = n6316 & n11486;
  assign n16799 = n16797 & ~n16798;
  assign n16800 = ~n16794 & n16799;
  assign n16801 = n16800 ^ x8;
  assign n16803 = n16802 ^ n16801;
  assign n16806 = n11957 & n16805;
  assign n16807 = n6309 & n11486;
  assign n16808 = n6316 & n11215;
  assign n16809 = ~n16807 & ~n16808;
  assign n16810 = x8 & n16809;
  assign n16811 = ~n11500 & n16810;
  assign n16812 = x7 & ~n16811;
  assign n16813 = ~n16806 & n16812;
  assign n16814 = ~n11957 & n16810;
  assign n16815 = n11500 & n16805;
  assign n16816 = ~x7 & ~n16815;
  assign n16817 = ~n16814 & n16816;
  assign n16818 = ~n16813 & ~n16817;
  assign n16821 = n16809 & ~n16820;
  assign n16822 = n16821 ^ x8;
  assign n16823 = ~n16818 & n16822;
  assign n16804 = n16728 ^ n16333;
  assign n16824 = n16823 ^ n16804;
  assign n16833 = n16725 ^ n16343;
  assign n16825 = n6306 & n11704;
  assign n16826 = n7168 & n11486;
  assign n16827 = n6309 & n11215;
  assign n16828 = n6316 & ~n10956;
  assign n16829 = ~n16827 & ~n16828;
  assign n16830 = ~n16826 & n16829;
  assign n16831 = ~n16825 & n16830;
  assign n16832 = n16831 ^ x8;
  assign n16834 = n16833 ^ n16832;
  assign n16843 = ~n12460 & n16805;
  assign n16836 = n6316 & ~n10663;
  assign n16837 = n6309 & ~n10956;
  assign n16838 = ~n16836 & ~n16837;
  assign n16839 = x8 & n16838;
  assign n16844 = ~n11215 & n16839;
  assign n16845 = ~n16843 & ~n16844;
  assign n16840 = n12460 & n16839;
  assign n16841 = n11215 & n16805;
  assign n16842 = ~n16840 & ~n16841;
  assign n16846 = n16845 ^ n16842;
  assign n16847 = ~x7 & n16846;
  assign n16848 = n16847 ^ n16845;
  assign n16849 = ~n16820 & n16838;
  assign n16850 = n16849 ^ x8;
  assign n16851 = n16848 & n16850;
  assign n16835 = n16722 ^ n16353;
  assign n16852 = n16851 ^ n16835;
  assign n16861 = n16719 ^ n16363;
  assign n16853 = n6306 & ~n10957;
  assign n16854 = n6309 & ~n10663;
  assign n16855 = n7168 & ~n10956;
  assign n16856 = n6316 & n10665;
  assign n16857 = ~n16855 & ~n16856;
  assign n16858 = ~n16854 & n16857;
  assign n16859 = ~n16853 & n16858;
  assign n16860 = n16859 ^ x8;
  assign n16862 = n16861 ^ n16860;
  assign n16871 = n16716 ^ n16373;
  assign n16863 = n6306 & ~n11694;
  assign n16864 = n7168 & ~n10663;
  assign n16865 = n6316 & n10680;
  assign n16866 = n6309 & n10665;
  assign n16867 = ~n16865 & ~n16866;
  assign n16868 = ~n16864 & n16867;
  assign n16869 = ~n16863 & n16868;
  assign n16870 = n16869 ^ x8;
  assign n16872 = n16871 ^ n16870;
  assign n16874 = n6306 & n12100;
  assign n16875 = n6309 & n10680;
  assign n16876 = n6316 & n10683;
  assign n16877 = ~n16875 & ~n16876;
  assign n16878 = n7168 & n10665;
  assign n16879 = n16877 & ~n16878;
  assign n16880 = ~n16874 & n16879;
  assign n16881 = n16880 ^ x8;
  assign n16873 = n16713 ^ n16383;
  assign n16882 = n16881 ^ n16873;
  assign n16884 = n6306 & n12524;
  assign n16885 = n7168 & n10680;
  assign n16886 = n6309 & n10683;
  assign n16887 = n6316 & n10694;
  assign n16888 = ~n16886 & ~n16887;
  assign n16889 = ~n16885 & n16888;
  assign n16890 = ~n16884 & n16889;
  assign n16891 = n16890 ^ x8;
  assign n16883 = n16710 ^ n16393;
  assign n16892 = n16891 ^ n16883;
  assign n16894 = n6306 & n11599;
  assign n16895 = n6309 & n10694;
  assign n16896 = n6316 & n10698;
  assign n16897 = ~n16895 & ~n16896;
  assign n16898 = n7168 & n10683;
  assign n16899 = n16897 & ~n16898;
  assign n16900 = ~n16894 & n16899;
  assign n16901 = n16900 ^ x8;
  assign n16893 = n16707 ^ n16403;
  assign n16902 = n16901 ^ n16893;
  assign n16904 = n12087 & n16805;
  assign n16905 = n6316 & n10715;
  assign n16906 = n6309 & n10698;
  assign n16907 = ~n16905 & ~n16906;
  assign n16908 = x8 & n16907;
  assign n16909 = ~n10694 & n16908;
  assign n16910 = x7 & ~n16909;
  assign n16911 = ~n16904 & n16910;
  assign n16912 = ~n12087 & n16908;
  assign n16913 = n10694 & n16805;
  assign n16914 = ~x7 & ~n16913;
  assign n16915 = ~n16912 & n16914;
  assign n16916 = ~n16911 & ~n16915;
  assign n16917 = ~n16820 & n16907;
  assign n16918 = n16917 ^ x8;
  assign n16919 = ~n16916 & n16918;
  assign n16903 = n16704 ^ n16413;
  assign n16920 = n16919 ^ n16903;
  assign n16922 = n12034 & n16805;
  assign n16923 = n6309 & n10715;
  assign n16924 = n6316 & n10718;
  assign n16925 = ~n16923 & ~n16924;
  assign n16926 = x8 & n16925;
  assign n16927 = ~n10698 & n16926;
  assign n16928 = ~n16922 & ~n16927;
  assign n16929 = x7 & n16928;
  assign n16930 = ~n12034 & n16926;
  assign n16931 = n10698 & n16805;
  assign n16932 = ~x7 & ~n16931;
  assign n16933 = ~n16930 & n16932;
  assign n16934 = ~n16929 & ~n16933;
  assign n16935 = ~n16820 & n16925;
  assign n16936 = n16935 ^ x8;
  assign n16937 = ~n16934 & n16936;
  assign n16921 = n16701 ^ n16423;
  assign n16938 = n16937 ^ n16921;
  assign n16940 = n12111 & n16805;
  assign n16941 = n6316 & ~n10736;
  assign n16942 = n6309 & n10718;
  assign n16943 = ~n16941 & ~n16942;
  assign n16944 = x8 & n16943;
  assign n16945 = ~n10715 & n16944;
  assign n16946 = x7 & ~n16945;
  assign n16947 = ~n16940 & n16946;
  assign n16948 = ~n12111 & n16944;
  assign n16949 = n10715 & n16805;
  assign n16950 = ~x7 & ~n16949;
  assign n16951 = ~n16948 & n16950;
  assign n16952 = ~n16947 & ~n16951;
  assign n16953 = ~n16820 & n16943;
  assign n16954 = n16953 ^ x8;
  assign n16955 = ~n16952 & n16954;
  assign n16939 = n16698 ^ n16433;
  assign n16956 = n16955 ^ n16939;
  assign n16958 = n12180 & n16805;
  assign n16959 = n6309 & ~n10736;
  assign n16960 = n6316 & n10738;
  assign n16961 = ~n16959 & ~n16960;
  assign n16962 = x8 & n16961;
  assign n16963 = ~n10718 & n16962;
  assign n16964 = ~n16958 & ~n16963;
  assign n16965 = x7 & n16964;
  assign n16966 = ~n12180 & n16962;
  assign n16967 = n10718 & n16805;
  assign n16968 = ~x7 & ~n16967;
  assign n16969 = ~n16966 & n16968;
  assign n16970 = ~n16965 & ~n16969;
  assign n16971 = ~n16820 & n16961;
  assign n16972 = n16971 ^ x8;
  assign n16973 = ~n16970 & n16972;
  assign n16957 = n16695 ^ n16443;
  assign n16974 = n16973 ^ n16957;
  assign n16976 = n6306 & ~n12596;
  assign n16977 = n7168 & ~n10736;
  assign n16978 = n6309 & n10738;
  assign n16979 = n6316 & n10740;
  assign n16980 = ~n16978 & ~n16979;
  assign n16981 = ~n16977 & n16980;
  assign n16982 = ~n16976 & n16981;
  assign n16983 = n16982 ^ x8;
  assign n16975 = n16692 ^ n16453;
  assign n16984 = n16983 ^ n16975;
  assign n16986 = n12194 & n16805;
  assign n16987 = n6309 & n10740;
  assign n16988 = n6316 & n10751;
  assign n16989 = ~n16987 & ~n16988;
  assign n16990 = x8 & n16989;
  assign n16991 = ~n10738 & n16990;
  assign n16992 = x7 & ~n16991;
  assign n16993 = ~n16986 & n16992;
  assign n16994 = ~n12194 & n16990;
  assign n16995 = n10738 & n16805;
  assign n16996 = ~x7 & ~n16995;
  assign n16997 = ~n16994 & n16996;
  assign n16998 = ~n16993 & ~n16997;
  assign n16999 = ~n16820 & n16989;
  assign n17000 = n16999 ^ x8;
  assign n17001 = ~n16998 & n17000;
  assign n16985 = n16689 ^ n16463;
  assign n17002 = n17001 ^ n16985;
  assign n17004 = n6306 & n13141;
  assign n17005 = n7168 & n10740;
  assign n17006 = n6309 & n10751;
  assign n17007 = n6316 & ~n10756;
  assign n17008 = ~n17006 & ~n17007;
  assign n17009 = ~n17005 & n17008;
  assign n17010 = ~n17004 & n17009;
  assign n17011 = n17010 ^ x8;
  assign n17003 = n16686 ^ n16473;
  assign n17012 = n17011 ^ n17003;
  assign n17014 = n6309 & ~n10756;
  assign n17015 = n6316 & n10757;
  assign n17016 = ~n17014 & ~n17015;
  assign n17017 = x8 & n17016;
  assign n17018 = ~n12940 & n17017;
  assign n17019 = n10751 & n16805;
  assign n17020 = ~n17018 & ~n17019;
  assign n17021 = ~x7 & ~n17020;
  assign n17022 = ~n16820 & n17016;
  assign n17023 = n17022 ^ x8;
  assign n17024 = ~n17021 & n17023;
  assign n17025 = n12940 & n16805;
  assign n17026 = ~n10751 & n17017;
  assign n17027 = ~n17025 & ~n17026;
  assign n17028 = x7 & ~n17027;
  assign n17029 = n17024 & ~n17028;
  assign n17013 = n16683 ^ n16491;
  assign n17030 = n17029 ^ n17013;
  assign n17031 = n16653 ^ n16544;
  assign n17033 = n6306 & ~n12832;
  assign n17034 = n7168 & ~n10777;
  assign n17035 = n6316 & ~n10789;
  assign n17036 = ~n17034 & ~n17035;
  assign n17037 = n6309 & n10785;
  assign n17038 = n17036 & ~n17037;
  assign n17039 = ~n17033 & n17038;
  assign n17040 = n17039 ^ x8;
  assign n17032 = n16650 ^ n16648;
  assign n17041 = n17040 ^ n17032;
  assign n17175 = n16635 ^ n16628;
  assign n17042 = n16617 ^ n16562;
  assign n17172 = n16626 ^ n16562;
  assign n17173 = ~n17042 & n17172;
  assign n17174 = n17173 ^ n16625;
  assign n17176 = n17175 ^ n17174;
  assign n17044 = n6306 & ~n13224;
  assign n17045 = n7168 & ~n10789;
  assign n17046 = n6316 & ~n10799;
  assign n17047 = ~n17045 & ~n17046;
  assign n17048 = n6309 & ~n10795;
  assign n17049 = n17047 & ~n17048;
  assign n17050 = ~n17044 & n17049;
  assign n17051 = n17050 ^ x8;
  assign n17043 = n17042 ^ n16626;
  assign n17052 = n17051 ^ n17043;
  assign n17055 = n6306 & ~n13239;
  assign n17056 = n7168 & ~n10795;
  assign n17057 = n6309 & ~n10799;
  assign n17058 = n6316 & ~n10800;
  assign n17059 = ~n17057 & ~n17058;
  assign n17060 = ~n17056 & n17059;
  assign n17061 = ~n17055 & n17060;
  assign n17062 = n17061 ^ x8;
  assign n17053 = n16614 ^ n16571;
  assign n17054 = n17053 ^ n16563;
  assign n17063 = n17062 ^ n17054;
  assign n17065 = n6306 & ~n13278;
  assign n17066 = n7168 & ~n10799;
  assign n17067 = n6309 & ~n10800;
  assign n17068 = n6316 & n10815;
  assign n17069 = ~n17067 & ~n17068;
  assign n17070 = ~n17066 & n17069;
  assign n17071 = ~n17065 & n17070;
  assign n17072 = n17071 ^ x8;
  assign n17064 = n16611 ^ n16590;
  assign n17073 = n17072 ^ n17064;
  assign n17076 = n6306 & ~n13341;
  assign n17077 = n7168 & ~n10800;
  assign n17078 = n6316 & n10819;
  assign n17079 = ~n17077 & ~n17078;
  assign n17080 = n6309 & n10815;
  assign n17081 = n17079 & ~n17080;
  assign n17082 = ~n17076 & n17081;
  assign n17083 = n17082 ^ x8;
  assign n17074 = n16601 ^ n16585;
  assign n17075 = n17074 ^ n16610;
  assign n17084 = n17083 ^ n17075;
  assign n17128 = ~n5812 & ~n10822;
  assign n17129 = n16600 & ~n17128;
  assign n17130 = n16599 & n17129;
  assign n17131 = x11 & n5812;
  assign n17132 = ~n14128 & n17131;
  assign n17133 = ~n16598 & ~n17132;
  assign n17134 = n5817 & n13532;
  assign n17135 = ~x11 & n5817;
  assign n17136 = ~n10822 & n17135;
  assign n17137 = ~n17134 & ~n17136;
  assign n17138 = ~n17133 & n17137;
  assign n17139 = ~n17130 & n17138;
  assign n17094 = n6306 & n13429;
  assign n17095 = n7168 & n10819;
  assign n17096 = n6309 & ~n10820;
  assign n17097 = n6316 & n10821;
  assign n17098 = ~n17096 & ~n17097;
  assign n17099 = ~n17095 & n17098;
  assign n17100 = ~n17094 & n17099;
  assign n17101 = n17100 ^ x8;
  assign n17085 = ~n5819 & ~n10822;
  assign n17086 = n8711 & ~n17085;
  assign n17087 = ~n8713 & ~n17086;
  assign n17088 = n10825 & ~n17087;
  assign n17089 = n5812 & n10825;
  assign n17090 = x10 & n17089;
  assign n17091 = n17090 ^ n5812;
  assign n17092 = ~n10822 & n17091;
  assign n17093 = ~n17088 & ~n17092;
  assign n17102 = n17101 ^ n17093;
  assign n17103 = n6306 & n10821;
  assign n17104 = ~n6316 & ~n17103;
  assign n17105 = n10825 & ~n17104;
  assign n17106 = n7168 & n10821;
  assign n17107 = ~n17105 & ~n17106;
  assign n17108 = n6306 & n16596;
  assign n17109 = n17107 & ~n17108;
  assign n17110 = x8 & n17109;
  assign n17111 = n6315 & n10825;
  assign n17112 = n17110 & ~n17111;
  assign n17113 = n6315 & ~n10822;
  assign n17114 = n17112 & ~n17113;
  assign n17115 = ~n17089 & ~n17114;
  assign n17116 = n6306 & ~n14111;
  assign n17117 = n7168 & ~n10820;
  assign n17118 = n6309 & n10821;
  assign n17119 = n6316 & ~n10822;
  assign n17120 = ~n17118 & ~n17119;
  assign n17121 = ~n17117 & n17120;
  assign n17122 = ~n17116 & n17121;
  assign n17123 = n17122 ^ x8;
  assign n17124 = ~n17115 & ~n17123;
  assign n17125 = n17124 ^ n17101;
  assign n17126 = ~n17102 & ~n17125;
  assign n17127 = n17126 ^ n17124;
  assign n17140 = n17139 ^ n17127;
  assign n17141 = n13387 & n16805;
  assign n17142 = n6309 & n10819;
  assign n17143 = n6316 & ~n10820;
  assign n17144 = ~n17142 & ~n17143;
  assign n17145 = x8 & n17144;
  assign n17146 = ~n10815 & n17145;
  assign n17147 = x7 & ~n17146;
  assign n17148 = ~n17141 & n17147;
  assign n17149 = ~n13387 & n17145;
  assign n17150 = n10815 & n16805;
  assign n17151 = ~x7 & ~n17150;
  assign n17152 = ~n17149 & n17151;
  assign n17153 = ~n17148 & ~n17152;
  assign n17154 = ~n16820 & n17144;
  assign n17155 = n17154 ^ x8;
  assign n17156 = ~n17153 & n17155;
  assign n17157 = n17156 ^ n17127;
  assign n17158 = n17140 & ~n17157;
  assign n17159 = n17158 ^ n17156;
  assign n17160 = n17159 ^ n17083;
  assign n17161 = ~n17084 & n17160;
  assign n17162 = n17161 ^ n17159;
  assign n17163 = n17162 ^ n17072;
  assign n17164 = n17073 & n17163;
  assign n17165 = n17164 ^ n17162;
  assign n17166 = n17165 ^ n17062;
  assign n17167 = n17063 & n17166;
  assign n17168 = n17167 ^ n17165;
  assign n17169 = n17168 ^ n17051;
  assign n17170 = ~n17052 & n17169;
  assign n17171 = n17170 ^ n17168;
  assign n17177 = n17176 ^ n17171;
  assign n17178 = n13197 & n16805;
  assign n17179 = n6316 & ~n10795;
  assign n17180 = n6309 & ~n10789;
  assign n17181 = ~n17179 & ~n17180;
  assign n17182 = x8 & n17181;
  assign n17183 = ~n10785 & n17182;
  assign n17184 = x7 & ~n17183;
  assign n17185 = ~n17178 & n17184;
  assign n17186 = ~n13197 & n17182;
  assign n17187 = n10785 & n16805;
  assign n17188 = ~x7 & ~n17187;
  assign n17189 = ~n17186 & n17188;
  assign n17190 = ~n17185 & ~n17189;
  assign n17191 = ~n16820 & n17181;
  assign n17192 = n17191 ^ x8;
  assign n17193 = ~n17190 & n17192;
  assign n17194 = n17193 ^ n17176;
  assign n17195 = ~n17177 & n17194;
  assign n17196 = n17195 ^ n17171;
  assign n17197 = n17196 ^ n17040;
  assign n17198 = n17041 & n17197;
  assign n17199 = n17198 ^ n17196;
  assign n17200 = ~n17031 & n17199;
  assign n17201 = n6306 & ~n13167;
  assign n17202 = n7168 & ~n10776;
  assign n17203 = n6316 & n10785;
  assign n17204 = n6309 & ~n10777;
  assign n17205 = ~n17203 & ~n17204;
  assign n17206 = ~n17202 & n17205;
  assign n17207 = ~n17201 & n17206;
  assign n17208 = n17207 ^ x8;
  assign n17209 = n16674 ^ n16658;
  assign n17210 = n6306 & n13155;
  assign n17211 = n7168 & n10773;
  assign n17212 = n6309 & ~n10776;
  assign n17213 = n6316 & ~n10777;
  assign n17214 = ~n17212 & ~n17213;
  assign n17215 = ~n17211 & n17214;
  assign n17216 = ~n17210 & n17215;
  assign n17217 = n17216 ^ n17207;
  assign n17218 = ~n17209 & n17217;
  assign n17219 = ~n17208 & n17218;
  assign n17220 = n17219 ^ n17208;
  assign n17221 = ~n17200 & ~n17220;
  assign n17222 = n17031 & ~n17199;
  assign n17223 = n17222 ^ n17209;
  assign n17224 = n17216 ^ x8;
  assign n17225 = n17224 ^ n17222;
  assign n17226 = n17223 & n17225;
  assign n17227 = n17226 ^ n17209;
  assign n17228 = ~n17221 & ~n17227;
  assign n17229 = n16677 ^ n16526;
  assign n17230 = n17228 & n17229;
  assign n17231 = n6306 & n12818;
  assign n17232 = n7168 & n10757;
  assign n17233 = n6316 & ~n10776;
  assign n17234 = ~n17232 & ~n17233;
  assign n17235 = n6309 & n10773;
  assign n17236 = n17234 & ~n17235;
  assign n17237 = ~n17231 & n17236;
  assign n17238 = ~n17230 & ~n17237;
  assign n17239 = ~n17228 & ~n17229;
  assign n17240 = ~n17238 & ~n17239;
  assign n17241 = n6306 & ~n12703;
  assign n17242 = n7168 & ~n10756;
  assign n17243 = n6309 & n10757;
  assign n17244 = n6316 & n10773;
  assign n17245 = ~n17243 & ~n17244;
  assign n17246 = ~n17242 & n17245;
  assign n17247 = ~n17241 & n17246;
  assign n17248 = n16680 ^ n16508;
  assign n17249 = n17247 & n17248;
  assign n17250 = ~n17240 & ~n17249;
  assign n17251 = ~n17247 & ~n17248;
  assign n17252 = ~x8 & ~n17251;
  assign n17253 = ~n17250 & n17252;
  assign n17254 = ~n17247 & n17248;
  assign n17255 = n17237 ^ n17229;
  assign n17256 = n17229 ^ n17228;
  assign n17257 = n17255 & n17256;
  assign n17258 = n17257 ^ n17228;
  assign n17259 = ~n17254 & ~n17258;
  assign n17260 = n17247 & ~n17248;
  assign n17261 = x8 & ~n17260;
  assign n17262 = ~n17259 & n17261;
  assign n17263 = ~n17253 & ~n17262;
  assign n17264 = n17263 ^ n17029;
  assign n17265 = n17030 & ~n17264;
  assign n17266 = n17265 ^ n17263;
  assign n17267 = n17266 ^ n17011;
  assign n17268 = ~n17012 & ~n17267;
  assign n17269 = n17268 ^ n17266;
  assign n17270 = n17269 ^ n17001;
  assign n17271 = ~n17002 & ~n17270;
  assign n17272 = n17271 ^ n17269;
  assign n17273 = n17272 ^ n16983;
  assign n17274 = ~n16984 & ~n17273;
  assign n17275 = n17274 ^ n17272;
  assign n17276 = n17275 ^ n16973;
  assign n17277 = n16974 & ~n17276;
  assign n17278 = n17277 ^ n17275;
  assign n17279 = n17278 ^ n16955;
  assign n17280 = n16956 & ~n17279;
  assign n17281 = n17280 ^ n17278;
  assign n17282 = n17281 ^ n16937;
  assign n17283 = ~n16938 & ~n17282;
  assign n17284 = n17283 ^ n17281;
  assign n17285 = n17284 ^ n16919;
  assign n17286 = n16920 & ~n17285;
  assign n17287 = n17286 ^ n17284;
  assign n17288 = n17287 ^ n16901;
  assign n17289 = ~n16902 & ~n17288;
  assign n17290 = n17289 ^ n17287;
  assign n17291 = n17290 ^ n16891;
  assign n17292 = ~n16892 & ~n17291;
  assign n17293 = n17292 ^ n17290;
  assign n17294 = n17293 ^ n16881;
  assign n17295 = ~n16882 & ~n17294;
  assign n17296 = n17295 ^ n17293;
  assign n17297 = n17296 ^ n16871;
  assign n17298 = ~n16872 & ~n17297;
  assign n17299 = n17298 ^ n17296;
  assign n17300 = n17299 ^ n16861;
  assign n17301 = ~n16862 & ~n17300;
  assign n17302 = n17301 ^ n17299;
  assign n17303 = n17302 ^ n16851;
  assign n17304 = ~n16852 & ~n17303;
  assign n17305 = n17304 ^ n17302;
  assign n17306 = n17305 ^ n16833;
  assign n17307 = n16834 & n17306;
  assign n17308 = n17307 ^ n17305;
  assign n17309 = n17308 ^ n16823;
  assign n17310 = ~n16824 & ~n17309;
  assign n17311 = n17310 ^ n17308;
  assign n17312 = n17311 ^ n16802;
  assign n17313 = n16803 & n17312;
  assign n17314 = n17313 ^ n17311;
  assign n17315 = n17314 ^ n16792;
  assign n17316 = n16793 & n17315;
  assign n17317 = n17316 ^ n17314;
  assign n17318 = n17317 ^ n16782;
  assign n17319 = n16783 & n17318;
  assign n17320 = n17319 ^ n17317;
  assign n17392 = n17391 ^ n17320;
  assign n17393 = n17317 ^ n16783;
  assign n17914 = n17314 ^ n16793;
  assign n17906 = n7515 & ~n11941;
  assign n17907 = n8029 & ~n11940;
  assign n17908 = n7518 & n11902;
  assign n17909 = n7520 & ~n11875;
  assign n17910 = ~n17908 & ~n17909;
  assign n17911 = ~n17907 & n17910;
  assign n17912 = ~n17906 & n17911;
  assign n17913 = n17912 ^ x5;
  assign n17915 = n17914 ^ n17913;
  assign n17415 = n17311 ^ n16803;
  assign n17396 = ~x5 & n7514;
  assign n17397 = n12504 & n17396;
  assign n17398 = n7518 & ~n11875;
  assign n17399 = n7520 & ~n11773;
  assign n17400 = ~n17398 & ~n17399;
  assign n17401 = x5 & n17400;
  assign n17402 = ~n11902 & n17401;
  assign n17403 = ~n17397 & ~n17402;
  assign n17404 = x4 & n17403;
  assign n17405 = ~n12504 & n17401;
  assign n17406 = n11902 & n17396;
  assign n17407 = ~x4 & ~n17406;
  assign n17408 = ~n17405 & n17407;
  assign n17409 = ~n17404 & ~n17408;
  assign n17410 = x5 & ~n7514;
  assign n17411 = n17410 ^ x5;
  assign n17412 = n17400 & ~n17411;
  assign n17413 = n17412 ^ x5;
  assign n17414 = ~n17409 & n17413;
  assign n17416 = n17415 ^ n17414;
  assign n17425 = n17308 ^ n16824;
  assign n17417 = n7515 & ~n12000;
  assign n17418 = n8029 & ~n11875;
  assign n17419 = n7518 & ~n11773;
  assign n17420 = n7520 & n11480;
  assign n17421 = ~n17419 & ~n17420;
  assign n17422 = ~n17418 & n17421;
  assign n17423 = ~n17417 & n17422;
  assign n17424 = n17423 ^ x5;
  assign n17426 = n17425 ^ n17424;
  assign n17435 = n17305 ^ n16834;
  assign n17427 = n7513 & n11776;
  assign n17428 = n17427 ^ n11773;
  assign n17429 = n7514 & ~n17428;
  assign n17430 = n7518 & n11480;
  assign n17431 = n7520 & n11500;
  assign n17432 = ~n17430 & ~n17431;
  assign n17433 = ~n17429 & n17432;
  assign n17434 = n17433 ^ x5;
  assign n17436 = n17435 ^ n17434;
  assign n17445 = n17302 ^ n16852;
  assign n17437 = n7515 & n11507;
  assign n17438 = n8029 & n11480;
  assign n17439 = n7518 & n11500;
  assign n17440 = ~n17438 & ~n17439;
  assign n17441 = n7520 & n11486;
  assign n17442 = n17440 & ~n17441;
  assign n17443 = ~n17437 & n17442;
  assign n17444 = n17443 ^ x5;
  assign n17446 = n17445 ^ n17444;
  assign n17447 = n17299 ^ n16862;
  assign n17448 = n7515 & n11957;
  assign n17449 = n8029 & n11500;
  assign n17450 = n7518 & n11486;
  assign n17451 = n7520 & n11215;
  assign n17452 = ~n17450 & ~n17451;
  assign n17453 = ~n17449 & n17452;
  assign n17454 = ~n17448 & n17453;
  assign n17455 = n17454 ^ x5;
  assign n17456 = ~n17447 & n17455;
  assign n17457 = n17447 & ~n17455;
  assign n17466 = n17296 ^ n16872;
  assign n17458 = n7515 & n11704;
  assign n17459 = n8029 & n11486;
  assign n17460 = n7518 & n11215;
  assign n17461 = n7520 & ~n10956;
  assign n17462 = ~n17460 & ~n17461;
  assign n17463 = ~n17459 & n17462;
  assign n17464 = ~n17458 & n17463;
  assign n17465 = n17464 ^ x5;
  assign n17467 = n17466 ^ n17465;
  assign n17468 = n17293 ^ n16882;
  assign n17469 = n7515 & ~n12460;
  assign n17470 = n8029 & n11215;
  assign n17471 = n7520 & ~n10663;
  assign n17472 = n7518 & ~n10956;
  assign n17473 = ~n17471 & ~n17472;
  assign n17474 = ~n17470 & n17473;
  assign n17475 = ~n17469 & n17474;
  assign n17476 = n17475 ^ x5;
  assign n17477 = ~n17468 & n17476;
  assign n17486 = n17290 ^ n16892;
  assign n17478 = n7515 & ~n10957;
  assign n17479 = n7518 & ~n10663;
  assign n17480 = n8029 & ~n10956;
  assign n17481 = n7520 & n10665;
  assign n17482 = ~n17480 & ~n17481;
  assign n17483 = ~n17479 & n17482;
  assign n17484 = ~n17478 & n17483;
  assign n17485 = n17484 ^ x5;
  assign n17487 = n17486 ^ n17485;
  assign n17870 = n17287 ^ n16902;
  assign n17488 = n17284 ^ n16920;
  assign n17497 = n17281 ^ n16938;
  assign n17489 = n7515 & n12524;
  assign n17490 = n8029 & n10680;
  assign n17491 = n7518 & n10683;
  assign n17492 = n7520 & n10694;
  assign n17493 = ~n17491 & ~n17492;
  assign n17494 = ~n17490 & n17493;
  assign n17495 = ~n17489 & n17494;
  assign n17496 = n17495 ^ x5;
  assign n17498 = n17497 ^ n17496;
  assign n17500 = n7515 & n11599;
  assign n17501 = n8029 & n10683;
  assign n17502 = n7518 & n10694;
  assign n17503 = ~n17501 & ~n17502;
  assign n17504 = n7520 & n10698;
  assign n17505 = n17503 & ~n17504;
  assign n17506 = ~n17500 & n17505;
  assign n17507 = n17506 ^ x5;
  assign n17499 = n17278 ^ n16956;
  assign n17508 = n17507 ^ n17499;
  assign n17510 = n7515 & n12087;
  assign n17511 = n8029 & n10694;
  assign n17512 = n7520 & n10715;
  assign n17513 = n7518 & n10698;
  assign n17514 = ~n17512 & ~n17513;
  assign n17515 = ~n17511 & n17514;
  assign n17516 = ~n17510 & n17515;
  assign n17517 = n17516 ^ x5;
  assign n17509 = n17275 ^ n16974;
  assign n17518 = n17517 ^ n17509;
  assign n17527 = n17272 ^ n16984;
  assign n17519 = n7513 & n12033;
  assign n17520 = n17519 ^ n10698;
  assign n17521 = n7514 & n17520;
  assign n17522 = n7518 & n10715;
  assign n17523 = n7520 & n10718;
  assign n17524 = ~n17522 & ~n17523;
  assign n17525 = ~n17521 & n17524;
  assign n17526 = n17525 ^ x5;
  assign n17528 = n17527 ^ n17526;
  assign n17530 = n12111 & n17396;
  assign n17531 = n7520 & ~n10736;
  assign n17532 = n7518 & n10718;
  assign n17533 = ~n17531 & ~n17532;
  assign n17534 = x5 & n17533;
  assign n17535 = ~n10715 & n17534;
  assign n17536 = x4 & ~n17535;
  assign n17537 = ~n17530 & n17536;
  assign n17538 = ~n12111 & n17534;
  assign n17539 = n10715 & n17396;
  assign n17540 = ~x4 & ~n17539;
  assign n17541 = ~n17538 & n17540;
  assign n17542 = ~n17537 & ~n17541;
  assign n17543 = ~n17411 & n17533;
  assign n17544 = n17543 ^ x5;
  assign n17545 = ~n17542 & n17544;
  assign n17529 = n17269 ^ n17002;
  assign n17546 = n17545 ^ n17529;
  assign n17548 = n7515 & n12180;
  assign n17549 = n7518 & ~n10736;
  assign n17550 = n7520 & n10738;
  assign n17551 = ~n17549 & ~n17550;
  assign n17552 = n8029 & n10718;
  assign n17553 = n17551 & ~n17552;
  assign n17554 = ~n17548 & n17553;
  assign n17555 = n17554 ^ x5;
  assign n17547 = n17266 ^ n17012;
  assign n17556 = n17555 ^ n17547;
  assign n17558 = n7515 & ~n12596;
  assign n17559 = n8029 & ~n10736;
  assign n17560 = n7518 & n10738;
  assign n17561 = n7520 & n10740;
  assign n17562 = ~n17560 & ~n17561;
  assign n17563 = ~n17559 & n17562;
  assign n17564 = ~n17558 & n17563;
  assign n17565 = n17564 ^ x5;
  assign n17557 = n17263 ^ n17030;
  assign n17566 = n17565 ^ n17557;
  assign n17573 = n7515 & n12194;
  assign n17574 = n8029 & n10738;
  assign n17575 = n7518 & n10740;
  assign n17576 = n7520 & n10751;
  assign n17577 = ~n17575 & ~n17576;
  assign n17578 = ~n17574 & n17577;
  assign n17579 = ~n17573 & n17578;
  assign n17580 = n17579 ^ x5;
  assign n17571 = n17248 ^ n17247;
  assign n17567 = n17229 ^ x8;
  assign n17568 = n17567 ^ n17237;
  assign n17569 = ~n17256 & n17568;
  assign n17570 = n17569 ^ n17237;
  assign n17572 = n17571 ^ n17570;
  assign n17581 = n17580 ^ n17572;
  assign n17584 = n7515 & n13141;
  assign n17585 = n8029 & n10740;
  assign n17586 = n7518 & n10751;
  assign n17587 = n7520 & ~n10756;
  assign n17588 = ~n17586 & ~n17587;
  assign n17589 = ~n17585 & n17588;
  assign n17590 = ~n17584 & n17589;
  assign n17591 = n17590 ^ x5;
  assign n17582 = n17255 ^ x8;
  assign n17583 = n17582 ^ n17228;
  assign n17592 = n17591 ^ n17583;
  assign n17599 = n7515 & n12940;
  assign n17600 = n8029 & n10751;
  assign n17601 = n7518 & ~n10756;
  assign n17602 = n7520 & n10757;
  assign n17603 = ~n17601 & ~n17602;
  assign n17604 = ~n17600 & n17603;
  assign n17605 = ~n17599 & n17604;
  assign n17606 = n17605 ^ x5;
  assign n17597 = n17216 ^ n17209;
  assign n17593 = n17199 ^ n17031;
  assign n17594 = n17208 ^ n17031;
  assign n17595 = n17593 & ~n17594;
  assign n17596 = n17595 ^ n17207;
  assign n17598 = n17597 ^ n17596;
  assign n17607 = n17606 ^ n17598;
  assign n17609 = n7515 & ~n12703;
  assign n17610 = n8029 & ~n10756;
  assign n17611 = n7518 & n10757;
  assign n17612 = n7520 & n10773;
  assign n17613 = ~n17611 & ~n17612;
  assign n17614 = ~n17610 & n17613;
  assign n17615 = ~n17609 & n17614;
  assign n17616 = n17615 ^ x5;
  assign n17608 = n17593 ^ n17208;
  assign n17617 = n17616 ^ n17608;
  assign n17619 = n7515 & n12818;
  assign n17620 = n7518 & n10773;
  assign n17621 = n8029 & n10757;
  assign n17622 = ~n17620 & ~n17621;
  assign n17623 = n7520 & ~n10776;
  assign n17624 = n17622 & ~n17623;
  assign n17625 = ~n17619 & n17624;
  assign n17626 = n17625 ^ x5;
  assign n17618 = n17196 ^ n17041;
  assign n17627 = n17626 ^ n17618;
  assign n17629 = n7515 & n13155;
  assign n17630 = n8029 & n10773;
  assign n17631 = n7518 & ~n10776;
  assign n17632 = n7520 & ~n10777;
  assign n17633 = ~n17631 & ~n17632;
  assign n17634 = ~n17630 & n17633;
  assign n17635 = ~n17629 & n17634;
  assign n17636 = n17635 ^ x5;
  assign n17628 = n17193 ^ n17177;
  assign n17637 = n17636 ^ n17628;
  assign n17639 = n7515 & ~n13167;
  assign n17640 = n8029 & ~n10776;
  assign n17641 = n7520 & n10785;
  assign n17642 = n7518 & ~n10777;
  assign n17643 = ~n17641 & ~n17642;
  assign n17644 = ~n17640 & n17643;
  assign n17645 = ~n17639 & n17644;
  assign n17646 = n17645 ^ x5;
  assign n17638 = n17168 ^ n17052;
  assign n17647 = n17646 ^ n17638;
  assign n17649 = n7515 & ~n12832;
  assign n17650 = n8029 & ~n10777;
  assign n17651 = n7520 & ~n10789;
  assign n17652 = ~n17650 & ~n17651;
  assign n17653 = n7518 & n10785;
  assign n17654 = n17652 & ~n17653;
  assign n17655 = ~n17649 & n17654;
  assign n17656 = n17655 ^ x5;
  assign n17648 = n17165 ^ n17063;
  assign n17657 = n17656 ^ n17648;
  assign n17659 = n7515 & n13197;
  assign n17660 = n8029 & n10785;
  assign n17661 = n7518 & ~n10789;
  assign n17662 = n7520 & ~n10795;
  assign n17663 = ~n17661 & ~n17662;
  assign n17664 = ~n17660 & n17663;
  assign n17665 = ~n17659 & n17664;
  assign n17666 = n17665 ^ x5;
  assign n17658 = n17162 ^ n17073;
  assign n17667 = n17666 ^ n17658;
  assign n17668 = n17156 ^ n17140;
  assign n17670 = n7515 & ~n13278;
  assign n17671 = n8029 & ~n10799;
  assign n17672 = n7518 & ~n10800;
  assign n17673 = n7520 & n10815;
  assign n17674 = ~n17672 & ~n17673;
  assign n17675 = ~n17671 & n17674;
  assign n17676 = ~n17670 & n17675;
  assign n17677 = n17676 ^ x5;
  assign n17669 = n17124 ^ n17102;
  assign n17678 = n17677 ^ n17669;
  assign n17688 = n7515 & ~n13341;
  assign n17689 = n8029 & ~n10800;
  assign n17690 = n7520 & n10819;
  assign n17691 = ~n17689 & ~n17690;
  assign n17692 = n7518 & n10815;
  assign n17693 = n17691 & ~n17692;
  assign n17694 = ~n17688 & n17693;
  assign n17695 = n17694 ^ x5;
  assign n17679 = ~n5812 & ~n17112;
  assign n17682 = n17110 & ~n17113;
  assign n17680 = n5812 & ~n6315;
  assign n17681 = n17110 & n17680;
  assign n17683 = n17682 ^ n17681;
  assign n17684 = n10825 & ~n17683;
  assign n17685 = n17684 ^ n17682;
  assign n17686 = ~n17679 & n17685;
  assign n17687 = n17686 ^ n17123;
  assign n17696 = n17695 ^ n17687;
  assign n17710 = n7515 & n13387;
  assign n17711 = n8029 & n10815;
  assign n17712 = n7518 & n10819;
  assign n17713 = n7520 & ~n10820;
  assign n17714 = ~n17712 & ~n17713;
  assign n17715 = ~n17711 & n17714;
  assign n17716 = ~n17710 & n17715;
  assign n17717 = n17716 ^ x5;
  assign n17697 = n17111 ^ n6305;
  assign n17698 = n10822 & n17697;
  assign n17699 = n17698 ^ n6305;
  assign n17700 = n17110 & n17699;
  assign n17701 = ~x8 & n6309;
  assign n17702 = ~n10822 & n17701;
  assign n17703 = ~n17700 & ~n17702;
  assign n17704 = n6309 & n13532;
  assign n17705 = n17109 & ~n17704;
  assign n17706 = x8 & n6305;
  assign n17707 = ~n14128 & n17706;
  assign n17708 = ~n17705 & ~n17707;
  assign n17709 = n17703 & ~n17708;
  assign n17718 = n17717 ^ n17709;
  assign n17727 = n7515 & n13429;
  assign n17728 = n8029 & n10819;
  assign n17729 = n7518 & ~n10820;
  assign n17730 = n7520 & n10821;
  assign n17731 = ~n17729 & ~n17730;
  assign n17732 = ~n17728 & n17731;
  assign n17733 = ~n17727 & n17732;
  assign n17734 = n17733 ^ x5;
  assign n17719 = ~n6313 & ~n10822;
  assign n17720 = n9197 & ~n17719;
  assign n17721 = ~n9195 & ~n17720;
  assign n17722 = n10825 & ~n17721;
  assign n17723 = x7 & n10825;
  assign n17724 = n6305 & ~n17723;
  assign n17725 = ~n10822 & n17724;
  assign n17726 = ~n17722 & ~n17725;
  assign n17735 = n17734 ^ n17726;
  assign n17736 = n7515 & ~n14111;
  assign n17737 = n8029 & ~n10820;
  assign n17738 = n7518 & n10821;
  assign n17739 = n7520 & ~n10822;
  assign n17740 = ~n17738 & ~n17739;
  assign n17741 = ~n17737 & n17740;
  assign n17742 = ~n17736 & n17741;
  assign n17743 = n7514 & ~n13532;
  assign n17744 = ~n8029 & ~n17743;
  assign n17745 = n10821 & ~n17744;
  assign n17746 = n7518 & ~n10822;
  assign n17747 = n7520 & n10825;
  assign n17748 = ~n17746 & ~n17747;
  assign n17749 = ~n17745 & n17748;
  assign n17750 = n7515 & n13533;
  assign n17751 = n17749 & ~n17750;
  assign n17752 = n7514 & ~n10822;
  assign n17753 = ~n7519 & n10825;
  assign n17754 = ~n17752 & ~n17753;
  assign n17755 = x5 & n17754;
  assign n17756 = n17751 & n17755;
  assign n17757 = ~n17742 & ~n17756;
  assign n17758 = n9236 & ~n17757;
  assign n17759 = n9220 & ~n17742;
  assign n17760 = ~n17758 & ~n17759;
  assign n17761 = n10825 & ~n17760;
  assign n17762 = n17742 & n17756;
  assign n17763 = ~n17761 & ~n17762;
  assign n17764 = n17763 ^ n17734;
  assign n17765 = ~n17735 & n17764;
  assign n17766 = n17765 ^ n17763;
  assign n17767 = n17766 ^ n17709;
  assign n17768 = n17718 & ~n17767;
  assign n17769 = n17768 ^ n17717;
  assign n17770 = n17769 ^ n17687;
  assign n17771 = n17696 & ~n17770;
  assign n17772 = n17771 ^ n17695;
  assign n17773 = n17772 ^ n17677;
  assign n17774 = n17678 & n17773;
  assign n17775 = n17774 ^ n17772;
  assign n17776 = ~n17668 & n17775;
  assign n17777 = n7515 & ~n13239;
  assign n17778 = n8029 & ~n10795;
  assign n17779 = n7518 & ~n10799;
  assign n17780 = n7520 & ~n10800;
  assign n17781 = ~n17779 & ~n17780;
  assign n17782 = ~n17778 & n17781;
  assign n17783 = ~n17777 & n17782;
  assign n17784 = n17783 ^ x5;
  assign n17785 = n17775 & n17784;
  assign n17786 = ~n17776 & ~n17785;
  assign n17787 = n7515 & ~n13224;
  assign n17788 = n8029 & ~n10789;
  assign n17789 = n7520 & ~n10799;
  assign n17790 = ~n17788 & ~n17789;
  assign n17791 = n7518 & ~n10795;
  assign n17792 = n17790 & ~n17791;
  assign n17793 = ~n17787 & n17792;
  assign n17794 = n17159 ^ n17084;
  assign n17795 = n17793 & n17794;
  assign n17796 = ~n17668 & n17783;
  assign n17797 = ~n17795 & ~n17796;
  assign n17798 = n17786 & n17797;
  assign n17799 = ~n17793 & ~n17794;
  assign n17800 = ~x5 & ~n17799;
  assign n17801 = ~n17798 & n17800;
  assign n17802 = ~n17793 & n17794;
  assign n17803 = ~n17668 & ~n17783;
  assign n17804 = ~n17802 & ~n17803;
  assign n17805 = n17786 & n17804;
  assign n17806 = n17793 & ~n17794;
  assign n17807 = x5 & ~n17806;
  assign n17808 = ~n17805 & n17807;
  assign n17809 = ~n17801 & ~n17808;
  assign n17810 = n17809 ^ n17658;
  assign n17811 = ~n17667 & ~n17810;
  assign n17812 = n17811 ^ n17666;
  assign n17813 = n17812 ^ n17648;
  assign n17814 = ~n17657 & n17813;
  assign n17815 = n17814 ^ n17656;
  assign n17816 = n17815 ^ n17646;
  assign n17817 = ~n17647 & n17816;
  assign n17818 = n17817 ^ n17815;
  assign n17819 = n17818 ^ n17628;
  assign n17820 = ~n17637 & n17819;
  assign n17821 = n17820 ^ n17636;
  assign n17822 = n17821 ^ n17618;
  assign n17823 = ~n17627 & n17822;
  assign n17824 = n17823 ^ n17626;
  assign n17825 = n17824 ^ n17616;
  assign n17826 = n17617 & n17825;
  assign n17827 = n17826 ^ n17824;
  assign n17828 = n17827 ^ n17606;
  assign n17829 = n17607 & n17828;
  assign n17830 = n17829 ^ n17827;
  assign n17831 = n17830 ^ n17591;
  assign n17832 = ~n17592 & n17831;
  assign n17833 = n17832 ^ n17830;
  assign n17834 = n17833 ^ n17580;
  assign n17835 = ~n17581 & n17834;
  assign n17836 = n17835 ^ n17833;
  assign n17837 = n17836 ^ n17565;
  assign n17838 = ~n17566 & n17837;
  assign n17839 = n17838 ^ n17836;
  assign n17840 = n17839 ^ n17555;
  assign n17841 = n17556 & n17840;
  assign n17842 = n17841 ^ n17839;
  assign n17843 = n17842 ^ n17529;
  assign n17844 = ~n17546 & n17843;
  assign n17845 = n17844 ^ n17545;
  assign n17846 = n17845 ^ n17527;
  assign n17847 = n17528 & ~n17846;
  assign n17848 = n17847 ^ n17845;
  assign n17849 = n17848 ^ n17517;
  assign n17850 = ~n17518 & n17849;
  assign n17851 = n17850 ^ n17848;
  assign n17852 = n17851 ^ n17507;
  assign n17853 = ~n17508 & n17852;
  assign n17854 = n17853 ^ n17851;
  assign n17855 = n17854 ^ n17497;
  assign n17856 = n17498 & ~n17855;
  assign n17857 = n17856 ^ n17854;
  assign n17858 = ~n17488 & ~n17857;
  assign n17859 = n17488 & n17857;
  assign n17860 = n7515 & n12100;
  assign n17861 = n7518 & n10680;
  assign n17862 = n7520 & n10683;
  assign n17863 = ~n17861 & ~n17862;
  assign n17864 = n8029 & n10665;
  assign n17865 = n17863 & ~n17864;
  assign n17866 = ~n17860 & n17865;
  assign n17867 = n17866 ^ x5;
  assign n17868 = ~n17859 & ~n17867;
  assign n17869 = ~n17858 & ~n17868;
  assign n17871 = n17870 ^ n17869;
  assign n17872 = n7515 & ~n11694;
  assign n17873 = n8029 & ~n10663;
  assign n17874 = n7520 & n10680;
  assign n17875 = n7518 & n10665;
  assign n17876 = ~n17874 & ~n17875;
  assign n17877 = ~n17873 & n17876;
  assign n17878 = ~n17872 & n17877;
  assign n17879 = n17878 ^ x5;
  assign n17880 = n17879 ^ n17869;
  assign n17881 = ~n17871 & ~n17880;
  assign n17882 = n17881 ^ n17870;
  assign n17883 = n17882 ^ n17486;
  assign n17884 = n17487 & n17883;
  assign n17885 = n17884 ^ n17882;
  assign n17886 = ~n17477 & n17885;
  assign n17887 = n17468 & ~n17476;
  assign n17888 = ~n17886 & ~n17887;
  assign n17889 = n17888 ^ n17466;
  assign n17890 = n17467 & ~n17889;
  assign n17891 = n17890 ^ n17888;
  assign n17892 = ~n17457 & n17891;
  assign n17893 = ~n17456 & ~n17892;
  assign n17894 = n17893 ^ n17444;
  assign n17895 = ~n17446 & n17894;
  assign n17896 = n17895 ^ n17445;
  assign n17897 = n17896 ^ n17435;
  assign n17898 = ~n17436 & ~n17897;
  assign n17899 = n17898 ^ n17896;
  assign n17900 = n17899 ^ n17425;
  assign n17901 = n17426 & n17900;
  assign n17902 = n17901 ^ n17899;
  assign n17903 = n17902 ^ n17415;
  assign n17904 = ~n17416 & ~n17903;
  assign n17905 = n17904 ^ n17902;
  assign n17916 = n17915 ^ n17905;
  assign n17394 = n9380 & n12019;
  assign n17395 = ~n12750 & ~n17394;
  assign n17917 = n17916 ^ n17395;
  assign n17928 = n17902 ^ n17416;
  assign n17918 = x2 & n17383;
  assign n17919 = x0 & ~n17918;
  assign n17920 = x1 & ~n17383;
  assign n17921 = n17919 & ~n17920;
  assign n17922 = x2 & n11940;
  assign n17923 = n9448 & n17922;
  assign n17924 = n12019 ^ x2;
  assign n17925 = n9378 & ~n17924;
  assign n17926 = ~n17923 & ~n17925;
  assign n17927 = ~n17921 & n17926;
  assign n17929 = n17928 ^ n17927;
  assign n17931 = n33 & ~n12013;
  assign n17932 = n17931 ^ x1;
  assign n17933 = ~n12019 & ~n17932;
  assign n17934 = x2 & n12019;
  assign n17935 = x0 & ~n17934;
  assign n17936 = ~n17933 & n17935;
  assign n17937 = n11940 ^ x2;
  assign n17938 = x1 & ~n17937;
  assign n17939 = n9346 & ~n11902;
  assign n17940 = ~x0 & ~n17939;
  assign n17941 = ~n17938 & n17940;
  assign n17942 = ~n17936 & ~n17941;
  assign n17930 = n17899 ^ n17426;
  assign n17943 = n17942 ^ n17930;
  assign n17944 = n33 & ~n11999;
  assign n17945 = n17944 ^ x1;
  assign n17946 = n17945 ^ n11875;
  assign n17947 = x0 & n17946;
  assign n17948 = n11773 ^ x2;
  assign n17949 = n9378 & n17948;
  assign n17950 = x2 & ~n11480;
  assign n17951 = n9448 & ~n17950;
  assign n17952 = ~n17949 & ~n17951;
  assign n17953 = ~n17947 & n17952;
  assign n18464 = n33 & ~n11776;
  assign n18465 = n18464 ^ x1;
  assign n18466 = n18465 ^ n11773;
  assign n18467 = x0 & n18466;
  assign n18468 = x2 & ~n11500;
  assign n18469 = n9448 & ~n18468;
  assign n18470 = n11480 ^ x2;
  assign n18471 = n9378 & ~n18470;
  assign n18472 = ~n18469 & ~n18471;
  assign n18473 = ~n18467 & n18472;
  assign n17964 = n17476 ^ n17468;
  assign n17965 = n17964 ^ n17885;
  assign n17954 = n33 & ~n11506;
  assign n17955 = n17954 ^ x1;
  assign n17956 = n17955 ^ n11480;
  assign n17957 = x0 & ~n17956;
  assign n17958 = n11500 ^ x2;
  assign n17959 = n9378 & ~n17958;
  assign n17960 = x2 & ~n11486;
  assign n17961 = n9448 & ~n17960;
  assign n17962 = ~n17959 & ~n17961;
  assign n17963 = ~n17957 & n17962;
  assign n17966 = n17965 ^ n17963;
  assign n17968 = n33 & ~n11956;
  assign n17969 = n17968 ^ x1;
  assign n17970 = n17969 ^ n11500;
  assign n17971 = x0 & n17970;
  assign n17972 = n11486 ^ x2;
  assign n17973 = n9378 & n17972;
  assign n17974 = x2 & ~n11215;
  assign n17975 = n9448 & n17974;
  assign n17976 = ~n17973 & ~n17975;
  assign n17977 = ~n17971 & n17976;
  assign n17967 = n17882 ^ n17487;
  assign n17978 = n17977 ^ n17967;
  assign n17986 = n33 & ~n11703;
  assign n17987 = n17986 ^ x1;
  assign n17988 = n17987 ^ n11486;
  assign n17989 = x0 & ~n17988;
  assign n17990 = n11215 ^ x2;
  assign n17991 = n9378 & ~n17990;
  assign n17992 = x2 & n10956;
  assign n17993 = n9448 & ~n17992;
  assign n17994 = ~n17991 & ~n17993;
  assign n17995 = ~n17989 & n17994;
  assign n17984 = n17878 ^ n17870;
  assign n17979 = n17857 ^ n17488;
  assign n17980 = n17488 ^ x5;
  assign n17981 = n17980 ^ n17866;
  assign n17982 = ~n17979 & n17981;
  assign n17983 = n17982 ^ n17866;
  assign n17985 = n17984 ^ n17983;
  assign n17996 = n17995 ^ n17985;
  assign n18008 = n17854 ^ n17498;
  assign n18014 = n33 & ~n10880;
  assign n18015 = n18014 ^ x1;
  assign n18016 = n18015 ^ n10956;
  assign n18010 = n10663 ^ x2;
  assign n18009 = x2 & ~n10665;
  assign n18011 = n18010 ^ n18009;
  assign n18012 = ~x1 & ~n18011;
  assign n18013 = n18012 ^ n18010;
  assign n18017 = n18016 ^ n18013;
  assign n18018 = ~x0 & n18017;
  assign n18019 = n18018 ^ n18016;
  assign n18020 = n18008 & ~n18019;
  assign n18021 = n33 & ~n11693;
  assign n18022 = n18021 ^ x1;
  assign n18023 = n18022 ^ n10663;
  assign n18024 = x0 & ~n18023;
  assign n18025 = n10665 ^ x2;
  assign n18026 = x1 & ~n18025;
  assign n18027 = n9431 & ~n10680;
  assign n18028 = ~n9378 & ~n18027;
  assign n18029 = ~n18026 & ~n18028;
  assign n18030 = ~n18024 & ~n18029;
  assign n18031 = n17851 ^ n17508;
  assign n18032 = ~n18030 & ~n18031;
  assign n18033 = ~n18020 & ~n18032;
  assign n18034 = n17848 ^ n17518;
  assign n18039 = n33 & ~n12099;
  assign n18040 = n18039 ^ x1;
  assign n18041 = n18040 ^ n10665;
  assign n18035 = n10680 ^ x2;
  assign n18036 = x1 & n18035;
  assign n18037 = n9346 & ~n10683;
  assign n18038 = ~n18036 & ~n18037;
  assign n18042 = n18041 ^ n18038;
  assign n18043 = ~x0 & ~n18042;
  assign n18044 = n18043 ^ n18041;
  assign n18045 = ~n18034 & n18044;
  assign n18427 = n33 & ~n11616;
  assign n18428 = n18427 ^ x1;
  assign n18429 = n18428 ^ n10680;
  assign n18430 = x0 & ~n18429;
  assign n18431 = x2 & ~n10694;
  assign n18432 = n9448 & ~n18431;
  assign n18433 = n10683 ^ x2;
  assign n18434 = n9378 & ~n18433;
  assign n18435 = ~n18432 & ~n18434;
  assign n18436 = ~n18430 & n18435;
  assign n18056 = n33 & ~n12033;
  assign n18057 = n18056 ^ x1;
  assign n18058 = n18057 ^ n10698;
  assign n18059 = x0 & ~n18058;
  assign n18060 = n10715 ^ x2;
  assign n18061 = x1 & n18060;
  assign n18062 = x2 & ~n10718;
  assign n18063 = ~x0 & ~n18062;
  assign n18064 = ~n9378 & ~n18063;
  assign n18065 = ~n18061 & ~n18064;
  assign n18066 = ~n18059 & ~n18065;
  assign n18067 = n17836 ^ n17566;
  assign n18068 = ~n18066 & n18067;
  assign n18079 = n33 & ~n12595;
  assign n18080 = n18079 ^ x1;
  assign n18081 = n18080 ^ n10736;
  assign n18082 = x0 & n18081;
  assign n18083 = n10738 ^ x2;
  assign n18084 = x1 & n18083;
  assign n18085 = x2 & ~n10740;
  assign n18086 = ~x0 & ~n18085;
  assign n18087 = ~n9378 & ~n18086;
  assign n18088 = ~n18084 & ~n18087;
  assign n18089 = ~n18082 & ~n18088;
  assign n18365 = n33 & ~n12193;
  assign n18366 = n18365 ^ x1;
  assign n18367 = n18366 ^ n10738;
  assign n18368 = x0 & ~n18367;
  assign n18351 = n10740 ^ x2;
  assign n18369 = n9378 & ~n18351;
  assign n18370 = x2 & ~n10751;
  assign n18371 = n9448 & ~n18370;
  assign n18372 = ~n18369 & ~n18371;
  assign n18373 = ~n18368 & n18372;
  assign n18348 = n10740 ^ x1;
  assign n18349 = n13140 & n18348;
  assign n18350 = x0 & ~n18349;
  assign n18352 = ~n13140 & n18351;
  assign n18353 = n18350 & ~n18352;
  assign n18354 = x2 & n10756;
  assign n18355 = n9448 & ~n18354;
  assign n18356 = n10751 ^ x2;
  assign n18357 = n9378 & ~n18356;
  assign n18358 = ~n18355 & ~n18357;
  assign n18359 = ~n18353 & n18358;
  assign n18324 = ~x2 & n10751;
  assign n18325 = x0 & n18324;
  assign n18330 = n10866 & n18325;
  assign n18331 = n10756 ^ x2;
  assign n18332 = ~x0 & ~n18331;
  assign n18333 = ~n18330 & ~n18332;
  assign n18334 = x0 & ~n10751;
  assign n18335 = ~x2 & ~n12939;
  assign n18336 = n18334 & ~n18335;
  assign n18337 = n18333 & ~n18336;
  assign n18338 = n10841 & n18324;
  assign n18339 = n18337 & ~n18338;
  assign n18326 = n8890 & ~n12940;
  assign n18327 = ~n18325 & ~n18326;
  assign n18328 = n9431 & ~n10757;
  assign n18329 = n18327 & ~n18328;
  assign n18340 = n18339 ^ n18329;
  assign n18341 = ~x1 & n18340;
  assign n18342 = n18341 ^ n18339;
  assign n18309 = n33 & ~n12702;
  assign n18310 = n18309 ^ x1;
  assign n18311 = n18310 ^ n10756;
  assign n18312 = x0 & n18311;
  assign n18313 = n10757 ^ x2;
  assign n18314 = x1 & n18313;
  assign n18315 = n9346 & ~n10773;
  assign n18316 = ~x0 & ~n18315;
  assign n18317 = ~n18314 & n18316;
  assign n18318 = ~n18312 & ~n18317;
  assign n18101 = n17812 ^ n17657;
  assign n18095 = n33 & ~n12817;
  assign n18096 = n18095 ^ x1;
  assign n18097 = n18096 ^ n10757;
  assign n18091 = n10773 ^ x2;
  assign n18090 = x2 & n10776;
  assign n18092 = n18091 ^ n18090;
  assign n18093 = ~x1 & n18092;
  assign n18094 = n18093 ^ n18091;
  assign n18098 = n18097 ^ n18094;
  assign n18099 = ~x0 & n18098;
  assign n18100 = n18099 ^ n18097;
  assign n18102 = n18101 ^ n18100;
  assign n18291 = n33 & ~n13154;
  assign n18292 = n18291 ^ x1;
  assign n18293 = n18292 ^ n10773;
  assign n18294 = x0 & ~n18293;
  assign n18295 = n10776 ^ x2;
  assign n18296 = n9378 & n18295;
  assign n18297 = x2 & n10777;
  assign n18298 = n9448 & ~n18297;
  assign n18299 = ~n18296 & ~n18298;
  assign n18300 = ~n18294 & n18299;
  assign n18271 = n33 & ~n13166;
  assign n18272 = n18271 ^ x1;
  assign n18273 = n18272 ^ n10776;
  assign n18274 = x0 & n18273;
  assign n18275 = x2 & ~n10785;
  assign n18276 = n9448 & ~n18275;
  assign n18277 = n10777 ^ x2;
  assign n18278 = n9378 & n18277;
  assign n18279 = ~n18276 & ~n18278;
  assign n18280 = ~n18274 & n18279;
  assign n18105 = n33 & ~n12831;
  assign n18106 = n18105 ^ x1;
  assign n18107 = n18106 ^ n10777;
  assign n18108 = x0 & ~n18107;
  assign n18109 = n10785 ^ x2;
  assign n18110 = n9378 & n18109;
  assign n18111 = x2 & n10789;
  assign n18112 = n9448 & n18111;
  assign n18113 = ~n18110 & ~n18112;
  assign n18114 = ~n18108 & n18113;
  assign n18103 = n17775 ^ n17668;
  assign n18104 = n18103 ^ n17784;
  assign n18115 = n18114 ^ n18104;
  assign n18126 = ~x1 & n10799;
  assign n18127 = ~n10800 & n18126;
  assign n18128 = ~x2 & ~n10799;
  assign n18129 = ~n10831 & ~n10855;
  assign n18130 = n18128 & ~n18129;
  assign n18131 = ~n18127 & ~n18130;
  assign n18132 = n10815 & n18131;
  assign n18133 = n10799 & n18129;
  assign n18134 = ~x2 & n18133;
  assign n18135 = ~x1 & n10800;
  assign n18136 = ~n10799 & n18135;
  assign n18137 = ~n10815 & ~n18136;
  assign n18138 = ~n18134 & n18137;
  assign n18139 = ~n18132 & ~n18138;
  assign n18140 = n10800 ^ n10799;
  assign n18141 = ~x2 & ~n18140;
  assign n18142 = n18129 ^ n10800;
  assign n18143 = n18140 & ~n18142;
  assign n18144 = ~x1 & n18143;
  assign n18145 = ~n18141 & ~n18144;
  assign n18146 = ~n18139 & n18145;
  assign n18147 = n18146 ^ n10795;
  assign n18148 = x0 & n18147;
  assign n18149 = n10799 ^ x2;
  assign n18150 = n9378 & n18149;
  assign n18151 = x2 & n10800;
  assign n18152 = n9448 & ~n18151;
  assign n18153 = ~n18150 & ~n18152;
  assign n18154 = ~n18148 & n18153;
  assign n18155 = n17766 ^ n17718;
  assign n18156 = n18154 & ~n18155;
  assign n18157 = n33 & ~n13277;
  assign n18158 = n18157 ^ x1;
  assign n18159 = n18158 ^ n10799;
  assign n18160 = x0 & ~n18159;
  assign n18161 = x2 & ~n10815;
  assign n18162 = n9448 & n18161;
  assign n18163 = n10800 ^ x2;
  assign n18164 = n9378 & ~n18163;
  assign n18165 = ~n18162 & ~n18164;
  assign n18166 = ~n18160 & n18165;
  assign n18177 = ~x6 & n10825;
  assign n18178 = n18177 ^ n17756;
  assign n18179 = ~x5 & ~n10825;
  assign n18180 = ~n18178 & ~n18179;
  assign n18181 = n18180 ^ n17742;
  assign n18171 = n33 & ~n13340;
  assign n18172 = n18171 ^ x1;
  assign n18173 = n18172 ^ n10800;
  assign n18167 = n10815 ^ x2;
  assign n18168 = x1 & n18167;
  assign n18169 = n9346 & ~n10819;
  assign n18170 = ~n18168 & ~n18169;
  assign n18174 = n18173 ^ n18170;
  assign n18175 = ~x0 & n18174;
  assign n18176 = n18175 ^ n18173;
  assign n18182 = n18181 ^ n18176;
  assign n18185 = n33 & ~n13386;
  assign n18186 = n18185 ^ x1;
  assign n18187 = n18186 ^ n10815;
  assign n18188 = x0 & ~n18187;
  assign n18189 = n10819 ^ x2;
  assign n18190 = x1 & n18189;
  assign n18191 = n9346 & n10820;
  assign n18192 = ~x0 & ~n18191;
  assign n18193 = ~n18190 & n18192;
  assign n18194 = ~n18188 & ~n18193;
  assign n18183 = x5 & ~n17754;
  assign n18184 = n18183 ^ n17751;
  assign n18195 = n18194 ^ n18184;
  assign n18196 = x2 & ~n10821;
  assign n18197 = ~n9431 & ~n18196;
  assign n18198 = ~n9448 & n13532;
  assign n18199 = n18198 ^ n10825;
  assign n18200 = ~n18197 & ~n18199;
  assign n18201 = n7514 & n10825;
  assign n18202 = ~n18200 & ~n18201;
  assign n18207 = n33 & ~n14110;
  assign n18208 = n18207 ^ x1;
  assign n18209 = n18208 ^ n10820;
  assign n18203 = n10821 ^ x2;
  assign n18204 = x1 & n18203;
  assign n18205 = n9346 & n10822;
  assign n18206 = ~n18204 & ~n18205;
  assign n18210 = n18209 ^ n18206;
  assign n18211 = ~x0 & n18210;
  assign n18212 = n18211 ^ n18209;
  assign n18213 = ~n18202 & ~n18212;
  assign n18214 = ~n9530 & ~n10822;
  assign n18215 = n9532 & ~n18214;
  assign n18216 = ~n9529 & ~n18215;
  assign n18217 = n10825 & ~n18216;
  assign n18218 = x4 & n10825;
  assign n18219 = n17752 & ~n18218;
  assign n18220 = ~n18217 & ~n18219;
  assign n18221 = ~n18213 & n18220;
  assign n18222 = n33 & ~n13428;
  assign n18223 = n18222 ^ x1;
  assign n18224 = n18223 ^ n10819;
  assign n18225 = x0 & ~n18224;
  assign n18226 = ~n18221 & ~n18225;
  assign n18227 = n10820 ^ x2;
  assign n18228 = n18227 ^ n18196;
  assign n18229 = x1 & ~n18228;
  assign n18230 = n18229 ^ n18196;
  assign n18231 = ~x0 & ~n18230;
  assign n18232 = n18226 & ~n18231;
  assign n18233 = n18213 & ~n18220;
  assign n18234 = ~n18232 & ~n18233;
  assign n18235 = n18234 ^ n18184;
  assign n18236 = ~n18195 & ~n18235;
  assign n18237 = n18236 ^ n18194;
  assign n18238 = n18237 ^ n18181;
  assign n18239 = n18182 & n18238;
  assign n18240 = n18239 ^ n18176;
  assign n18241 = ~n18166 & ~n18240;
  assign n18242 = ~n18156 & ~n18241;
  assign n18243 = n18166 & n18240;
  assign n18244 = n17763 ^ n17735;
  assign n18245 = ~n18243 & ~n18244;
  assign n18246 = n18242 & ~n18245;
  assign n18247 = n33 & ~n13223;
  assign n18248 = n18247 ^ x1;
  assign n18249 = n18248 ^ n10789;
  assign n18250 = x0 & ~n18249;
  assign n18251 = n10795 ^ x2;
  assign n18252 = n9378 & ~n18251;
  assign n18253 = n9431 & n18126;
  assign n18254 = ~n18252 & ~n18253;
  assign n18255 = ~n18250 & n18254;
  assign n18256 = n17769 ^ n17696;
  assign n18257 = n18255 & n18256;
  assign n18258 = ~n18154 & n18155;
  assign n18259 = ~n18257 & ~n18258;
  assign n18260 = ~n18246 & n18259;
  assign n18261 = ~n18255 & ~n18256;
  assign n18262 = ~n18260 & ~n18261;
  assign n18116 = n33 & ~n13196;
  assign n18117 = n18116 ^ x1;
  assign n18118 = n18117 ^ n10785;
  assign n18119 = x0 & ~n18118;
  assign n18120 = x2 & n10795;
  assign n18121 = n9448 & ~n18120;
  assign n18122 = n10789 ^ x2;
  assign n18123 = n9378 & n18122;
  assign n18124 = ~n18121 & ~n18123;
  assign n18125 = ~n18119 & n18124;
  assign n18263 = n18262 ^ n18125;
  assign n18264 = n17772 ^ n17678;
  assign n18265 = n18264 ^ n18125;
  assign n18266 = ~n18263 & ~n18265;
  assign n18267 = n18266 ^ n18262;
  assign n18268 = n18267 ^ n18104;
  assign n18269 = ~n18115 & n18268;
  assign n18270 = n18269 ^ n18114;
  assign n18281 = n18280 ^ n18270;
  assign n18286 = n17794 ^ n17793;
  assign n18282 = n17668 ^ x5;
  assign n18283 = n18282 ^ n17783;
  assign n18284 = n18103 & ~n18283;
  assign n18285 = n18284 ^ n17783;
  assign n18287 = n18286 ^ n18285;
  assign n18288 = n18287 ^ n18280;
  assign n18289 = ~n18281 & n18288;
  assign n18290 = n18289 ^ n18270;
  assign n18301 = n18300 ^ n18290;
  assign n18302 = n17809 ^ n17667;
  assign n18303 = n18302 ^ n18300;
  assign n18304 = ~n18301 & n18303;
  assign n18305 = n18304 ^ n18290;
  assign n18306 = n18305 ^ n18101;
  assign n18307 = n18102 & n18306;
  assign n18308 = n18307 ^ n18100;
  assign n18319 = n18318 ^ n18308;
  assign n18320 = n17815 ^ n17647;
  assign n18321 = n18320 ^ n18318;
  assign n18322 = n18319 & n18321;
  assign n18323 = n18322 ^ n18308;
  assign n18343 = n18342 ^ n18323;
  assign n18344 = n17818 ^ n17637;
  assign n18345 = n18344 ^ n18323;
  assign n18346 = ~n18343 & ~n18345;
  assign n18347 = n18346 ^ n18342;
  assign n18360 = n18359 ^ n18347;
  assign n18361 = n17821 ^ n17627;
  assign n18362 = n18361 ^ n18359;
  assign n18363 = ~n18360 & ~n18362;
  assign n18364 = n18363 ^ n18347;
  assign n18374 = n18373 ^ n18364;
  assign n18375 = n17824 ^ n17617;
  assign n18376 = n18375 ^ n18373;
  assign n18377 = ~n18374 & ~n18376;
  assign n18378 = n18377 ^ n18364;
  assign n18379 = n18089 & ~n18378;
  assign n18380 = n17827 ^ n17607;
  assign n18381 = ~n18379 & ~n18380;
  assign n18382 = ~n18089 & n18378;
  assign n18383 = n33 & ~n12179;
  assign n18384 = n18383 ^ x1;
  assign n18385 = n18384 ^ n10718;
  assign n18386 = x0 & ~n18385;
  assign n18387 = n10736 ^ x2;
  assign n18388 = x1 & ~n18387;
  assign n18389 = n9346 & ~n10738;
  assign n18390 = ~x0 & ~n18389;
  assign n18391 = ~n18388 & n18390;
  assign n18392 = ~n18386 & ~n18391;
  assign n18393 = n17830 ^ n17592;
  assign n18394 = ~n18392 & n18393;
  assign n18395 = ~n18382 & ~n18394;
  assign n18396 = ~n18381 & n18395;
  assign n18397 = n18392 & ~n18393;
  assign n18398 = ~n18396 & ~n18397;
  assign n18073 = n33 & ~n12110;
  assign n18074 = n18073 ^ x1;
  assign n18075 = n18074 ^ n10715;
  assign n18069 = n10718 ^ x2;
  assign n18070 = x1 & n18069;
  assign n18071 = n9346 & n10736;
  assign n18072 = ~n18070 & ~n18071;
  assign n18076 = n18075 ^ n18072;
  assign n18077 = ~x0 & ~n18076;
  assign n18078 = n18077 ^ n18075;
  assign n18399 = n18398 ^ n18078;
  assign n18400 = n17833 ^ n17581;
  assign n18401 = n18400 ^ n18078;
  assign n18402 = ~n18399 & n18401;
  assign n18403 = n18402 ^ n18398;
  assign n18404 = ~n18068 & ~n18403;
  assign n18405 = n17839 ^ n17556;
  assign n18410 = n33 & ~n12086;
  assign n18411 = n18410 ^ x1;
  assign n18412 = n18411 ^ n10694;
  assign n18406 = n10698 ^ x2;
  assign n18407 = x1 & n18406;
  assign n18408 = n9346 & ~n10715;
  assign n18409 = ~n18407 & ~n18408;
  assign n18413 = n18412 ^ n18409;
  assign n18414 = ~x0 & ~n18413;
  assign n18415 = n18414 ^ n18412;
  assign n18416 = n18405 & n18415;
  assign n18417 = n18066 & ~n18067;
  assign n18418 = ~n18416 & ~n18417;
  assign n18419 = ~n18404 & n18418;
  assign n18420 = ~n18405 & ~n18415;
  assign n18421 = ~n18419 & ~n18420;
  assign n18046 = n33 & ~n11598;
  assign n18047 = n18046 ^ x1;
  assign n18048 = n18047 ^ n10683;
  assign n18049 = x0 & ~n18048;
  assign n18050 = n10694 ^ x2;
  assign n18051 = x1 & n18050;
  assign n18052 = n9346 & ~n10698;
  assign n18053 = ~x0 & ~n18052;
  assign n18054 = ~n18051 & n18053;
  assign n18055 = ~n18049 & ~n18054;
  assign n18422 = n18421 ^ n18055;
  assign n18423 = n17842 ^ n17546;
  assign n18424 = n18423 ^ n18055;
  assign n18425 = n18422 & ~n18424;
  assign n18426 = n18425 ^ n18421;
  assign n18437 = n18436 ^ n18426;
  assign n18438 = n17845 ^ n17528;
  assign n18439 = n18438 ^ n18436;
  assign n18440 = n18437 & ~n18439;
  assign n18441 = n18440 ^ n18426;
  assign n18442 = ~n18045 & ~n18441;
  assign n18443 = n18030 & n18031;
  assign n18444 = n18034 & ~n18044;
  assign n18445 = ~n18443 & ~n18444;
  assign n18446 = ~n18442 & n18445;
  assign n18447 = n18033 & ~n18446;
  assign n18448 = ~n18008 & n18019;
  assign n18449 = ~n18447 & ~n18448;
  assign n17997 = n11226 ^ n10956;
  assign n17998 = n33 & n17997;
  assign n17999 = n17998 ^ x1;
  assign n18000 = n17999 ^ n11215;
  assign n18001 = x0 & n18000;
  assign n18002 = x2 & n10663;
  assign n18003 = n9448 & n18002;
  assign n18004 = n10956 ^ x2;
  assign n18005 = n9378 & ~n18004;
  assign n18006 = ~n18003 & ~n18005;
  assign n18007 = ~n18001 & n18006;
  assign n18450 = n18449 ^ n18007;
  assign n18451 = n17979 ^ n17867;
  assign n18452 = n18451 ^ n18007;
  assign n18453 = ~n18450 & ~n18452;
  assign n18454 = n18453 ^ n18449;
  assign n18455 = n18454 ^ n17985;
  assign n18456 = n17996 & ~n18455;
  assign n18457 = n18456 ^ n17995;
  assign n18458 = n18457 ^ n17977;
  assign n18459 = ~n17978 & ~n18458;
  assign n18460 = n18459 ^ n18457;
  assign n18461 = n18460 ^ n17965;
  assign n18462 = n17966 & ~n18461;
  assign n18463 = n18462 ^ n18460;
  assign n18474 = n18473 ^ n18463;
  assign n18475 = n17888 ^ n17467;
  assign n18476 = n18475 ^ n18473;
  assign n18477 = n18474 & ~n18476;
  assign n18478 = n18477 ^ n18463;
  assign n18479 = ~n17953 & ~n18478;
  assign n18480 = n17446 & ~n17893;
  assign n18481 = ~n17446 & ~n17891;
  assign n18482 = ~n17455 & n18481;
  assign n18483 = ~n18480 & ~n18482;
  assign n18484 = n18479 & ~n18483;
  assign n18485 = n17953 & n18478;
  assign n18486 = n17455 ^ n17447;
  assign n18487 = ~n17891 & n18486;
  assign n18488 = n17892 ^ n17456;
  assign n18489 = ~n17446 & ~n18488;
  assign n18490 = n18489 ^ n17456;
  assign n18491 = ~n18487 & n18490;
  assign n18492 = ~n18485 & n18491;
  assign n18493 = ~n18484 & ~n18492;
  assign n18494 = n17896 ^ n17436;
  assign n18495 = ~n18493 & ~n18494;
  assign n18496 = x2 & ~n18495;
  assign n18500 = n33 & n11907;
  assign n18501 = n18500 ^ n11940;
  assign n18497 = x1 & n11902;
  assign n18498 = n9346 & ~n11875;
  assign n18499 = ~n18497 & ~n18498;
  assign n18502 = n18501 ^ n18499;
  assign n18503 = ~x0 & n18502;
  assign n18504 = n18503 ^ n18501;
  assign n18505 = n18504 ^ n18494;
  assign n18506 = ~n17456 & n18481;
  assign n18507 = n17891 & n18486;
  assign n18508 = n17446 & ~n17457;
  assign n18509 = ~n18507 & ~n18508;
  assign n18510 = ~n18506 & n18509;
  assign n18511 = ~n18479 & n18510;
  assign n18512 = n17455 & n17891;
  assign n18513 = n18512 ^ n17893;
  assign n18514 = ~n17446 & n18513;
  assign n18515 = n18514 ^ n17893;
  assign n18516 = n18485 & n18515;
  assign n18517 = ~n18511 & ~n18516;
  assign n18518 = n33 & n12504;
  assign n18519 = ~n33 & n11902;
  assign n18520 = x0 & ~n18519;
  assign n18521 = ~n18518 & n18520;
  assign n18522 = n9378 & n11875;
  assign n18523 = ~n18521 & ~n18522;
  assign n18524 = x2 & ~n11773;
  assign n18525 = n9448 & ~n18524;
  assign n18526 = n18523 & ~n18525;
  assign n18527 = n18517 & ~n18526;
  assign n18528 = n18493 & ~n18527;
  assign n18529 = n18528 ^ n18494;
  assign n18530 = n18505 & n18529;
  assign n18531 = n18530 ^ n18528;
  assign n18532 = ~n18496 & ~n18531;
  assign n18533 = n18517 & n18526;
  assign n18534 = n18493 & ~n18533;
  assign n18535 = n18494 & n18534;
  assign n18536 = x2 & ~n18535;
  assign n18537 = ~n18494 & n18533;
  assign n18538 = n18504 & ~n18537;
  assign n18539 = n18536 & ~n18538;
  assign n18540 = ~n18532 & ~n18539;
  assign n18541 = n18540 ^ n17942;
  assign n18542 = n17943 & n18541;
  assign n18543 = n18542 ^ n18540;
  assign n18544 = n18543 ^ n17928;
  assign n18545 = n17929 & n18544;
  assign n18546 = n18545 ^ n18543;
  assign n18547 = n18546 ^ n17916;
  assign n18548 = n17917 & n18547;
  assign n18549 = n18548 ^ n18546;
  assign n18550 = ~n17393 & n18549;
  assign n18551 = n17392 & n18550;
  assign n18552 = n17393 & ~n18549;
  assign n18553 = n7513 & n12013;
  assign n18554 = n7514 & ~n12019;
  assign n18555 = ~n18553 & n18554;
  assign n18556 = n7518 & ~n11940;
  assign n18557 = n7520 & n11902;
  assign n18558 = ~n18556 & ~n18557;
  assign n18559 = ~n18555 & n18558;
  assign n18560 = n18559 ^ x5;
  assign n18561 = n18560 ^ n12750;
  assign n18562 = n17914 ^ n17905;
  assign n18563 = ~n17915 & ~n18562;
  assign n18564 = n18563 ^ n17905;
  assign n18565 = n18564 ^ n18560;
  assign n18566 = n18564 ^ n17392;
  assign n18567 = n18565 & n18566;
  assign n18568 = n18561 & n18567;
  assign n18569 = n18568 ^ n17392;
  assign n18570 = ~n18552 & n18569;
  assign n18571 = ~n18551 & ~n18570;
  assign n18572 = ~n17392 & ~n18550;
  assign n18573 = n18560 & ~n18564;
  assign n18574 = ~n18560 & n18564;
  assign n18575 = ~n12750 & ~n18574;
  assign n18576 = ~n18573 & ~n18575;
  assign n18577 = ~n18572 & n18576;
  assign n18578 = n18571 & ~n18577;
  assign n18579 = n17390 ^ n17320;
  assign n18580 = ~n17391 & ~n18579;
  assign n18581 = n18580 ^ n17320;
  assign n18582 = n18578 & ~n18581;
  assign n18615 = n6306 & ~n11941;
  assign n18616 = n7168 & ~n11940;
  assign n18617 = n6309 & n11902;
  assign n18618 = n6316 & ~n11875;
  assign n18619 = ~n18617 & ~n18618;
  assign n18620 = ~n18616 & n18619;
  assign n18621 = ~n18615 & n18620;
  assign n18622 = n18621 ^ x8;
  assign n18605 = n5814 & ~n11777;
  assign n18606 = n6295 & ~n11773;
  assign n18607 = n5817 & n11480;
  assign n18608 = n5824 & n11500;
  assign n18609 = ~n18607 & ~n18608;
  assign n18610 = ~n18606 & n18609;
  assign n18611 = ~n18605 & n18610;
  assign n18612 = n18611 ^ x11;
  assign n18603 = n15330 ^ n15316;
  assign n18600 = n17344 ^ n17329;
  assign n18601 = n17331 & n18600;
  assign n18602 = n18601 ^ n17344;
  assign n18604 = n18603 ^ n18602;
  assign n18613 = n18612 ^ n18604;
  assign n18597 = n17361 ^ n17326;
  assign n18598 = n17362 & ~n18597;
  assign n18599 = n18598 ^ n17326;
  assign n18614 = n18613 ^ n18599;
  assign n18623 = n18622 ^ n18614;
  assign n18583 = x4 & ~x5;
  assign n18584 = n17934 & n18583;
  assign n18585 = ~x2 & x5;
  assign n18586 = ~n18584 & ~n18585;
  assign n18587 = x3 & ~n18586;
  assign n18588 = x5 & n12019;
  assign n18589 = ~x4 & n9530;
  assign n18590 = ~n18588 & n18589;
  assign n18591 = n9528 ^ x2;
  assign n18592 = x4 & ~n18591;
  assign n18593 = n18592 ^ x2;
  assign n18594 = x5 & n18593;
  assign n18595 = ~n18590 & ~n18594;
  assign n18596 = ~n18587 & n18595;
  assign n18624 = n18623 ^ n18596;
  assign n18625 = n17363 ^ n17323;
  assign n18626 = n17380 & ~n18625;
  assign n18627 = n18626 ^ n17379;
  assign n18628 = n18627 ^ n18623;
  assign n18629 = n18624 & n18628;
  assign n18630 = n18629 ^ n18627;
  assign n18631 = ~n18582 & ~n18630;
  assign n18641 = n6304 & n12013;
  assign n18642 = n6305 & ~n12019;
  assign n18643 = ~n18641 & n18642;
  assign n18644 = n6309 & ~n11940;
  assign n18645 = n6316 & n11902;
  assign n18646 = ~n18644 & ~n18645;
  assign n18647 = ~n18643 & n18646;
  assign n18648 = n18647 ^ x8;
  assign n18639 = n15343 ^ n15335;
  assign n18636 = n18612 ^ n18603;
  assign n18637 = n18604 & ~n18636;
  assign n18638 = n18637 ^ n18612;
  assign n18640 = n18639 ^ n18638;
  assign n18649 = n18648 ^ n18640;
  assign n18632 = n18622 ^ n18599;
  assign n18633 = ~n18614 & ~n18632;
  assign n18634 = n18633 ^ n18622;
  assign n18635 = n18634 ^ n12756;
  assign n18650 = n18649 ^ n18635;
  assign n18651 = ~n18631 & n18650;
  assign n18652 = ~n18578 & n18581;
  assign n18653 = ~n18596 & n18623;
  assign n18654 = n18627 & n18653;
  assign n18655 = ~n18650 & ~n18654;
  assign n18656 = n18596 & ~n18623;
  assign n18657 = ~n18627 & n18656;
  assign n18658 = ~n18655 & ~n18657;
  assign n18659 = ~n18652 & n18658;
  assign n18660 = n18582 & n18630;
  assign n18661 = ~n18659 & ~n18660;
  assign n18662 = ~n18651 & n18661;
  assign n18663 = n18649 ^ n18634;
  assign n18664 = ~n18635 & n18663;
  assign n18665 = n18664 ^ n18649;
  assign n18666 = n18648 ^ n18639;
  assign n18667 = ~n18640 & n18666;
  assign n18668 = n18667 ^ n18648;
  assign n18669 = ~n18665 & ~n18668;
  assign n18670 = n15367 ^ n15366;
  assign n18671 = n18669 & n18670;
  assign n18672 = n6306 & n17383;
  assign n18673 = n6316 & ~n11940;
  assign n18674 = n6309 & ~n12019;
  assign n18675 = ~n7168 & ~n18674;
  assign n18676 = ~n18673 & n18675;
  assign n18677 = ~n18672 & n18676;
  assign n18678 = n18677 ^ x8;
  assign n18679 = n15356 ^ n15355;
  assign n18680 = ~n18678 & n18679;
  assign n18681 = ~n18671 & ~n18680;
  assign n18682 = ~n18662 & n18681;
  assign n18683 = n18678 & ~n18679;
  assign n18684 = n18683 ^ n18669;
  assign n18685 = n18683 ^ n18670;
  assign n18686 = ~n18684 & n18685;
  assign n18687 = n18686 ^ n18669;
  assign n18688 = ~n18682 & n18687;
  assign n18689 = n18670 & ~n18683;
  assign n18690 = ~n18662 & ~n18689;
  assign n18691 = n18665 & n18668;
  assign n18692 = ~n18670 & ~n18680;
  assign n18693 = ~n18691 & ~n18692;
  assign n18694 = ~n18690 & n18693;
  assign n18695 = ~n18688 & ~n18694;
  assign n18696 = n18695 ^ n15371;
  assign n18697 = n15372 & ~n18696;
  assign n18698 = n18697 ^ n18695;
  assign n18699 = ~n14994 & n18698;
  assign n18700 = n14305 & n14993;
  assign n18701 = n5814 & n17383;
  assign n18702 = n5824 & ~n11940;
  assign n18703 = n5817 & ~n12019;
  assign n18704 = ~n6295 & ~n18703;
  assign n18705 = ~n18702 & n18704;
  assign n18706 = ~n18701 & n18705;
  assign n18707 = n18706 ^ x11;
  assign n18708 = n14634 ^ n14625;
  assign n18709 = ~n14626 & n18708;
  assign n18710 = n18709 ^ n14634;
  assign n18711 = ~n18707 & ~n18710;
  assign n18712 = ~n18700 & n18711;
  assign n18713 = n14298 ^ n14020;
  assign n18714 = ~n18700 & n18713;
  assign n18715 = ~n18712 & ~n18714;
  assign n18716 = ~n18699 & ~n18715;
  assign n18717 = n18711 & n18713;
  assign n18718 = ~n18716 & ~n18717;
  assign n18719 = n18698 & ~n18714;
  assign n18720 = n18707 & n18710;
  assign n18721 = ~n14994 & ~n18713;
  assign n18722 = ~n18720 & ~n18721;
  assign n18723 = ~n18719 & n18722;
  assign n18724 = n18718 & ~n18723;
  assign n18725 = n18724 ^ n14303;
  assign n18726 = ~n14304 & n18725;
  assign n18727 = n18726 ^ n18724;
  assign n18728 = ~n14011 & ~n18727;
  assign n18729 = n5752 & ~n11940;
  assign n18730 = ~n5746 & ~n12019;
  assign n18731 = ~n18729 & ~n18730;
  assign n18732 = n6048 ^ x14;
  assign n18733 = n18731 & n18732;
  assign n18734 = n18733 ^ x14;
  assign n18735 = n7860 ^ n5796;
  assign n18736 = n17383 & n18735;
  assign n18737 = n18736 ^ n5796;
  assign n18738 = ~n18734 & ~n18737;
  assign n18739 = n13715 ^ n13699;
  assign n18740 = n18738 & ~n18739;
  assign n18741 = ~n14006 & ~n14009;
  assign n18742 = ~n13758 & ~n18741;
  assign n18743 = ~n18740 & ~n18742;
  assign n18744 = ~n18728 & n18743;
  assign n18745 = ~n18727 & ~n18741;
  assign n18746 = ~n18738 & n18739;
  assign n18747 = ~n13758 & ~n18746;
  assign n18748 = ~n14010 & ~n18747;
  assign n18749 = ~n18745 & n18748;
  assign n18750 = ~n18744 & ~n18749;
  assign n18751 = n13758 & n18746;
  assign n18752 = n18750 & ~n18751;
  assign n18753 = n13752 ^ n13734;
  assign n18754 = n13736 & n18753;
  assign n18755 = n18754 ^ n13752;
  assign n18756 = n18752 & ~n18755;
  assign n18757 = n13757 & n18756;
  assign n18783 = n18782 ^ n18760;
  assign n18784 = ~n13087 & ~n13756;
  assign n18785 = n11578 & ~n18784;
  assign n18786 = ~n13757 & ~n18785;
  assign n18787 = n18783 & ~n18786;
  assign n18788 = ~n18757 & ~n18787;
  assign n18789 = ~n18783 & ~n18785;
  assign n18790 = n18756 & ~n18789;
  assign n18791 = ~n18752 & n18755;
  assign n18792 = n13756 ^ n13087;
  assign n18793 = n13087 ^ n11578;
  assign n18794 = n18783 ^ n11578;
  assign n18795 = ~n18793 & n18794;
  assign n18796 = ~n18792 & n18795;
  assign n18797 = n18796 ^ n18783;
  assign n18798 = ~n18791 & n18797;
  assign n18799 = ~n18790 & ~n18798;
  assign n18800 = n18788 & n18799;
  assign n18801 = n18764 ^ n18763;
  assign n18802 = ~n18773 & n18801;
  assign n18803 = n18802 ^ n18772;
  assign n18832 = n18800 & n18803;
  assign n19097 = n18831 & n18832;
  assign n18804 = ~n18800 & ~n18803;
  assign n18822 = ~n18805 & ~n18816;
  assign n18823 = n18820 & n18822;
  assign n19098 = ~n18804 & n18823;
  assign n19099 = ~n19097 & ~n19098;
  assign n18817 = n18805 & n18816;
  assign n18821 = n18817 & ~n18820;
  assign n19100 = n18821 & ~n18832;
  assign n19101 = n18804 & ~n18831;
  assign n19102 = ~n19100 & ~n19101;
  assign n19103 = n19099 & n19102;
  assign n12685 = n4672 & n12013;
  assign n12686 = n4671 & ~n12019;
  assign n12687 = ~n12685 & n12686;
  assign n12688 = n4685 & ~n11940;
  assign n12689 = ~n4681 & n11902;
  assign n12690 = ~n12688 & ~n12689;
  assign n12691 = ~n12687 & n12690;
  assign n12692 = n12691 ^ x20;
  assign n12438 = n4478 & ~n12000;
  assign n12439 = n4487 & ~n11875;
  assign n12440 = n4484 & ~n11773;
  assign n12441 = n4480 & n11480;
  assign n12442 = ~n12440 & ~n12441;
  assign n12443 = ~n12439 & n12442;
  assign n12444 = ~n12438 & n12443;
  assign n12445 = n12444 ^ x23;
  assign n12418 = n11957 & n12417;
  assign n12419 = n3435 & n11486;
  assign n12420 = ~n3440 & n11215;
  assign n12421 = ~n12419 & ~n12420;
  assign n12422 = x26 & n12421;
  assign n12423 = ~n11500 & n12422;
  assign n12424 = x25 & ~n12423;
  assign n12425 = ~n12418 & n12424;
  assign n12426 = ~n11957 & n12422;
  assign n12427 = n11500 & n12417;
  assign n12428 = ~x25 & ~n12427;
  assign n12429 = ~n12426 & n12428;
  assign n12430 = ~n12425 & ~n12429;
  assign n12433 = n12421 & ~n12432;
  assign n12434 = n12433 ^ x26;
  assign n12435 = ~n12430 & n12434;
  assign n12407 = n44 & ~n10957;
  assign n12408 = n3277 & ~n10663;
  assign n12409 = n3280 & ~n10956;
  assign n12410 = n3275 & n10665;
  assign n12411 = ~n12409 & ~n12410;
  assign n12412 = ~n12408 & n12411;
  assign n12413 = ~n12407 & n12412;
  assign n12414 = n12413 ^ x29;
  assign n12398 = x31 & n11616;
  assign n12399 = n12398 ^ n10680;
  assign n12400 = n41 & n12399;
  assign n12401 = x31 & n11604;
  assign n12402 = ~n3673 & n10683;
  assign n12403 = ~n12401 & ~n12402;
  assign n12404 = ~n12400 & n12403;
  assign n11638 = n3469 & n3713;
  assign n11639 = n1164 & n2038;
  assign n11640 = n3163 & n4388;
  assign n11641 = n11639 & n11640;
  assign n11642 = ~n326 & ~n800;
  assign n11643 = ~n4086 & n11642;
  assign n11644 = n949 & n1197;
  assign n11645 = n11643 & n11644;
  assign n11646 = n11641 & n11645;
  assign n11647 = ~n417 & n1561;
  assign n11648 = n1312 & n2957;
  assign n11649 = n11647 & n11648;
  assign n11650 = n11646 & n11649;
  assign n11651 = ~n170 & ~n443;
  assign n11652 = ~n409 & n11651;
  assign n11653 = n5033 & n11652;
  assign n11654 = n11650 & n11653;
  assign n11655 = n2891 & n4245;
  assign n11656 = n11654 & n11655;
  assign n11657 = n732 & n11656;
  assign n11658 = n11638 & n11657;
  assign n12397 = n11658 ^ n11554;
  assign n12405 = n12404 ^ n12397;
  assign n11611 = n11610 ^ n11596;
  assign n11612 = n11597 & ~n11611;
  assign n11613 = n11612 ^ n11610;
  assign n12406 = n12405 ^ n11613;
  assign n12415 = n12414 ^ n12406;
  assign n12394 = n12371 ^ n12358;
  assign n12395 = n12380 & ~n12394;
  assign n12396 = n12395 ^ n12379;
  assign n12416 = n12415 ^ n12396;
  assign n12436 = n12435 ^ n12416;
  assign n12391 = n12390 ^ n12357;
  assign n12392 = n12382 & ~n12391;
  assign n12393 = n12392 ^ n12390;
  assign n12437 = n12436 ^ n12393;
  assign n12683 = n12445 ^ n12437;
  assign n12680 = n12665 ^ n12656;
  assign n12681 = n12657 & ~n12680;
  assign n12682 = n12681 ^ n12665;
  assign n12684 = n12683 ^ n12682;
  assign n12693 = n12692 ^ n12684;
  assign n12676 = n12675 ^ n12652;
  assign n12677 = n12667 & n12676;
  assign n12678 = n12677 ^ n12675;
  assign n11675 = ~n4966 & ~n11674;
  assign n12679 = n12678 ^ n11675;
  assign n18824 = n12693 ^ n12679;
  assign n19104 = n19103 ^ n18824;
  assign n19105 = n11578 & n13757;
  assign n19106 = ~n18791 & n19105;
  assign n19107 = n18756 & n18785;
  assign n19108 = ~n19106 & ~n19107;
  assign n19109 = ~n13087 & n18755;
  assign n19110 = ~n13756 & n19109;
  assign n19111 = ~n18752 & n19110;
  assign n19112 = ~n18757 & ~n19111;
  assign n19113 = n19108 & n19112;
  assign n19114 = n18755 ^ n13087;
  assign n19115 = n18755 ^ n13756;
  assign n19116 = n19114 & ~n19115;
  assign n19117 = n19116 ^ n13756;
  assign n19118 = ~n18752 & ~n19117;
  assign n19119 = ~n19110 & ~n19118;
  assign n19120 = ~n11578 & ~n19119;
  assign n19121 = n19113 & ~n19120;
  assign n19122 = n19121 ^ n18783;
  assign n19129 = ~n18678 & ~n18691;
  assign n19130 = ~n18669 & ~n19129;
  assign n19131 = n18679 & ~n19130;
  assign n19132 = n18669 & ~n18678;
  assign n19133 = n18683 & n18691;
  assign n19134 = ~n19132 & ~n19133;
  assign n19135 = ~n19131 & n19134;
  assign n19123 = n18678 ^ n18668;
  assign n19126 = n18679 ^ n18678;
  assign n19127 = ~n19123 & n19126;
  assign n19124 = n19123 ^ n18679;
  assign n19125 = n18665 & n19124;
  assign n19128 = n19127 ^ n19125;
  assign n19136 = n19135 ^ n19128;
  assign n19137 = ~n18662 & ~n19136;
  assign n19138 = n19137 ^ n19135;
  assign n19139 = n19138 ^ n18670;
  assign n19140 = n19126 ^ n18668;
  assign n19141 = n19140 ^ n18665;
  assign n19142 = n19141 ^ n18662;
  assign n19143 = n18549 & ~n18560;
  assign n19144 = n17393 & ~n18564;
  assign n19145 = ~n12750 & n19144;
  assign n19146 = ~n19143 & n19145;
  assign n19147 = ~n18549 & n18560;
  assign n19148 = ~n17393 & n18564;
  assign n19149 = n12750 & n19148;
  assign n19150 = ~n19147 & n19149;
  assign n19151 = ~n19146 & ~n19150;
  assign n19152 = n12750 & ~n19144;
  assign n19153 = n19143 & n19152;
  assign n19154 = n19151 & ~n19153;
  assign n19155 = n19147 & ~n19152;
  assign n19156 = n19155 ^ n19143;
  assign n19157 = n19148 & n19156;
  assign n19158 = n19157 ^ n19155;
  assign n19159 = n19154 & ~n19158;
  assign n19160 = n19159 ^ n17392;
  assign n19161 = n18540 ^ n17943;
  assign n19162 = n18546 ^ n17917;
  assign n19163 = n19160 & ~n19162;
  assign n19164 = n18534 ^ n18528;
  assign n19165 = x2 & ~n19164;
  assign n19166 = n19165 ^ n18528;
  assign n19167 = n19166 ^ n18505;
  assign n19169 = n18493 & n18517;
  assign n19168 = n18526 ^ x2;
  assign n19170 = n19169 ^ n19168;
  assign n19171 = n18486 ^ n17891;
  assign n19172 = n19171 ^ n17953;
  assign n19173 = n19172 ^ n18478;
  assign n19174 = n18475 ^ n18474;
  assign n19175 = n18460 ^ n17966;
  assign n19176 = n19174 & ~n19175;
  assign n19177 = ~n19173 & ~n19176;
  assign n19178 = n19170 & ~n19177;
  assign n19179 = n19167 & ~n19178;
  assign n19180 = ~n19161 & ~n19179;
  assign n19183 = n17964 ^ n17963;
  assign n19184 = ~n17885 & ~n19183;
  assign n19181 = n17963 ^ n17476;
  assign n19182 = n17964 & n19181;
  assign n19185 = n19184 ^ n19182;
  assign n19186 = n19185 ^ n17467;
  assign n19187 = n19186 ^ n18473;
  assign n19188 = n18457 ^ n17978;
  assign n19189 = ~n19187 & ~n19188;
  assign n19190 = ~n19175 & ~n19189;
  assign n19191 = ~n19174 & ~n19190;
  assign n19192 = n19173 & ~n19191;
  assign n19193 = ~n19170 & ~n19192;
  assign n19194 = ~n19167 & ~n19193;
  assign n19195 = ~n19180 & ~n19194;
  assign n19196 = n19163 & ~n19195;
  assign n19197 = n18560 ^ n17393;
  assign n19198 = n19197 ^ n12750;
  assign n19199 = n19198 ^ n18564;
  assign n19200 = n19199 ^ n18549;
  assign n19201 = n18543 ^ n17929;
  assign n19202 = n19200 & ~n19201;
  assign n19203 = ~n19196 & ~n19202;
  assign n19204 = ~n19161 & ~n19203;
  assign n19205 = ~n19160 & n19162;
  assign n19206 = n19200 & ~n19205;
  assign n19207 = ~n19195 & n19202;
  assign n19208 = ~n19206 & ~n19207;
  assign n19209 = n19163 & ~n19201;
  assign n19210 = n19208 & ~n19209;
  assign n19211 = ~n19204 & n19210;
  assign n19212 = ~n19160 & n19211;
  assign n19213 = n18627 ^ n18624;
  assign n19214 = n19213 ^ n18581;
  assign n19215 = n19214 ^ n18578;
  assign n19216 = ~n19212 & ~n19215;
  assign n19217 = ~n19142 & n19216;
  assign n19218 = n18654 ^ n18630;
  assign n19219 = ~n18652 & ~n19218;
  assign n19220 = n19219 ^ n18630;
  assign n19221 = n18657 ^ n18630;
  assign n19222 = ~n18582 & n19221;
  assign n19223 = n19222 ^ n18630;
  assign n19224 = n19220 & ~n19223;
  assign n19225 = n19224 ^ n18650;
  assign n19226 = ~n19217 & n19225;
  assign n19227 = n19160 & ~n19211;
  assign n19228 = n19215 & ~n19227;
  assign n19229 = n19142 & n19228;
  assign n19230 = ~n19226 & ~n19229;
  assign n19231 = n19142 & ~n19230;
  assign n19232 = n19139 & ~n19231;
  assign n19233 = n18695 ^ n15372;
  assign n19234 = ~n19232 & ~n19233;
  assign n19235 = n18707 ^ n14305;
  assign n19236 = n19235 ^ n18710;
  assign n19237 = n19236 ^ n14993;
  assign n19238 = n19237 ^ n18698;
  assign n19239 = ~n19234 & ~n19238;
  assign n19242 = n18700 & ~n18711;
  assign n19243 = ~n14994 & n18720;
  assign n19244 = ~n19242 & ~n19243;
  assign n19240 = n14994 & ~n18720;
  assign n19241 = ~n18712 & ~n19240;
  assign n19245 = n19244 ^ n19241;
  assign n19246 = ~n18698 & n19245;
  assign n19247 = n19246 ^ n19244;
  assign n19248 = n18710 ^ n14993;
  assign n19249 = n18710 ^ n14305;
  assign n19250 = ~n19235 & ~n19249;
  assign n19251 = ~n19248 & n19250;
  assign n19252 = n19247 & ~n19251;
  assign n19253 = n19252 ^ n18713;
  assign n19254 = ~n19239 & ~n19253;
  assign n19255 = n18724 ^ n14304;
  assign n19256 = ~n19254 & ~n19255;
  assign n19257 = n18739 ^ n18738;
  assign n19258 = n19257 ^ n14009;
  assign n19259 = n19258 ^ n14006;
  assign n19260 = n19259 ^ n18727;
  assign n19261 = ~n19256 & ~n19260;
  assign n19267 = n14006 & ~n18746;
  assign n19268 = ~n18740 & ~n19267;
  assign n19269 = n14009 & ~n19268;
  assign n19270 = n14006 & n18740;
  assign n19271 = n18741 & n18746;
  assign n19272 = ~n19270 & ~n19271;
  assign n19273 = ~n19269 & n19272;
  assign n19262 = n18738 ^ n14009;
  assign n19264 = n19262 ^ n18739;
  assign n19265 = ~n14006 & ~n19264;
  assign n19263 = n19257 & ~n19262;
  assign n19266 = n19265 ^ n19263;
  assign n19274 = n19273 ^ n19266;
  assign n19275 = ~n18727 & ~n19274;
  assign n19276 = n19275 ^ n19266;
  assign n19277 = n19276 ^ n13758;
  assign n19278 = ~n19261 & n19277;
  assign n19279 = n18793 ^ n18755;
  assign n19280 = n19279 ^ n13756;
  assign n19281 = n19280 ^ n18752;
  assign n19282 = ~n19278 & n19281;
  assign n19283 = n19122 & ~n19282;
  assign n19284 = n18828 ^ n18803;
  assign n19285 = n19284 ^ n18820;
  assign n19286 = n19285 ^ n18800;
  assign n19287 = ~n19283 & n19286;
  assign n19288 = n19104 & ~n19287;
  assign n19577 = ~n19142 & ~n19226;
  assign n19578 = ~n19139 & ~n19577;
  assign n19579 = n19233 & ~n19578;
  assign n19580 = n19238 & ~n19579;
  assign n19581 = n19253 & ~n19580;
  assign n19582 = n19255 & ~n19581;
  assign n19583 = n19260 & ~n19582;
  assign n19584 = ~n19277 & ~n19583;
  assign n19585 = ~n19281 & ~n19584;
  assign n19586 = ~n19122 & ~n19585;
  assign n19587 = ~n19286 & ~n19586;
  assign n19588 = ~n19104 & ~n19587;
  assign n21683 = ~n19288 & ~n19588;
  assign n18839 = n4673 & n17383;
  assign n18840 = ~n4681 & ~n11940;
  assign n18841 = n4685 & ~n12019;
  assign n18842 = ~n4688 & ~n18841;
  assign n18843 = ~n18840 & n18842;
  assign n18844 = ~n18839 & n18843;
  assign n18845 = n18844 ^ x20;
  assign n12505 = n12502 & n12504;
  assign n12506 = n4484 & ~n11875;
  assign n12507 = n4480 & ~n11773;
  assign n12508 = ~n12506 & ~n12507;
  assign n12509 = x23 & n12508;
  assign n12510 = ~n11902 & n12509;
  assign n12511 = ~n12505 & ~n12510;
  assign n12512 = x22 & n12511;
  assign n12513 = ~n12504 & n12509;
  assign n12514 = n11902 & n12502;
  assign n12515 = ~x22 & ~n12514;
  assign n12516 = ~n12513 & n12515;
  assign n12517 = ~n12512 & ~n12516;
  assign n12520 = n12508 & ~n12519;
  assign n12521 = n12520 ^ x23;
  assign n12522 = ~n12517 & n12521;
  assign n12481 = n12404 & n12414;
  assign n12482 = ~n11658 & n12481;
  assign n12483 = n11613 & ~n12482;
  assign n12484 = n11554 & ~n12483;
  assign n12485 = n12404 ^ n11658;
  assign n12486 = n12414 ^ n12404;
  assign n12487 = n12485 & n12486;
  assign n12488 = n12487 ^ n12414;
  assign n12489 = n12484 & n12488;
  assign n11614 = ~n11554 & n11613;
  assign n12490 = n11614 & ~n12488;
  assign n12491 = ~n11613 & n12482;
  assign n11680 = n11554 & ~n11613;
  assign n11684 = n11658 & ~n11680;
  assign n12492 = ~n12404 & ~n12414;
  assign n12493 = n11684 & n12492;
  assign n12494 = ~n12491 & ~n12493;
  assign n12495 = ~n12490 & n12494;
  assign n12496 = ~n12489 & n12495;
  assign n10969 = ~n327 & ~n373;
  assign n10970 = ~n797 & n10969;
  assign n10971 = ~n652 & n3113;
  assign n10972 = n10970 & n10971;
  assign n10973 = n10968 & n10972;
  assign n10974 = n187 & n4078;
  assign n10975 = n2202 & n10974;
  assign n10976 = n10973 & n10975;
  assign n11008 = ~n156 & ~n758;
  assign n11659 = n58 & n11008;
  assign n11660 = n526 & n3007;
  assign n11661 = n11659 & n11660;
  assign n11662 = ~n336 & ~n410;
  assign n11663 = n801 & n11662;
  assign n11664 = n441 & n2180;
  assign n11665 = n11663 & n11664;
  assign n11666 = n11661 & n11665;
  assign n11667 = n783 & n960;
  assign n11668 = n4618 & n11667;
  assign n11669 = n11666 & n11668;
  assign n11670 = n10976 & n11669;
  assign n11671 = n1340 & n11411;
  assign n11672 = n11670 & n11671;
  assign n11673 = n4748 & n11672;
  assign n11676 = n11675 ^ n11673;
  assign n11685 = n11676 ^ n11658;
  assign n11615 = n10680 & n11606;
  assign n11617 = n41 & n11616;
  assign n11618 = ~n11615 & ~n11617;
  assign n11619 = ~n10665 & ~n11618;
  assign n11620 = x31 & ~n11619;
  assign n11621 = ~n54 & n10875;
  assign n11622 = n10665 & n11621;
  assign n11623 = ~n91 & ~n11622;
  assign n11624 = ~n10680 & ~n11623;
  assign n11625 = n11620 & ~n11624;
  assign n11627 = ~n91 & n10665;
  assign n11628 = n11626 & n11627;
  assign n11629 = ~n54 & ~n11223;
  assign n11630 = ~n11628 & n11629;
  assign n11631 = ~n10683 & ~n11630;
  assign n11632 = n11625 & ~n11631;
  assign n11633 = n54 & ~n10680;
  assign n11634 = n3640 & ~n11633;
  assign n11635 = ~n54 & ~n10665;
  assign n11636 = n11634 & ~n11635;
  assign n11637 = ~n11632 & ~n11636;
  assign n12480 = n11685 ^ n11637;
  assign n12497 = n12496 ^ n12480;
  assign n12469 = ~n12460 & n12466;
  assign n12461 = n3275 & ~n10663;
  assign n12462 = n3277 & ~n10956;
  assign n12463 = ~n12461 & ~n12462;
  assign n12464 = x29 & n12463;
  assign n12470 = ~n11215 & n12464;
  assign n12471 = ~n12469 & ~n12470;
  assign n12465 = n12460 & n12464;
  assign n12467 = n11215 & n12466;
  assign n12468 = ~n12465 & ~n12467;
  assign n12472 = n12471 ^ n12468;
  assign n12473 = ~x28 & n12472;
  assign n12474 = n12473 ^ n12471;
  assign n12477 = n12463 & ~n12476;
  assign n12478 = n12477 ^ x29;
  assign n12479 = n12474 & n12478;
  assign n12498 = n12497 ^ n12479;
  assign n12452 = n3285 & n11507;
  assign n12453 = n3435 & n11500;
  assign n12454 = ~n3440 & n11486;
  assign n12455 = ~n12453 & ~n12454;
  assign n12456 = n3437 & n11480;
  assign n12457 = n12455 & ~n12456;
  assign n12458 = ~n12452 & n12457;
  assign n12459 = n12458 ^ x26;
  assign n12499 = n12498 ^ n12459;
  assign n12449 = n12435 ^ n12415;
  assign n12450 = ~n12416 & n12449;
  assign n12451 = n12450 ^ n12435;
  assign n12500 = n12499 ^ n12451;
  assign n12446 = n12445 ^ n12436;
  assign n12447 = ~n12437 & n12446;
  assign n12448 = n12447 ^ n12445;
  assign n12501 = n12500 ^ n12448;
  assign n12523 = n12522 ^ n12501;
  assign n19289 = n18845 ^ n12523;
  assign n12698 = n12692 ^ n12683;
  assign n12699 = ~n12684 & n12698;
  assign n12700 = n12699 ^ n12692;
  assign n19290 = n19289 ^ n12700;
  assign n12694 = n12693 ^ n12678;
  assign n12695 = n12679 & n12694;
  assign n12696 = n12695 ^ n12693;
  assign n19291 = n19290 ^ n12696;
  assign n18825 = ~n18823 & n18824;
  assign n18826 = ~n18821 & ~n18825;
  assign n18827 = ~n18804 & n18826;
  assign n18833 = n18832 ^ n18831;
  assign n18834 = n18831 ^ n18824;
  assign n18835 = n18833 & n18834;
  assign n18836 = n18835 ^ n18832;
  assign n18837 = ~n18827 & ~n18836;
  assign n19292 = n19291 ^ n18837;
  assign n21684 = n21683 ^ n19292;
  assign n21867 = n5814 & n21684;
  assign n21868 = n6295 & n19292;
  assign n21869 = n5817 & n19104;
  assign n21870 = n5824 & ~n19286;
  assign n21871 = ~n21869 & ~n21870;
  assign n21872 = ~n21868 & n21871;
  assign n21873 = ~n21867 & n21872;
  assign n21874 = n21873 ^ x11;
  assign n19695 = ~n19254 & ~n19581;
  assign n19696 = n19695 ^ n19255;
  assign n21340 = n4963 & ~n19696;
  assign n21341 = n4972 & ~n19255;
  assign n21342 = n4976 & n19253;
  assign n21343 = n4970 & ~n19238;
  assign n21344 = ~n21342 & ~n21343;
  assign n21345 = ~n21341 & n21344;
  assign n21346 = ~n21340 & n21345;
  assign n21347 = n21346 ^ x17;
  assign n20293 = ~n19232 & ~n19578;
  assign n20294 = n20293 ^ n19233;
  assign n21330 = n4673 & n20294;
  assign n21331 = n4688 & n19233;
  assign n21332 = n4685 & n19139;
  assign n21333 = ~n4681 & ~n19142;
  assign n21334 = ~n21332 & ~n21333;
  assign n21335 = ~n21331 & n21334;
  assign n21336 = ~n21330 & n21335;
  assign n21337 = n21336 ^ x20;
  assign n20209 = ~n19216 & ~n19228;
  assign n20210 = n20209 ^ n19225;
  assign n21320 = n12502 & ~n20210;
  assign n21313 = n4480 & n19160;
  assign n21314 = n4484 & ~n19215;
  assign n21315 = ~n21313 & ~n21314;
  assign n21316 = x23 & n21315;
  assign n21321 = n19225 & n21316;
  assign n21322 = ~n21320 & ~n21321;
  assign n21317 = n20210 & n21316;
  assign n21318 = n12502 & ~n19225;
  assign n21319 = ~n21317 & ~n21318;
  assign n21323 = n21322 ^ n21319;
  assign n21324 = ~x22 & n21323;
  assign n21325 = n21324 ^ n21322;
  assign n21326 = ~n12519 & n21315;
  assign n21327 = n21326 ^ x23;
  assign n21328 = n21325 & n21327;
  assign n19810 = n19161 & ~n19194;
  assign n19811 = ~n19201 & ~n19810;
  assign n19812 = n19162 & ~n19811;
  assign n19813 = ~n19180 & n19201;
  assign n19814 = ~n19162 & ~n19813;
  assign n19815 = ~n19812 & ~n19814;
  assign n19816 = n19815 ^ n19200;
  assign n21302 = n3285 & n19816;
  assign n21303 = n3437 & n19200;
  assign n21304 = n3435 & ~n19162;
  assign n21305 = ~n3440 & ~n19201;
  assign n21306 = ~n21304 & ~n21305;
  assign n21307 = ~n21303 & n21306;
  assign n21308 = ~n21302 & n21307;
  assign n21309 = n21308 ^ x26;
  assign n19798 = ~n19179 & ~n19194;
  assign n19799 = n19798 ^ n19161;
  assign n21292 = n44 & ~n19799;
  assign n21293 = n3280 & ~n19161;
  assign n21294 = n3277 & ~n19167;
  assign n21295 = n3275 & n19170;
  assign n21296 = ~n21294 & ~n21295;
  assign n21297 = ~n21293 & n21296;
  assign n21298 = ~n21292 & n21297;
  assign n21299 = n21298 ^ x29;
  assign n19719 = n19190 ^ n19174;
  assign n19720 = n19719 ^ n19173;
  assign n21279 = n41 & n19720;
  assign n21280 = n91 & n19174;
  assign n21281 = n54 & ~n19175;
  assign n21282 = x31 & ~n21281;
  assign n21283 = ~n21280 & n21282;
  assign n21284 = ~n21279 & n21283;
  assign n21285 = n41 & n19173;
  assign n21286 = n54 & n19174;
  assign n21287 = ~x31 & ~n21286;
  assign n21288 = ~n21285 & n21287;
  assign n21289 = ~n21284 & ~n21288;
  assign n21261 = ~n443 & ~n463;
  assign n21262 = n4040 & n21261;
  assign n21263 = n4065 & n21262;
  assign n21264 = n2199 & n21263;
  assign n21265 = ~n500 & n635;
  assign n21266 = ~n152 & ~n424;
  assign n21267 = ~n117 & ~n222;
  assign n21268 = n21266 & n21267;
  assign n21269 = n21265 & n21268;
  assign n21270 = n520 & n3515;
  assign n21271 = n441 & ~n691;
  assign n21272 = n21270 & n21271;
  assign n21273 = n21269 & n21272;
  assign n21274 = n21264 & n21273;
  assign n21275 = n3728 & n21274;
  assign n21276 = n4203 & n21275;
  assign n21277 = n2747 & n21276;
  assign n21278 = n367 & n21277;
  assign n21290 = n21289 ^ n21278;
  assign n20691 = n41 & ~n19175;
  assign n20693 = n5636 & n19188;
  assign n20692 = x31 & n19188;
  assign n20694 = n20693 ^ n20692;
  assign n20695 = n20691 & ~n20694;
  assign n20696 = n20695 ^ n20693;
  assign n20697 = ~n576 & n1301;
  assign n20698 = n2104 & n20697;
  assign n20699 = n2622 & n20698;
  assign n20700 = n13418 & n20699;
  assign n20701 = n3572 & n4522;
  assign n20702 = n12302 & n20701;
  assign n20703 = n2209 & n2607;
  assign n20704 = n1238 & n2240;
  assign n20705 = n20703 & n20704;
  assign n20706 = n20702 & n20705;
  assign n20707 = n20700 & n20706;
  assign n20708 = ~n504 & ~n929;
  assign n20709 = ~n535 & n20708;
  assign n20710 = n13184 & n20709;
  assign n20711 = n10092 & n20710;
  assign n20712 = n551 & n2138;
  assign n20713 = ~n206 & n3515;
  assign n20714 = n20712 & n20713;
  assign n20715 = n20711 & n20714;
  assign n20716 = n20707 & n20715;
  assign n20717 = n1043 & n1312;
  assign n20718 = n12145 & n20717;
  assign n20719 = ~n471 & ~n797;
  assign n20720 = ~n514 & ~n617;
  assign n20721 = n20719 & n20720;
  assign n20722 = n20718 & n20721;
  assign n20723 = n10218 & n12072;
  assign n20724 = n20722 & n20723;
  assign n20725 = n1855 & n2166;
  assign n20726 = n3953 & n3964;
  assign n20727 = n20725 & n20726;
  assign n20728 = n20724 & n20727;
  assign n20729 = n20716 & n20728;
  assign n20730 = n13300 & n20729;
  assign n20842 = n20696 & ~n20730;
  assign n20825 = n3710 & n11588;
  assign n20826 = n2335 & n20825;
  assign n20827 = n4129 & n20826;
  assign n20828 = n2633 & n20827;
  assign n20829 = n2997 & n11523;
  assign n20830 = n1314 & n2239;
  assign n20831 = n20829 & n20830;
  assign n20832 = n191 & n3059;
  assign n20833 = ~n243 & ~n266;
  assign n20834 = ~n51 & ~n525;
  assign n20835 = n20833 & n20834;
  assign n20836 = n20832 & n20835;
  assign n20837 = n20831 & n20836;
  assign n20838 = n3695 & n20837;
  assign n20839 = n20828 & n20838;
  assign n20840 = n5528 & n20839;
  assign n20841 = n13301 & n20840;
  assign n20843 = n20842 ^ n20841;
  assign n19987 = ~n19174 & ~n19188;
  assign n20844 = n11234 & ~n19987;
  assign n20845 = n5636 & ~n19175;
  assign n20846 = ~n20844 & n20845;
  assign n19729 = ~n19175 & ~n19188;
  assign n20847 = x31 & n19729;
  assign n20848 = n41 & ~n20847;
  assign n20849 = n19174 & n20848;
  assign n20850 = n3669 & n19188;
  assign n20851 = ~n20849 & ~n20850;
  assign n20852 = ~n20846 & n20851;
  assign n21258 = n20852 ^ n20842;
  assign n21259 = n20843 & ~n21258;
  assign n21260 = n21259 ^ n20852;
  assign n21291 = n21290 ^ n21260;
  assign n21300 = n21299 ^ n21291;
  assign n19760 = ~n19178 & ~n19193;
  assign n19761 = n19760 ^ n19167;
  assign n20854 = n44 & ~n19761;
  assign n20855 = n3280 & ~n19167;
  assign n20856 = n3277 & n19170;
  assign n20857 = n3275 & n19173;
  assign n20858 = ~n20856 & ~n20857;
  assign n20859 = ~n20855 & n20858;
  assign n20860 = ~n20854 & n20859;
  assign n20861 = n20860 ^ x29;
  assign n20853 = n20852 ^ n20843;
  assign n20862 = n20861 ^ n20853;
  assign n20245 = n44 & n19720;
  assign n20246 = n3280 & n19173;
  assign n20247 = n3277 & n19174;
  assign n20248 = n3275 & ~n19175;
  assign n20249 = ~n20247 & ~n20248;
  assign n20250 = ~n20246 & n20249;
  assign n20251 = ~n20245 & n20250;
  assign n20252 = n20251 ^ x29;
  assign n19988 = n44 & n19987;
  assign n19989 = ~n3277 & ~n19988;
  assign n19990 = ~n19175 & ~n19989;
  assign n19991 = n44 & ~n19729;
  assign n19992 = ~n3280 & ~n19991;
  assign n19993 = n19174 & ~n19992;
  assign n19994 = n3275 & n19188;
  assign n19995 = ~n19993 & ~n19994;
  assign n19996 = ~n19990 & n19995;
  assign n19933 = n42 & ~n19175;
  assign n19984 = n6179 & n19188;
  assign n19985 = ~n19933 & ~n19984;
  assign n20253 = x29 & n19985;
  assign n20254 = n19996 & n20253;
  assign n20259 = n41 & n19188;
  assign n20732 = ~n20254 & ~n20259;
  assign n20733 = ~n20252 & ~n20732;
  assign n20731 = n20730 ^ n20696;
  assign n20734 = n20733 ^ n20731;
  assign n19747 = ~n19177 & ~n19192;
  assign n19748 = n19747 ^ n19170;
  assign n20735 = ~x28 & n19748;
  assign n20736 = x28 & n19170;
  assign n20737 = x29 & ~n20736;
  assign n20738 = ~n20735 & n20737;
  assign n20739 = ~n12475 & ~n20738;
  assign n20740 = n3277 & n19173;
  assign n20741 = n3275 & n19174;
  assign n20742 = ~n20740 & ~n20741;
  assign n20743 = ~n20739 & n20742;
  assign n20744 = x28 & ~n6475;
  assign n20745 = ~n6177 & n20744;
  assign n20746 = n19748 & n20745;
  assign n20747 = ~x28 & n42;
  assign n20748 = n19170 & n20747;
  assign n20749 = n20742 & ~n20748;
  assign n20750 = ~n20746 & n20749;
  assign n20751 = ~x29 & ~n20750;
  assign n20752 = ~n20743 & ~n20751;
  assign n20822 = n20752 ^ n20733;
  assign n20823 = n20734 & ~n20822;
  assign n20824 = n20823 ^ n20752;
  assign n21255 = n20853 ^ n20824;
  assign n21256 = ~n20862 & n21255;
  assign n21257 = n21256 ^ n20861;
  assign n21301 = n21300 ^ n21257;
  assign n21310 = n21309 ^ n21301;
  assign n19827 = ~n19811 & ~n19813;
  assign n19828 = n19827 ^ n19162;
  assign n20864 = n3285 & ~n19828;
  assign n20865 = n3437 & ~n19162;
  assign n20866 = n3435 & ~n19201;
  assign n20867 = ~n3440 & ~n19161;
  assign n20868 = ~n20866 & ~n20867;
  assign n20869 = ~n20865 & n20868;
  assign n20870 = ~n20864 & n20869;
  assign n20871 = n20870 ^ x26;
  assign n20863 = n20862 ^ n20824;
  assign n20872 = n20871 ^ n20863;
  assign n19839 = ~n19180 & ~n19810;
  assign n19840 = n19839 ^ n19201;
  assign n20754 = n3285 & ~n19840;
  assign n20755 = n3437 & ~n19201;
  assign n20756 = n3435 & ~n19161;
  assign n20757 = ~n3440 & ~n19167;
  assign n20758 = ~n20756 & ~n20757;
  assign n20759 = ~n20755 & n20758;
  assign n20760 = ~n20754 & n20759;
  assign n20761 = n20760 ^ x26;
  assign n20753 = n20752 ^ n20734;
  assign n20762 = n20761 ^ n20753;
  assign n20263 = n3285 & ~n19799;
  assign n20264 = n3437 & ~n19161;
  assign n20265 = n3435 & ~n19167;
  assign n20266 = ~n3440 & n19170;
  assign n20267 = ~n20265 & ~n20266;
  assign n20268 = ~n20264 & n20267;
  assign n20269 = ~n20263 & n20268;
  assign n20270 = n20269 ^ x26;
  assign n20255 = n20254 ^ n20252;
  assign n20256 = n91 & n20251;
  assign n20257 = ~n54 & n19188;
  assign n20258 = ~n20256 & n20257;
  assign n20260 = n20259 ^ n20258;
  assign n20261 = n20255 & ~n20260;
  assign n20262 = n20261 ^ n20259;
  assign n20271 = n20270 ^ n20262;
  assign n19998 = n3285 & ~n19761;
  assign n19999 = n3437 & ~n19167;
  assign n20000 = n3435 & n19170;
  assign n20001 = ~n3440 & n19173;
  assign n20002 = ~n20000 & ~n20001;
  assign n20003 = ~n19999 & n20002;
  assign n20004 = ~n19998 & n20003;
  assign n20005 = n20004 ^ x26;
  assign n19986 = x29 & ~n19985;
  assign n19997 = n19996 ^ n19986;
  assign n20006 = n20005 ^ n19997;
  assign n19789 = n3285 & n19720;
  assign n19790 = n3437 & n19173;
  assign n19791 = n3435 & n19174;
  assign n19792 = ~n3440 & ~n19175;
  assign n19793 = ~n19791 & ~n19792;
  assign n19794 = ~n19790 & n19793;
  assign n19795 = ~n19789 & n19794;
  assign n19796 = n19795 ^ x26;
  assign n19785 = n42 & n19188;
  assign n19730 = n19729 ^ n19174;
  assign n19774 = n3285 & n19730;
  assign n19775 = n3437 & n19174;
  assign n19776 = n3435 & ~n19175;
  assign n19777 = ~n3440 & n19188;
  assign n19778 = ~n19776 & ~n19777;
  assign n19779 = ~n19775 & n19778;
  assign n19780 = ~n19774 & n19779;
  assign n19713 = n735 & ~n19175;
  assign n19771 = ~n6509 & n19188;
  assign n19772 = ~n19713 & ~n19771;
  assign n19786 = x26 & n19772;
  assign n19787 = n19780 & n19786;
  assign n19940 = ~n19785 & ~n19787;
  assign n19941 = ~n19796 & ~n19940;
  assign n19934 = x28 & n19188;
  assign n19935 = n19933 & ~n19934;
  assign n19936 = n14428 & ~n19175;
  assign n19937 = n6476 & n19188;
  assign n19938 = ~n19936 & n19937;
  assign n19939 = ~n19935 & ~n19938;
  assign n19942 = n19941 ^ n19939;
  assign n19943 = n3285 & n19748;
  assign n19944 = n3437 & n19170;
  assign n19945 = n3435 & n19173;
  assign n19946 = ~n3440 & n19174;
  assign n19947 = ~n19945 & ~n19946;
  assign n19948 = ~n19944 & n19947;
  assign n19949 = ~n19943 & n19948;
  assign n19950 = n19949 ^ x26;
  assign n19981 = n19950 ^ n19941;
  assign n19982 = n19942 & ~n19981;
  assign n19983 = n19982 ^ n19950;
  assign n20242 = n19997 ^ n19983;
  assign n20243 = n20006 & ~n20242;
  assign n20244 = n20243 ^ n20005;
  assign n20688 = n20270 ^ n20244;
  assign n20689 = ~n20271 & n20688;
  assign n20690 = n20689 ^ n20244;
  assign n20819 = n20761 ^ n20690;
  assign n20820 = n20762 & n20819;
  assign n20821 = n20820 ^ n20690;
  assign n21252 = n20871 ^ n20821;
  assign n21253 = n20872 & n21252;
  assign n21254 = n21253 ^ n20821;
  assign n21311 = n21310 ^ n21254;
  assign n20873 = n20872 ^ n20821;
  assign n19963 = n19814 ^ n19812;
  assign n19964 = ~n19200 & n19963;
  assign n19965 = n19964 ^ n19812;
  assign n19966 = n19965 ^ n19160;
  assign n20767 = n4478 & n19966;
  assign n20768 = n4487 & n19160;
  assign n20769 = n4484 & n19200;
  assign n20770 = n4480 & ~n19162;
  assign n20771 = ~n20769 & ~n20770;
  assign n20772 = ~n20768 & n20771;
  assign n20773 = ~n20767 & n20772;
  assign n20774 = n20773 ^ x23;
  assign n20273 = n4478 & n19816;
  assign n20274 = n4487 & n19200;
  assign n20275 = n4484 & ~n19162;
  assign n20276 = n4480 & ~n19201;
  assign n20277 = ~n20275 & ~n20276;
  assign n20278 = ~n20274 & n20277;
  assign n20279 = ~n20273 & n20278;
  assign n20280 = n20279 ^ x23;
  assign n20272 = n20271 ^ n20244;
  assign n20281 = n20280 ^ n20272;
  assign n20008 = n4478 & ~n19828;
  assign n20009 = n4487 & ~n19162;
  assign n20010 = n4484 & ~n19201;
  assign n20011 = n4480 & ~n19161;
  assign n20012 = ~n20010 & ~n20011;
  assign n20013 = ~n20009 & n20012;
  assign n20014 = ~n20008 & n20013;
  assign n20015 = n20014 ^ x23;
  assign n20007 = n20006 ^ n19983;
  assign n20016 = n20015 ^ n20007;
  assign n19952 = n4478 & ~n19840;
  assign n19953 = n4487 & ~n19201;
  assign n19954 = n4484 & ~n19161;
  assign n19955 = n4480 & ~n19167;
  assign n19956 = ~n19954 & ~n19955;
  assign n19957 = ~n19953 & n19956;
  assign n19958 = ~n19952 & n19957;
  assign n19959 = n19958 ^ x23;
  assign n19951 = n19950 ^ n19942;
  assign n19960 = n19959 ^ n19951;
  assign n19800 = n4478 & ~n19799;
  assign n19801 = n4487 & ~n19161;
  assign n19802 = n4484 & ~n19167;
  assign n19803 = n4480 & n19170;
  assign n19804 = ~n19802 & ~n19803;
  assign n19805 = ~n19801 & n19804;
  assign n19806 = ~n19800 & n19805;
  assign n19807 = n19806 ^ x23;
  assign n19788 = n19787 ^ n19785;
  assign n19797 = n19796 ^ n19788;
  assign n19808 = n19807 ^ n19797;
  assign n19762 = n4478 & ~n19761;
  assign n19763 = n4487 & ~n19167;
  assign n19764 = n4484 & n19170;
  assign n19765 = n4480 & n19173;
  assign n19766 = ~n19764 & ~n19765;
  assign n19767 = ~n19763 & n19766;
  assign n19768 = ~n19762 & n19767;
  assign n19769 = n19768 ^ x23;
  assign n19721 = n4478 & n19720;
  assign n19722 = n4487 & n19173;
  assign n19723 = n4484 & n19174;
  assign n19724 = n4480 & ~n19175;
  assign n19725 = ~n19723 & ~n19724;
  assign n19726 = ~n19722 & n19725;
  assign n19727 = ~n19721 & n19726;
  assign n19728 = n19727 ^ x23;
  assign n19731 = n4478 & n19730;
  assign n19732 = n4487 & n19174;
  assign n19733 = n4484 & ~n19175;
  assign n19734 = n4480 & n19188;
  assign n19735 = ~n19733 & ~n19734;
  assign n19736 = ~n19732 & n19735;
  assign n19737 = ~n19731 & n19736;
  assign n19738 = n4476 & ~n19175;
  assign n19739 = n38 & n19188;
  assign n19740 = ~n19738 & ~n19739;
  assign n19741 = x23 & n19740;
  assign n19742 = n19737 & n19741;
  assign n19743 = n735 & n19188;
  assign n19744 = ~n19742 & ~n19743;
  assign n19745 = ~n19728 & ~n19744;
  assign n19715 = n6715 & n19188;
  assign n19714 = x25 & n19188;
  assign n19716 = n19715 ^ n19714;
  assign n19717 = n19713 & ~n19716;
  assign n19718 = n19717 ^ n19715;
  assign n19746 = n19745 ^ n19718;
  assign n19749 = n4478 & n19748;
  assign n19750 = n4487 & n19170;
  assign n19751 = n4484 & n19173;
  assign n19752 = n4480 & n19174;
  assign n19753 = ~n19751 & ~n19752;
  assign n19754 = ~n19750 & n19753;
  assign n19755 = ~n19749 & n19754;
  assign n19756 = n19755 ^ x23;
  assign n19757 = n19756 ^ n19745;
  assign n19758 = ~n19746 & ~n19757;
  assign n19759 = n19758 ^ n19756;
  assign n19770 = n19769 ^ n19759;
  assign n19773 = x26 & ~n19772;
  assign n19781 = n19780 ^ n19773;
  assign n19782 = n19781 ^ n19769;
  assign n19783 = n19770 & ~n19782;
  assign n19784 = n19783 ^ n19759;
  assign n19930 = n19807 ^ n19784;
  assign n19931 = ~n19808 & n19930;
  assign n19932 = n19931 ^ n19784;
  assign n19978 = n19959 ^ n19932;
  assign n19979 = n19960 & n19978;
  assign n19980 = n19979 ^ n19932;
  assign n20239 = n20015 ^ n19980;
  assign n20240 = ~n20016 & n20239;
  assign n20241 = n20240 ^ n19980;
  assign n20764 = n20280 ^ n20241;
  assign n20765 = ~n20281 & n20764;
  assign n20766 = n20765 ^ n20241;
  assign n20775 = n20774 ^ n20766;
  assign n20763 = n20762 ^ n20690;
  assign n20816 = n20766 ^ n20763;
  assign n20817 = n20775 & n20816;
  assign n20818 = n20817 ^ n20774;
  assign n20874 = n20873 ^ n20818;
  assign n20019 = n19215 ^ n19160;
  assign n20020 = n20019 ^ n19211;
  assign n20875 = n4478 & n20020;
  assign n20876 = n4484 & n19160;
  assign n20877 = n4487 & ~n19215;
  assign n20878 = n4480 & n19200;
  assign n20879 = ~n20877 & ~n20878;
  assign n20880 = ~n20876 & n20879;
  assign n20881 = ~n20875 & n20880;
  assign n20882 = n20881 ^ x23;
  assign n21249 = n20882 ^ n20818;
  assign n21250 = n20874 & n21249;
  assign n21251 = n21250 ^ n20882;
  assign n21312 = n21311 ^ n21251;
  assign n21329 = n21328 ^ n21312;
  assign n21338 = n21337 ^ n21329;
  assign n20030 = n19230 ^ n19142;
  assign n20031 = n20030 ^ n19139;
  assign n20884 = n4673 & ~n20031;
  assign n20885 = n4688 & n19139;
  assign n20886 = n4685 & ~n19142;
  assign n20887 = ~n4681 & ~n19225;
  assign n20888 = ~n20886 & ~n20887;
  assign n20889 = ~n20885 & n20888;
  assign n20890 = ~n20884 & n20889;
  assign n20891 = n20890 ^ x20;
  assign n20883 = n20882 ^ n20874;
  assign n20892 = n20891 ^ n20883;
  assign n20776 = n20775 ^ n20763;
  assign n20282 = n20281 ^ n20241;
  assign n20017 = n20016 ^ n19980;
  assign n19961 = n19960 ^ n19932;
  assign n19817 = n4673 & n19816;
  assign n19818 = n4688 & n19200;
  assign n19819 = n4685 & ~n19162;
  assign n19820 = ~n4681 & ~n19201;
  assign n19821 = ~n19819 & ~n19820;
  assign n19822 = ~n19818 & n19821;
  assign n19823 = ~n19817 & n19822;
  assign n19824 = n19823 ^ x20;
  assign n19809 = n19808 ^ n19784;
  assign n19825 = n19824 ^ n19809;
  assign n19829 = n4673 & ~n19828;
  assign n19830 = n4688 & ~n19162;
  assign n19831 = n4685 & ~n19201;
  assign n19832 = ~n4681 & ~n19161;
  assign n19833 = ~n19831 & ~n19832;
  assign n19834 = ~n19830 & n19833;
  assign n19835 = ~n19829 & n19834;
  assign n19836 = n19835 ^ x20;
  assign n19826 = n19781 ^ n19770;
  assign n19837 = n19836 ^ n19826;
  assign n19841 = n4673 & ~n19840;
  assign n19842 = n4688 & ~n19201;
  assign n19843 = n4685 & ~n19161;
  assign n19844 = ~n4681 & ~n19167;
  assign n19845 = ~n19843 & ~n19844;
  assign n19846 = ~n19842 & n19845;
  assign n19847 = ~n19841 & n19846;
  assign n19848 = n19847 ^ x20;
  assign n19838 = n19756 ^ n19746;
  assign n19849 = n19848 ^ n19838;
  assign n19852 = n4673 & ~n19799;
  assign n19853 = n4688 & ~n19161;
  assign n19854 = n4685 & ~n19167;
  assign n19855 = ~n4681 & n19170;
  assign n19856 = ~n19854 & ~n19855;
  assign n19857 = ~n19853 & n19856;
  assign n19858 = ~n19852 & n19857;
  assign n19859 = n19858 ^ x20;
  assign n19850 = n19743 ^ n19742;
  assign n19851 = n19850 ^ n19728;
  assign n19860 = n19859 ^ n19851;
  assign n19904 = x23 & ~n19740;
  assign n19905 = n19904 ^ n19737;
  assign n19866 = n4673 & n19174;
  assign n19867 = n4681 & ~n19866;
  assign n19868 = n19188 & ~n19867;
  assign n19869 = n4688 & n19174;
  assign n19870 = ~n19868 & ~n19869;
  assign n19871 = ~n19174 & ~n19729;
  assign n19872 = ~n19176 & ~n19871;
  assign n19873 = n4673 & n19872;
  assign n19874 = n19870 & ~n19873;
  assign n19875 = n19175 & ~n19188;
  assign n19876 = ~n7059 & ~n19875;
  assign n19877 = n19874 & ~n19876;
  assign n19878 = n4476 & n19188;
  assign n19879 = ~n19877 & ~n19878;
  assign n19880 = n4673 & n19720;
  assign n19881 = n4688 & n19173;
  assign n19882 = n4685 & n19174;
  assign n19883 = ~n4681 & ~n19175;
  assign n19884 = ~n19882 & ~n19883;
  assign n19885 = ~n19881 & n19884;
  assign n19886 = ~n19880 & n19885;
  assign n19887 = x20 & ~n19886;
  assign n19888 = ~n19879 & ~n19887;
  assign n19889 = n19878 & ~n19886;
  assign n19890 = ~x20 & ~n19889;
  assign n19891 = n19888 & ~n19890;
  assign n19862 = x22 & n19188;
  assign n19861 = n7030 & n19188;
  assign n19863 = n19862 ^ n19861;
  assign n19864 = ~n19738 & ~n19863;
  assign n19865 = n19864 ^ n19862;
  assign n19892 = n19891 ^ n19865;
  assign n19893 = n4673 & n19748;
  assign n19894 = n4688 & n19170;
  assign n19895 = n4685 & n19173;
  assign n19896 = ~n4681 & n19174;
  assign n19897 = ~n19895 & ~n19896;
  assign n19898 = ~n19894 & n19897;
  assign n19899 = ~n19893 & n19898;
  assign n19900 = n19899 ^ x20;
  assign n19901 = n19900 ^ n19891;
  assign n19902 = n19892 & ~n19901;
  assign n19903 = n19902 ^ n19900;
  assign n19906 = n19905 ^ n19903;
  assign n19907 = n4673 & ~n19761;
  assign n19908 = n4688 & ~n19167;
  assign n19909 = n4685 & n19170;
  assign n19910 = ~n4681 & n19173;
  assign n19911 = ~n19909 & ~n19910;
  assign n19912 = ~n19908 & n19911;
  assign n19913 = ~n19907 & n19912;
  assign n19914 = n19913 ^ x20;
  assign n19915 = n19914 ^ n19905;
  assign n19916 = n19906 & ~n19915;
  assign n19917 = n19916 ^ n19903;
  assign n19918 = n19917 ^ n19859;
  assign n19919 = ~n19860 & n19918;
  assign n19920 = n19919 ^ n19917;
  assign n19921 = n19920 ^ n19848;
  assign n19922 = ~n19849 & n19921;
  assign n19923 = n19922 ^ n19920;
  assign n19924 = n19923 ^ n19836;
  assign n19925 = ~n19837 & n19924;
  assign n19926 = n19925 ^ n19923;
  assign n19927 = n19926 ^ n19809;
  assign n19928 = n19825 & ~n19927;
  assign n19929 = n19928 ^ n19824;
  assign n19962 = n19961 ^ n19929;
  assign n19967 = n4673 & n19966;
  assign n19968 = n4688 & n19160;
  assign n19969 = n4685 & n19200;
  assign n19970 = ~n4681 & ~n19162;
  assign n19971 = ~n19969 & ~n19970;
  assign n19972 = ~n19968 & n19971;
  assign n19973 = ~n19967 & n19972;
  assign n19974 = n19973 ^ x20;
  assign n19975 = n19974 ^ n19929;
  assign n19976 = n19962 & n19975;
  assign n19977 = n19976 ^ n19974;
  assign n20018 = n20017 ^ n19977;
  assign n20021 = n4673 & n20020;
  assign n20022 = n4685 & n19160;
  assign n20023 = n4688 & ~n19215;
  assign n20024 = ~n4681 & n19200;
  assign n20025 = ~n20023 & ~n20024;
  assign n20026 = ~n20022 & n20025;
  assign n20027 = ~n20021 & n20026;
  assign n20028 = n20027 ^ x20;
  assign n20236 = n20028 ^ n19977;
  assign n20237 = ~n20018 & n20236;
  assign n20238 = n20237 ^ n20028;
  assign n20283 = n20282 ^ n20238;
  assign n20284 = n4673 & ~n20210;
  assign n20285 = n4688 & ~n19225;
  assign n20286 = ~n4681 & n19160;
  assign n20287 = n4685 & ~n19215;
  assign n20288 = ~n20286 & ~n20287;
  assign n20289 = ~n20285 & n20288;
  assign n20290 = ~n20284 & n20289;
  assign n20291 = n20290 ^ x20;
  assign n20685 = n20291 ^ n20238;
  assign n20686 = ~n20283 & n20685;
  assign n20687 = n20686 ^ n20291;
  assign n20777 = n20776 ^ n20687;
  assign n20042 = n19228 ^ n19216;
  assign n20043 = ~n19225 & n20042;
  assign n20044 = n20043 ^ n19216;
  assign n20045 = n20044 ^ n19142;
  assign n20669 = n13653 & ~n20045;
  assign n20670 = n4685 & ~n19225;
  assign n20671 = ~n4681 & ~n19215;
  assign n20672 = ~n20670 & ~n20671;
  assign n20673 = x20 & n20672;
  assign n20674 = n19142 & n20673;
  assign n20675 = x19 & ~n20674;
  assign n20676 = ~n20669 & n20675;
  assign n20677 = n20045 & n20673;
  assign n20678 = n13653 & ~n19142;
  assign n20679 = ~x19 & ~n20678;
  assign n20680 = ~n20677 & n20679;
  assign n20681 = ~n20676 & ~n20680;
  assign n20682 = ~n13668 & n20672;
  assign n20683 = n20682 ^ x20;
  assign n20684 = ~n20681 & n20683;
  assign n20813 = n20776 ^ n20684;
  assign n20814 = ~n20777 & n20813;
  assign n20815 = n20814 ^ n20687;
  assign n21246 = n20891 ^ n20815;
  assign n21247 = n20892 & n21246;
  assign n21248 = n21247 ^ n20815;
  assign n21339 = n21338 ^ n21248;
  assign n21348 = n21347 ^ n21339;
  assign n20307 = ~n19239 & ~n19580;
  assign n20308 = n20307 ^ n19253;
  assign n20894 = n4963 & n20308;
  assign n20895 = n4972 & n19253;
  assign n20896 = n4976 & ~n19238;
  assign n20897 = n4970 & n19233;
  assign n20898 = ~n20896 & ~n20897;
  assign n20899 = ~n20895 & n20898;
  assign n20900 = ~n20894 & n20899;
  assign n20901 = n20900 ^ x17;
  assign n20893 = n20892 ^ n20815;
  assign n20902 = n20901 ^ n20893;
  assign n20327 = ~n19234 & ~n19579;
  assign n20328 = n20327 ^ n19238;
  assign n20779 = n4963 & ~n20328;
  assign n20780 = n4972 & ~n19238;
  assign n20781 = n4976 & n19233;
  assign n20782 = n4970 & n19139;
  assign n20783 = ~n20781 & ~n20782;
  assign n20784 = ~n20780 & n20783;
  assign n20785 = ~n20779 & n20784;
  assign n20786 = n20785 ^ x17;
  assign n20778 = n20777 ^ n20684;
  assign n20787 = n20786 ^ n20778;
  assign n20295 = n4963 & n20294;
  assign n20296 = n4972 & n19233;
  assign n20297 = n4976 & n19139;
  assign n20298 = n4970 & ~n19142;
  assign n20299 = ~n20297 & ~n20298;
  assign n20300 = ~n20296 & n20299;
  assign n20301 = ~n20295 & n20300;
  assign n20302 = n20301 ^ x17;
  assign n20292 = n20291 ^ n20283;
  assign n20303 = n20302 ^ n20292;
  assign n20032 = n4963 & ~n20031;
  assign n20033 = n4972 & n19139;
  assign n20034 = n4976 & ~n19142;
  assign n20035 = n4970 & ~n19225;
  assign n20036 = ~n20034 & ~n20035;
  assign n20037 = ~n20033 & n20036;
  assign n20038 = ~n20032 & n20037;
  assign n20039 = n20038 ^ x17;
  assign n20029 = n20028 ^ n20018;
  assign n20040 = n20039 ^ n20029;
  assign n20046 = n5771 & ~n20045;
  assign n20047 = n4976 & ~n19225;
  assign n20048 = n4970 & ~n19215;
  assign n20049 = ~n20047 & ~n20048;
  assign n20050 = x17 & n20049;
  assign n20051 = n19142 & n20050;
  assign n20052 = x16 & ~n20051;
  assign n20053 = ~n20046 & n20052;
  assign n20054 = n20045 & n20050;
  assign n20055 = n5771 & ~n19142;
  assign n20056 = ~x16 & ~n20055;
  assign n20057 = ~n20054 & n20056;
  assign n20058 = ~n20053 & ~n20057;
  assign n20059 = ~n5786 & n20049;
  assign n20060 = n20059 ^ x17;
  assign n20061 = ~n20058 & n20060;
  assign n20041 = n19974 ^ n19962;
  assign n20062 = n20061 ^ n20041;
  assign n20207 = n19926 ^ n19825;
  assign n20194 = n19923 ^ n19837;
  assign n20181 = n4963 & n19966;
  assign n20182 = n4972 & n19160;
  assign n20183 = n4976 & n19200;
  assign n20184 = n4970 & ~n19162;
  assign n20185 = ~n20183 & ~n20184;
  assign n20186 = ~n20182 & n20185;
  assign n20187 = ~n20181 & n20186;
  assign n20188 = n20187 ^ x17;
  assign n20064 = n4963 & n19816;
  assign n20065 = n4972 & n19200;
  assign n20066 = n4976 & ~n19162;
  assign n20067 = n4970 & ~n19201;
  assign n20068 = ~n20066 & ~n20067;
  assign n20069 = ~n20065 & n20068;
  assign n20070 = ~n20064 & n20069;
  assign n20071 = n20070 ^ x17;
  assign n20063 = n19917 ^ n19860;
  assign n20072 = n20071 ^ n20063;
  assign n20074 = n4963 & ~n19828;
  assign n20075 = n4972 & ~n19162;
  assign n20076 = n4976 & ~n19201;
  assign n20077 = n4970 & ~n19161;
  assign n20078 = ~n20076 & ~n20077;
  assign n20079 = ~n20075 & n20078;
  assign n20080 = ~n20074 & n20079;
  assign n20081 = n20080 ^ x17;
  assign n20073 = n19914 ^ n19906;
  assign n20082 = n20081 ^ n20073;
  assign n20084 = n4963 & ~n19840;
  assign n20085 = n4972 & ~n19201;
  assign n20086 = n4976 & ~n19161;
  assign n20087 = n4970 & ~n19167;
  assign n20088 = ~n20086 & ~n20087;
  assign n20089 = ~n20085 & n20088;
  assign n20090 = ~n20084 & n20089;
  assign n20091 = n20090 ^ x17;
  assign n20083 = n19900 ^ n19892;
  assign n20092 = n20091 ^ n20083;
  assign n20096 = n4963 & ~n19799;
  assign n20097 = n4972 & ~n19161;
  assign n20098 = n4976 & ~n19167;
  assign n20099 = n4970 & n19170;
  assign n20100 = ~n20098 & ~n20099;
  assign n20101 = ~n20097 & n20100;
  assign n20102 = ~n20096 & n20101;
  assign n20103 = n20102 ^ x17;
  assign n20094 = x20 & ~n19877;
  assign n20093 = n19886 ^ n19878;
  assign n20095 = n20094 ^ n20093;
  assign n20104 = n20103 ^ n20095;
  assign n20116 = n4963 & ~n19761;
  assign n20117 = n4972 & ~n19167;
  assign n20118 = n4976 & n19170;
  assign n20119 = n4970 & n19173;
  assign n20120 = ~n20118 & ~n20119;
  assign n20121 = ~n20117 & n20120;
  assign n20122 = ~n20116 & n20121;
  assign n20123 = n20122 ^ x17;
  assign n20105 = n7366 & ~n19875;
  assign n20106 = ~n4671 & ~n19175;
  assign n20107 = n20105 & ~n20106;
  assign n20108 = n4685 & ~n19175;
  assign n20109 = ~x20 & n20108;
  assign n20110 = ~n20107 & ~n20109;
  assign n20111 = n19874 & ~n20110;
  assign n20112 = n4685 & n19729;
  assign n20113 = ~n20111 & ~n20112;
  assign n20114 = ~n19874 & ~n20105;
  assign n20115 = n20113 & ~n20114;
  assign n20124 = n20123 ^ n20115;
  assign n20131 = n4963 & n19720;
  assign n20132 = n4972 & n19173;
  assign n20133 = n4976 & n19174;
  assign n20134 = n4970 & ~n19175;
  assign n20135 = ~n20133 & ~n20134;
  assign n20136 = ~n20132 & n20135;
  assign n20137 = ~n20131 & n20136;
  assign n20138 = n20137 ^ x17;
  assign n20139 = n4963 & n19730;
  assign n20140 = n4972 & n19174;
  assign n20141 = n4976 & ~n19175;
  assign n20142 = n4970 & n19188;
  assign n20143 = ~n20141 & ~n20142;
  assign n20144 = ~n20140 & n20143;
  assign n20145 = ~n20139 & n20144;
  assign n20146 = n4961 & ~n19175;
  assign n20147 = n4969 & n19188;
  assign n20148 = ~n20146 & ~n20147;
  assign n20149 = x17 & n20148;
  assign n20150 = n20145 & n20149;
  assign n20151 = n4671 & n19188;
  assign n20152 = ~n20150 & ~n20151;
  assign n20153 = ~n20138 & ~n20152;
  assign n20125 = n4671 & ~n19175;
  assign n20126 = n15624 & n19188;
  assign n20127 = ~n20125 & ~n20126;
  assign n20128 = n15622 & n19188;
  assign n20129 = ~n19175 & n20128;
  assign n20130 = ~n20127 & ~n20129;
  assign n20154 = n20153 ^ n20130;
  assign n20155 = n4963 & n19748;
  assign n20156 = n4972 & n19170;
  assign n20157 = n4976 & n19173;
  assign n20158 = n4970 & n19174;
  assign n20159 = ~n20157 & ~n20158;
  assign n20160 = ~n20156 & n20159;
  assign n20161 = ~n20155 & n20160;
  assign n20162 = n20161 ^ x17;
  assign n20163 = n20162 ^ n20153;
  assign n20164 = ~n20154 & ~n20163;
  assign n20165 = n20164 ^ n20162;
  assign n20166 = n20165 ^ n20115;
  assign n20167 = n20124 & ~n20166;
  assign n20168 = n20167 ^ n20123;
  assign n20169 = n20168 ^ n20103;
  assign n20170 = ~n20104 & n20169;
  assign n20171 = n20170 ^ n20168;
  assign n20172 = n20171 ^ n20091;
  assign n20173 = n20092 & n20172;
  assign n20174 = n20173 ^ n20171;
  assign n20175 = n20174 ^ n20081;
  assign n20176 = ~n20082 & n20175;
  assign n20177 = n20176 ^ n20174;
  assign n20178 = n20177 ^ n20071;
  assign n20179 = ~n20072 & n20178;
  assign n20180 = n20179 ^ n20177;
  assign n20189 = n20188 ^ n20180;
  assign n20190 = n19920 ^ n19849;
  assign n20191 = n20190 ^ n20180;
  assign n20192 = n20189 & ~n20191;
  assign n20193 = n20192 ^ n20188;
  assign n20195 = n20194 ^ n20193;
  assign n20196 = n4963 & n20020;
  assign n20197 = n4976 & n19160;
  assign n20198 = n4972 & ~n19215;
  assign n20199 = n4970 & n19200;
  assign n20200 = ~n20198 & ~n20199;
  assign n20201 = ~n20197 & n20200;
  assign n20202 = ~n20196 & n20201;
  assign n20203 = n20202 ^ x17;
  assign n20204 = n20203 ^ n20193;
  assign n20205 = ~n20195 & n20204;
  assign n20206 = n20205 ^ n20203;
  assign n20208 = n20207 ^ n20206;
  assign n20218 = n5771 & ~n20210;
  assign n20211 = n4970 & n19160;
  assign n20212 = n4976 & ~n19215;
  assign n20213 = ~n20211 & ~n20212;
  assign n20214 = x17 & n20213;
  assign n20219 = n19225 & n20214;
  assign n20220 = ~n20218 & ~n20219;
  assign n20215 = n20210 & n20214;
  assign n20216 = n5771 & ~n19225;
  assign n20217 = ~n20215 & ~n20216;
  assign n20221 = n20220 ^ n20217;
  assign n20222 = ~x16 & n20221;
  assign n20223 = n20222 ^ n20220;
  assign n20224 = ~n5786 & n20213;
  assign n20225 = n20224 ^ x17;
  assign n20226 = n20223 & n20225;
  assign n20227 = n20226 ^ n20206;
  assign n20228 = ~n20208 & n20227;
  assign n20229 = n20228 ^ n20226;
  assign n20230 = n20229 ^ n20061;
  assign n20231 = n20062 & n20230;
  assign n20232 = n20231 ^ n20229;
  assign n20233 = n20232 ^ n20039;
  assign n20234 = ~n20040 & n20233;
  assign n20235 = n20234 ^ n20232;
  assign n20666 = n20302 ^ n20235;
  assign n20667 = ~n20303 & n20666;
  assign n20668 = n20667 ^ n20235;
  assign n20810 = n20786 ^ n20668;
  assign n20811 = n20787 & n20810;
  assign n20812 = n20811 ^ n20668;
  assign n21243 = n20901 ^ n20812;
  assign n21244 = n20902 & n21243;
  assign n21245 = n21244 ^ n20812;
  assign n21349 = n21348 ^ n21245;
  assign n20907 = ~n19278 & ~n19584;
  assign n20908 = n20907 ^ n19281;
  assign n21227 = n6033 & ~n20908;
  assign n21228 = ~n5746 & n19277;
  assign n21229 = n5752 & n19260;
  assign n21230 = ~n21228 & ~n21229;
  assign n21231 = x14 & n21230;
  assign n21232 = n19281 & n21231;
  assign n21233 = x13 & ~n21232;
  assign n21234 = ~n21227 & n21233;
  assign n21235 = n20908 & n21231;
  assign n21236 = n6033 & ~n19281;
  assign n21237 = ~x13 & ~n21236;
  assign n21238 = ~n21235 & n21237;
  assign n21239 = ~n21234 & ~n21238;
  assign n21240 = ~n7589 & n21230;
  assign n21241 = n21240 ^ x14;
  assign n21242 = ~n21239 & n21241;
  assign n21350 = n21349 ^ n21242;
  assign n20903 = n20902 ^ n20812;
  assign n20792 = ~n19261 & ~n19583;
  assign n20793 = n20792 ^ n19277;
  assign n20794 = n6033 & n20793;
  assign n20795 = ~n5746 & n19260;
  assign n20796 = n5752 & ~n19255;
  assign n20797 = ~n20795 & ~n20796;
  assign n20798 = x14 & n20797;
  assign n20799 = ~n19277 & n20798;
  assign n20800 = x13 & ~n20799;
  assign n20801 = ~n20794 & n20800;
  assign n20802 = ~n20793 & n20798;
  assign n20803 = n6033 & n19277;
  assign n20804 = ~x13 & ~n20803;
  assign n20805 = ~n20802 & n20804;
  assign n20806 = ~n20801 & ~n20805;
  assign n20807 = ~n7589 & n20797;
  assign n20808 = n20807 ^ x14;
  assign n20809 = ~n20806 & n20808;
  assign n20904 = n20903 ^ n20809;
  assign n20656 = ~n19256 & ~n19582;
  assign n20657 = n5749 & n20656;
  assign n20658 = n20657 ^ n19260;
  assign n20659 = n5748 & n20658;
  assign n20660 = ~n5746 & ~n19255;
  assign n20661 = n5752 & n19253;
  assign n20662 = ~n20660 & ~n20661;
  assign n20663 = ~n20659 & n20662;
  assign n20664 = n20663 ^ x14;
  assign n20304 = n20303 ^ n20235;
  assign n19697 = n6033 & ~n19696;
  assign n19698 = ~n5746 & n19253;
  assign n19699 = n5752 & ~n19238;
  assign n19700 = ~n19698 & ~n19699;
  assign n19701 = x14 & n19700;
  assign n19702 = n19255 & n19701;
  assign n19703 = x13 & ~n19702;
  assign n19704 = ~n19697 & n19703;
  assign n19705 = n19696 & n19701;
  assign n19706 = n6033 & ~n19255;
  assign n19707 = ~x13 & ~n19706;
  assign n19708 = ~n19705 & n19707;
  assign n19709 = ~n19704 & ~n19708;
  assign n19710 = ~n7589 & n19700;
  assign n19711 = n19710 ^ x14;
  assign n19712 = ~n19709 & n19711;
  assign n20305 = n20304 ^ n19712;
  assign n20309 = n6033 & n20308;
  assign n20310 = ~n5746 & ~n19238;
  assign n20311 = n5752 & n19233;
  assign n20312 = ~n20310 & ~n20311;
  assign n20313 = x14 & n20312;
  assign n20314 = ~n19253 & n20313;
  assign n20315 = x13 & ~n20314;
  assign n20316 = ~n20309 & n20315;
  assign n20317 = ~n20308 & n20313;
  assign n20318 = n6033 & n19253;
  assign n20319 = ~x13 & ~n20318;
  assign n20320 = ~n20317 & n20319;
  assign n20321 = ~n20316 & ~n20320;
  assign n20322 = ~n7589 & n20312;
  assign n20323 = n20322 ^ x14;
  assign n20324 = ~n20321 & n20323;
  assign n20306 = n20232 ^ n20040;
  assign n20325 = n20324 ^ n20306;
  assign n20336 = n6033 & ~n20328;
  assign n20329 = ~n5746 & n19233;
  assign n20330 = n5752 & n19139;
  assign n20331 = ~n20329 & ~n20330;
  assign n20332 = x14 & n20331;
  assign n20337 = n19238 & n20332;
  assign n20338 = ~n20336 & ~n20337;
  assign n20333 = n20328 & n20332;
  assign n20334 = n6033 & ~n19238;
  assign n20335 = ~n20333 & ~n20334;
  assign n20339 = n20338 ^ n20335;
  assign n20340 = ~x13 & n20339;
  assign n20341 = n20340 ^ n20338;
  assign n20342 = ~n7589 & n20331;
  assign n20343 = n20342 ^ x14;
  assign n20344 = n20341 & n20343;
  assign n20326 = n20229 ^ n20062;
  assign n20345 = n20344 ^ n20326;
  assign n20354 = n6033 & n20294;
  assign n20347 = ~n5746 & n19139;
  assign n20348 = n5752 & ~n19142;
  assign n20349 = ~n20347 & ~n20348;
  assign n20350 = x14 & n20349;
  assign n20355 = ~n19233 & n20350;
  assign n20356 = ~n20354 & ~n20355;
  assign n20351 = ~n20294 & n20350;
  assign n20352 = n6033 & n19233;
  assign n20353 = ~n20351 & ~n20352;
  assign n20357 = n20356 ^ n20353;
  assign n20358 = ~x13 & n20357;
  assign n20359 = n20358 ^ n20356;
  assign n20360 = ~n7589 & n20349;
  assign n20361 = n20360 ^ x14;
  assign n20362 = n20359 & n20361;
  assign n20346 = n20226 ^ n20208;
  assign n20363 = n20362 ^ n20346;
  assign n20365 = n5749 & n20030;
  assign n20366 = n20365 ^ x13;
  assign n20367 = n20366 ^ n19139;
  assign n20368 = n5748 & n20367;
  assign n20369 = n13989 & ~n19142;
  assign n20370 = x12 & ~n20369;
  assign n20371 = n13719 & n19225;
  assign n20372 = n20370 & ~n20371;
  assign n20373 = ~x13 & ~n19225;
  assign n20374 = n14928 & ~n19142;
  assign n20375 = ~n20373 & ~n20374;
  assign n20376 = ~x12 & n20375;
  assign n20377 = ~n20372 & ~n20376;
  assign n20378 = ~n14941 & n19142;
  assign n20379 = ~n5742 & ~n5745;
  assign n20380 = ~n20378 & ~n20379;
  assign n20381 = ~n7559 & ~n20380;
  assign n20382 = ~n20377 & ~n20381;
  assign n20383 = ~n20368 & ~n20382;
  assign n20364 = n20203 ^ n20195;
  assign n20384 = n20383 ^ n20364;
  assign n20386 = n6033 & ~n20045;
  assign n20387 = ~n5746 & ~n19225;
  assign n20388 = n5752 & ~n19215;
  assign n20389 = ~n20387 & ~n20388;
  assign n20390 = x14 & n20389;
  assign n20391 = n19142 & n20390;
  assign n20392 = x13 & ~n20391;
  assign n20393 = ~n20386 & n20392;
  assign n20394 = n20045 & n20390;
  assign n20395 = n6033 & ~n19142;
  assign n20396 = ~x13 & ~n20395;
  assign n20397 = ~n20394 & n20396;
  assign n20398 = ~n20393 & ~n20397;
  assign n20399 = ~n7589 & n20389;
  assign n20400 = n20399 ^ x14;
  assign n20401 = ~n20398 & n20400;
  assign n20385 = n20190 ^ n20189;
  assign n20402 = n20401 ^ n20385;
  assign n20404 = x13 & n20209;
  assign n20405 = n20404 ^ n19225;
  assign n20406 = n6033 & ~n20405;
  assign n20407 = ~x13 & n20210;
  assign n20408 = x13 & n19225;
  assign n20409 = n7860 & ~n20408;
  assign n20410 = ~n20407 & n20409;
  assign n20411 = n5752 & n19160;
  assign n20412 = ~n5746 & ~n19215;
  assign n20413 = ~n20411 & ~n20412;
  assign n20414 = n20413 ^ x14;
  assign n20415 = ~n20410 & ~n20414;
  assign n20416 = ~n20406 & ~n20415;
  assign n20403 = n20177 ^ n20072;
  assign n20417 = n20416 ^ n20403;
  assign n20615 = n20174 ^ n20082;
  assign n20595 = n20171 ^ n20092;
  assign n20419 = n6033 & n19816;
  assign n20420 = ~n5746 & ~n19162;
  assign n20421 = n5752 & ~n19201;
  assign n20422 = ~n20420 & ~n20421;
  assign n20423 = x14 & n20422;
  assign n20424 = ~n19200 & n20423;
  assign n20425 = x13 & ~n20424;
  assign n20426 = ~n20419 & n20425;
  assign n20427 = ~n19816 & n20423;
  assign n20428 = n6033 & n19200;
  assign n20429 = ~x13 & ~n20428;
  assign n20430 = ~n20427 & n20429;
  assign n20431 = ~n20426 & ~n20430;
  assign n20432 = ~n7589 & n20422;
  assign n20433 = n20432 ^ x14;
  assign n20434 = ~n20431 & n20433;
  assign n20418 = n20168 ^ n20104;
  assign n20435 = n20434 ^ n20418;
  assign n20437 = n6033 & ~n19828;
  assign n20438 = ~n5746 & ~n19201;
  assign n20439 = n5752 & ~n19161;
  assign n20440 = ~n20438 & ~n20439;
  assign n20441 = x14 & n20440;
  assign n20442 = n19162 & n20441;
  assign n20443 = ~n20437 & ~n20442;
  assign n20444 = x13 & n20443;
  assign n20445 = n19828 & n20441;
  assign n20446 = n6033 & ~n19162;
  assign n20447 = ~x13 & ~n20446;
  assign n20448 = ~n20445 & n20447;
  assign n20449 = ~n20444 & ~n20448;
  assign n20450 = ~n7589 & n20440;
  assign n20451 = n20450 ^ x14;
  assign n20452 = ~n20449 & n20451;
  assign n20436 = n20165 ^ n20124;
  assign n20453 = n20452 ^ n20436;
  assign n20455 = ~n5746 & ~n19161;
  assign n20456 = n5752 & ~n19167;
  assign n20457 = ~n20455 & ~n20456;
  assign n20458 = x14 & n20457;
  assign n20459 = n19839 & n20458;
  assign n20460 = ~n6033 & ~n20459;
  assign n20461 = x13 & n19839;
  assign n20462 = ~n19201 & ~n20461;
  assign n20463 = ~n20460 & n20462;
  assign n20464 = n6033 & n19839;
  assign n20465 = ~n20458 & ~n20464;
  assign n20466 = ~x13 & n19839;
  assign n20467 = ~n20465 & ~n20466;
  assign n20468 = n19201 & n20467;
  assign n20469 = ~n20463 & ~n20468;
  assign n20470 = ~n7589 & n20457;
  assign n20471 = n20470 ^ x14;
  assign n20472 = n20469 & n20471;
  assign n20454 = n20162 ^ n20154;
  assign n20473 = n20472 ^ n20454;
  assign n20476 = n19180 & ~n19194;
  assign n20477 = ~x13 & n19798;
  assign n20478 = ~n6033 & ~n19161;
  assign n20479 = ~n20477 & ~n20478;
  assign n20480 = n20479 ^ x13;
  assign n20481 = ~n20476 & ~n20480;
  assign n20482 = n20481 ^ x13;
  assign n20486 = n19161 & ~n19798;
  assign n20487 = n5748 & ~n20486;
  assign n20483 = ~n5746 & ~n19167;
  assign n20484 = n5752 & n19170;
  assign n20485 = ~n20483 & ~n20484;
  assign n20488 = n20487 ^ n20485;
  assign n20489 = x14 & n20488;
  assign n20490 = n20489 ^ n20487;
  assign n20491 = ~n20482 & n20490;
  assign n20492 = x14 & ~n20485;
  assign n20493 = ~n7559 & n20485;
  assign n20494 = ~n20492 & ~n20493;
  assign n20495 = ~n20491 & ~n20494;
  assign n20474 = n20151 ^ n20150;
  assign n20475 = n20474 ^ n20138;
  assign n20496 = n20495 ^ n20475;
  assign n20499 = n6033 & ~n19761;
  assign n20500 = ~n5746 & n19170;
  assign n20501 = n5752 & n19173;
  assign n20502 = ~n20500 & ~n20501;
  assign n20503 = x14 & n20502;
  assign n20504 = n19167 & n20503;
  assign n20505 = x13 & ~n20504;
  assign n20506 = ~n20499 & n20505;
  assign n20507 = n19761 & n20503;
  assign n20508 = n6033 & ~n19167;
  assign n20509 = ~x13 & ~n20508;
  assign n20510 = ~n20507 & n20509;
  assign n20511 = ~n20506 & ~n20510;
  assign n20512 = ~n7589 & n20502;
  assign n20513 = n20512 ^ x14;
  assign n20514 = ~n20511 & n20513;
  assign n20497 = x17 & ~n20148;
  assign n20498 = n20497 ^ n20145;
  assign n20515 = n20514 ^ n20498;
  assign n20521 = n6033 & n19720;
  assign n20522 = ~n5746 & n19174;
  assign n20523 = n5752 & ~n19175;
  assign n20524 = ~n20522 & ~n20523;
  assign n20525 = x14 & n20524;
  assign n20526 = ~n19173 & n20525;
  assign n20527 = ~n20521 & ~n20526;
  assign n20528 = x13 & n20527;
  assign n20529 = ~n19720 & n20525;
  assign n20530 = n6033 & n19173;
  assign n20531 = ~x13 & ~n20530;
  assign n20532 = ~n20529 & n20531;
  assign n20533 = ~n20528 & ~n20532;
  assign n20534 = ~n7589 & n20524;
  assign n20535 = n20534 ^ x14;
  assign n20536 = ~n20533 & n20535;
  assign n20537 = n6033 & ~n19871;
  assign n20538 = n19174 & ~n19729;
  assign n20539 = ~n5746 & ~n19175;
  assign n20540 = n5752 & n19188;
  assign n20541 = ~n20539 & ~n20540;
  assign n20542 = x14 & n20541;
  assign n20543 = ~n20538 & n20542;
  assign n20544 = ~n20537 & ~n20543;
  assign n20545 = n19174 ^ x13;
  assign n20546 = n19729 & ~n20545;
  assign n20547 = ~n20544 & ~n20546;
  assign n20548 = ~n7589 & n20541;
  assign n20549 = n20548 ^ x14;
  assign n20550 = ~n20547 & n20549;
  assign n20551 = n5748 & ~n19175;
  assign n20552 = n5746 & ~n5748;
  assign n20553 = n19188 & ~n20552;
  assign n20554 = x14 & ~n20553;
  assign n20555 = ~n20551 & n20554;
  assign n20556 = ~n20550 & n20555;
  assign n20557 = n4961 & n19188;
  assign n20558 = ~n20556 & ~n20557;
  assign n20559 = ~n20536 & ~n20558;
  assign n20517 = x16 & n19188;
  assign n20516 = n16092 & n19188;
  assign n20518 = n20517 ^ n20516;
  assign n20519 = ~n20146 & ~n20518;
  assign n20520 = n20519 ^ n20517;
  assign n20560 = n20559 ^ n20520;
  assign n20561 = n6033 & n19748;
  assign n20562 = ~n5746 & n19173;
  assign n20563 = n5752 & n19174;
  assign n20564 = ~n20562 & ~n20563;
  assign n20565 = x14 & n20564;
  assign n20566 = ~n19170 & n20565;
  assign n20567 = x13 & ~n20566;
  assign n20568 = ~n20561 & n20567;
  assign n20569 = ~n19748 & n20565;
  assign n20570 = n6033 & n19170;
  assign n20571 = ~x13 & ~n20570;
  assign n20572 = ~n20569 & n20571;
  assign n20573 = ~n20568 & ~n20572;
  assign n20574 = ~n7589 & n20564;
  assign n20575 = n20574 ^ x14;
  assign n20576 = ~n20573 & n20575;
  assign n20577 = n20576 ^ n20559;
  assign n20578 = n20560 & ~n20577;
  assign n20579 = n20578 ^ n20576;
  assign n20580 = n20579 ^ n20498;
  assign n20581 = n20515 & ~n20580;
  assign n20582 = n20581 ^ n20514;
  assign n20583 = n20582 ^ n20475;
  assign n20584 = n20496 & ~n20583;
  assign n20585 = n20584 ^ n20495;
  assign n20586 = n20585 ^ n20472;
  assign n20587 = ~n20473 & n20586;
  assign n20588 = n20587 ^ n20585;
  assign n20589 = n20588 ^ n20452;
  assign n20590 = ~n20453 & n20589;
  assign n20591 = n20590 ^ n20588;
  assign n20592 = n20591 ^ n20434;
  assign n20593 = ~n20435 & n20592;
  assign n20594 = n20593 ^ n20591;
  assign n20596 = n20595 ^ n20594;
  assign n20597 = n13989 & ~n19966;
  assign n20598 = n14928 & ~n19160;
  assign n20599 = ~n5746 & n19200;
  assign n20600 = n5752 & ~n19162;
  assign n20601 = ~n20599 & ~n20600;
  assign n20602 = ~n7559 & n20601;
  assign n20603 = ~n20598 & n20602;
  assign n20604 = ~n20597 & n20603;
  assign n20605 = x14 & ~n20601;
  assign n20606 = ~n20604 & ~n20605;
  assign n20607 = x13 & ~n19966;
  assign n20608 = ~x13 & ~n19160;
  assign n20609 = n6033 & ~n20608;
  assign n20610 = ~n20607 & n20609;
  assign n20611 = ~n20606 & ~n20610;
  assign n20612 = n20611 ^ n20594;
  assign n20613 = n20596 & n20612;
  assign n20614 = n20613 ^ n20611;
  assign n20616 = n20615 ^ n20614;
  assign n20617 = n13989 & ~n20020;
  assign n20618 = ~n5746 & n19160;
  assign n20619 = n5752 & n19200;
  assign n20620 = ~n20618 & ~n20619;
  assign n20621 = ~n7559 & n20620;
  assign n20622 = n14928 & n19215;
  assign n20623 = n20621 & ~n20622;
  assign n20624 = ~n20617 & n20623;
  assign n20625 = x14 & ~n20620;
  assign n20626 = ~n20624 & ~n20625;
  assign n20627 = x13 & ~n20020;
  assign n20628 = ~x13 & n19215;
  assign n20629 = n6033 & ~n20628;
  assign n20630 = ~n20627 & n20629;
  assign n20631 = ~n20626 & ~n20630;
  assign n20632 = n20631 ^ n20614;
  assign n20633 = ~n20616 & n20632;
  assign n20634 = n20633 ^ n20631;
  assign n20635 = n20634 ^ n20403;
  assign n20636 = n20417 & ~n20635;
  assign n20637 = n20636 ^ n20416;
  assign n20638 = n20637 ^ n20401;
  assign n20639 = ~n20402 & n20638;
  assign n20640 = n20639 ^ n20637;
  assign n20641 = n20640 ^ n20383;
  assign n20642 = ~n20384 & n20641;
  assign n20643 = n20642 ^ n20640;
  assign n20644 = n20643 ^ n20362;
  assign n20645 = ~n20363 & n20644;
  assign n20646 = n20645 ^ n20643;
  assign n20647 = n20646 ^ n20344;
  assign n20648 = n20345 & n20647;
  assign n20649 = n20648 ^ n20646;
  assign n20650 = n20649 ^ n20324;
  assign n20651 = ~n20325 & n20650;
  assign n20652 = n20651 ^ n20649;
  assign n20653 = n20652 ^ n20304;
  assign n20654 = ~n20305 & n20653;
  assign n20655 = n20654 ^ n20652;
  assign n20665 = n20664 ^ n20655;
  assign n20788 = n20787 ^ n20668;
  assign n20789 = n20788 ^ n20664;
  assign n20790 = n20665 & n20789;
  assign n20791 = n20790 ^ n20655;
  assign n21224 = n20903 ^ n20791;
  assign n21225 = n20904 & ~n21224;
  assign n21226 = n21225 ^ n20791;
  assign n21351 = n21350 ^ n21226;
  assign n21214 = ~n19287 & ~n19587;
  assign n21215 = n21214 ^ n19104;
  assign n21216 = n5814 & n21215;
  assign n21217 = n6295 & n19104;
  assign n21218 = n5824 & n19122;
  assign n21219 = n5817 & ~n19286;
  assign n21220 = ~n21218 & ~n21219;
  assign n21221 = ~n21217 & n21220;
  assign n21222 = ~n21216 & n21221;
  assign n21223 = n21222 ^ x11;
  assign n21352 = n21351 ^ n21223;
  assign n20905 = n20904 ^ n20791;
  assign n19677 = ~n19283 & ~n19586;
  assign n19678 = n19677 ^ n19286;
  assign n19679 = n7536 & ~n19678;
  assign n19680 = n5817 & n19122;
  assign n19681 = n5824 & ~n19281;
  assign n19682 = ~n19680 & ~n19681;
  assign n19683 = x11 & n19682;
  assign n19684 = n19286 & n19683;
  assign n19685 = ~n19679 & ~n19684;
  assign n19686 = x10 & n19685;
  assign n19687 = n19678 & n19683;
  assign n19688 = n7536 & ~n19286;
  assign n19689 = ~x10 & ~n19688;
  assign n19690 = ~n19687 & n19689;
  assign n19691 = ~n19686 & ~n19690;
  assign n19692 = ~n7551 & n19682;
  assign n19693 = n19692 ^ x11;
  assign n19694 = ~n19691 & n19693;
  assign n20906 = n20905 ^ n19694;
  assign n21188 = ~n19282 & ~n19585;
  assign n21189 = n21188 ^ n19122;
  assign n21190 = n7536 & n21189;
  assign n21191 = n5817 & ~n19281;
  assign n21192 = n5824 & n19277;
  assign n21193 = ~n21191 & ~n21192;
  assign n21194 = x11 & n21193;
  assign n21195 = ~n19122 & n21194;
  assign n21196 = x10 & ~n21195;
  assign n21197 = ~n21190 & n21196;
  assign n21198 = ~n21189 & n21194;
  assign n21199 = n7536 & n19122;
  assign n21200 = ~x10 & ~n21199;
  assign n21201 = ~n21198 & n21200;
  assign n21202 = ~n21197 & ~n21201;
  assign n21203 = ~n7551 & n21193;
  assign n21204 = n21203 ^ x11;
  assign n21205 = ~n21202 & n21204;
  assign n20917 = n20652 ^ n20305;
  assign n20909 = n5814 & ~n20908;
  assign n20910 = n6295 & ~n19281;
  assign n20911 = n5817 & n19277;
  assign n20912 = n5824 & n19260;
  assign n20913 = ~n20911 & ~n20912;
  assign n20914 = ~n20910 & n20913;
  assign n20915 = ~n20909 & n20914;
  assign n20916 = n20915 ^ x11;
  assign n20918 = n20917 ^ n20916;
  assign n20927 = n20649 ^ n20325;
  assign n20919 = n5814 & n20793;
  assign n20920 = n6295 & n19277;
  assign n20921 = n5817 & n19260;
  assign n20922 = n5824 & ~n19255;
  assign n20923 = ~n20921 & ~n20922;
  assign n20924 = ~n20920 & n20923;
  assign n20925 = ~n20919 & n20924;
  assign n20926 = n20925 ^ x11;
  assign n20928 = n20927 ^ n20926;
  assign n20946 = n20646 ^ n20345;
  assign n20929 = n20656 ^ n19260;
  assign n20930 = n7536 & n20929;
  assign n20931 = n5817 & ~n19255;
  assign n20932 = n5824 & n19253;
  assign n20933 = ~n20931 & ~n20932;
  assign n20934 = x11 & n20933;
  assign n20935 = ~n19260 & n20934;
  assign n20936 = x10 & ~n20935;
  assign n20937 = ~n20930 & n20936;
  assign n20938 = ~n20929 & n20934;
  assign n20939 = n7536 & n19260;
  assign n20940 = ~x10 & ~n20939;
  assign n20941 = ~n20938 & n20940;
  assign n20942 = ~n20937 & ~n20941;
  assign n20943 = ~n7551 & n20933;
  assign n20944 = n20943 ^ x11;
  assign n20945 = ~n20942 & n20944;
  assign n20947 = n20946 ^ n20945;
  assign n20956 = n20643 ^ n20363;
  assign n20948 = n5814 & ~n19696;
  assign n20949 = n6295 & ~n19255;
  assign n20950 = n5817 & n19253;
  assign n20951 = n5824 & ~n19238;
  assign n20952 = ~n20950 & ~n20951;
  assign n20953 = ~n20949 & n20952;
  assign n20954 = ~n20948 & n20953;
  assign n20955 = n20954 ^ x11;
  assign n20957 = n20956 ^ n20955;
  assign n20966 = n20640 ^ n20384;
  assign n20958 = n5814 & n20308;
  assign n20959 = n6295 & n19253;
  assign n20960 = n5817 & ~n19238;
  assign n20961 = n5824 & n19233;
  assign n20962 = ~n20960 & ~n20961;
  assign n20963 = ~n20959 & n20962;
  assign n20964 = ~n20958 & n20963;
  assign n20965 = n20964 ^ x11;
  assign n20967 = n20966 ^ n20965;
  assign n20969 = n5814 & ~n20328;
  assign n20970 = n6295 & ~n19238;
  assign n20971 = n5817 & n19233;
  assign n20972 = n5824 & n19139;
  assign n20973 = ~n20971 & ~n20972;
  assign n20974 = ~n20970 & n20973;
  assign n20975 = ~n20969 & n20974;
  assign n20976 = n20975 ^ x11;
  assign n20968 = n20637 ^ n20402;
  assign n20977 = n20976 ^ n20968;
  assign n20979 = n5814 & n20294;
  assign n20980 = n6295 & n19233;
  assign n20981 = n5817 & n19139;
  assign n20982 = n5824 & ~n19142;
  assign n20983 = ~n20981 & ~n20982;
  assign n20984 = ~n20980 & n20983;
  assign n20985 = ~n20979 & n20984;
  assign n20986 = n20985 ^ x11;
  assign n20978 = n20634 ^ n20417;
  assign n20987 = n20986 ^ n20978;
  assign n20989 = n5814 & ~n20031;
  assign n20990 = n6295 & n19139;
  assign n20991 = n5817 & ~n19142;
  assign n20992 = n5824 & ~n19225;
  assign n20993 = ~n20991 & ~n20992;
  assign n20994 = ~n20990 & n20993;
  assign n20995 = ~n20989 & n20994;
  assign n20996 = n20995 ^ x11;
  assign n20988 = n20631 ^ n20616;
  assign n20997 = n20996 ^ n20988;
  assign n20999 = n5814 & ~n20045;
  assign n21000 = n6295 & ~n19142;
  assign n21001 = n5824 & ~n19215;
  assign n21002 = ~n21000 & ~n21001;
  assign n21003 = n5817 & ~n19225;
  assign n21004 = n21002 & ~n21003;
  assign n21005 = ~n20999 & n21004;
  assign n21006 = n21005 ^ x11;
  assign n20998 = n20611 ^ n20596;
  assign n21007 = n21006 ^ n20998;
  assign n21140 = n20591 ^ n20435;
  assign n21127 = n5814 & n20020;
  assign n21128 = n5817 & n19160;
  assign n21129 = n6295 & ~n19215;
  assign n21130 = n5824 & n19200;
  assign n21131 = ~n21129 & ~n21130;
  assign n21132 = ~n21128 & n21131;
  assign n21133 = ~n21127 & n21132;
  assign n21134 = n21133 ^ x11;
  assign n21114 = n5814 & n19966;
  assign n21115 = n6295 & n19160;
  assign n21116 = n5817 & n19200;
  assign n21117 = n5824 & ~n19162;
  assign n21118 = ~n21116 & ~n21117;
  assign n21119 = ~n21115 & n21118;
  assign n21120 = ~n21114 & n21119;
  assign n21121 = n21120 ^ x11;
  assign n21009 = n5814 & n19816;
  assign n21010 = n6295 & n19200;
  assign n21011 = n5817 & ~n19162;
  assign n21012 = n5824 & ~n19201;
  assign n21013 = ~n21011 & ~n21012;
  assign n21014 = ~n21010 & n21013;
  assign n21015 = ~n21009 & n21014;
  assign n21016 = n21015 ^ x11;
  assign n21008 = n20582 ^ n20496;
  assign n21017 = n21016 ^ n21008;
  assign n21019 = n5814 & ~n19828;
  assign n21020 = n6295 & ~n19162;
  assign n21021 = n5817 & ~n19201;
  assign n21022 = n5824 & ~n19161;
  assign n21023 = ~n21021 & ~n21022;
  assign n21024 = ~n21020 & n21023;
  assign n21025 = ~n21019 & n21024;
  assign n21026 = n21025 ^ x11;
  assign n21018 = n20579 ^ n20515;
  assign n21027 = n21026 ^ n21018;
  assign n21029 = n5814 & ~n19840;
  assign n21030 = n6295 & ~n19201;
  assign n21031 = n5817 & ~n19161;
  assign n21032 = n5824 & ~n19167;
  assign n21033 = ~n21031 & ~n21032;
  assign n21034 = ~n21030 & n21033;
  assign n21035 = ~n21029 & n21034;
  assign n21036 = n21035 ^ x11;
  assign n21028 = n20576 ^ n20560;
  assign n21037 = n21036 ^ n21028;
  assign n21040 = n5814 & ~n19799;
  assign n21041 = n6295 & ~n19161;
  assign n21042 = n5817 & ~n19167;
  assign n21043 = n5824 & n19170;
  assign n21044 = ~n21042 & ~n21043;
  assign n21045 = ~n21041 & n21044;
  assign n21046 = ~n21040 & n21045;
  assign n21047 = n21046 ^ x11;
  assign n21038 = n20557 ^ n20556;
  assign n21039 = n21038 ^ n20536;
  assign n21048 = n21047 ^ n21039;
  assign n21089 = n20555 ^ n20550;
  assign n21056 = n5814 & n19872;
  assign n21057 = n6295 & n19174;
  assign n21058 = ~n21056 & ~n21057;
  assign n21059 = n5814 & n19174;
  assign n21060 = ~n5824 & ~n21059;
  assign n21061 = n19188 & ~n21060;
  assign n21062 = n21058 & ~n21061;
  assign n21063 = x11 & n21062;
  assign n21064 = n5823 & ~n19875;
  assign n21065 = n21063 & ~n21064;
  assign n21066 = n5748 & n19188;
  assign n21067 = ~n21065 & ~n21066;
  assign n21068 = n5814 & n19720;
  assign n21069 = n6295 & n19173;
  assign n21070 = n5817 & n19174;
  assign n21071 = n5824 & ~n19175;
  assign n21072 = ~n21070 & ~n21071;
  assign n21073 = ~n21069 & n21072;
  assign n21074 = ~n21068 & n21073;
  assign n21075 = n21074 ^ x11;
  assign n21076 = ~n21067 & ~n21075;
  assign n21049 = ~n5744 & ~n19175;
  assign n21050 = n8210 & ~n21049;
  assign n21051 = ~n5743 & ~n21050;
  assign n21052 = n19188 & ~n21051;
  assign n21053 = x13 & n19188;
  assign n21054 = n20551 & ~n21053;
  assign n21055 = ~n21052 & ~n21054;
  assign n21077 = n21076 ^ n21055;
  assign n21078 = n5814 & n19748;
  assign n21079 = n6295 & n19170;
  assign n21080 = n5817 & n19173;
  assign n21081 = n5824 & n19174;
  assign n21082 = ~n21080 & ~n21081;
  assign n21083 = ~n21079 & n21082;
  assign n21084 = ~n21078 & n21083;
  assign n21085 = n21084 ^ x11;
  assign n21086 = n21085 ^ n21076;
  assign n21087 = n21077 & ~n21086;
  assign n21088 = n21087 ^ n21085;
  assign n21090 = n21089 ^ n21088;
  assign n21091 = n5814 & ~n19761;
  assign n21092 = n6295 & ~n19167;
  assign n21093 = n5817 & n19170;
  assign n21094 = n5824 & n19173;
  assign n21095 = ~n21093 & ~n21094;
  assign n21096 = ~n21092 & n21095;
  assign n21097 = ~n21091 & n21096;
  assign n21098 = n21097 ^ x11;
  assign n21099 = n21098 ^ n21088;
  assign n21100 = ~n21090 & n21099;
  assign n21101 = n21100 ^ n21098;
  assign n21102 = n21101 ^ n21047;
  assign n21103 = ~n21048 & n21102;
  assign n21104 = n21103 ^ n21101;
  assign n21105 = n21104 ^ n21036;
  assign n21106 = n21037 & n21105;
  assign n21107 = n21106 ^ n21104;
  assign n21108 = n21107 ^ n21026;
  assign n21109 = ~n21027 & n21108;
  assign n21110 = n21109 ^ n21107;
  assign n21111 = n21110 ^ n21016;
  assign n21112 = ~n21017 & n21111;
  assign n21113 = n21112 ^ n21110;
  assign n21122 = n21121 ^ n21113;
  assign n21123 = n20585 ^ n20473;
  assign n21124 = n21123 ^ n21113;
  assign n21125 = n21122 & ~n21124;
  assign n21126 = n21125 ^ n21121;
  assign n21135 = n21134 ^ n21126;
  assign n21136 = n20588 ^ n20453;
  assign n21137 = n21136 ^ n21126;
  assign n21138 = n21135 & ~n21137;
  assign n21139 = n21138 ^ n21134;
  assign n21141 = n21140 ^ n21139;
  assign n21149 = n7536 & ~n20210;
  assign n21142 = n5824 & n19160;
  assign n21143 = n5817 & ~n19215;
  assign n21144 = ~n21142 & ~n21143;
  assign n21145 = x11 & n21144;
  assign n21150 = n19225 & n21145;
  assign n21151 = ~n21149 & ~n21150;
  assign n21146 = n20210 & n21145;
  assign n21147 = n7536 & ~n19225;
  assign n21148 = ~n21146 & ~n21147;
  assign n21152 = n21151 ^ n21148;
  assign n21153 = ~x10 & n21152;
  assign n21154 = n21153 ^ n21151;
  assign n21155 = ~n7551 & n21144;
  assign n21156 = n21155 ^ x11;
  assign n21157 = n21154 & n21156;
  assign n21158 = n21157 ^ n21139;
  assign n21159 = ~n21141 & n21158;
  assign n21160 = n21159 ^ n21157;
  assign n21161 = n21160 ^ n21006;
  assign n21162 = n21007 & n21161;
  assign n21163 = n21162 ^ n21160;
  assign n21164 = n21163 ^ n20996;
  assign n21165 = ~n20997 & n21164;
  assign n21166 = n21165 ^ n21163;
  assign n21167 = n21166 ^ n20986;
  assign n21168 = ~n20987 & n21167;
  assign n21169 = n21168 ^ n21166;
  assign n21170 = n21169 ^ n20976;
  assign n21171 = ~n20977 & n21170;
  assign n21172 = n21171 ^ n21169;
  assign n21173 = n21172 ^ n20966;
  assign n21174 = ~n20967 & n21173;
  assign n21175 = n21174 ^ n21172;
  assign n21176 = n21175 ^ n20956;
  assign n21177 = ~n20957 & n21176;
  assign n21178 = n21177 ^ n21175;
  assign n21179 = n21178 ^ n20946;
  assign n21180 = n20947 & ~n21179;
  assign n21181 = n21180 ^ n21178;
  assign n21182 = n21181 ^ n20927;
  assign n21183 = ~n20928 & n21182;
  assign n21184 = n21183 ^ n21181;
  assign n21185 = n21184 ^ n20917;
  assign n21186 = ~n20918 & n21185;
  assign n21187 = n21186 ^ n21184;
  assign n21206 = n21205 ^ n21187;
  assign n21207 = n20788 ^ n20665;
  assign n21208 = n21207 ^ n21205;
  assign n21209 = n21206 & n21208;
  assign n21210 = n21209 ^ n21187;
  assign n21211 = n21210 ^ n20905;
  assign n21212 = n20906 & ~n21211;
  assign n21213 = n21212 ^ n21210;
  assign n21864 = n21351 ^ n21213;
  assign n21865 = n21352 & ~n21864;
  assign n21866 = n21865 ^ n21213;
  assign n21875 = n21874 ^ n21866;
  assign n21850 = n4673 & ~n20328;
  assign n21851 = n4688 & ~n19238;
  assign n21852 = n4685 & n19233;
  assign n21853 = ~n4681 & n19139;
  assign n21854 = ~n21852 & ~n21853;
  assign n21855 = ~n21851 & n21854;
  assign n21856 = ~n21850 & n21855;
  assign n21857 = n21856 ^ x20;
  assign n21832 = n12502 & ~n20045;
  assign n21833 = n4484 & ~n19225;
  assign n21834 = n4480 & ~n19215;
  assign n21835 = ~n21833 & ~n21834;
  assign n21836 = x23 & n21835;
  assign n21837 = n19142 & n21836;
  assign n21838 = x22 & ~n21837;
  assign n21839 = ~n21832 & n21838;
  assign n21840 = n20045 & n21836;
  assign n21841 = n12502 & ~n19142;
  assign n21842 = ~x22 & ~n21841;
  assign n21843 = ~n21840 & n21842;
  assign n21844 = ~n21839 & ~n21843;
  assign n21845 = ~n12519 & n21835;
  assign n21846 = n21845 ^ x23;
  assign n21847 = ~n21844 & n21846;
  assign n21820 = n44 & ~n19840;
  assign n21821 = n3280 & ~n19201;
  assign n21822 = n3277 & ~n19161;
  assign n21823 = n3275 & ~n19167;
  assign n21824 = ~n21822 & ~n21823;
  assign n21825 = ~n21821 & n21824;
  assign n21826 = ~n21820 & n21825;
  assign n21827 = n21826 ^ x29;
  assign n21808 = n41 & n19748;
  assign n21809 = n91 & n19173;
  assign n21810 = x31 & ~n21286;
  assign n21811 = ~n21809 & n21810;
  assign n21812 = ~n21808 & n21811;
  assign n21813 = n41 & n19170;
  assign n21814 = n54 & n19173;
  assign n21815 = ~x31 & ~n21814;
  assign n21816 = ~n21813 & n21815;
  assign n21817 = ~n21812 & ~n21816;
  assign n11968 = n236 & n3263;
  assign n11969 = n986 & n11968;
  assign n11971 = n4077 & n4736;
  assign n11972 = n11970 & n11971;
  assign n11973 = ~n319 & ~n370;
  assign n11974 = ~n659 & n11973;
  assign n11975 = n1723 & n3064;
  assign n11976 = n11974 & n11975;
  assign n11977 = n11972 & n11976;
  assign n11978 = n11969 & n11977;
  assign n11002 = n1274 & n11001;
  assign n11003 = n1205 & n11002;
  assign n11004 = ~n248 & ~n303;
  assign n11005 = n5449 & n11004;
  assign n11006 = n5384 & n11005;
  assign n11007 = n11003 & n11006;
  assign n21793 = ~n301 & ~n313;
  assign n21794 = ~n155 & n21793;
  assign n21795 = ~n202 & ~n417;
  assign n21796 = n1688 & n21795;
  assign n21797 = n21794 & n21796;
  assign n21798 = ~n64 & ~n104;
  assign n21799 = n12229 & n21798;
  assign n21800 = n437 & n2202;
  assign n21801 = n21799 & n21800;
  assign n21802 = n21797 & n21801;
  assign n10978 = ~n517 & ~n710;
  assign n10979 = ~n193 & ~n378;
  assign n10980 = n10978 & n10979;
  assign n10981 = ~n323 & ~n582;
  assign n10982 = n3039 & n10981;
  assign n10983 = n10980 & n10982;
  assign n21803 = n10983 & n13270;
  assign n21804 = n21802 & n21803;
  assign n21805 = n11007 & n21804;
  assign n21806 = n11978 & n21805;
  assign n21807 = n13366 & n21806;
  assign n21818 = n21817 ^ n21807;
  assign n21790 = n21289 ^ n21260;
  assign n21791 = n21290 & ~n21790;
  assign n21792 = n21791 ^ n21260;
  assign n21819 = n21818 ^ n21792;
  assign n21828 = n21827 ^ n21819;
  assign n21787 = n21291 ^ n21257;
  assign n21788 = ~n21300 & n21787;
  assign n21789 = n21788 ^ n21299;
  assign n21829 = n21828 ^ n21789;
  assign n21784 = n21309 ^ n21254;
  assign n21785 = n21310 & n21784;
  assign n21786 = n21785 ^ n21254;
  assign n21830 = n21829 ^ n21786;
  assign n21776 = n3285 & n19966;
  assign n21777 = n3437 & n19160;
  assign n21778 = n3435 & n19200;
  assign n21779 = ~n3440 & ~n19162;
  assign n21780 = ~n21778 & ~n21779;
  assign n21781 = ~n21777 & n21780;
  assign n21782 = ~n21776 & n21781;
  assign n21783 = n21782 ^ x26;
  assign n21831 = n21830 ^ n21783;
  assign n21848 = n21847 ^ n21831;
  assign n21773 = n21328 ^ n21251;
  assign n21774 = n21312 & n21773;
  assign n21775 = n21774 ^ n21328;
  assign n21849 = n21848 ^ n21775;
  assign n21858 = n21857 ^ n21849;
  assign n21770 = n21337 ^ n21248;
  assign n21771 = n21338 & n21770;
  assign n21772 = n21771 ^ n21248;
  assign n21859 = n21858 ^ n21772;
  assign n21754 = n5771 & n20929;
  assign n21755 = n4976 & ~n19255;
  assign n21756 = n4970 & n19253;
  assign n21757 = ~n21755 & ~n21756;
  assign n21758 = x17 & n21757;
  assign n21759 = ~n19260 & n21758;
  assign n21760 = x16 & ~n21759;
  assign n21761 = ~n21754 & n21760;
  assign n21762 = ~n20929 & n21758;
  assign n21763 = n5771 & n19260;
  assign n21764 = ~x16 & ~n21763;
  assign n21765 = ~n21762 & n21764;
  assign n21766 = ~n21761 & ~n21765;
  assign n21767 = ~n5786 & n21757;
  assign n21768 = n21767 ^ x17;
  assign n21769 = ~n21766 & n21768;
  assign n21860 = n21859 ^ n21769;
  assign n21751 = n21347 ^ n21245;
  assign n21752 = n21348 & n21751;
  assign n21753 = n21752 ^ n21245;
  assign n21861 = n21860 ^ n21753;
  assign n21736 = ~x13 & n21189;
  assign n21737 = x13 & n19122;
  assign n21738 = x14 & ~n21737;
  assign n21739 = ~n21736 & n21738;
  assign n21740 = ~n5746 & ~n19281;
  assign n21741 = n5752 & n19277;
  assign n21742 = ~n21740 & ~n21741;
  assign n21743 = ~n7559 & n21742;
  assign n21744 = ~n21739 & n21743;
  assign n21745 = x14 & ~n21742;
  assign n21746 = ~n21744 & ~n21745;
  assign n21747 = x13 & n21188;
  assign n21748 = n21747 ^ n19122;
  assign n21749 = n6033 & n21748;
  assign n21750 = ~n21746 & ~n21749;
  assign n21862 = n21861 ^ n21750;
  assign n21733 = n21349 ^ n21226;
  assign n21734 = n21350 & ~n21733;
  assign n21735 = n21734 ^ n21226;
  assign n21863 = n21862 ^ n21735;
  assign n21876 = n21875 ^ n21863;
  assign n19079 = n18837 ^ n12696;
  assign n19080 = n12696 ^ n12523;
  assign n19081 = ~n19079 & ~n19080;
  assign n19082 = n19081 ^ n18837;
  assign n19083 = n18845 & ~n19082;
  assign n18909 = n12523 & n12696;
  assign n19084 = ~n18837 & n18909;
  assign n19085 = n12700 & ~n19084;
  assign n19086 = ~n19083 & n19085;
  assign n19087 = ~n18845 & n19082;
  assign n12697 = ~n12523 & ~n12696;
  assign n19088 = n12697 & n18837;
  assign n19089 = ~n12700 & ~n19088;
  assign n19090 = ~n19087 & n19089;
  assign n19091 = ~n19086 & ~n19090;
  assign n18906 = ~n18837 & n18845;
  assign n19092 = n18906 & n18909;
  assign n18908 = n18837 & ~n18845;
  assign n19093 = n12697 & n18908;
  assign n19094 = ~n19092 & ~n19093;
  assign n19095 = ~n19091 & n19094;
  assign n18884 = ~x22 & ~n11941;
  assign n18885 = x22 & ~n11940;
  assign n18886 = x23 & ~n18885;
  assign n18887 = ~n18884 & n18886;
  assign n18888 = ~n12518 & ~n18887;
  assign n18889 = n4484 & n11902;
  assign n18890 = n4480 & ~n11875;
  assign n18891 = ~n18889 & ~n18890;
  assign n18892 = ~n18888 & n18891;
  assign n18893 = ~n11941 & n14738;
  assign n18894 = ~n11940 & n14740;
  assign n18895 = n18891 & ~n18894;
  assign n18896 = ~n18893 & n18895;
  assign n18897 = ~x23 & ~n18896;
  assign n18898 = ~n18892 & ~n18897;
  assign n18870 = ~n12479 & n12497;
  assign n18871 = ~n12480 & ~n12493;
  assign n18872 = ~n12490 & n18871;
  assign n18873 = n11680 & n12492;
  assign n18874 = n12480 & ~n18873;
  assign n18875 = n11680 ^ n11658;
  assign n18876 = ~n11614 & ~n18875;
  assign n18877 = ~n12481 & n18876;
  assign n18878 = n18874 & ~n18877;
  assign n18879 = ~n18872 & ~n18878;
  assign n18880 = ~n18870 & ~n18879;
  assign n11689 = n11675 ^ n11658;
  assign n11690 = ~n11676 & n11689;
  assign n11691 = n11690 ^ n11658;
  assign n11677 = ~n11658 & ~n11676;
  assign n11678 = n11637 & ~n11677;
  assign n11679 = n11614 & ~n11678;
  assign n11681 = n11658 & n11676;
  assign n11682 = ~n11680 & n11681;
  assign n11683 = n11637 & ~n11682;
  assign n11686 = ~n11684 & n11685;
  assign n11687 = ~n11683 & ~n11686;
  assign n11688 = ~n11679 & ~n11687;
  assign n18867 = n11691 ^ n11688;
  assign n10984 = n10977 & n10983;
  assign n10985 = n679 & n1792;
  assign n10987 = n1116 & n10986;
  assign n10988 = n10985 & n10987;
  assign n10989 = ~n189 & ~n750;
  assign n10990 = ~n396 & n10989;
  assign n10991 = n1650 & n10990;
  assign n10992 = n10988 & n10991;
  assign n10993 = n10984 & n10992;
  assign n10994 = ~n141 & ~n1135;
  assign n10995 = n3938 & n10994;
  assign n10996 = n1273 & n2013;
  assign n10997 = n10995 & n10996;
  assign n10998 = n10993 & n10997;
  assign n10999 = n10976 & n10998;
  assign n11000 = n1372 & n10999;
  assign n11009 = ~n567 & ~n928;
  assign n11010 = n11008 & n11009;
  assign n11011 = n459 & n11010;
  assign n11012 = n813 & n4064;
  assign n11013 = n11011 & n11012;
  assign n11014 = ~n403 & ~n755;
  assign n11015 = ~n346 & n11014;
  assign n11017 = n884 & n11016;
  assign n11018 = n11015 & n11017;
  assign n11019 = n11013 & n11018;
  assign n11020 = n11007 & n11019;
  assign n11021 = n11000 & n11020;
  assign n18868 = n18867 ^ n11021;
  assign n11705 = n44 & n11704;
  assign n11706 = n3280 & n11486;
  assign n11707 = n3277 & n11215;
  assign n11708 = n3275 & ~n10956;
  assign n11709 = ~n11707 & ~n11708;
  assign n11710 = ~n11706 & n11709;
  assign n11711 = ~n11705 & n11710;
  assign n11712 = n11711 ^ x29;
  assign n11695 = n41 & n11694;
  assign n11696 = ~n11633 & ~n11695;
  assign n11697 = x31 & ~n11696;
  assign n11698 = ~n91 & ~n10663;
  assign n11699 = n5358 & ~n11698;
  assign n11700 = ~n5354 & ~n10665;
  assign n11701 = ~n11699 & ~n11700;
  assign n11702 = ~n11697 & n11701;
  assign n11713 = n11712 ^ n11702;
  assign n18869 = n18868 ^ n11713;
  assign n18881 = n18880 ^ n18869;
  assign n18859 = n3285 & ~n11777;
  assign n18860 = n3437 & ~n11773;
  assign n18861 = ~n3440 & n11500;
  assign n18862 = n3435 & n11480;
  assign n18863 = ~n18861 & ~n18862;
  assign n18864 = ~n18860 & n18863;
  assign n18865 = ~n18859 & n18864;
  assign n18866 = n18865 ^ x26;
  assign n18882 = n18881 ^ n18866;
  assign n18856 = n12498 ^ n12451;
  assign n18857 = ~n12499 & n18856;
  assign n18858 = n18857 ^ n12451;
  assign n18883 = n18882 ^ n18858;
  assign n18899 = n18898 ^ n18883;
  assign n18850 = x20 & n12019;
  assign n18851 = n4676 & ~n18850;
  assign n18852 = n4680 & n12019;
  assign n18853 = ~n7366 & ~n18852;
  assign n18854 = ~n18851 & n18853;
  assign n18847 = n12522 ^ n12448;
  assign n18848 = ~n12501 & n18847;
  assign n18849 = n18848 ^ n12522;
  assign n18855 = n18854 ^ n18849;
  assign n18900 = n18899 ^ n18855;
  assign n19096 = n19095 ^ n18900;
  assign n19293 = ~n19288 & ~n19292;
  assign n19294 = n19096 & ~n19293;
  assign n18968 = n4477 & n12013;
  assign n18969 = n4476 & ~n12019;
  assign n18970 = ~n18968 & n18969;
  assign n18971 = n4484 & ~n11940;
  assign n18972 = n4480 & n11902;
  assign n18973 = ~n18971 & ~n18972;
  assign n18974 = ~n18970 & n18973;
  assign n18975 = n18974 ^ x23;
  assign n18950 = ~n12000 & n12417;
  assign n18951 = n3435 & ~n11773;
  assign n18952 = ~n3440 & n11480;
  assign n18953 = ~n18951 & ~n18952;
  assign n18954 = x26 & n18953;
  assign n18955 = n11875 & n18954;
  assign n18956 = x25 & ~n18955;
  assign n18957 = ~n18950 & n18956;
  assign n18958 = n12000 & n18954;
  assign n18959 = ~n11875 & n12417;
  assign n18960 = ~x25 & ~n18959;
  assign n18961 = ~n18958 & n18960;
  assign n18962 = ~n18957 & ~n18961;
  assign n18963 = ~n12432 & n18953;
  assign n18964 = n18963 ^ x26;
  assign n18965 = ~n18962 & n18964;
  assign n18933 = n11702 ^ n11688;
  assign n18934 = ~n18867 & ~n18933;
  assign n18935 = n18934 ^ n11702;
  assign n18936 = n11712 & ~n18935;
  assign n18937 = ~n11021 & ~n18936;
  assign n11692 = n11688 & n11691;
  assign n18938 = n11692 & ~n11702;
  assign n18939 = n18937 & ~n18938;
  assign n18940 = ~n11712 & n18935;
  assign n11725 = ~n11688 & ~n11691;
  assign n18941 = n11702 & n11725;
  assign n18942 = n11021 & ~n18941;
  assign n18943 = ~n18940 & n18942;
  assign n18944 = ~n18939 & ~n18943;
  assign n18945 = ~n18938 & ~n18941;
  assign n18946 = n11713 & ~n18945;
  assign n18947 = ~n18944 & ~n18946;
  assign n11037 = ~n553 & n2755;
  assign n11038 = ~n218 & ~n245;
  assign n11039 = n11037 & n11038;
  assign n11041 = n584 & n11040;
  assign n11042 = n413 & n1153;
  assign n11043 = n11041 & n11042;
  assign n11044 = n11039 & n11043;
  assign n11045 = n2592 & n11044;
  assign n11046 = ~n278 & ~n449;
  assign n11047 = ~n248 & n11046;
  assign n11048 = n2145 & n2160;
  assign n11049 = n11047 & n11048;
  assign n11050 = n2043 & n5557;
  assign n11051 = n11049 & n11050;
  assign n11052 = n11045 & n11051;
  assign n11053 = n1876 & n11052;
  assign n11054 = n11036 & n11053;
  assign n11055 = n4135 & n11054;
  assign n11715 = n11055 ^ n11021;
  assign n10958 = n41 & n10957;
  assign n10959 = n54 & ~n10665;
  assign n10960 = x31 & ~n10959;
  assign n10961 = ~n10958 & n10960;
  assign n10962 = n3671 & ~n10663;
  assign n10963 = ~n10961 & ~n10962;
  assign n10964 = n3676 & ~n10956;
  assign n10965 = n10963 & ~n10964;
  assign n10966 = n91 & n10663;
  assign n10967 = ~n10965 & ~n10966;
  assign n11716 = n11715 ^ n10967;
  assign n18948 = n18947 ^ n11716;
  assign n18925 = n44 & n11957;
  assign n18926 = n3280 & n11500;
  assign n18927 = n3277 & n11486;
  assign n18928 = n3275 & n11215;
  assign n18929 = ~n18927 & ~n18928;
  assign n18930 = ~n18926 & n18929;
  assign n18931 = ~n18925 & n18930;
  assign n18932 = n18931 ^ x29;
  assign n18949 = n18948 ^ n18932;
  assign n18966 = n18965 ^ n18949;
  assign n18922 = n18869 ^ n18866;
  assign n18923 = n18881 & ~n18922;
  assign n18924 = n18923 ^ n18880;
  assign n18967 = n18966 ^ n18924;
  assign n18976 = n18975 ^ n18967;
  assign n11058 = x19 ^ x18;
  assign n11059 = ~n4672 & ~n11058;
  assign n11060 = ~n4671 & n11059;
  assign n11061 = n11060 ^ x20;
  assign n19295 = n18976 ^ n11061;
  assign n18977 = n18898 ^ n18858;
  assign n18978 = ~n18883 & n18977;
  assign n18979 = n18978 ^ n18898;
  assign n19296 = n19295 ^ n18979;
  assign n18916 = n18899 ^ n18849;
  assign n18917 = n18855 & n18916;
  assign n18918 = n18917 ^ n18899;
  assign n19297 = n19296 ^ n18918;
  assign n18838 = n18837 ^ n12700;
  assign n18846 = n18845 ^ n12700;
  assign n18901 = n18900 ^ n18845;
  assign n18902 = ~n18846 & ~n18901;
  assign n18903 = n18838 & n18902;
  assign n18904 = n18903 ^ n18900;
  assign n18905 = ~n12697 & ~n18904;
  assign n18907 = ~n12700 & ~n18906;
  assign n18910 = n18900 & ~n18909;
  assign n18911 = ~n18908 & ~n18910;
  assign n18912 = ~n18907 & n18911;
  assign n18913 = ~n18900 & n18909;
  assign n18914 = ~n18912 & ~n18913;
  assign n18915 = ~n18905 & n18914;
  assign n19298 = n19297 ^ n18915;
  assign n19299 = ~n19294 & ~n19298;
  assign n19589 = n19292 & ~n19588;
  assign n19590 = ~n19096 & ~n19589;
  assign n19591 = n19298 & ~n19590;
  assign n21714 = ~n19299 & ~n19591;
  assign n19064 = n18979 ^ n18976;
  assign n19065 = n18979 ^ n18915;
  assign n19066 = ~n19064 & ~n19065;
  assign n19067 = n19066 ^ n18915;
  assign n19068 = ~n18918 & n19067;
  assign n18980 = ~n18976 & ~n18979;
  assign n19069 = n18915 & n18980;
  assign n19070 = n11061 & ~n19069;
  assign n19071 = n19068 & ~n19070;
  assign n18921 = n11061 & n18918;
  assign n19072 = n18921 & ~n19067;
  assign n19073 = ~n11061 & n19069;
  assign n18919 = ~n11061 & ~n18918;
  assign n18920 = ~n18915 & ~n18919;
  assign n19020 = n18976 & n18979;
  assign n19074 = n18920 & n19020;
  assign n19075 = ~n19073 & ~n19074;
  assign n19076 = ~n19072 & n19075;
  assign n19077 = ~n19071 & n19076;
  assign n18995 = n12417 & n12504;
  assign n18996 = n3435 & ~n11875;
  assign n18997 = ~n3440 & ~n11773;
  assign n18998 = ~n18996 & ~n18997;
  assign n18999 = x26 & n18998;
  assign n19000 = ~n11902 & n18999;
  assign n19001 = ~n18995 & ~n19000;
  assign n19002 = x25 & n19001;
  assign n19003 = ~n12504 & n18999;
  assign n19004 = n11902 & n12417;
  assign n19005 = ~x25 & ~n19004;
  assign n19006 = ~n19003 & n19005;
  assign n19007 = ~n19002 & ~n19006;
  assign n19008 = ~n12432 & n18998;
  assign n19009 = n19008 ^ x26;
  assign n19010 = ~n19007 & n19009;
  assign n11714 = n11702 ^ n11021;
  assign n11717 = n11716 ^ n11021;
  assign n11718 = ~n11714 & ~n11717;
  assign n11719 = n11713 & n11718;
  assign n11720 = n11719 ^ n11716;
  assign n11721 = ~n11692 & ~n11720;
  assign n11722 = n11702 & ~n11712;
  assign n11723 = ~n11021 & ~n11722;
  assign n11724 = ~n11702 & n11712;
  assign n11726 = n11716 & ~n11725;
  assign n11727 = ~n11724 & ~n11726;
  assign n11728 = ~n11723 & n11727;
  assign n11729 = ~n11716 & n11725;
  assign n11730 = ~n11728 & ~n11729;
  assign n11731 = ~n11721 & n11730;
  assign n11508 = n44 & n11507;
  assign n11509 = n3280 & n11480;
  assign n11510 = n3277 & n11500;
  assign n11511 = ~n11509 & ~n11510;
  assign n11512 = n3275 & n11486;
  assign n11513 = n11511 & ~n11512;
  assign n11514 = ~n11508 & n11513;
  assign n11515 = n11514 ^ x29;
  assign n11228 = n10956 & n11227;
  assign n11229 = n3667 & n11228;
  assign n11230 = n3676 & n11215;
  assign n11231 = n3669 & ~n10663;
  assign n11232 = ~n11230 & ~n11231;
  assign n11233 = ~n11229 & n11232;
  assign n11235 = n11227 & n11234;
  assign n11236 = n5636 & ~n10956;
  assign n11237 = ~n11235 & n11236;
  assign n11238 = n11233 & ~n11237;
  assign n11062 = n584 & n1160;
  assign n11063 = n100 & n11062;
  assign n11064 = n191 & n4040;
  assign n11065 = n11063 & n11064;
  assign n11067 = n1333 & n11066;
  assign n11068 = n11065 & n11067;
  assign n11069 = ~n265 & n1611;
  assign n11070 = ~n244 & ~n812;
  assign n11071 = ~n656 & n11070;
  assign n11072 = n11069 & n11071;
  assign n11073 = n251 & n3163;
  assign n11074 = n11072 & n11073;
  assign n11075 = n2446 & n11074;
  assign n11076 = n11068 & n11075;
  assign n11077 = ~n336 & ~n418;
  assign n11078 = ~n612 & n11077;
  assign n11079 = n3538 & n11078;
  assign n11080 = n285 & ~n588;
  assign n11081 = n1037 & n11080;
  assign n11082 = n11079 & n11081;
  assign n11083 = n274 & n498;
  assign n11085 = n925 & n11084;
  assign n11086 = n11083 & n11085;
  assign n11087 = n11082 & n11086;
  assign n11088 = n1291 & n2667;
  assign n11089 = n11087 & n11088;
  assign n11090 = n11076 & n11089;
  assign n11091 = n2103 & n11090;
  assign n11092 = n11091 ^ n11061;
  assign n11239 = n11238 ^ n11092;
  assign n11022 = n11021 ^ n10967;
  assign n11056 = n11055 ^ n10967;
  assign n11057 = n11022 & n11056;
  assign n11240 = n11239 ^ n11057;
  assign n11516 = n11515 ^ n11240;
  assign n18994 = n11731 ^ n11516;
  assign n19011 = n19010 ^ n18994;
  assign n18991 = n18965 ^ n18948;
  assign n18992 = ~n18949 & n18991;
  assign n18993 = n18992 ^ n18965;
  assign n19012 = n19011 ^ n18993;
  assign n18984 = n4478 & n17383;
  assign n18985 = n4480 & ~n11940;
  assign n18986 = n4484 & ~n12019;
  assign n18987 = ~n4487 & ~n18986;
  assign n18988 = ~n18985 & n18987;
  assign n18989 = ~n18984 & n18988;
  assign n18990 = n18989 ^ x23;
  assign n19013 = n19012 ^ n18990;
  assign n18981 = n18975 ^ n18966;
  assign n18982 = ~n18967 & n18981;
  assign n18983 = n18982 ^ n18975;
  assign n19014 = n19013 ^ n18983;
  assign n19078 = n19077 ^ n19014;
  assign n21715 = n21714 ^ n19078;
  assign n21716 = ~x7 & ~n21715;
  assign n21717 = x7 & ~n19078;
  assign n21718 = x8 & ~n21717;
  assign n21719 = ~n21716 & n21718;
  assign n21720 = ~n16819 & ~n21719;
  assign n21721 = n6316 & n19096;
  assign n21722 = n6309 & n19298;
  assign n21723 = ~n21721 & ~n21722;
  assign n21724 = ~n21720 & n21723;
  assign n21725 = x7 & n21715;
  assign n21726 = ~x7 & n19078;
  assign n21727 = n16805 & ~n21726;
  assign n21728 = ~n21725 & n21727;
  assign n21729 = ~x8 & ~n21723;
  assign n21730 = ~n21728 & ~n21729;
  assign n21731 = ~n21724 & n21730;
  assign n21353 = n21352 ^ n21213;
  assign n19667 = ~n19294 & ~n19590;
  assign n19668 = n19667 ^ n19298;
  assign n19669 = n6306 & n19668;
  assign n19670 = n7168 & n19298;
  assign n19671 = n6316 & n19292;
  assign n19672 = ~n19670 & ~n19671;
  assign n19673 = n6309 & n19096;
  assign n19674 = n19672 & ~n19673;
  assign n19675 = ~n19669 & n19674;
  assign n19676 = n19675 ^ x8;
  assign n21354 = n21353 ^ n19676;
  assign n21696 = n21210 ^ n20906;
  assign n21681 = n21207 ^ n21206;
  assign n21363 = n21184 ^ n20918;
  assign n21355 = n6306 & n21215;
  assign n21356 = n7168 & n19104;
  assign n21357 = n6316 & n19122;
  assign n21358 = n6309 & ~n19286;
  assign n21359 = ~n21357 & ~n21358;
  assign n21360 = ~n21356 & n21359;
  assign n21361 = ~n21355 & n21360;
  assign n21362 = n21361 ^ x8;
  assign n21364 = n21363 ^ n21362;
  assign n21373 = n21181 ^ n20928;
  assign n21365 = n6306 & ~n19678;
  assign n21366 = n6309 & n19122;
  assign n21367 = n7168 & ~n19286;
  assign n21368 = n6316 & ~n19281;
  assign n21369 = ~n21367 & ~n21368;
  assign n21370 = ~n21366 & n21369;
  assign n21371 = ~n21365 & n21370;
  assign n21372 = n21371 ^ x8;
  assign n21374 = n21373 ^ n21372;
  assign n21375 = n21175 ^ n20957;
  assign n21384 = n21172 ^ n20967;
  assign n21376 = n6306 & n20793;
  assign n21377 = n7168 & n19277;
  assign n21378 = n6309 & n19260;
  assign n21379 = n6316 & ~n19255;
  assign n21380 = ~n21378 & ~n21379;
  assign n21381 = ~n21377 & n21380;
  assign n21382 = ~n21376 & n21381;
  assign n21383 = n21382 ^ x8;
  assign n21385 = n21384 ^ n21383;
  assign n21394 = n21169 ^ n20977;
  assign n21386 = n6306 & n20929;
  assign n21387 = n7168 & n19260;
  assign n21388 = n6309 & ~n19255;
  assign n21389 = n6316 & n19253;
  assign n21390 = ~n21388 & ~n21389;
  assign n21391 = ~n21387 & n21390;
  assign n21392 = ~n21386 & n21391;
  assign n21393 = n21392 ^ x8;
  assign n21395 = n21394 ^ n21393;
  assign n21412 = n21166 ^ n20987;
  assign n21396 = n16805 & ~n19696;
  assign n21397 = n6309 & n19253;
  assign n21398 = n6316 & ~n19238;
  assign n21399 = ~n21397 & ~n21398;
  assign n21400 = x8 & n21399;
  assign n21401 = n19255 & n21400;
  assign n21402 = x7 & ~n21401;
  assign n21403 = ~n21396 & n21402;
  assign n21404 = n19696 & n21400;
  assign n21405 = n16805 & ~n19255;
  assign n21406 = ~x7 & ~n21405;
  assign n21407 = ~n21404 & n21406;
  assign n21408 = ~n21403 & ~n21407;
  assign n21409 = ~n16820 & n21399;
  assign n21410 = n21409 ^ x8;
  assign n21411 = ~n21408 & n21410;
  assign n21413 = n21412 ^ n21411;
  assign n21422 = n21163 ^ n20997;
  assign n21414 = n6306 & n20308;
  assign n21415 = n7168 & n19253;
  assign n21416 = n6309 & ~n19238;
  assign n21417 = n6316 & n19233;
  assign n21418 = ~n21416 & ~n21417;
  assign n21419 = ~n21415 & n21418;
  assign n21420 = ~n21414 & n21419;
  assign n21421 = n21420 ^ x8;
  assign n21423 = n21422 ^ n21421;
  assign n21432 = n21160 ^ n21007;
  assign n21424 = n6306 & ~n20328;
  assign n21425 = n7168 & ~n19238;
  assign n21426 = n6309 & n19233;
  assign n21427 = n6316 & n19139;
  assign n21428 = ~n21426 & ~n21427;
  assign n21429 = ~n21425 & n21428;
  assign n21430 = ~n21424 & n21429;
  assign n21431 = n21430 ^ x8;
  assign n21433 = n21432 ^ n21431;
  assign n21435 = n6306 & n20294;
  assign n21436 = n7168 & n19233;
  assign n21437 = n6309 & n19139;
  assign n21438 = n6316 & ~n19142;
  assign n21439 = ~n21437 & ~n21438;
  assign n21440 = ~n21436 & n21439;
  assign n21441 = ~n21435 & n21440;
  assign n21442 = n21441 ^ x8;
  assign n21434 = n21157 ^ n21141;
  assign n21443 = n21442 ^ n21434;
  assign n21445 = n6306 & ~n20031;
  assign n21446 = n7168 & n19139;
  assign n21447 = n6309 & ~n19142;
  assign n21448 = n6316 & ~n19225;
  assign n21449 = ~n21447 & ~n21448;
  assign n21450 = ~n21446 & n21449;
  assign n21451 = ~n21445 & n21450;
  assign n21452 = n21451 ^ x8;
  assign n21444 = n21136 ^ n21135;
  assign n21453 = n21452 ^ n21444;
  assign n21455 = n6306 & ~n20045;
  assign n21456 = n7168 & ~n19142;
  assign n21457 = n6316 & ~n19215;
  assign n21458 = ~n21456 & ~n21457;
  assign n21459 = n6309 & ~n19225;
  assign n21460 = n21458 & ~n21459;
  assign n21461 = ~n21455 & n21460;
  assign n21462 = n21461 ^ x8;
  assign n21454 = n21123 ^ n21122;
  assign n21463 = n21462 ^ n21454;
  assign n21609 = n6306 & ~n20210;
  assign n21610 = n7168 & ~n19225;
  assign n21611 = n6316 & n19160;
  assign n21612 = n6309 & ~n19215;
  assign n21613 = ~n21611 & ~n21612;
  assign n21614 = ~n21610 & n21613;
  assign n21615 = ~n21609 & n21614;
  assign n21616 = n21615 ^ x8;
  assign n21596 = n21107 ^ n21027;
  assign n21583 = n21104 ^ n21037;
  assign n21472 = n21101 ^ n21048;
  assign n21464 = n6306 & n19816;
  assign n21465 = n7168 & n19200;
  assign n21466 = n6309 & ~n19162;
  assign n21467 = n6316 & ~n19201;
  assign n21468 = ~n21466 & ~n21467;
  assign n21469 = ~n21465 & n21468;
  assign n21470 = ~n21464 & n21469;
  assign n21471 = n21470 ^ x8;
  assign n21473 = n21472 ^ n21471;
  assign n21482 = n21098 ^ n21090;
  assign n21474 = n6306 & ~n19828;
  assign n21475 = n7168 & ~n19162;
  assign n21476 = n6309 & ~n19201;
  assign n21477 = n6316 & ~n19161;
  assign n21478 = ~n21476 & ~n21477;
  assign n21479 = ~n21475 & n21478;
  assign n21480 = ~n21474 & n21479;
  assign n21481 = n21480 ^ x8;
  assign n21483 = n21482 ^ n21481;
  assign n21485 = n6306 & ~n19840;
  assign n21486 = n7168 & ~n19201;
  assign n21487 = n6309 & ~n19161;
  assign n21488 = n6316 & ~n19167;
  assign n21489 = ~n21487 & ~n21488;
  assign n21490 = ~n21486 & n21489;
  assign n21491 = ~n21485 & n21490;
  assign n21492 = n21491 ^ x8;
  assign n21484 = n21085 ^ n21077;
  assign n21493 = n21492 ^ n21484;
  assign n21560 = n6306 & ~n19799;
  assign n21561 = n7168 & ~n19161;
  assign n21562 = n6309 & ~n19167;
  assign n21563 = n6316 & n19170;
  assign n21564 = ~n21562 & ~n21563;
  assign n21565 = ~n21561 & n21564;
  assign n21566 = ~n21560 & n21565;
  assign n21567 = n21566 ^ x8;
  assign n21537 = n5817 & ~n19175;
  assign n21538 = n21062 & ~n21537;
  assign n21539 = ~x11 & ~n21538;
  assign n21540 = ~n21062 & ~n21064;
  assign n21541 = n5817 & n19729;
  assign n21542 = ~n21540 & ~n21541;
  assign n21543 = ~n21539 & n21542;
  assign n21544 = ~n5812 & ~n19175;
  assign n21545 = n21064 & ~n21544;
  assign n21546 = n21063 & n21545;
  assign n21547 = n21543 & ~n21546;
  assign n21503 = n6306 & n19720;
  assign n21504 = n7168 & n19173;
  assign n21505 = n6309 & n19174;
  assign n21506 = n6316 & ~n19175;
  assign n21507 = ~n21505 & ~n21506;
  assign n21508 = ~n21504 & n21507;
  assign n21509 = ~n21503 & n21508;
  assign n21510 = n21509 ^ x8;
  assign n21498 = n5812 & n19188;
  assign n21511 = n6306 & n19730;
  assign n21512 = n7168 & n19174;
  assign n21513 = n6309 & ~n19175;
  assign n21514 = n6316 & n19188;
  assign n21515 = ~n21513 & ~n21514;
  assign n21516 = ~n21512 & n21515;
  assign n21517 = ~n21511 & n21516;
  assign n21518 = n6305 & ~n19175;
  assign n21519 = ~n19188 & ~n21518;
  assign n21520 = n6315 & ~n21519;
  assign n21521 = x8 & ~n21520;
  assign n21522 = n21517 & n21521;
  assign n21523 = ~n21498 & ~n21522;
  assign n21524 = ~n21510 & ~n21523;
  assign n21494 = ~n5819 & ~n19175;
  assign n21495 = n8711 & ~n21494;
  assign n21496 = ~n8713 & ~n21495;
  assign n21497 = n19188 & ~n21496;
  assign n21499 = x10 & n21498;
  assign n21500 = n21499 ^ n5812;
  assign n21501 = ~n19175 & n21500;
  assign n21502 = ~n21497 & ~n21501;
  assign n21525 = n21524 ^ n21502;
  assign n21526 = n6306 & n19748;
  assign n21527 = n7168 & n19170;
  assign n21528 = n6309 & n19173;
  assign n21529 = n6316 & n19174;
  assign n21530 = ~n21528 & ~n21529;
  assign n21531 = ~n21527 & n21530;
  assign n21532 = ~n21526 & n21531;
  assign n21533 = n21532 ^ x8;
  assign n21534 = n21533 ^ n21524;
  assign n21535 = n21525 & ~n21534;
  assign n21536 = n21535 ^ n21533;
  assign n21548 = n21547 ^ n21536;
  assign n21549 = n6306 & ~n19761;
  assign n21550 = n7168 & ~n19167;
  assign n21551 = n6309 & n19170;
  assign n21552 = n6316 & n19173;
  assign n21553 = ~n21551 & ~n21552;
  assign n21554 = ~n21550 & n21553;
  assign n21555 = ~n21549 & n21554;
  assign n21556 = n21555 ^ x8;
  assign n21557 = n21556 ^ n21547;
  assign n21558 = n21548 & ~n21557;
  assign n21559 = n21558 ^ n21536;
  assign n21568 = n21567 ^ n21559;
  assign n21569 = n21075 ^ n21066;
  assign n21570 = n21569 ^ n21065;
  assign n21571 = n21570 ^ n21567;
  assign n21572 = n21568 & ~n21571;
  assign n21573 = n21572 ^ n21559;
  assign n21574 = n21573 ^ n21484;
  assign n21575 = ~n21493 & n21574;
  assign n21576 = n21575 ^ n21492;
  assign n21577 = n21576 ^ n21482;
  assign n21578 = ~n21483 & n21577;
  assign n21579 = n21578 ^ n21576;
  assign n21580 = n21579 ^ n21472;
  assign n21581 = ~n21473 & n21580;
  assign n21582 = n21581 ^ n21579;
  assign n21584 = n21583 ^ n21582;
  assign n21585 = n6306 & n19966;
  assign n21586 = n7168 & n19160;
  assign n21587 = n6309 & n19200;
  assign n21588 = n6316 & ~n19162;
  assign n21589 = ~n21587 & ~n21588;
  assign n21590 = ~n21586 & n21589;
  assign n21591 = ~n21585 & n21590;
  assign n21592 = n21591 ^ x8;
  assign n21593 = n21592 ^ n21583;
  assign n21594 = ~n21584 & n21593;
  assign n21595 = n21594 ^ n21582;
  assign n21597 = n21596 ^ n21595;
  assign n21598 = n6306 & n20020;
  assign n21599 = n6309 & n19160;
  assign n21600 = n7168 & ~n19215;
  assign n21601 = n6316 & n19200;
  assign n21602 = ~n21600 & ~n21601;
  assign n21603 = ~n21599 & n21602;
  assign n21604 = ~n21598 & n21603;
  assign n21605 = n21604 ^ x8;
  assign n21606 = n21605 ^ n21595;
  assign n21607 = ~n21597 & n21606;
  assign n21608 = n21607 ^ n21605;
  assign n21617 = n21616 ^ n21608;
  assign n21618 = n21110 ^ n21017;
  assign n21619 = n21618 ^ n21608;
  assign n21620 = n21617 & ~n21619;
  assign n21621 = n21620 ^ n21616;
  assign n21622 = n21621 ^ n21462;
  assign n21623 = ~n21463 & n21622;
  assign n21624 = n21623 ^ n21621;
  assign n21625 = n21624 ^ n21452;
  assign n21626 = ~n21453 & n21625;
  assign n21627 = n21626 ^ n21624;
  assign n21628 = n21627 ^ n21442;
  assign n21629 = ~n21443 & n21628;
  assign n21630 = n21629 ^ n21627;
  assign n21631 = n21630 ^ n21432;
  assign n21632 = n21433 & ~n21631;
  assign n21633 = n21632 ^ n21630;
  assign n21634 = n21633 ^ n21422;
  assign n21635 = ~n21423 & n21634;
  assign n21636 = n21635 ^ n21633;
  assign n21637 = n21636 ^ n21412;
  assign n21638 = ~n21413 & n21637;
  assign n21639 = n21638 ^ n21636;
  assign n21640 = n21639 ^ n21394;
  assign n21641 = ~n21395 & n21640;
  assign n21642 = n21641 ^ n21639;
  assign n21643 = n21642 ^ n21384;
  assign n21644 = ~n21385 & n21643;
  assign n21645 = n21644 ^ n21642;
  assign n21646 = ~n21375 & ~n21645;
  assign n21647 = n21178 ^ n20947;
  assign n21648 = ~n21646 & ~n21647;
  assign n21649 = n6306 & n21189;
  assign n21650 = n7168 & n19122;
  assign n21651 = n6309 & ~n19281;
  assign n21652 = n6316 & n19277;
  assign n21653 = ~n21651 & ~n21652;
  assign n21654 = ~n21650 & n21653;
  assign n21655 = ~n21649 & n21654;
  assign n21656 = n21655 ^ x8;
  assign n21657 = ~n21648 & ~n21656;
  assign n21658 = n21375 & n21645;
  assign n21659 = n6306 & ~n20908;
  assign n21660 = n7168 & ~n19281;
  assign n21661 = n6309 & n19277;
  assign n21662 = n6316 & n19260;
  assign n21663 = ~n21661 & ~n21662;
  assign n21664 = ~n21660 & n21663;
  assign n21665 = ~n21659 & n21664;
  assign n21666 = n21665 ^ x8;
  assign n21667 = n21665 ^ n21655;
  assign n21668 = ~n21647 & n21667;
  assign n21669 = ~n21666 & n21668;
  assign n21670 = n21669 ^ n21666;
  assign n21671 = ~n21658 & ~n21670;
  assign n21672 = n21646 & n21647;
  assign n21673 = ~n21671 & ~n21672;
  assign n21674 = ~n21657 & n21673;
  assign n21675 = n21674 ^ n21373;
  assign n21676 = ~n21374 & n21675;
  assign n21677 = n21676 ^ n21674;
  assign n21678 = n21677 ^ n21363;
  assign n21679 = ~n21364 & n21678;
  assign n21680 = n21679 ^ n21677;
  assign n21682 = n21681 ^ n21680;
  assign n21685 = n6306 & n21684;
  assign n21686 = n7168 & n19292;
  assign n21687 = n6309 & n19104;
  assign n21688 = n6316 & ~n19286;
  assign n21689 = ~n21687 & ~n21688;
  assign n21690 = ~n21686 & n21689;
  assign n21691 = ~n21685 & n21690;
  assign n21692 = n21691 ^ x8;
  assign n21693 = n21692 ^ n21681;
  assign n21694 = ~n21682 & n21693;
  assign n21695 = n21694 ^ n21680;
  assign n21697 = n21696 ^ n21695;
  assign n21698 = ~n19293 & ~n19589;
  assign n21699 = n21698 ^ n19096;
  assign n21700 = n6306 & n21699;
  assign n21701 = n7168 & n19096;
  assign n21702 = n6309 & n19292;
  assign n21703 = n6316 & n19104;
  assign n21704 = ~n21702 & ~n21703;
  assign n21705 = ~n21701 & n21704;
  assign n21706 = ~n21700 & n21705;
  assign n21707 = n21706 ^ x8;
  assign n21708 = n21707 ^ n21696;
  assign n21709 = ~n21697 & n21708;
  assign n21710 = n21709 ^ n21695;
  assign n21711 = n21710 ^ n21353;
  assign n21712 = n21354 & ~n21711;
  assign n21713 = n21712 ^ n21710;
  assign n21732 = n21731 ^ n21713;
  assign n22046 = n21876 ^ n21732;
  assign n19015 = ~n18980 & n19014;
  assign n19016 = ~n18921 & ~n19015;
  assign n19017 = ~n18920 & n19016;
  assign n19018 = ~n18921 & ~n19014;
  assign n19019 = ~n18915 & ~n19018;
  assign n19021 = ~n18919 & n19014;
  assign n19022 = ~n19020 & ~n19021;
  assign n19023 = ~n19019 & n19022;
  assign n19024 = ~n19017 & ~n19023;
  assign n19025 = n18980 & ~n19014;
  assign n19026 = n19024 & ~n19025;
  assign n19027 = n19012 ^ n18983;
  assign n19028 = ~n19013 & n19027;
  assign n19029 = n19028 ^ n18983;
  assign n19030 = ~n19026 & ~n19029;
  assign n11942 = n3285 & ~n11941;
  assign n11943 = n3437 & ~n11940;
  assign n11944 = n3435 & n11902;
  assign n11945 = ~n3440 & ~n11875;
  assign n11946 = ~n11944 & ~n11945;
  assign n11947 = ~n11943 & n11946;
  assign n11948 = ~n11942 & n11947;
  assign n11949 = n11948 ^ x26;
  assign n11820 = ~n10967 & n11055;
  assign n11821 = ~n11092 & ~n11238;
  assign n11822 = n11820 & ~n11821;
  assign n11823 = n11092 & n11238;
  assign n11824 = n11021 & ~n11823;
  assign n11825 = ~n11822 & n11824;
  assign n11826 = n10967 & ~n11055;
  assign n11827 = n11826 ^ n11238;
  assign n11828 = ~n11021 & n11092;
  assign n11829 = n11828 ^ n11238;
  assign n11830 = ~n11827 & n11829;
  assign n11831 = n11830 ^ n11826;
  assign n11832 = ~n11825 & ~n11831;
  assign n11803 = n2085 & n2143;
  assign n11804 = n3128 & n11803;
  assign n11805 = n1261 & n11804;
  assign n11806 = n11802 & n11805;
  assign n11807 = ~n136 & ~n424;
  assign n11808 = ~n83 & ~n640;
  assign n11809 = n11807 & n11808;
  assign n11810 = n11024 & n11809;
  assign n11811 = ~n524 & ~n549;
  assign n11812 = n883 & n11811;
  assign n11813 = n4783 & n11812;
  assign n11814 = n11810 & n11813;
  assign n11815 = n11806 & n11814;
  assign n11816 = n11138 & n11815;
  assign n11817 = n2283 & n11816;
  assign n11797 = n11061 ^ n11021;
  assign n11798 = n11092 & ~n11797;
  assign n11799 = n11798 ^ n11021;
  assign n11818 = n11817 ^ n11799;
  assign n11789 = n41 & ~n11704;
  assign n11790 = n91 & ~n11215;
  assign n11791 = n54 & n10956;
  assign n11792 = ~n11790 & ~n11791;
  assign n11793 = ~n11789 & n11792;
  assign n11786 = n41 & n11486;
  assign n11787 = n54 & n11215;
  assign n11788 = ~n11786 & ~n11787;
  assign n11794 = n11793 ^ n11788;
  assign n11795 = ~x31 & ~n11794;
  assign n11796 = n11795 ^ n11793;
  assign n11819 = n11818 ^ n11796;
  assign n11833 = n11832 ^ n11819;
  assign n11778 = n44 & ~n11777;
  assign n11779 = n3280 & ~n11773;
  assign n11780 = n3275 & n11500;
  assign n11781 = n3277 & n11480;
  assign n11782 = ~n11780 & ~n11781;
  assign n11783 = ~n11779 & n11782;
  assign n11784 = ~n11778 & n11783;
  assign n11785 = n11784 ^ x29;
  assign n11834 = n11833 ^ n11785;
  assign n11732 = n11731 ^ n11515;
  assign n11733 = ~n11516 & n11732;
  assign n11734 = n11733 ^ n11731;
  assign n11835 = n11834 ^ n11734;
  assign n19031 = n11949 ^ n11835;
  assign n19032 = x22 & ~x23;
  assign n19033 = n18850 & n19032;
  assign n19034 = ~x20 & x23;
  assign n19035 = ~n19033 & ~n19034;
  assign n19036 = x21 & ~n19035;
  assign n19037 = x23 & n12019;
  assign n19038 = n35 & ~n19037;
  assign n19039 = ~x20 & ~x22;
  assign n19040 = x23 & ~n19039;
  assign n19041 = ~n37 & n19040;
  assign n19042 = ~n19038 & ~n19041;
  assign n19043 = ~n19036 & n19042;
  assign n19044 = n19031 & ~n19043;
  assign n19045 = n18994 ^ n18993;
  assign n19046 = n19011 & ~n19045;
  assign n19047 = n19046 ^ n19010;
  assign n19048 = n19044 & n19047;
  assign n19049 = ~n19030 & n19048;
  assign n19050 = n19026 & n19029;
  assign n19051 = n19043 ^ n19031;
  assign n19052 = n19047 ^ n19031;
  assign n19053 = n19051 & n19052;
  assign n19054 = n19053 ^ n19047;
  assign n19055 = n19050 & n19054;
  assign n19056 = ~n19049 & ~n19055;
  assign n19057 = ~n19031 & n19043;
  assign n19058 = ~n19047 & n19057;
  assign n19059 = ~n19050 & n19058;
  assign n19060 = n19030 & ~n19054;
  assign n19061 = ~n19059 & ~n19060;
  assign n19062 = n19056 & n19061;
  assign n12014 = n643 & n12013;
  assign n12020 = n735 & ~n12019;
  assign n12021 = ~n12014 & n12020;
  assign n12022 = n3435 & ~n11940;
  assign n12023 = ~n3440 & n11902;
  assign n12024 = ~n12022 & ~n12023;
  assign n12025 = ~n12021 & n12024;
  assign n12026 = n12025 ^ x26;
  assign n12001 = n44 & ~n12000;
  assign n12002 = n3280 & ~n11875;
  assign n12003 = n3277 & ~n11773;
  assign n12004 = n3275 & n11480;
  assign n12005 = ~n12003 & ~n12004;
  assign n12006 = ~n12002 & n12005;
  assign n12007 = ~n12001 & n12006;
  assign n12008 = n12007 ^ x29;
  assign n11992 = n11799 & n11817;
  assign n11993 = ~n11796 & n11992;
  assign n11994 = ~n11799 & ~n11817;
  assign n11995 = n11796 & n11994;
  assign n11996 = ~n11993 & ~n11995;
  assign n11979 = n713 & n11304;
  assign n11980 = n875 & n11979;
  assign n11981 = n1422 & n5403;
  assign n11982 = ~n343 & n3074;
  assign n11983 = n11981 & n11982;
  assign n11984 = n11980 & n11983;
  assign n11985 = n4622 & n11984;
  assign n11986 = n11978 & n11985;
  assign n11987 = n11020 & n11986;
  assign n11988 = n1996 & n3291;
  assign n11989 = n3123 & n11988;
  assign n11990 = n11987 & n11989;
  assign n11991 = n4379 & n11990;
  assign n11997 = n11996 ^ n11991;
  assign n11958 = n41 & n11957;
  assign n11959 = n91 & n11486;
  assign n11960 = x31 & ~n11787;
  assign n11961 = ~n11959 & n11960;
  assign n11962 = ~n11958 & n11961;
  assign n11963 = n41 & n11500;
  assign n11964 = n54 & n11486;
  assign n11965 = ~x31 & ~n11964;
  assign n11966 = ~n11963 & n11965;
  assign n11967 = ~n11962 & ~n11966;
  assign n11998 = n11997 ^ n11967;
  assign n12009 = n12008 ^ n11998;
  assign n11953 = n11819 ^ n11785;
  assign n11954 = n11833 & ~n11953;
  assign n11955 = n11954 ^ n11832;
  assign n12010 = n12009 ^ n11955;
  assign n12027 = n12026 ^ n12010;
  assign n11950 = n11949 ^ n11734;
  assign n11951 = ~n11835 & n11950;
  assign n11952 = n11951 ^ n11949;
  assign n12028 = n12027 ^ n11952;
  assign n39 = ~x23 & n38;
  assign n40 = n39 ^ n37;
  assign n12029 = n12028 ^ n40;
  assign n19063 = n19062 ^ n12029;
  assign n19300 = ~n19078 & ~n19299;
  assign n19301 = n19051 ^ n19047;
  assign n19302 = n19301 ^ n19029;
  assign n19303 = n19302 ^ n19026;
  assign n19304 = ~n19300 & ~n19303;
  assign n19305 = n19063 & ~n19304;
  assign n19592 = n19078 & ~n19591;
  assign n19593 = n19303 & ~n19592;
  assign n19594 = ~n19063 & ~n19593;
  assign n22036 = ~n19305 & ~n19594;
  assign n19365 = ~n12029 & ~n19060;
  assign n19366 = ~n19059 & n19365;
  assign n19367 = n19056 & ~n19366;
  assign n19355 = n3285 & n17383;
  assign n19356 = ~n3440 & ~n11940;
  assign n19357 = n3435 & ~n12019;
  assign n19358 = ~n3437 & ~n19357;
  assign n19359 = ~n19356 & n19358;
  assign n19360 = ~n19355 & n19359;
  assign n19361 = n19360 ^ x26;
  assign n19345 = n44 & n12504;
  assign n19346 = n3280 & n11902;
  assign n19347 = n3277 & ~n11875;
  assign n19348 = n3275 & ~n11773;
  assign n19349 = ~n19347 & ~n19348;
  assign n19350 = ~n19346 & n19349;
  assign n19351 = ~n19345 & n19350;
  assign n19352 = n19351 ^ x29;
  assign n19333 = n41 & n11507;
  assign n19334 = x31 & ~n11964;
  assign n19335 = ~n19333 & n19334;
  assign n19336 = n54 & n11500;
  assign n19337 = ~x31 & ~n19336;
  assign n19338 = n41 & n11480;
  assign n19339 = n19337 & ~n19338;
  assign n19340 = ~n19335 & ~n19339;
  assign n19341 = n3672 & n11500;
  assign n19342 = ~n19340 & ~n19341;
  assign n19318 = n4781 & n12275;
  assign n19319 = n13492 & n19318;
  assign n19320 = n3218 & n3697;
  assign n19321 = ~n185 & ~n238;
  assign n19322 = ~n280 & n19321;
  assign n19323 = n2392 & n3936;
  assign n19324 = n19322 & n19323;
  assign n19325 = n1091 & n19324;
  assign n19326 = n19320 & n19325;
  assign n19327 = n4098 & n12057;
  assign n19328 = n641 & n19327;
  assign n19329 = n19326 & n19328;
  assign n19330 = n11533 & n19329;
  assign n19331 = n19319 & n19330;
  assign n19332 = n19331 ^ n40;
  assign n19343 = n19342 ^ n19332;
  assign n19315 = n11995 ^ n11993;
  assign n19316 = ~n11991 & n19315;
  assign n19317 = n19316 ^ n11993;
  assign n19344 = n19343 ^ n19317;
  assign n19353 = n19352 ^ n19344;
  assign n19312 = n12008 ^ n11997;
  assign n19313 = ~n11998 & ~n19312;
  assign n19314 = n19313 ^ n12008;
  assign n19354 = n19353 ^ n19314;
  assign n19362 = n19361 ^ n19354;
  assign n19309 = n12026 ^ n12009;
  assign n19310 = ~n12010 & n19309;
  assign n19311 = n19310 ^ n12026;
  assign n19363 = n19362 ^ n19311;
  assign n19306 = n11952 ^ n40;
  assign n19307 = n12028 & n19306;
  assign n19308 = n19307 ^ n12027;
  assign n19364 = n19363 ^ n19308;
  assign n19368 = n19367 ^ n19364;
  assign n22037 = n22036 ^ n19368;
  assign n22038 = n7515 & ~n22037;
  assign n22039 = n8029 & ~n19368;
  assign n22040 = n7518 & n19063;
  assign n22041 = n7520 & n19303;
  assign n22042 = ~n22040 & ~n22041;
  assign n22043 = ~n22039 & n22042;
  assign n22044 = ~n22038 & n22043;
  assign n22045 = n22044 ^ x5;
  assign n22047 = n22046 ^ n22045;
  assign n22048 = n21710 ^ n21354;
  assign n19657 = ~n19300 & ~n19592;
  assign n19658 = n19657 ^ n19303;
  assign n22426 = n7515 & n19658;
  assign n22427 = n7518 & ~n19078;
  assign n22428 = n8029 & n19303;
  assign n22429 = n7520 & n19298;
  assign n22430 = ~n22428 & ~n22429;
  assign n22431 = ~n22427 & n22430;
  assign n22432 = ~n22426 & n22431;
  assign n22433 = n22432 ^ x5;
  assign n22065 = n21692 ^ n21682;
  assign n22049 = n7520 & n19096;
  assign n22050 = n7518 & n19298;
  assign n22051 = ~n22049 & ~n22050;
  assign n22052 = x5 & n22051;
  assign n22053 = n21715 & n22052;
  assign n22054 = n17396 & ~n19078;
  assign n22055 = ~n22053 & ~n22054;
  assign n22056 = ~x4 & ~n22055;
  assign n22057 = ~n17411 & n22051;
  assign n22058 = n22057 ^ x5;
  assign n22059 = ~n22056 & n22058;
  assign n22060 = n17396 & ~n21715;
  assign n22061 = n19078 & n22052;
  assign n22062 = ~n22060 & ~n22061;
  assign n22063 = x4 & ~n22062;
  assign n22064 = n22059 & ~n22063;
  assign n22066 = n22065 ^ n22064;
  assign n22075 = n21677 ^ n21364;
  assign n22067 = n7515 & n19668;
  assign n22068 = n7518 & n19096;
  assign n22069 = n7520 & n19292;
  assign n22070 = ~n22068 & ~n22069;
  assign n22071 = n8029 & n19298;
  assign n22072 = n22070 & ~n22071;
  assign n22073 = ~n22067 & n22072;
  assign n22074 = n22073 ^ x5;
  assign n22076 = n22075 ^ n22074;
  assign n22085 = n21674 ^ n21374;
  assign n22077 = n7515 & n21699;
  assign n22078 = n8029 & n19096;
  assign n22079 = n7518 & n19292;
  assign n22080 = n7520 & n19104;
  assign n22081 = ~n22079 & ~n22080;
  assign n22082 = ~n22078 & n22081;
  assign n22083 = ~n22077 & n22082;
  assign n22084 = n22083 ^ x5;
  assign n22086 = n22085 ^ n22084;
  assign n22094 = n7515 & n21684;
  assign n22095 = n8029 & n19292;
  assign n22096 = n7518 & n19104;
  assign n22097 = n7520 & ~n19286;
  assign n22098 = ~n22096 & ~n22097;
  assign n22099 = ~n22095 & n22098;
  assign n22100 = ~n22094 & n22099;
  assign n22101 = n22100 ^ x5;
  assign n22092 = n21655 ^ n21647;
  assign n22087 = n21645 ^ n21375;
  assign n22088 = n21375 ^ x8;
  assign n22089 = n22088 ^ n21665;
  assign n22090 = ~n22087 & n22089;
  assign n22091 = n22090 ^ n21665;
  assign n22093 = n22092 ^ n22091;
  assign n22102 = n22101 ^ n22093;
  assign n22104 = n7515 & n21215;
  assign n22105 = n8029 & n19104;
  assign n22106 = n7520 & n19122;
  assign n22107 = n7518 & ~n19286;
  assign n22108 = ~n22106 & ~n22107;
  assign n22109 = ~n22105 & n22108;
  assign n22110 = ~n22104 & n22109;
  assign n22111 = n22110 ^ x5;
  assign n22103 = n22087 ^ n21666;
  assign n22112 = n22111 ^ n22103;
  assign n22121 = n21642 ^ n21385;
  assign n22113 = n7515 & ~n19678;
  assign n22114 = n7518 & n19122;
  assign n22115 = n8029 & ~n19286;
  assign n22116 = n7520 & ~n19281;
  assign n22117 = ~n22115 & ~n22116;
  assign n22118 = ~n22114 & n22117;
  assign n22119 = ~n22113 & n22118;
  assign n22120 = n22119 ^ x5;
  assign n22122 = n22121 ^ n22120;
  assign n22131 = n21639 ^ n21395;
  assign n22123 = n7515 & n21189;
  assign n22124 = n8029 & n19122;
  assign n22125 = n7518 & ~n19281;
  assign n22126 = n7520 & n19277;
  assign n22127 = ~n22125 & ~n22126;
  assign n22128 = ~n22124 & n22127;
  assign n22129 = ~n22123 & n22128;
  assign n22130 = n22129 ^ x5;
  assign n22132 = n22131 ^ n22130;
  assign n22141 = n21636 ^ n21413;
  assign n22133 = n7515 & ~n20908;
  assign n22134 = n8029 & ~n19281;
  assign n22135 = n7518 & n19277;
  assign n22136 = n7520 & n19260;
  assign n22137 = ~n22135 & ~n22136;
  assign n22138 = ~n22134 & n22137;
  assign n22139 = ~n22133 & n22138;
  assign n22140 = n22139 ^ x5;
  assign n22142 = n22141 ^ n22140;
  assign n22151 = n21633 ^ n21423;
  assign n22143 = n7515 & n20793;
  assign n22144 = n8029 & n19277;
  assign n22145 = n7518 & n19260;
  assign n22146 = n7520 & ~n19255;
  assign n22147 = ~n22145 & ~n22146;
  assign n22148 = ~n22144 & n22147;
  assign n22149 = ~n22143 & n22148;
  assign n22150 = n22149 ^ x5;
  assign n22152 = n22151 ^ n22150;
  assign n22161 = n21630 ^ n21433;
  assign n22153 = n7515 & n20929;
  assign n22154 = n8029 & n19260;
  assign n22155 = n7518 & ~n19255;
  assign n22156 = n7520 & n19253;
  assign n22157 = ~n22155 & ~n22156;
  assign n22158 = ~n22154 & n22157;
  assign n22159 = ~n22153 & n22158;
  assign n22160 = n22159 ^ x5;
  assign n22162 = n22161 ^ n22160;
  assign n22164 = n7515 & ~n19696;
  assign n22165 = n8029 & ~n19255;
  assign n22166 = n7518 & n19253;
  assign n22167 = n7520 & ~n19238;
  assign n22168 = ~n22166 & ~n22167;
  assign n22169 = ~n22165 & n22168;
  assign n22170 = ~n22164 & n22169;
  assign n22171 = n22170 ^ x5;
  assign n22163 = n21627 ^ n21443;
  assign n22172 = n22171 ^ n22163;
  assign n22174 = n7515 & n20308;
  assign n22175 = n8029 & n19253;
  assign n22176 = n7518 & ~n19238;
  assign n22177 = n7520 & n19233;
  assign n22178 = ~n22176 & ~n22177;
  assign n22179 = ~n22175 & n22178;
  assign n22180 = ~n22174 & n22179;
  assign n22181 = n22180 ^ x5;
  assign n22173 = n21624 ^ n21453;
  assign n22182 = n22181 ^ n22173;
  assign n22184 = n7515 & ~n20328;
  assign n22185 = n8029 & ~n19238;
  assign n22186 = n7518 & n19233;
  assign n22187 = n7520 & n19139;
  assign n22188 = ~n22186 & ~n22187;
  assign n22189 = ~n22185 & n22188;
  assign n22190 = ~n22184 & n22189;
  assign n22191 = n22190 ^ x5;
  assign n22183 = n21621 ^ n21463;
  assign n22192 = n22191 ^ n22183;
  assign n22201 = n21618 ^ n21617;
  assign n22193 = n7513 & n20293;
  assign n22194 = n22193 ^ n19233;
  assign n22195 = n7514 & n22194;
  assign n22196 = n7518 & n19139;
  assign n22197 = n7520 & ~n19142;
  assign n22198 = ~n22196 & ~n22197;
  assign n22199 = ~n22195 & n22198;
  assign n22200 = n22199 ^ x5;
  assign n22202 = n22201 ^ n22200;
  assign n22204 = n7513 & ~n20030;
  assign n22205 = n22204 ^ n19139;
  assign n22206 = n7514 & n22205;
  assign n22207 = n7520 & ~n19225;
  assign n22208 = n7518 & ~n19142;
  assign n22209 = ~n22207 & ~n22208;
  assign n22210 = ~n22206 & n22209;
  assign n22211 = n22210 ^ x5;
  assign n22203 = n21605 ^ n21597;
  assign n22212 = n22211 ^ n22203;
  assign n22214 = n7515 & ~n20045;
  assign n22215 = n8029 & ~n19142;
  assign n22216 = n7518 & ~n19225;
  assign n22217 = ~n22215 & ~n22216;
  assign n22218 = n7520 & ~n19215;
  assign n22219 = n22217 & ~n22218;
  assign n22220 = ~n22214 & n22219;
  assign n22221 = n22220 ^ x5;
  assign n22213 = n21592 ^ n21584;
  assign n22222 = n22221 ^ n22213;
  assign n22224 = n7515 & ~n20210;
  assign n22225 = n8029 & ~n19225;
  assign n22226 = n7520 & n19160;
  assign n22227 = n7518 & ~n19215;
  assign n22228 = ~n22226 & ~n22227;
  assign n22229 = ~n22225 & n22228;
  assign n22230 = ~n22224 & n22229;
  assign n22231 = n22230 ^ x5;
  assign n22223 = n21579 ^ n21473;
  assign n22232 = n22231 ^ n22223;
  assign n22362 = n7515 & n20020;
  assign n22363 = n7518 & n19160;
  assign n22364 = n8029 & ~n19215;
  assign n22365 = n7520 & n19200;
  assign n22366 = ~n22364 & ~n22365;
  assign n22367 = ~n22363 & n22366;
  assign n22368 = ~n22362 & n22367;
  assign n22369 = n22368 ^ x5;
  assign n22241 = n21573 ^ n21493;
  assign n22233 = n7515 & n19966;
  assign n22234 = n8029 & n19160;
  assign n22235 = n7518 & n19200;
  assign n22236 = n7520 & ~n19162;
  assign n22237 = ~n22235 & ~n22236;
  assign n22238 = ~n22234 & n22237;
  assign n22239 = ~n22233 & n22238;
  assign n22240 = n22239 ^ x5;
  assign n22242 = n22241 ^ n22240;
  assign n22251 = n21570 ^ n21568;
  assign n22243 = n7515 & n19816;
  assign n22244 = n8029 & n19200;
  assign n22245 = n7518 & ~n19162;
  assign n22246 = n7520 & ~n19201;
  assign n22247 = ~n22245 & ~n22246;
  assign n22248 = ~n22244 & n22247;
  assign n22249 = ~n22243 & n22248;
  assign n22250 = n22249 ^ x5;
  assign n22252 = n22251 ^ n22250;
  assign n22254 = n7515 & ~n19828;
  assign n22255 = n8029 & ~n19162;
  assign n22256 = n7518 & ~n19201;
  assign n22257 = n7520 & ~n19161;
  assign n22258 = ~n22256 & ~n22257;
  assign n22259 = ~n22255 & n22258;
  assign n22260 = ~n22254 & n22259;
  assign n22261 = n22260 ^ x5;
  assign n22253 = n21556 ^ n21548;
  assign n22262 = n22261 ^ n22253;
  assign n22264 = n7515 & ~n19840;
  assign n22265 = n8029 & ~n19201;
  assign n22266 = n7518 & ~n19161;
  assign n22267 = n7520 & ~n19167;
  assign n22268 = ~n22266 & ~n22267;
  assign n22269 = ~n22265 & n22268;
  assign n22270 = ~n22264 & n22269;
  assign n22271 = n22270 ^ x5;
  assign n22263 = n21533 ^ n21525;
  assign n22272 = n22271 ^ n22263;
  assign n22275 = n7515 & ~n19799;
  assign n22276 = n8029 & ~n19161;
  assign n22277 = n7518 & ~n19167;
  assign n22278 = n7520 & n19170;
  assign n22279 = ~n22277 & ~n22278;
  assign n22280 = ~n22276 & n22279;
  assign n22281 = ~n22275 & n22280;
  assign n22282 = n22281 ^ x5;
  assign n22273 = n21522 ^ n21498;
  assign n22274 = n22273 ^ n21510;
  assign n22283 = n22282 ^ n22274;
  assign n22284 = n7515 & n19720;
  assign n22285 = n8029 & n19173;
  assign n22286 = n7518 & n19174;
  assign n22287 = n7520 & ~n19175;
  assign n22288 = ~n22286 & ~n22287;
  assign n22289 = ~n22285 & n22288;
  assign n22290 = ~n22284 & n22289;
  assign n22291 = n22290 ^ x5;
  assign n22292 = n7514 & ~n19175;
  assign n22293 = ~n19174 & n22292;
  assign n22294 = ~n19188 & ~n22293;
  assign n22295 = ~n7519 & n19188;
  assign n22296 = n7513 & ~n22295;
  assign n22297 = ~n22294 & n22296;
  assign n22298 = n7514 & ~n19729;
  assign n22299 = ~n8029 & ~n22298;
  assign n22300 = n19174 & ~n22299;
  assign n22301 = n7518 & ~n19175;
  assign n22302 = ~n22300 & ~n22301;
  assign n22303 = ~n22297 & n22302;
  assign n22304 = ~n22292 & ~n22295;
  assign n22305 = x5 & n22304;
  assign n22306 = n22303 & n22305;
  assign n22307 = n6305 & n19188;
  assign n22308 = ~n22306 & ~n22307;
  assign n22309 = ~n22291 & ~n22308;
  assign n22310 = ~n6313 & ~n19175;
  assign n22311 = n9197 & ~n22310;
  assign n22312 = ~n9195 & ~n22311;
  assign n22313 = x7 & n19188;
  assign n22314 = n21518 & ~n22313;
  assign n22315 = n22312 & ~n22314;
  assign n22316 = ~n21519 & ~n22315;
  assign n22317 = ~n22309 & ~n22316;
  assign n22318 = n7515 & n19748;
  assign n22319 = n8029 & n19170;
  assign n22320 = n7518 & n19173;
  assign n22321 = n7520 & n19174;
  assign n22322 = ~n22320 & ~n22321;
  assign n22323 = ~n22319 & n22322;
  assign n22324 = ~n22318 & n22323;
  assign n22325 = n22324 ^ x5;
  assign n22326 = n15363 & ~n21519;
  assign n22327 = n22326 ^ n21517;
  assign n22328 = n7515 & ~n19761;
  assign n22329 = n8029 & ~n19167;
  assign n22330 = n7518 & n19170;
  assign n22331 = n7520 & n19173;
  assign n22332 = ~n22330 & ~n22331;
  assign n22333 = ~n22329 & n22332;
  assign n22334 = ~n22328 & n22333;
  assign n22335 = n22334 ^ n22324;
  assign n22336 = n22327 & n22335;
  assign n22337 = ~n22325 & n22336;
  assign n22338 = n22337 ^ n22325;
  assign n22339 = ~n22317 & ~n22338;
  assign n22340 = n22334 ^ x5;
  assign n22341 = n22340 ^ n22327;
  assign n22342 = n22309 & n22316;
  assign n22343 = n22342 ^ n22340;
  assign n22344 = n22341 & n22343;
  assign n22345 = n22344 ^ n22327;
  assign n22346 = ~n22339 & n22345;
  assign n22347 = n22346 ^ n22282;
  assign n22348 = ~n22283 & n22347;
  assign n22349 = n22348 ^ n22346;
  assign n22350 = n22349 ^ n22271;
  assign n22351 = n22272 & n22350;
  assign n22352 = n22351 ^ n22349;
  assign n22353 = n22352 ^ n22261;
  assign n22354 = ~n22262 & n22353;
  assign n22355 = n22354 ^ n22352;
  assign n22356 = n22355 ^ n22251;
  assign n22357 = ~n22252 & n22356;
  assign n22358 = n22357 ^ n22355;
  assign n22359 = n22358 ^ n22241;
  assign n22360 = n22242 & ~n22359;
  assign n22361 = n22360 ^ n22358;
  assign n22370 = n22369 ^ n22361;
  assign n22371 = n21576 ^ n21483;
  assign n22372 = n22371 ^ n22361;
  assign n22373 = n22370 & ~n22372;
  assign n22374 = n22373 ^ n22369;
  assign n22375 = n22374 ^ n22223;
  assign n22376 = n22232 & ~n22375;
  assign n22377 = n22376 ^ n22231;
  assign n22378 = n22377 ^ n22221;
  assign n22379 = n22222 & n22378;
  assign n22380 = n22379 ^ n22377;
  assign n22381 = n22380 ^ n22203;
  assign n22382 = n22212 & ~n22381;
  assign n22383 = n22382 ^ n22211;
  assign n22384 = n22383 ^ n22201;
  assign n22385 = ~n22202 & n22384;
  assign n22386 = n22385 ^ n22383;
  assign n22387 = n22386 ^ n22191;
  assign n22388 = ~n22192 & n22387;
  assign n22389 = n22388 ^ n22386;
  assign n22390 = n22389 ^ n22181;
  assign n22391 = ~n22182 & n22390;
  assign n22392 = n22391 ^ n22389;
  assign n22393 = n22392 ^ n22171;
  assign n22394 = ~n22172 & n22393;
  assign n22395 = n22394 ^ n22392;
  assign n22396 = n22395 ^ n22161;
  assign n22397 = n22162 & ~n22396;
  assign n22398 = n22397 ^ n22395;
  assign n22399 = n22398 ^ n22151;
  assign n22400 = ~n22152 & n22399;
  assign n22401 = n22400 ^ n22398;
  assign n22402 = n22401 ^ n22141;
  assign n22403 = ~n22142 & n22402;
  assign n22404 = n22403 ^ n22401;
  assign n22405 = n22404 ^ n22131;
  assign n22406 = ~n22132 & n22405;
  assign n22407 = n22406 ^ n22404;
  assign n22408 = n22407 ^ n22121;
  assign n22409 = ~n22122 & n22408;
  assign n22410 = n22409 ^ n22407;
  assign n22411 = n22410 ^ n22111;
  assign n22412 = ~n22112 & n22411;
  assign n22413 = n22412 ^ n22410;
  assign n22414 = n22413 ^ n22101;
  assign n22415 = n22102 & n22414;
  assign n22416 = n22415 ^ n22413;
  assign n22417 = n22416 ^ n22085;
  assign n22418 = ~n22086 & n22417;
  assign n22419 = n22418 ^ n22416;
  assign n22420 = n22419 ^ n22075;
  assign n22421 = ~n22076 & n22420;
  assign n22422 = n22421 ^ n22419;
  assign n22423 = n22422 ^ n22065;
  assign n22424 = n22066 & ~n22423;
  assign n22425 = n22424 ^ n22422;
  assign n22434 = n22433 ^ n22425;
  assign n22435 = n21707 ^ n21697;
  assign n22436 = n22435 ^ n22433;
  assign n22437 = n22434 & n22436;
  assign n22438 = n22437 ^ n22425;
  assign n22439 = ~n22048 & n22438;
  assign n22440 = ~n19304 & ~n19593;
  assign n22441 = n22440 ^ n19063;
  assign n22442 = n7515 & n22441;
  assign n22443 = n8029 & n19063;
  assign n22444 = n7520 & ~n19078;
  assign n22445 = n7518 & n19303;
  assign n22446 = ~n22444 & ~n22445;
  assign n22447 = ~n22443 & n22446;
  assign n22448 = ~n22442 & n22447;
  assign n22449 = n22448 ^ x5;
  assign n22450 = ~n22439 & ~n22449;
  assign n22451 = n22048 & ~n22438;
  assign n22452 = ~n22450 & ~n22451;
  assign n22469 = n22047 & ~n22452;
  assign n22470 = ~n22047 & n22449;
  assign n22471 = ~n22048 & n22470;
  assign n22472 = ~n22469 & ~n22471;
  assign n22951 = n22435 ^ n22434;
  assign n22484 = n22422 ^ n22066;
  assign n22478 = n33 & ~n22036;
  assign n22479 = n22478 ^ x1;
  assign n22480 = n22479 ^ n19368;
  assign n22474 = n19063 ^ x2;
  assign n22473 = x2 & ~n19303;
  assign n22475 = n22474 ^ n22473;
  assign n22476 = ~x1 & n22475;
  assign n22477 = n22476 ^ n22474;
  assign n22481 = n22480 ^ n22477;
  assign n22482 = ~x0 & ~n22481;
  assign n22483 = n22482 ^ n22480;
  assign n22485 = n22484 ^ n22483;
  assign n22931 = n22419 ^ n22076;
  assign n22916 = n33 & ~n19657;
  assign n22917 = n22916 ^ x1;
  assign n22918 = n22917 ^ n19303;
  assign n22919 = x0 & ~n22918;
  assign n22920 = n19078 ^ x2;
  assign n22921 = n9378 & n22920;
  assign n22922 = x2 & ~n19298;
  assign n22923 = n9448 & ~n22922;
  assign n22924 = ~n22921 & ~n22923;
  assign n22925 = ~n22919 & n22924;
  assign n22901 = n33 & ~n21714;
  assign n22902 = n22901 ^ x1;
  assign n22903 = n22902 ^ n19078;
  assign n22904 = x0 & n22903;
  assign n22905 = n19298 ^ x2;
  assign n22906 = x1 & n22905;
  assign n22907 = n9346 & ~n19096;
  assign n22908 = ~x0 & ~n22907;
  assign n22909 = ~n22906 & n22908;
  assign n22910 = ~n22904 & ~n22909;
  assign n22885 = n22410 ^ n22112;
  assign n22870 = n33 & ~n21698;
  assign n22871 = n22870 ^ x1;
  assign n22872 = n22871 ^ n19096;
  assign n22873 = x0 & ~n22872;
  assign n22874 = n19292 ^ x2;
  assign n22875 = x1 & n22874;
  assign n22876 = n9346 & ~n19104;
  assign n22877 = ~x0 & ~n22876;
  assign n22878 = ~n22875 & n22877;
  assign n22879 = ~n22873 & ~n22878;
  assign n22855 = n22404 ^ n22132;
  assign n22835 = n22398 ^ n22152;
  assign n22820 = n22395 ^ n22162;
  assign n22497 = n33 & ~n20293;
  assign n22498 = n22497 ^ x1;
  assign n22499 = n22498 ^ n19233;
  assign n22500 = x0 & ~n22499;
  assign n22501 = n19139 ^ x2;
  assign n22502 = n9378 & ~n22501;
  assign n22503 = x2 & n19142;
  assign n22504 = n9448 & ~n22503;
  assign n22505 = ~n22502 & ~n22504;
  assign n22506 = ~n22500 & n22505;
  assign n22507 = n22374 ^ n22232;
  assign n22508 = n22506 & ~n22507;
  assign n22520 = n9378 & ~n19225;
  assign n22521 = ~x1 & ~n19215;
  assign n22522 = n9431 & ~n22521;
  assign n22523 = ~n22520 & ~n22522;
  assign n22524 = n8886 & ~n19225;
  assign n22525 = ~n22523 & ~n22524;
  assign n22526 = n33 & ~n20044;
  assign n22527 = n22526 ^ x1;
  assign n22528 = n22527 ^ n19142;
  assign n22529 = x0 & ~n22528;
  assign n22530 = ~n22525 & ~n22529;
  assign n22519 = n22358 ^ n22242;
  assign n22531 = n22530 ^ n22519;
  assign n22542 = n22355 ^ n22252;
  assign n22536 = n33 & ~n20209;
  assign n22537 = n22536 ^ x1;
  assign n22538 = n22537 ^ n19225;
  assign n22532 = n19215 ^ x2;
  assign n22533 = x1 & ~n22532;
  assign n22534 = n9346 & ~n19160;
  assign n22535 = ~n22533 & ~n22534;
  assign n22539 = n22538 ^ n22535;
  assign n22540 = ~x0 & n22539;
  assign n22541 = n22540 ^ n22538;
  assign n22543 = n22542 ^ n22541;
  assign n22696 = n20020 ^ n19215;
  assign n22697 = n19215 ^ x1;
  assign n22698 = n22697 ^ x2;
  assign n22699 = n22698 ^ n20020;
  assign n22700 = n22696 & ~n22699;
  assign n22701 = n22700 ^ n22697;
  assign n22692 = n19160 ^ x2;
  assign n22691 = x2 & ~n19200;
  assign n22693 = n22692 ^ n22691;
  assign n22694 = ~x1 & n22693;
  assign n22695 = n22694 ^ n22692;
  assign n22702 = n22701 ^ n22695;
  assign n22703 = ~x0 & ~n22702;
  assign n22704 = n22703 ^ n22701;
  assign n22545 = n19200 ^ x2;
  assign n22546 = n9378 & ~n22545;
  assign n22547 = x2 & n19162;
  assign n22548 = n9448 & ~n22547;
  assign n22549 = ~n22546 & ~n22548;
  assign n22550 = n33 & ~n19965;
  assign n22551 = n22550 ^ x1;
  assign n22552 = n22551 ^ n19160;
  assign n22553 = x0 & ~n22552;
  assign n22554 = n22549 & ~n22553;
  assign n22544 = n22349 ^ n22272;
  assign n22555 = n22554 ^ n22544;
  assign n22566 = n22346 ^ n22283;
  assign n22560 = n33 & ~n19815;
  assign n22561 = n22560 ^ x1;
  assign n22562 = n22561 ^ n19200;
  assign n22556 = n19162 ^ x2;
  assign n22557 = x1 & ~n22556;
  assign n22558 = n9346 & n19201;
  assign n22559 = ~n22557 & ~n22558;
  assign n22563 = n22562 ^ n22559;
  assign n22564 = ~x0 & ~n22563;
  assign n22565 = n22564 ^ n22562;
  assign n22567 = n22566 ^ n22565;
  assign n22665 = n33 & ~n19827;
  assign n22666 = n22665 ^ x1;
  assign n22667 = n22666 ^ n19162;
  assign n22668 = x0 & ~n22667;
  assign n22669 = n9378 & ~n19201;
  assign n22670 = ~x1 & ~n19161;
  assign n22671 = n9431 & ~n22670;
  assign n22672 = ~n22669 & ~n22671;
  assign n22673 = n8886 & ~n19201;
  assign n22674 = ~n22672 & ~n22673;
  assign n22675 = ~n22668 & ~n22674;
  assign n22589 = n22306 ^ n22291;
  assign n22590 = n22589 ^ n22307;
  assign n22583 = n33 & ~n19798;
  assign n22584 = n22583 ^ x1;
  assign n22585 = n22584 ^ n19161;
  assign n22579 = n19167 ^ x2;
  assign n22580 = x1 & ~n22579;
  assign n22581 = n9346 & ~n19170;
  assign n22582 = ~n22580 & ~n22581;
  assign n22586 = n22585 ^ n22582;
  assign n22587 = ~x0 & n22586;
  assign n22588 = n22587 ^ n22585;
  assign n22591 = n22590 ^ n22588;
  assign n22592 = n33 & n19761;
  assign n22593 = ~n33 & n19167;
  assign n22594 = x0 & ~n22593;
  assign n22595 = ~n22592 & n22594;
  assign n22596 = n9378 & n19170;
  assign n22597 = n9380 & n19173;
  assign n22598 = ~n22596 & ~n22597;
  assign n22599 = ~n22595 & n22598;
  assign n22600 = n22599 ^ x2;
  assign n22601 = x5 & ~n22304;
  assign n22602 = n22601 ^ n22303;
  assign n22603 = n22600 & n22602;
  assign n22604 = n33 & ~n19748;
  assign n22605 = ~n33 & ~n19170;
  assign n22606 = x0 & ~n22605;
  assign n22607 = ~n22604 & n22606;
  assign n22608 = n9378 & n19173;
  assign n22609 = n9380 & n19174;
  assign n22610 = ~n22608 & ~n22609;
  assign n22611 = ~n22607 & n22610;
  assign n22612 = n22611 ^ x2;
  assign n22613 = ~n9530 & ~n19175;
  assign n22614 = n9532 & ~n22613;
  assign n22615 = ~n9529 & ~n22614;
  assign n22616 = n19188 & ~n22615;
  assign n22617 = x4 & n19188;
  assign n22618 = n22292 & ~n22617;
  assign n22619 = ~n22616 & ~n22618;
  assign n22620 = n22612 & n22619;
  assign n22621 = x2 & ~x3;
  assign n22622 = n33 & ~n19720;
  assign n22623 = ~n33 & ~n19173;
  assign n22624 = x0 & ~n22623;
  assign n22625 = ~n22622 & n22624;
  assign n22626 = n9378 & n19174;
  assign n22627 = n9380 & ~n19175;
  assign n22628 = ~n22626 & ~n22627;
  assign n22629 = ~n22625 & n22628;
  assign n22630 = ~n22621 & n22629;
  assign n22631 = n19188 & ~n22630;
  assign n22632 = ~x2 & x3;
  assign n22633 = ~n22629 & ~n22632;
  assign n22634 = n22631 & ~n22633;
  assign n22635 = ~n9448 & n19174;
  assign n22636 = x2 & n19875;
  assign n22637 = ~n22635 & n22636;
  assign n22638 = ~n22625 & n22637;
  assign n22639 = ~n22634 & ~n22638;
  assign n22640 = ~n22620 & ~n22639;
  assign n22641 = ~n22603 & n22640;
  assign n22642 = ~n22611 & ~n22619;
  assign n22643 = ~n22602 & n22642;
  assign n22644 = n22599 & ~n22643;
  assign n22645 = n22602 & ~n22642;
  assign n22646 = ~x2 & ~n22645;
  assign n22647 = ~n22644 & n22646;
  assign n22648 = n22611 & ~n22619;
  assign n22649 = ~n22602 & n22648;
  assign n22650 = ~n22599 & ~n22649;
  assign n22651 = n22602 & ~n22648;
  assign n22652 = x2 & ~n22651;
  assign n22653 = ~n22650 & n22652;
  assign n22654 = ~n22647 & ~n22653;
  assign n22655 = ~n22641 & n22654;
  assign n22656 = n22655 ^ n22590;
  assign n22657 = n22591 & ~n22656;
  assign n22658 = n22657 ^ n22588;
  assign n22573 = n33 & ~n19839;
  assign n22574 = n22573 ^ x1;
  assign n22575 = n22574 ^ n19201;
  assign n22569 = n19161 ^ x2;
  assign n22568 = x2 & n19167;
  assign n22570 = n22569 ^ n22568;
  assign n22571 = ~x1 & ~n22570;
  assign n22572 = n22571 ^ n22569;
  assign n22576 = n22575 ^ n22572;
  assign n22577 = ~x0 & n22576;
  assign n22578 = n22577 ^ n22575;
  assign n22659 = n22658 ^ n22578;
  assign n22660 = n22316 ^ n22309;
  assign n22661 = n22660 ^ n22325;
  assign n22662 = n22661 ^ n22578;
  assign n22663 = n22659 & ~n22662;
  assign n22664 = n22663 ^ n22658;
  assign n22676 = n22675 ^ n22664;
  assign n22680 = n22334 ^ n22327;
  assign n22677 = n22325 ^ n22316;
  assign n22678 = ~n22660 & ~n22677;
  assign n22679 = n22678 ^ n22324;
  assign n22681 = n22680 ^ n22679;
  assign n22682 = n22681 ^ n22675;
  assign n22683 = n22676 & ~n22682;
  assign n22684 = n22683 ^ n22664;
  assign n22685 = n22684 ^ n22566;
  assign n22686 = ~n22567 & ~n22685;
  assign n22687 = n22686 ^ n22565;
  assign n22688 = n22687 ^ n22544;
  assign n22689 = n22555 & ~n22688;
  assign n22690 = n22689 ^ n22554;
  assign n22705 = n22704 ^ n22690;
  assign n22706 = n22352 ^ n22262;
  assign n22707 = n22706 ^ n22690;
  assign n22708 = ~n22705 & n22707;
  assign n22709 = n22708 ^ n22704;
  assign n22710 = n22709 ^ n22542;
  assign n22711 = n22543 & ~n22710;
  assign n22712 = n22711 ^ n22541;
  assign n22713 = n22712 ^ n22519;
  assign n22714 = ~n22531 & n22713;
  assign n22715 = n22714 ^ n22530;
  assign n22513 = n33 & n20030;
  assign n22514 = n22513 ^ x1;
  assign n22515 = n22514 ^ n19139;
  assign n22509 = n19142 ^ x2;
  assign n22510 = x1 & ~n22509;
  assign n22511 = n9346 & n19225;
  assign n22512 = ~n22510 & ~n22511;
  assign n22516 = n22515 ^ n22512;
  assign n22517 = ~x0 & ~n22516;
  assign n22518 = n22517 ^ n22515;
  assign n22716 = n22715 ^ n22518;
  assign n22717 = n22371 ^ n22369;
  assign n22718 = n22717 ^ n22361;
  assign n22719 = n22718 ^ n22518;
  assign n22720 = ~n22716 & n22719;
  assign n22721 = n22720 ^ n22715;
  assign n22722 = ~n22508 & n22721;
  assign n22723 = n22377 ^ n22222;
  assign n22729 = n33 & ~n20327;
  assign n22730 = n22729 ^ x1;
  assign n22731 = n22730 ^ n19238;
  assign n22725 = n19233 ^ x2;
  assign n22724 = x2 & ~n19139;
  assign n22726 = n22725 ^ n22724;
  assign n22727 = ~x1 & n22726;
  assign n22728 = n22727 ^ n22725;
  assign n22732 = n22731 ^ n22728;
  assign n22733 = ~x0 & ~n22732;
  assign n22734 = n22733 ^ n22731;
  assign n22735 = ~n22723 & n22734;
  assign n22736 = ~n22506 & n22507;
  assign n22737 = ~n22735 & ~n22736;
  assign n22738 = ~n22722 & n22737;
  assign n22739 = n22723 & ~n22734;
  assign n22740 = ~n22738 & ~n22739;
  assign n22741 = n22380 ^ n22212;
  assign n22742 = ~n22740 & ~n22741;
  assign n22748 = n33 & ~n19695;
  assign n22749 = n22748 ^ x1;
  assign n22750 = n22749 ^ n19255;
  assign n22744 = n19253 ^ x2;
  assign n22743 = x2 & n19238;
  assign n22745 = n22744 ^ n22743;
  assign n22746 = ~x1 & n22745;
  assign n22747 = n22746 ^ n22744;
  assign n22751 = n22750 ^ n22747;
  assign n22752 = x0 & ~n22751;
  assign n22753 = n22752 ^ n22747;
  assign n22754 = ~n22742 & ~n22753;
  assign n22755 = n22383 ^ n22202;
  assign n22756 = ~n22754 & ~n22755;
  assign n22757 = n22740 & n22741;
  assign n22758 = n19238 ^ x2;
  assign n22759 = n9378 & n22758;
  assign n22760 = x2 & ~n19233;
  assign n22761 = n9448 & ~n22760;
  assign n22762 = ~n22759 & ~n22761;
  assign n22763 = n33 & ~n20307;
  assign n22764 = n22763 ^ x1;
  assign n22765 = n22764 ^ n19253;
  assign n22766 = x0 & ~n22765;
  assign n22767 = n22762 & ~n22766;
  assign n22768 = ~n22755 & n22767;
  assign n22769 = ~n22753 & ~n22768;
  assign n22770 = ~n22757 & ~n22769;
  assign n22771 = ~n22756 & ~n22770;
  assign n22772 = ~n22742 & ~n22767;
  assign n22773 = n22755 & n22772;
  assign n22774 = ~n22771 & ~n22773;
  assign n22775 = n22386 ^ n22192;
  assign n22780 = n33 & ~n20656;
  assign n22781 = n22780 ^ x1;
  assign n22782 = n22781 ^ n19260;
  assign n22776 = n19255 ^ x2;
  assign n22777 = x1 & ~n22776;
  assign n22778 = n9346 & ~n19253;
  assign n22779 = ~n22777 & ~n22778;
  assign n22783 = n22782 ^ n22779;
  assign n22784 = ~x0 & ~n22783;
  assign n22785 = n22784 ^ n22782;
  assign n22786 = ~n22775 & n22785;
  assign n22787 = ~n22774 & ~n22786;
  assign n22788 = n22389 ^ n22182;
  assign n22789 = n33 & ~n20792;
  assign n22790 = n22789 ^ x1;
  assign n22791 = n22790 ^ n19277;
  assign n22792 = x0 & ~n22791;
  assign n22793 = n19260 ^ x2;
  assign n22794 = x1 & n22793;
  assign n22795 = n9346 & n19255;
  assign n22796 = ~x0 & ~n22795;
  assign n22797 = ~n22794 & n22796;
  assign n22798 = ~n22792 & ~n22797;
  assign n22799 = n22788 & ~n22798;
  assign n22800 = n22775 & ~n22785;
  assign n22801 = ~n22799 & ~n22800;
  assign n22802 = ~n22787 & n22801;
  assign n22803 = ~n22788 & n22798;
  assign n22804 = ~n22802 & ~n22803;
  assign n22496 = n22392 ^ n22172;
  assign n22805 = n22804 ^ n22496;
  assign n22811 = n33 & ~n20907;
  assign n22812 = n22811 ^ x1;
  assign n22813 = n22812 ^ n19281;
  assign n22807 = n19277 ^ x2;
  assign n22806 = x2 & ~n19260;
  assign n22808 = n22807 ^ n22806;
  assign n22809 = ~x1 & n22808;
  assign n22810 = n22809 ^ n22807;
  assign n22814 = n22813 ^ n22810;
  assign n22815 = ~x0 & ~n22814;
  assign n22816 = n22815 ^ n22813;
  assign n22817 = n22816 ^ n22496;
  assign n22818 = n22805 & ~n22817;
  assign n22819 = n22818 ^ n22804;
  assign n22821 = n22820 ^ n22819;
  assign n22822 = n33 & ~n21188;
  assign n22823 = n22822 ^ x1;
  assign n22824 = n22823 ^ n19122;
  assign n22825 = x0 & ~n22824;
  assign n22826 = n19281 ^ x2;
  assign n22827 = x1 & ~n22826;
  assign n22828 = n9346 & ~n19277;
  assign n22829 = ~x0 & ~n22828;
  assign n22830 = ~n22827 & n22829;
  assign n22831 = ~n22825 & ~n22830;
  assign n22832 = n22831 ^ n22820;
  assign n22833 = ~n22821 & ~n22832;
  assign n22834 = n22833 ^ n22819;
  assign n22836 = n22835 ^ n22834;
  assign n22841 = n33 & ~n19677;
  assign n22842 = n22841 ^ x1;
  assign n22843 = n22842 ^ n19286;
  assign n22837 = n19122 ^ x2;
  assign n22838 = x1 & n22837;
  assign n22839 = n9346 & n19281;
  assign n22840 = ~n22838 & ~n22839;
  assign n22844 = n22843 ^ n22840;
  assign n22845 = ~x0 & n22844;
  assign n22846 = n22845 ^ n22843;
  assign n22847 = n22846 ^ n22835;
  assign n22848 = n22836 & ~n22847;
  assign n22849 = n22848 ^ n22834;
  assign n22490 = n33 & ~n21214;
  assign n22491 = n22490 ^ x1;
  assign n22492 = n22491 ^ n19104;
  assign n22486 = n19286 ^ x2;
  assign n22487 = x1 & ~n22486;
  assign n22488 = n9346 & ~n19122;
  assign n22489 = ~n22487 & ~n22488;
  assign n22493 = n22492 ^ n22489;
  assign n22494 = ~x0 & ~n22493;
  assign n22495 = n22494 ^ n22492;
  assign n22850 = n22849 ^ n22495;
  assign n22851 = n22401 ^ n22142;
  assign n22852 = n22851 ^ n22495;
  assign n22853 = ~n22850 & n22852;
  assign n22854 = n22853 ^ n22849;
  assign n22856 = n22855 ^ n22854;
  assign n22861 = n33 & ~n21683;
  assign n22862 = n22861 ^ x1;
  assign n22863 = n22862 ^ n19292;
  assign n22857 = n19104 ^ x2;
  assign n22858 = x1 & n22857;
  assign n22859 = n9346 & n19286;
  assign n22860 = ~n22858 & ~n22859;
  assign n22864 = n22863 ^ n22860;
  assign n22865 = ~x0 & ~n22864;
  assign n22866 = n22865 ^ n22863;
  assign n22867 = n22866 ^ n22855;
  assign n22868 = n22856 & n22867;
  assign n22869 = n22868 ^ n22854;
  assign n22880 = n22879 ^ n22869;
  assign n22881 = n22407 ^ n22122;
  assign n22882 = n22881 ^ n22879;
  assign n22883 = ~n22880 & n22882;
  assign n22884 = n22883 ^ n22869;
  assign n22886 = n22885 ^ n22884;
  assign n22892 = n33 & ~n19667;
  assign n22893 = n22892 ^ x1;
  assign n22894 = n22893 ^ n19298;
  assign n22888 = n19096 ^ x2;
  assign n22887 = x2 & ~n19292;
  assign n22889 = n22888 ^ n22887;
  assign n22890 = ~x1 & n22889;
  assign n22891 = n22890 ^ n22888;
  assign n22895 = n22894 ^ n22891;
  assign n22896 = ~x0 & n22895;
  assign n22897 = n22896 ^ n22894;
  assign n22898 = n22897 ^ n22885;
  assign n22899 = n22886 & n22898;
  assign n22900 = n22899 ^ n22884;
  assign n22911 = n22910 ^ n22900;
  assign n22912 = n22413 ^ n22102;
  assign n22913 = n22912 ^ n22910;
  assign n22914 = ~n22911 & ~n22913;
  assign n22915 = n22914 ^ n22900;
  assign n22926 = n22925 ^ n22915;
  assign n22927 = n22416 ^ n22086;
  assign n22928 = n22927 ^ n22925;
  assign n22929 = ~n22926 & n22928;
  assign n22930 = n22929 ^ n22915;
  assign n22932 = n22931 ^ n22930;
  assign n22933 = n33 & ~n22440;
  assign n22934 = n22933 ^ x1;
  assign n22935 = n22934 ^ n19063;
  assign n22936 = x0 & n22935;
  assign n22937 = x2 & n19078;
  assign n22938 = ~x1 & ~n22937;
  assign n22939 = ~x0 & ~n22938;
  assign n22940 = n8886 ^ x2;
  assign n22941 = n19303 & ~n22940;
  assign n22942 = n22941 ^ x2;
  assign n22943 = n22939 & n22942;
  assign n22944 = ~n22936 & ~n22943;
  assign n22945 = n22944 ^ n22931;
  assign n22946 = n22932 & ~n22945;
  assign n22947 = n22946 ^ n22930;
  assign n22948 = n22947 ^ n22483;
  assign n22949 = ~n22485 & ~n22948;
  assign n22950 = n22949 ^ n22484;
  assign n22952 = n22951 ^ n22950;
  assign n22953 = ~x1 & n19063;
  assign n22954 = n9431 & ~n22953;
  assign n22955 = n9378 & ~n19368;
  assign n22956 = ~n22954 & ~n22955;
  assign n22957 = n8886 & ~n19368;
  assign n22958 = ~n22956 & ~n22957;
  assign n19369 = ~n19305 & n19368;
  assign n19595 = ~n19368 & ~n19594;
  assign n22456 = ~n19369 & ~n19595;
  assign n22959 = n33 & ~n22456;
  assign n22960 = n22959 ^ x1;
  assign n19429 = n119 & n12019;
  assign n19431 = x26 & n12019;
  assign n19430 = x26 & ~n690;
  assign n19432 = n19431 ^ n19430;
  assign n19433 = ~n5451 & ~n19432;
  assign n19434 = n19433 ^ n19431;
  assign n19435 = ~n19429 & n19434;
  assign n19426 = n19344 ^ n19314;
  assign n19427 = ~n19353 & n19426;
  assign n19428 = n19427 ^ n19352;
  assign n19436 = n19435 ^ n19428;
  assign n19417 = n44 & ~n11941;
  assign n19418 = n3280 & ~n11940;
  assign n19419 = n3277 & n11902;
  assign n19420 = n3275 & ~n11875;
  assign n19421 = ~n19419 & ~n19420;
  assign n19422 = ~n19418 & n19421;
  assign n19423 = ~n19417 & n19422;
  assign n19424 = n19423 ^ x29;
  assign n19403 = n19332 & n19342;
  assign n19404 = n11995 & ~n19403;
  assign n19405 = ~n19332 & ~n19342;
  assign n19406 = ~n11991 & ~n19405;
  assign n19407 = ~n19404 & n19406;
  assign n19408 = n19342 ^ n11993;
  assign n19409 = n11991 & ~n19332;
  assign n19410 = n19409 ^ n19342;
  assign n19411 = n19408 & ~n19410;
  assign n19412 = n19411 ^ n11993;
  assign n19413 = ~n19407 & ~n19412;
  assign n19389 = n2477 & n2584;
  assign n19390 = n1498 & n19389;
  assign n19391 = ~n206 & n1902;
  assign n19392 = n19390 & n19391;
  assign n19393 = n3251 & n19392;
  assign n19394 = ~n278 & ~n518;
  assign n19395 = ~n850 & n19394;
  assign n19396 = n2038 & n19395;
  assign n19397 = n3290 & n4902;
  assign n19398 = n19396 & n19397;
  assign n19399 = n5598 & n19398;
  assign n19400 = n11744 & n19399;
  assign n19401 = n19393 & n19400;
  assign n19402 = n3161 & n19401;
  assign n19414 = n19413 ^ n19402;
  assign n19379 = n41 & ~n11777;
  assign n19380 = x31 & ~n19336;
  assign n19381 = n91 & n11480;
  assign n19382 = n19380 & ~n19381;
  assign n19383 = ~n19379 & n19382;
  assign n19384 = n41 & ~n11773;
  assign n19385 = n54 & n11480;
  assign n19386 = ~x31 & ~n19385;
  assign n19387 = ~n19384 & n19386;
  assign n19388 = ~n19383 & ~n19387;
  assign n19415 = n19414 ^ n19388;
  assign n19376 = n11991 ^ n40;
  assign n19377 = ~n19332 & n19376;
  assign n19378 = n19377 ^ n11991;
  assign n19416 = n19415 ^ n19378;
  assign n19425 = n19424 ^ n19416;
  assign n19437 = n19436 ^ n19425;
  assign n19373 = n19361 ^ n19311;
  assign n19374 = n19362 & n19373;
  assign n19375 = n19374 ^ n19311;
  assign n19438 = n19437 ^ n19375;
  assign n19370 = n19367 ^ n19308;
  assign n19371 = n19364 & ~n19370;
  assign n19372 = n19371 ^ n19367;
  assign n19439 = n19438 ^ n19372;
  assign n22961 = n22960 ^ n19439;
  assign n22962 = x0 & n22961;
  assign n22963 = ~n22958 & ~n22962;
  assign n22964 = n22963 ^ n22950;
  assign n22965 = n22952 & n22964;
  assign n22966 = n22965 ^ n22951;
  assign n19440 = ~n19369 & n19439;
  assign n19596 = ~n19439 & ~n19595;
  assign n22971 = ~n19440 & ~n19596;
  assign n22972 = n33 & ~n22971;
  assign n22973 = n22972 ^ x1;
  assign n19492 = n19375 & ~n19425;
  assign n19493 = n19372 & ~n19492;
  assign n19494 = ~n19375 & n19425;
  assign n19495 = n19494 ^ n19435;
  assign n19496 = ~n19436 & ~n19495;
  assign n19497 = n19496 ^ n19428;
  assign n19498 = n19493 & ~n19497;
  assign n19499 = ~n19428 & n19435;
  assign n19500 = n19425 ^ n19375;
  assign n19501 = n19428 & ~n19435;
  assign n19502 = n19501 ^ n19425;
  assign n19503 = ~n19500 & n19502;
  assign n19504 = n19503 ^ n19375;
  assign n19505 = ~n19499 & n19504;
  assign n19506 = ~n19372 & n19505;
  assign n19507 = ~n19492 & ~n19499;
  assign n19508 = ~n19494 & ~n19501;
  assign n19509 = ~n19507 & ~n19508;
  assign n19510 = ~n19506 & ~n19509;
  assign n19511 = ~n19498 & n19510;
  assign n19472 = n19378 & ~n19388;
  assign n19473 = ~n19402 & n19413;
  assign n19474 = n19473 ^ n19414;
  assign n19475 = n19424 & ~n19474;
  assign n19476 = n19475 ^ n19414;
  assign n19477 = ~n19472 & ~n19476;
  assign n19482 = ~n19378 & n19388;
  assign n19483 = n19473 ^ n19402;
  assign n19484 = ~n19482 & n19483;
  assign n19485 = n19484 ^ n19402;
  assign n19478 = n19388 ^ n19378;
  assign n19479 = n19402 & ~n19413;
  assign n19480 = n19479 ^ n19378;
  assign n19481 = n19478 & ~n19480;
  assign n19486 = n19485 ^ n19481;
  assign n19487 = n19424 & n19486;
  assign n19488 = n19487 ^ n19485;
  assign n19489 = ~n19477 & ~n19488;
  assign n19461 = n41 & ~n12000;
  assign n19462 = n91 & ~n11773;
  assign n19463 = x31 & ~n19385;
  assign n19464 = ~n19462 & n19463;
  assign n19465 = ~n19461 & n19464;
  assign n19466 = n41 & ~n11875;
  assign n19467 = n54 & ~n11773;
  assign n19468 = ~x31 & ~n19467;
  assign n19469 = ~n19466 & n19468;
  assign n19470 = ~n19465 & ~n19469;
  assign n19451 = ~n226 & ~n593;
  assign n19452 = ~n347 & ~n709;
  assign n19453 = n19451 & n19452;
  assign n19454 = n1440 & n12864;
  assign n19455 = n19453 & n19454;
  assign n19456 = n999 & n19455;
  assign n19457 = n3305 & n19456;
  assign n19458 = n3397 & n19457;
  assign n19459 = n11745 & n19458;
  assign n19460 = n3245 & n19459;
  assign n19471 = n19470 ^ n19460;
  assign n19490 = n19489 ^ n19471;
  assign n19442 = n43 & n12013;
  assign n19443 = n42 & ~n12019;
  assign n19444 = ~n19442 & n19443;
  assign n19445 = n3277 & ~n11940;
  assign n19446 = n3275 & n11902;
  assign n19447 = ~n19445 & ~n19446;
  assign n19448 = ~n19444 & n19447;
  assign n19449 = n19448 ^ x29;
  assign n19441 = ~n5451 & ~n19430;
  assign n19450 = n19449 ^ n19441;
  assign n19491 = n19490 ^ n19450;
  assign n19512 = n19511 ^ n19491;
  assign n22974 = n22973 ^ n19512;
  assign n22967 = n19439 ^ x2;
  assign n22968 = x1 & n22967;
  assign n22969 = n9346 & n19368;
  assign n22970 = ~n22968 & ~n22969;
  assign n22975 = n22974 ^ n22970;
  assign n22976 = ~x0 & n22975;
  assign n22977 = n22976 ^ n22974;
  assign n22978 = n22966 & ~n22977;
  assign n22979 = ~n22472 & n22978;
  assign n22980 = ~n22966 & n22977;
  assign n22981 = n22451 ^ n22450;
  assign n22982 = n22047 & ~n22981;
  assign n22983 = n22982 ^ n22450;
  assign n22984 = ~n22980 & ~n22983;
  assign n22985 = n22438 ^ n22048;
  assign n22986 = n22449 & n22985;
  assign n22987 = n22984 & ~n22986;
  assign n22988 = ~n22979 & ~n22987;
  assign n19513 = ~n19440 & n19512;
  assign n19597 = ~n19512 & ~n19596;
  assign n22989 = ~n19513 & ~n19597;
  assign n22990 = n33 & ~n22989;
  assign n22991 = n22990 ^ x1;
  assign n19566 = ~n19491 & ~n19501;
  assign n19567 = ~n19494 & ~n19566;
  assign n19568 = ~n19493 & n19567;
  assign n19569 = ~n19491 & ~n19492;
  assign n19570 = ~n19499 & ~n19569;
  assign n19571 = ~n19372 & n19570;
  assign n19572 = n19491 & n19497;
  assign n19573 = ~n19571 & ~n19572;
  assign n19574 = ~n19568 & n19573;
  assign n19549 = n19413 & ~n19424;
  assign n19550 = ~n19471 & ~n19549;
  assign n19551 = ~n19472 & ~n19550;
  assign n19552 = ~n19413 & n19424;
  assign n19553 = ~n19471 & ~n19482;
  assign n19554 = ~n19552 & ~n19553;
  assign n19555 = ~n19551 & ~n19554;
  assign n19556 = n19402 & ~n19555;
  assign n19557 = ~n19402 & ~n19471;
  assign n19558 = ~n19552 & n19557;
  assign n19559 = ~n19482 & ~n19558;
  assign n19560 = ~n19472 & n19557;
  assign n19561 = ~n19549 & ~n19560;
  assign n19562 = ~n19559 & ~n19561;
  assign n19563 = ~n19556 & ~n19562;
  assign n19534 = ~x29 & n17383;
  assign n19535 = n42 & ~n574;
  assign n19536 = ~n19534 & n19535;
  assign n19537 = n6177 & ~n11940;
  assign n19538 = x29 & n6475;
  assign n19539 = ~x28 & ~n19538;
  assign n19540 = ~n19537 & n19539;
  assign n19541 = ~x26 & x29;
  assign n19542 = x28 & ~n19541;
  assign n19543 = ~n19540 & ~n19542;
  assign n19544 = ~n1507 & ~n6178;
  assign n19545 = ~x29 & ~n19544;
  assign n19546 = ~n19543 & ~n19545;
  assign n19547 = ~n19536 & n19546;
  assign n19526 = n3667 & n12504;
  assign n19527 = n3676 & n11902;
  assign n19528 = ~n54 & ~n3672;
  assign n19529 = ~n11875 & ~n19528;
  assign n19530 = ~n19527 & ~n19529;
  assign n19531 = ~n19526 & n19530;
  assign n19519 = n3424 & n3873;
  assign n19520 = ~n79 & n19519;
  assign n19521 = ~n709 & n1240;
  assign n19522 = n19520 & n19521;
  assign n19523 = n3384 & n19522;
  assign n19524 = n3391 & n19523;
  assign n19525 = n19524 ^ n19441;
  assign n19532 = n19531 ^ n19525;
  assign n19517 = n19470 ^ n19402;
  assign n19518 = n19471 & n19517;
  assign n19533 = n19532 ^ n19518;
  assign n19548 = n19547 ^ n19533;
  assign n19564 = n19563 ^ n19548;
  assign n19514 = n19490 ^ n19449;
  assign n19515 = n19450 & ~n19514;
  assign n19516 = n19515 ^ n19490;
  assign n19565 = n19564 ^ n19516;
  assign n19575 = n19574 ^ n19565;
  assign n22992 = n22991 ^ n19575;
  assign n22993 = x0 & n22992;
  assign n22994 = n19512 ^ x2;
  assign n22995 = x1 & ~n22994;
  assign n22996 = ~x0 & ~n22995;
  assign n22997 = n9346 & ~n19439;
  assign n22998 = n22996 & ~n22997;
  assign n22999 = ~n22993 & ~n22998;
  assign n23000 = ~n22988 & n22999;
  assign n23001 = n22048 & ~n22449;
  assign n23002 = ~n22047 & ~n23001;
  assign n23003 = n22980 & ~n23002;
  assign n23004 = ~n22469 & n23003;
  assign n23005 = n22047 & ~n22439;
  assign n23006 = ~n22449 & n22985;
  assign n23007 = ~n23005 & ~n23006;
  assign n23008 = ~n22978 & n23007;
  assign n23009 = ~n22451 & n22470;
  assign n23010 = n23008 & ~n23009;
  assign n23011 = ~n23004 & ~n23010;
  assign n23012 = ~n22999 & ~n23011;
  assign n23013 = ~n23000 & ~n23012;
  assign n22457 = n22456 ^ n19439;
  assign n22458 = n7515 & n22457;
  assign n22459 = n8029 & n19439;
  assign n22460 = n7518 & ~n19368;
  assign n22461 = n7520 & n19063;
  assign n22462 = ~n22460 & ~n22461;
  assign n22463 = ~n22459 & n22462;
  assign n22464 = ~n22458 & n22463;
  assign n22465 = n22464 ^ x5;
  assign n22453 = n22452 ^ n22046;
  assign n22454 = n22047 & ~n22453;
  assign n22455 = n22454 ^ n22452;
  assign n22466 = n22465 ^ n22455;
  assign n22024 = n5814 & n21699;
  assign n22025 = n6295 & n19096;
  assign n22026 = n5817 & n19292;
  assign n22027 = n5824 & n19104;
  assign n22028 = ~n22026 & ~n22027;
  assign n22029 = ~n22025 & n22028;
  assign n22030 = ~n22024 & n22029;
  assign n22031 = n22030 ^ x11;
  assign n22021 = n21874 ^ n21863;
  assign n22022 = n21875 & n22021;
  assign n22023 = n22022 ^ n21866;
  assign n22032 = n22031 ^ n22023;
  assign n21934 = n21775 & n21847;
  assign n21974 = n3285 & n20020;
  assign n21975 = n3435 & n19160;
  assign n21976 = n3437 & ~n19215;
  assign n21977 = ~n3440 & n19200;
  assign n21978 = ~n21976 & ~n21977;
  assign n21979 = ~n21975 & n21978;
  assign n21980 = ~n21974 & n21979;
  assign n21981 = n21980 ^ x26;
  assign n21964 = n44 & ~n19828;
  assign n21965 = n3280 & ~n19162;
  assign n21966 = n3277 & ~n19201;
  assign n21967 = n3275 & ~n19161;
  assign n21968 = ~n21966 & ~n21967;
  assign n21969 = ~n21965 & n21968;
  assign n21970 = ~n21964 & n21969;
  assign n21971 = n21970 ^ x29;
  assign n21955 = n41 & ~n19761;
  assign n21956 = ~n21814 & ~n21955;
  assign n21957 = x31 & ~n21956;
  assign n21958 = n3676 & ~n19167;
  assign n21959 = ~n3673 & n19170;
  assign n21960 = ~n21958 & ~n21959;
  assign n21961 = ~n21957 & n21960;
  assign n21941 = n4048 & n12216;
  assign n21942 = n1273 & n3039;
  assign n21943 = n21941 & n21942;
  assign n21944 = n11649 & n21943;
  assign n21945 = n4757 & n21944;
  assign n21946 = n294 & ~n558;
  assign n21947 = n4744 & n21946;
  assign n21948 = ~n369 & n1514;
  assign n21949 = n1590 & n21948;
  assign n21950 = n21947 & n21949;
  assign n21951 = n3513 & n21950;
  assign n21952 = n21945 & n21951;
  assign n21953 = n4400 & n21952;
  assign n21954 = n11535 & n21953;
  assign n21962 = n21961 ^ n21954;
  assign n21938 = n21807 ^ n21792;
  assign n21939 = ~n21818 & ~n21938;
  assign n21940 = n21939 ^ n21817;
  assign n21963 = n21962 ^ n21940;
  assign n21972 = n21971 ^ n21963;
  assign n21935 = n21827 ^ n21789;
  assign n21936 = n21828 & n21935;
  assign n21937 = n21936 ^ n21789;
  assign n21973 = n21972 ^ n21937;
  assign n21982 = n21981 ^ n21973;
  assign n21984 = n21786 & ~n21829;
  assign n21985 = ~n21783 & ~n21984;
  assign n21986 = ~n21786 & n21829;
  assign n21987 = ~n21985 & ~n21986;
  assign n21983 = ~n21783 & n21829;
  assign n21988 = n21987 ^ n21983;
  assign n21989 = ~n21982 & n21988;
  assign n21990 = n21989 ^ n21987;
  assign n21991 = n21934 & n21990;
  assign n21992 = ~n21775 & ~n21847;
  assign n21996 = n21783 & n21984;
  assign n21993 = n21783 & ~n21829;
  assign n21994 = ~n21831 & n21993;
  assign n21995 = n21994 ^ n21831;
  assign n21997 = n21996 ^ n21995;
  assign n21998 = n21982 & ~n21997;
  assign n21999 = n21998 ^ n21995;
  assign n22000 = ~n21992 & ~n21999;
  assign n22001 = ~n21991 & ~n22000;
  assign n22002 = n21982 & ~n21987;
  assign n22003 = ~n21982 & n21993;
  assign n22004 = ~n22002 & ~n22003;
  assign n22005 = n21992 & ~n22004;
  assign n22006 = n21783 & n21830;
  assign n22007 = n21986 ^ n21985;
  assign n22008 = n21982 & ~n22007;
  assign n22009 = n22008 ^ n21985;
  assign n22010 = ~n22006 & ~n22009;
  assign n22011 = ~n21934 & n22010;
  assign n22012 = ~n22005 & ~n22011;
  assign n22013 = n22001 & n22012;
  assign n21926 = n4478 & ~n20031;
  assign n21927 = n4487 & n19139;
  assign n21928 = n4484 & ~n19142;
  assign n21929 = n4480 & ~n19225;
  assign n21930 = ~n21928 & ~n21929;
  assign n21931 = ~n21927 & n21930;
  assign n21932 = ~n21926 & n21931;
  assign n21933 = n21932 ^ x23;
  assign n22014 = n22013 ^ n21933;
  assign n21918 = n4673 & n20308;
  assign n21919 = n4688 & n19253;
  assign n21920 = n4685 & ~n19238;
  assign n21921 = ~n4681 & n19233;
  assign n21922 = ~n21920 & ~n21921;
  assign n21923 = ~n21919 & n21922;
  assign n21924 = ~n21918 & n21923;
  assign n21925 = n21924 ^ x20;
  assign n22015 = n22014 ^ n21925;
  assign n21915 = n21857 ^ n21772;
  assign n21916 = n21858 & n21915;
  assign n21917 = n21916 ^ n21772;
  assign n22016 = n22015 ^ n21917;
  assign n21907 = n4963 & n20793;
  assign n21908 = n4972 & n19277;
  assign n21909 = n4976 & n19260;
  assign n21910 = n4970 & ~n19255;
  assign n21911 = ~n21909 & ~n21910;
  assign n21912 = ~n21908 & n21911;
  assign n21913 = ~n21907 & n21912;
  assign n21914 = n21913 ^ x17;
  assign n22017 = n22016 ^ n21914;
  assign n21904 = n21859 ^ n21753;
  assign n21905 = n21860 & ~n21904;
  assign n21906 = n21905 ^ n21753;
  assign n22018 = n22017 ^ n21906;
  assign n21883 = ~x13 & n19122;
  assign n21884 = n13719 & ~n19281;
  assign n21885 = n5742 & ~n21884;
  assign n21886 = ~n21883 & n21885;
  assign n21887 = n13989 & ~n19281;
  assign n21888 = n5744 & ~n21887;
  assign n21889 = ~n21737 & n21888;
  assign n21890 = ~n21886 & ~n21889;
  assign n21891 = ~x14 & n21890;
  assign n21892 = ~n19286 & n21891;
  assign n21893 = n7860 & n19678;
  assign n21894 = ~n21892 & ~n21893;
  assign n21895 = ~x13 & n21894;
  assign n21896 = ~n19678 & n21891;
  assign n21897 = n7860 & n19286;
  assign n21898 = x13 & ~n21897;
  assign n21899 = ~n21896 & n21898;
  assign n21900 = ~n21895 & ~n21899;
  assign n21901 = n18732 & n21890;
  assign n21902 = n21901 ^ x14;
  assign n21903 = ~n21900 & ~n21902;
  assign n22019 = n22018 ^ n21903;
  assign n21880 = n21861 ^ n21735;
  assign n21881 = n21862 & ~n21880;
  assign n21882 = n21881 ^ n21735;
  assign n22020 = n22019 ^ n21882;
  assign n22033 = n22032 ^ n22020;
  assign n21877 = n21876 ^ n21731;
  assign n21878 = n21732 & n21877;
  assign n21879 = n21878 ^ n21713;
  assign n22034 = n22033 ^ n21879;
  assign n19659 = n6306 & n19658;
  assign n19660 = n6309 & ~n19078;
  assign n19661 = n7168 & n19303;
  assign n19662 = n6316 & n19298;
  assign n19663 = ~n19661 & ~n19662;
  assign n19664 = ~n19660 & n19663;
  assign n19665 = ~n19659 & n19664;
  assign n19666 = n19665 ^ x8;
  assign n22035 = n22034 ^ n19666;
  assign n22467 = n22466 ^ n22035;
  assign n19633 = n19516 & n19574;
  assign n19634 = ~n19533 & ~n19547;
  assign n19635 = n19563 & n19634;
  assign n19636 = ~n19633 & n19635;
  assign n19637 = ~n19516 & ~n19574;
  assign n19638 = n19533 & n19547;
  assign n19639 = ~n19563 & n19638;
  assign n19640 = ~n19637 & n19639;
  assign n19641 = ~n19636 & ~n19640;
  assign n19642 = n19574 ^ n19516;
  assign n19643 = n19563 ^ n19547;
  assign n19644 = ~n19548 & ~n19643;
  assign n19645 = n19644 ^ n19563;
  assign n19646 = n19645 ^ n19516;
  assign n19647 = ~n19642 & n19646;
  assign n19648 = n19641 & ~n19647;
  assign n19618 = n19460 & ~n19470;
  assign n19619 = n19525 & ~n19531;
  assign n19620 = n19618 & ~n19619;
  assign n19621 = ~n19525 & n19531;
  assign n19622 = n19402 & ~n19621;
  assign n19623 = ~n19620 & n19622;
  assign n19624 = ~n19460 & n19470;
  assign n19625 = n19624 ^ n19531;
  assign n19626 = ~n19402 & ~n19525;
  assign n19627 = n19626 ^ n19531;
  assign n19628 = ~n19625 & n19627;
  assign n19629 = n19628 ^ n19624;
  assign n19630 = ~n19623 & ~n19629;
  assign n19616 = x29 & n6179;
  assign n19617 = n19616 ^ n6178;
  assign n19631 = n19630 ^ n19617;
  assign n19608 = n11906 & ~n11940;
  assign n19609 = ~n19467 & ~n19608;
  assign n19610 = x31 & ~n19609;
  assign n19611 = n3676 & ~n11940;
  assign n19612 = ~n3673 & n11902;
  assign n19613 = ~n19611 & ~n19612;
  assign n19614 = ~n19610 & n19613;
  assign n19605 = n3871 & n19520;
  assign n19606 = n3364 & n19605;
  assign n19602 = n19441 ^ n19402;
  assign n19603 = ~n19525 & n19602;
  assign n19604 = n19603 ^ n19402;
  assign n19607 = n19606 ^ n19604;
  assign n19615 = n19614 ^ n19607;
  assign n19632 = n19631 ^ n19615;
  assign n19649 = n19648 ^ n19632;
  assign n19576 = ~n19513 & ~n19575;
  assign n19598 = n19575 & ~n19597;
  assign n19599 = ~n19576 & ~n19598;
  assign n19600 = n33 & ~n19599;
  assign n19601 = n19600 ^ x1;
  assign n19650 = n19649 ^ n19601;
  assign n19651 = x0 & n19650;
  assign n19652 = n19575 ^ x2;
  assign n19653 = n9378 & ~n19652;
  assign n19654 = n9380 & n19512;
  assign n19655 = ~n19653 & ~n19654;
  assign n19656 = ~n19651 & n19655;
  assign n22468 = n22467 ^ n19656;
  assign n23014 = n23013 ^ n22468;
  assign n23239 = n21932 & n22013;
  assign n23240 = n22012 ^ n22001;
  assign n23241 = x23 & n23240;
  assign n23242 = n23241 ^ n22001;
  assign n23243 = ~n23239 & n23242;
  assign n23231 = n4478 & n20294;
  assign n23232 = n4487 & n19233;
  assign n23233 = n4484 & n19139;
  assign n23234 = n4480 & ~n19142;
  assign n23235 = ~n23233 & ~n23234;
  assign n23236 = ~n23232 & n23235;
  assign n23237 = ~n23231 & n23236;
  assign n23221 = n12417 & ~n20210;
  assign n23214 = ~n3440 & n19160;
  assign n23215 = n3435 & ~n19215;
  assign n23216 = ~n23214 & ~n23215;
  assign n23217 = x26 & n23216;
  assign n23222 = n19225 & n23217;
  assign n23223 = ~n23221 & ~n23222;
  assign n23218 = n20210 & n23217;
  assign n23219 = n12417 & ~n19225;
  assign n23220 = ~n23218 & ~n23219;
  assign n23224 = n23223 ^ n23220;
  assign n23225 = ~x25 & n23224;
  assign n23226 = n23225 ^ n23223;
  assign n23227 = ~n12432 & n23216;
  assign n23228 = n23227 ^ x26;
  assign n23229 = n23226 & n23228;
  assign n23186 = ~n54 & n19761;
  assign n23187 = ~n19170 & ~n23186;
  assign n23188 = ~n19167 & ~n23187;
  assign n23189 = n41 & n19179;
  assign n23190 = ~n23188 & ~n23189;
  assign n23191 = ~n19161 & ~n23190;
  assign n23192 = n19167 & ~n19760;
  assign n23193 = n19161 & n23192;
  assign n23194 = ~n54 & ~n23193;
  assign n23195 = ~n91 & n19170;
  assign n23196 = ~n23194 & n23195;
  assign n23197 = ~n23191 & ~n23196;
  assign n23198 = ~n54 & ~n19170;
  assign n23199 = ~n19761 & n23198;
  assign n23200 = n19161 & n23199;
  assign n23201 = ~n91 & ~n23200;
  assign n23202 = ~n19167 & ~n23201;
  assign n23203 = x31 & ~n23202;
  assign n23204 = n23197 & n23203;
  assign n23205 = n41 & ~n19161;
  assign n23206 = n54 & ~n19167;
  assign n23207 = ~x31 & ~n23206;
  assign n23208 = ~n23205 & n23207;
  assign n23209 = ~n23204 & ~n23208;
  assign n23168 = ~n323 & ~n920;
  assign n23169 = ~n1005 & n23168;
  assign n23170 = n4762 & n23169;
  assign n23171 = n1029 & n12226;
  assign n23172 = n857 & n1192;
  assign n23173 = n23171 & n23172;
  assign n23174 = n23170 & n23173;
  assign n23175 = n5657 & n23174;
  assign n23176 = n2228 & n3064;
  assign n23177 = n2895 & n3606;
  assign n23178 = n1273 & n23177;
  assign n23179 = n23176 & n23178;
  assign n23180 = n5501 & n23179;
  assign n23181 = n23175 & n23180;
  assign n23182 = n848 & n23181;
  assign n23183 = n3018 & n12248;
  assign n23184 = n23182 & n23183;
  assign n23165 = n21954 ^ n21940;
  assign n23166 = n21962 & n23165;
  assign n23167 = n23166 ^ n21961;
  assign n23185 = n23184 ^ n23167;
  assign n23210 = n23209 ^ n23185;
  assign n23162 = n21963 ^ n21937;
  assign n23163 = ~n21972 & n23162;
  assign n23164 = n23163 ^ n21971;
  assign n23211 = n23210 ^ n23164;
  assign n23154 = n44 & n19816;
  assign n23155 = n3280 & n19200;
  assign n23156 = n3277 & ~n19162;
  assign n23157 = n3275 & ~n19201;
  assign n23158 = ~n23156 & ~n23157;
  assign n23159 = ~n23155 & n23158;
  assign n23160 = ~n23154 & n23159;
  assign n23161 = n23160 ^ x29;
  assign n23212 = n23211 ^ n23161;
  assign n23151 = n21987 ^ n21973;
  assign n23152 = ~n21982 & n23151;
  assign n23153 = n23152 ^ n21981;
  assign n23213 = n23212 ^ n23153;
  assign n23230 = n23229 ^ n23213;
  assign n23238 = n23237 ^ n23230;
  assign n23244 = n23243 ^ n23238;
  assign n23143 = n4673 & ~n19696;
  assign n23144 = n4688 & ~n19255;
  assign n23145 = n4685 & n19253;
  assign n23146 = ~n4681 & ~n19238;
  assign n23147 = ~n23145 & ~n23146;
  assign n23148 = ~n23144 & n23147;
  assign n23149 = ~n23143 & n23148;
  assign n23150 = n23149 ^ x20;
  assign n23245 = n23244 ^ n23150;
  assign n23140 = n22014 ^ n21917;
  assign n23141 = ~n22015 & n23140;
  assign n23142 = n23141 ^ n21917;
  assign n23246 = n23245 ^ n23142;
  assign n23132 = n4963 & ~n20908;
  assign n23133 = n4972 & ~n19281;
  assign n23134 = n4976 & n19277;
  assign n23135 = n4970 & n19260;
  assign n23136 = ~n23134 & ~n23135;
  assign n23137 = ~n23133 & n23136;
  assign n23138 = ~n23132 & n23137;
  assign n23139 = n23138 ^ x17;
  assign n23247 = n23246 ^ n23139;
  assign n23129 = n22016 ^ n21906;
  assign n23130 = ~n22017 & n23129;
  assign n23131 = n23130 ^ n21906;
  assign n23248 = n23247 ^ n23131;
  assign n23114 = n13989 & ~n21215;
  assign n23115 = n14928 & ~n19104;
  assign n23116 = ~n7559 & ~n23115;
  assign n23117 = ~n23114 & n23116;
  assign n23118 = n5752 & n19122;
  assign n23119 = ~n5746 & ~n19286;
  assign n23120 = ~n23118 & ~n23119;
  assign n23121 = ~n23117 & n23120;
  assign n23122 = x13 & ~n21215;
  assign n23123 = ~x13 & ~n19104;
  assign n23124 = n6033 & ~n23123;
  assign n23125 = ~n23122 & n23124;
  assign n23126 = ~x14 & ~n23120;
  assign n23127 = ~n23125 & ~n23126;
  assign n23128 = ~n23121 & n23127;
  assign n23249 = n23248 ^ n23128;
  assign n23111 = n22018 ^ n21882;
  assign n23112 = ~n22019 & n23111;
  assign n23113 = n23112 ^ n21882;
  assign n23250 = n23249 ^ n23113;
  assign n23108 = n22031 ^ n22020;
  assign n23109 = n22032 & ~n23108;
  assign n23110 = n23109 ^ n22023;
  assign n23251 = n23250 ^ n23110;
  assign n23092 = n7536 & n19668;
  assign n23093 = n5817 & n19096;
  assign n23094 = n5824 & n19292;
  assign n23095 = ~n23093 & ~n23094;
  assign n23096 = x11 & n23095;
  assign n23097 = ~n19298 & n23096;
  assign n23098 = ~n23092 & ~n23097;
  assign n23099 = x10 & n23098;
  assign n23100 = ~n19668 & n23096;
  assign n23101 = n7536 & n19298;
  assign n23102 = ~x10 & ~n23101;
  assign n23103 = ~n23100 & n23102;
  assign n23104 = ~n23099 & ~n23103;
  assign n23105 = ~n7551 & n23095;
  assign n23106 = n23105 ^ x11;
  assign n23107 = ~n23104 & n23106;
  assign n23252 = n23251 ^ n23107;
  assign n23089 = n22033 ^ n19666;
  assign n23090 = n22034 & ~n23089;
  assign n23091 = n23090 ^ n21879;
  assign n23253 = n23252 ^ n23091;
  assign n23081 = n6306 & n22441;
  assign n23082 = n7168 & n19063;
  assign n23083 = n6316 & ~n19078;
  assign n23084 = n6309 & n19303;
  assign n23085 = ~n23083 & ~n23084;
  assign n23086 = ~n23082 & n23085;
  assign n23087 = ~n23081 & n23086;
  assign n23088 = n23087 ^ x8;
  assign n23254 = n23253 ^ n23088;
  assign n23064 = n22971 ^ n19512;
  assign n23065 = ~x4 & ~n23064;
  assign n23066 = x4 & ~n19512;
  assign n23067 = x5 & ~n23066;
  assign n23068 = ~n23065 & n23067;
  assign n23069 = ~n17410 & ~n23068;
  assign n23070 = n7518 & n19439;
  assign n23071 = n7520 & ~n19368;
  assign n23072 = ~n23070 & ~n23071;
  assign n23073 = ~n23069 & n23072;
  assign n23074 = x4 & n23064;
  assign n23075 = ~x4 & n19512;
  assign n23076 = n17396 & ~n23075;
  assign n23077 = ~n23074 & n23076;
  assign n23078 = ~x5 & ~n23072;
  assign n23079 = ~n23077 & ~n23078;
  assign n23080 = ~n23073 & n23079;
  assign n23255 = n23254 ^ n23080;
  assign n23061 = n22465 ^ n22035;
  assign n23062 = n22466 & ~n23061;
  assign n23063 = n23062 ^ n22455;
  assign n23256 = n23255 ^ n23063;
  assign n23046 = n19632 & ~n19637;
  assign n23047 = n19645 & ~n23046;
  assign n23048 = n19632 & ~n19635;
  assign n23049 = ~n19639 & ~n23048;
  assign n23050 = ~n19633 & n23049;
  assign n23051 = ~n23047 & ~n23050;
  assign n23039 = n19604 & n19614;
  assign n23040 = n19606 & n23039;
  assign n23041 = ~n19604 & ~n19614;
  assign n23042 = ~n19606 & n23041;
  assign n23043 = ~n23040 & ~n23042;
  assign n23038 = n3422 & n3874;
  assign n23044 = n23043 ^ n23038;
  assign n23032 = x31 & ~n13863;
  assign n23033 = n3669 & ~n11902;
  assign n23034 = ~n91 & ~n23033;
  assign n23035 = ~n23032 & n23034;
  assign n23036 = n23035 ^ n19617;
  assign n23029 = n19617 ^ n19615;
  assign n23030 = n19631 & n23029;
  assign n23031 = n23030 ^ n19630;
  assign n23037 = n23036 ^ n23031;
  assign n23045 = n23044 ^ n23037;
  assign n23052 = n23051 ^ n23045;
  assign n23024 = ~n19576 & ~n19649;
  assign n23025 = ~n19598 & n19649;
  assign n23026 = ~n23024 & ~n23025;
  assign n23027 = n33 & ~n23026;
  assign n23028 = n23027 ^ x1;
  assign n23053 = n23052 ^ n23028;
  assign n23054 = x0 & ~n23053;
  assign n23055 = n19649 ^ x2;
  assign n23056 = n9378 & ~n23055;
  assign n23057 = x2 & n19575;
  assign n23058 = n9448 & ~n23057;
  assign n23059 = ~n23056 & ~n23058;
  assign n23060 = ~n23054 & n23059;
  assign n23257 = n23256 ^ n23060;
  assign n23015 = n22988 & ~n22999;
  assign n23016 = n23011 & ~n23015;
  assign n23021 = n23016 ^ n19656;
  assign n23022 = n22468 & n23021;
  assign n23023 = n23022 ^ n22467;
  assign n23258 = n23257 ^ n23023;
  assign n23017 = n22468 & n23016;
  assign n23018 = ~n22468 & ~n23000;
  assign n23019 = ~n23012 & ~n23018;
  assign n23020 = ~n23017 & n23019;
  assign n23259 = n23258 ^ n23020;
  assign n23468 = n22989 ^ n19575;
  assign n23469 = n17396 & ~n23468;
  assign n23470 = n7518 & ~n19512;
  assign n23471 = n7520 & n19439;
  assign n23472 = ~n23470 & ~n23471;
  assign n23473 = x5 & n23472;
  assign n23474 = n19575 & n23473;
  assign n23475 = ~n23469 & ~n23474;
  assign n23476 = x4 & n23475;
  assign n23477 = n23468 & n23473;
  assign n23478 = n17396 & ~n19575;
  assign n23479 = ~x4 & ~n23478;
  assign n23480 = ~n23477 & n23479;
  assign n23481 = ~n23476 & ~n23480;
  assign n23482 = ~n17411 & n23472;
  assign n23483 = n23482 ^ x5;
  assign n23484 = ~n23481 & n23483;
  assign n23465 = n23254 ^ n23063;
  assign n23466 = ~n23255 & n23465;
  assign n23467 = n23466 ^ n23063;
  assign n23485 = n23484 ^ n23467;
  assign n23453 = n5814 & ~n21715;
  assign n23454 = n6295 & ~n19078;
  assign n23455 = n5817 & n19298;
  assign n23456 = n5824 & n19096;
  assign n23457 = ~n23455 & ~n23456;
  assign n23458 = ~n23454 & n23457;
  assign n23459 = ~n23453 & n23458;
  assign n23460 = n23459 ^ x11;
  assign n23450 = n23250 ^ n23107;
  assign n23451 = n23251 & ~n23450;
  assign n23452 = n23451 ^ n23110;
  assign n23461 = n23460 ^ n23452;
  assign n23428 = n21932 & n22012;
  assign n23429 = ~n23230 & n23237;
  assign n23430 = n22001 & ~n23429;
  assign n23431 = ~n23428 & n23430;
  assign n23432 = n23230 & ~n23237;
  assign n23433 = ~x23 & ~n23432;
  assign n23434 = ~n23431 & n23433;
  assign n23435 = ~n21932 & n22012;
  assign n23436 = ~n23230 & ~n23237;
  assign n23437 = n22001 & ~n23436;
  assign n23438 = ~n23435 & n23437;
  assign n23439 = n23230 & n23237;
  assign n23440 = x23 & ~n23439;
  assign n23441 = ~n23438 & n23440;
  assign n23442 = ~n23434 & ~n23441;
  assign n23409 = n12417 & ~n20045;
  assign n23410 = n3435 & ~n19225;
  assign n23411 = ~n3440 & ~n19215;
  assign n23412 = ~n23410 & ~n23411;
  assign n23413 = x26 & n23412;
  assign n23414 = n19142 & n23413;
  assign n23415 = x25 & ~n23414;
  assign n23416 = ~n23409 & n23415;
  assign n23417 = n20045 & n23413;
  assign n23418 = n12417 & ~n19142;
  assign n23419 = ~x25 & ~n23418;
  assign n23420 = ~n23417 & n23419;
  assign n23421 = ~n23416 & ~n23420;
  assign n23422 = ~n12432 & n23412;
  assign n23423 = n23422 ^ x26;
  assign n23424 = ~n23421 & n23423;
  assign n23399 = n44 & n19966;
  assign n23400 = n3280 & n19160;
  assign n23401 = n3277 & n19200;
  assign n23402 = n3275 & ~n19162;
  assign n23403 = ~n23401 & ~n23402;
  assign n23404 = ~n23400 & n23403;
  assign n23405 = ~n23399 & n23404;
  assign n23406 = n23405 ^ x29;
  assign n23396 = n23210 ^ n23161;
  assign n23397 = ~n23211 & n23396;
  assign n23398 = n23397 ^ n23164;
  assign n23407 = n23406 ^ n23398;
  assign n23387 = x31 & n19839;
  assign n23388 = n23387 ^ n19201;
  assign n23389 = n41 & ~n23388;
  assign n23390 = ~n3673 & ~n19161;
  assign n23391 = x31 & n23206;
  assign n23392 = ~n23390 & ~n23391;
  assign n23393 = ~n23389 & n23392;
  assign n23370 = n2060 & n11567;
  assign n23371 = n2392 & n3808;
  assign n23372 = n175 & n437;
  assign n23373 = n23371 & n23372;
  assign n23374 = n2943 & n12864;
  assign n23375 = n1889 & n23374;
  assign n23376 = n23373 & n23375;
  assign n23377 = n23370 & n23376;
  assign n23378 = ~n409 & ~n680;
  assign n23379 = ~n93 & n23378;
  assign n23380 = n267 & n2595;
  assign n23381 = n23379 & n23380;
  assign n23382 = n1715 & n23381;
  assign n23383 = n3556 & n23382;
  assign n23384 = n23377 & n23383;
  assign n23385 = n3581 & n23384;
  assign n23386 = n1797 & n23385;
  assign n23394 = n23393 ^ n23386;
  assign n23367 = n23209 ^ n23167;
  assign n23368 = ~n23185 & ~n23367;
  assign n23369 = n23368 ^ n23209;
  assign n23395 = n23394 ^ n23369;
  assign n23408 = n23407 ^ n23395;
  assign n23425 = n23424 ^ n23408;
  assign n23364 = n23229 ^ n23153;
  assign n23365 = n23213 & n23364;
  assign n23366 = n23365 ^ n23229;
  assign n23426 = n23425 ^ n23366;
  assign n23356 = n4478 & ~n20328;
  assign n23357 = n4487 & ~n19238;
  assign n23358 = n4484 & n19233;
  assign n23359 = n4480 & n19139;
  assign n23360 = ~n23358 & ~n23359;
  assign n23361 = ~n23357 & n23360;
  assign n23362 = ~n23356 & n23361;
  assign n23363 = n23362 ^ x23;
  assign n23427 = n23426 ^ n23363;
  assign n23443 = n23442 ^ n23427;
  assign n23348 = n4673 & n20929;
  assign n23349 = n4688 & n19260;
  assign n23350 = n4685 & ~n19255;
  assign n23351 = ~n4681 & n19253;
  assign n23352 = ~n23350 & ~n23351;
  assign n23353 = ~n23349 & n23352;
  assign n23354 = ~n23348 & n23353;
  assign n23355 = n23354 ^ x20;
  assign n23444 = n23443 ^ n23355;
  assign n23345 = n23244 ^ n23142;
  assign n23346 = ~n23245 & n23345;
  assign n23347 = n23346 ^ n23142;
  assign n23445 = n23444 ^ n23347;
  assign n23337 = n4963 & n21189;
  assign n23338 = n4972 & n19122;
  assign n23339 = n4976 & ~n19281;
  assign n23340 = n4970 & n19277;
  assign n23341 = ~n23339 & ~n23340;
  assign n23342 = ~n23338 & n23341;
  assign n23343 = ~n23337 & n23342;
  assign n23344 = n23343 ^ x17;
  assign n23446 = n23445 ^ n23344;
  assign n23334 = n23246 ^ n23131;
  assign n23335 = ~n23247 & n23334;
  assign n23336 = n23335 ^ n23131;
  assign n23447 = n23446 ^ n23336;
  assign n23318 = n6033 & n21684;
  assign n23319 = ~n5746 & n19104;
  assign n23320 = n5752 & ~n19286;
  assign n23321 = ~n23319 & ~n23320;
  assign n23322 = x14 & n23321;
  assign n23323 = ~n19292 & n23322;
  assign n23324 = ~n23318 & ~n23323;
  assign n23325 = x13 & n23324;
  assign n23326 = ~n21684 & n23322;
  assign n23327 = n6033 & n19292;
  assign n23328 = ~x13 & ~n23327;
  assign n23329 = ~n23326 & n23328;
  assign n23330 = ~n23325 & ~n23329;
  assign n23331 = ~n7589 & n23321;
  assign n23332 = n23331 ^ x14;
  assign n23333 = ~n23330 & n23332;
  assign n23448 = n23447 ^ n23333;
  assign n23315 = n23248 ^ n23113;
  assign n23316 = ~n23249 & n23315;
  assign n23317 = n23316 ^ n23113;
  assign n23449 = n23448 ^ n23317;
  assign n23462 = n23461 ^ n23449;
  assign n23307 = n6306 & ~n22037;
  assign n23308 = n7168 & ~n19368;
  assign n23309 = n6309 & n19063;
  assign n23310 = n6316 & n19303;
  assign n23311 = ~n23309 & ~n23310;
  assign n23312 = ~n23308 & n23311;
  assign n23313 = ~n23307 & n23312;
  assign n23314 = n23313 ^ x8;
  assign n23463 = n23462 ^ n23314;
  assign n23304 = n23252 ^ n23088;
  assign n23305 = n23253 & ~n23304;
  assign n23306 = n23305 ^ n23091;
  assign n23464 = n23463 ^ n23306;
  assign n23486 = n23485 ^ n23464;
  assign n23301 = n23256 ^ n23023;
  assign n23302 = n23257 & n23301;
  assign n23303 = n23302 ^ n23023;
  assign n23487 = n23486 ^ n23303;
  assign n23274 = n23035 ^ n23031;
  assign n23275 = n23051 ^ n23031;
  assign n23276 = n23274 & ~n23275;
  assign n23277 = n23276 ^ n23051;
  assign n23278 = n19617 & ~n23277;
  assign n23279 = n23031 & ~n23035;
  assign n23280 = ~n23051 & n23279;
  assign n23281 = n23044 & ~n23280;
  assign n23282 = n23278 & ~n23281;
  assign n23283 = ~n19617 & n23044;
  assign n23284 = n23277 & n23283;
  assign n23285 = ~n23044 & n23280;
  assign n23286 = ~n23031 & n23035;
  assign n23287 = n23051 & n23286;
  assign n23288 = ~n19617 & n23287;
  assign n23289 = ~n23285 & ~n23288;
  assign n23290 = ~n23284 & n23289;
  assign n23291 = ~n23282 & n23290;
  assign n23267 = n3428 & n23040;
  assign n23268 = ~n3428 & ~n23039;
  assign n23269 = n23038 & ~n23268;
  assign n23270 = ~n23267 & n23269;
  assign n23271 = ~n23038 & ~n23042;
  assign n23272 = ~n23270 & ~n23271;
  assign n23266 = n19617 ^ n12591;
  assign n23273 = n23272 ^ n23266;
  assign n23292 = n23291 ^ n23273;
  assign n23261 = n23025 ^ n23024;
  assign n23262 = ~n23052 & n23261;
  assign n23263 = n23262 ^ n23024;
  assign n23264 = n33 & ~n23263;
  assign n23265 = n23264 ^ x1;
  assign n23293 = n23292 ^ n23265;
  assign n23294 = x0 & ~n23293;
  assign n23295 = n23052 ^ x2;
  assign n23296 = x1 & ~n23295;
  assign n23297 = n9431 & ~n19649;
  assign n23298 = ~n9378 & ~n23297;
  assign n23299 = ~n23296 & ~n23298;
  assign n23300 = ~n23294 & ~n23299;
  assign n23488 = n23487 ^ n23300;
  assign n23260 = n23020 & n23258;
  assign n23489 = n23488 ^ n23260;
  assign n23657 = ~x25 & ~n20030;
  assign n23658 = n19139 & ~n23657;
  assign n23659 = n12417 & n20030;
  assign n23660 = n23658 & ~n23659;
  assign n23661 = n735 & ~n23660;
  assign n23662 = ~n3440 & ~n19225;
  assign n23663 = n3435 & ~n19142;
  assign n23664 = ~n23662 & ~n23663;
  assign n23665 = x26 & n23664;
  assign n23666 = n23665 ^ x25;
  assign n23667 = n20030 & n23666;
  assign n23668 = n23667 ^ x25;
  assign n23669 = ~n19139 & ~n23668;
  assign n23670 = n23661 & ~n23669;
  assign n23671 = ~n12431 & n23664;
  assign n23672 = ~n23670 & n23671;
  assign n23673 = x26 & ~n23664;
  assign n23674 = ~n23672 & ~n23673;
  assign n23648 = n44 & n20020;
  assign n23649 = n3277 & n19160;
  assign n23650 = n3280 & ~n19215;
  assign n23651 = n3275 & n19200;
  assign n23652 = ~n23650 & ~n23651;
  assign n23653 = ~n23649 & n23652;
  assign n23654 = ~n23648 & n23653;
  assign n23655 = n23654 ^ x29;
  assign n23634 = n41 & n19828;
  assign n23635 = n91 & n19201;
  assign n23636 = n54 & n19161;
  assign n23637 = x31 & ~n23636;
  assign n23638 = ~n23635 & n23637;
  assign n23639 = ~n23634 & n23638;
  assign n23640 = ~n54 & n19162;
  assign n23641 = n54 & n19201;
  assign n23642 = n3640 & ~n23641;
  assign n23643 = ~n23640 & n23642;
  assign n23644 = ~n23639 & ~n23643;
  assign n23620 = ~n319 & n3510;
  assign n23621 = n11170 & n23620;
  assign n23622 = n2036 & n2137;
  assign n23623 = n23621 & n23622;
  assign n23624 = n302 & n2975;
  assign n23625 = n949 & n23624;
  assign n23626 = n23623 & n23625;
  assign n23627 = n766 & n4411;
  assign n23628 = n4761 & n23627;
  assign n23629 = n13190 & n23628;
  assign n23630 = n23626 & n23629;
  assign n23631 = n1437 & n23630;
  assign n23632 = n5681 & n23631;
  assign n23633 = n5608 & n23632;
  assign n23645 = n23644 ^ n23633;
  assign n23617 = n23393 ^ n23369;
  assign n23618 = ~n23394 & ~n23617;
  assign n23619 = n23618 ^ n23369;
  assign n23646 = n23645 ^ n23619;
  assign n23614 = n23398 ^ n23395;
  assign n23615 = n23407 & n23614;
  assign n23616 = n23615 ^ n23406;
  assign n23647 = n23646 ^ n23616;
  assign n23656 = n23655 ^ n23647;
  assign n23675 = n23674 ^ n23656;
  assign n23611 = n23424 ^ n23366;
  assign n23612 = n23425 & n23611;
  assign n23613 = n23612 ^ n23366;
  assign n23676 = n23675 ^ n23613;
  assign n23603 = n4478 & n20308;
  assign n23604 = n4487 & n19253;
  assign n23605 = n4484 & ~n19238;
  assign n23606 = n4480 & n19233;
  assign n23607 = ~n23605 & ~n23606;
  assign n23608 = ~n23604 & n23607;
  assign n23609 = ~n23603 & n23608;
  assign n23610 = n23609 ^ x23;
  assign n23677 = n23676 ^ n23610;
  assign n23600 = n23442 ^ n23426;
  assign n23601 = n23427 & n23600;
  assign n23602 = n23601 ^ n23442;
  assign n23678 = n23677 ^ n23602;
  assign n23592 = n4673 & n20793;
  assign n23593 = n4688 & n19277;
  assign n23594 = n4685 & n19260;
  assign n23595 = ~n4681 & ~n19255;
  assign n23596 = ~n23594 & ~n23595;
  assign n23597 = ~n23593 & n23596;
  assign n23598 = ~n23592 & n23597;
  assign n23599 = n23598 ^ x20;
  assign n23679 = n23678 ^ n23599;
  assign n23589 = n23443 ^ n23347;
  assign n23590 = ~n23444 & n23589;
  assign n23591 = n23590 ^ n23347;
  assign n23680 = n23679 ^ n23591;
  assign n23581 = n4963 & ~n19678;
  assign n23582 = n4976 & n19122;
  assign n23583 = n4972 & ~n19286;
  assign n23584 = n4970 & ~n19281;
  assign n23585 = ~n23583 & ~n23584;
  assign n23586 = ~n23582 & n23585;
  assign n23587 = ~n23581 & n23586;
  assign n23588 = n23587 ^ x17;
  assign n23681 = n23680 ^ n23588;
  assign n23578 = n23445 ^ n23336;
  assign n23579 = ~n23446 & n23578;
  assign n23580 = n23579 ^ n23336;
  assign n23682 = n23681 ^ n23580;
  assign n23564 = x13 & n21698;
  assign n23565 = ~n6033 & ~n21698;
  assign n23566 = ~n23564 & ~n23565;
  assign n23562 = n5749 & ~n21698;
  assign n23563 = n23562 ^ x13;
  assign n23567 = n23566 ^ n23563;
  assign n23568 = n19096 & n23567;
  assign n23569 = n23568 ^ n23563;
  assign n23570 = n5748 & ~n23569;
  assign n23571 = ~n5746 & n19292;
  assign n23572 = n5752 & n19104;
  assign n23573 = ~n23571 & ~n23572;
  assign n23574 = ~n6048 & n23573;
  assign n23575 = ~n23570 & n23574;
  assign n23576 = ~x14 & ~n23573;
  assign n23577 = ~n23575 & ~n23576;
  assign n23683 = n23682 ^ n23577;
  assign n23559 = n23447 ^ n23317;
  assign n23560 = ~n23448 & n23559;
  assign n23561 = n23560 ^ n23317;
  assign n23684 = n23683 ^ n23561;
  assign n23556 = n23460 ^ n23449;
  assign n23557 = n23461 & ~n23556;
  assign n23558 = n23557 ^ n23452;
  assign n23685 = n23684 ^ n23558;
  assign n23548 = n5814 & n19658;
  assign n23549 = n5817 & ~n19078;
  assign n23550 = n6295 & n19303;
  assign n23551 = n5824 & n19298;
  assign n23552 = ~n23550 & ~n23551;
  assign n23553 = ~n23549 & n23552;
  assign n23554 = ~n23548 & n23553;
  assign n23555 = n23554 ^ x11;
  assign n23686 = n23685 ^ n23555;
  assign n23545 = n23462 ^ n23306;
  assign n23546 = ~n23463 & n23545;
  assign n23547 = n23546 ^ n23306;
  assign n23687 = n23686 ^ n23547;
  assign n23537 = n6306 & n22457;
  assign n23538 = n7168 & n19439;
  assign n23539 = n6309 & ~n19368;
  assign n23540 = n6316 & n19063;
  assign n23541 = ~n23539 & ~n23540;
  assign n23542 = ~n23538 & n23541;
  assign n23543 = ~n23537 & n23542;
  assign n23544 = n23543 ^ x8;
  assign n23688 = n23687 ^ n23544;
  assign n23520 = n19649 ^ n19599;
  assign n23521 = n17396 & n23520;
  assign n23522 = n7520 & ~n19512;
  assign n23523 = n7518 & ~n19575;
  assign n23524 = ~n23522 & ~n23523;
  assign n23525 = x5 & n23524;
  assign n23526 = ~n19649 & n23525;
  assign n23527 = x4 & ~n23526;
  assign n23528 = ~n23521 & n23527;
  assign n23529 = ~n23520 & n23525;
  assign n23530 = n17396 & n19649;
  assign n23531 = ~x4 & ~n23530;
  assign n23532 = ~n23529 & n23531;
  assign n23533 = ~n23528 & ~n23532;
  assign n23534 = ~n17411 & n23524;
  assign n23535 = n23534 ^ x5;
  assign n23536 = ~n23533 & n23535;
  assign n23689 = n23688 ^ n23536;
  assign n23517 = n23484 ^ n23464;
  assign n23518 = n23485 & ~n23517;
  assign n23519 = n23518 ^ n23467;
  assign n23690 = n23689 ^ n23519;
  assign n23514 = n23486 ^ n23300;
  assign n23515 = n23487 & ~n23514;
  assign n23516 = n23515 ^ n23303;
  assign n23691 = n23690 ^ n23516;
  assign n23512 = n23260 & ~n23488;
  assign n23490 = ~n23025 & ~n23052;
  assign n23491 = ~n23292 & ~n23490;
  assign n23492 = n23024 & n23052;
  assign n23493 = ~n23491 & ~n23492;
  assign n23494 = ~x2 & n23493;
  assign n23495 = ~n23052 & n23292;
  assign n23496 = x2 & ~n23495;
  assign n23497 = x0 & ~n23496;
  assign n23498 = ~n23494 & n23497;
  assign n23499 = n9431 & ~n23292;
  assign n23500 = ~n23498 & ~n23499;
  assign n23501 = x1 & ~n23500;
  assign n23502 = ~x1 & ~n23495;
  assign n23503 = ~x0 & n23292;
  assign n23504 = ~n23502 & ~n23503;
  assign n23505 = ~x2 & ~n23504;
  assign n23506 = ~x1 & n8890;
  assign n23507 = n23493 & n23506;
  assign n23508 = n9448 & n23052;
  assign n23509 = ~n23507 & ~n23508;
  assign n23510 = ~n23505 & n23509;
  assign n23511 = ~n23501 & n23510;
  assign n23513 = n23512 ^ n23511;
  assign n23692 = n23691 ^ n23513;
  assign n23841 = n3285 & n20294;
  assign n23842 = n3437 & n19233;
  assign n23843 = n3435 & n19139;
  assign n23844 = ~n3440 & ~n19142;
  assign n23845 = ~n23843 & ~n23844;
  assign n23846 = ~n23842 & n23845;
  assign n23847 = ~n23841 & n23846;
  assign n23848 = n23847 ^ x26;
  assign n23831 = n44 & ~n20210;
  assign n23832 = n3280 & ~n19225;
  assign n23833 = n3275 & n19160;
  assign n23834 = n3277 & ~n19215;
  assign n23835 = ~n23833 & ~n23834;
  assign n23836 = ~n23832 & n23835;
  assign n23837 = ~n23831 & n23836;
  assign n23838 = n23837 ^ x29;
  assign n23828 = n23655 ^ n23616;
  assign n23829 = n23647 & n23828;
  assign n23830 = n23829 ^ n23655;
  assign n23839 = n23838 ^ n23830;
  assign n23816 = n41 & ~n19816;
  assign n23817 = n91 & n19162;
  assign n23818 = x31 & ~n23641;
  assign n23819 = ~n23817 & n23818;
  assign n23820 = ~n23816 & n23819;
  assign n23821 = ~n54 & ~n19200;
  assign n23822 = n54 & n19162;
  assign n23823 = n3640 & ~n23822;
  assign n23824 = ~n23821 & n23823;
  assign n23825 = ~n23820 & ~n23824;
  assign n23793 = n4273 & ~n13178;
  assign n23794 = n2615 & n23793;
  assign n23795 = n1295 & n1567;
  assign n23796 = n118 & n3087;
  assign n23797 = n23795 & n23796;
  assign n23798 = n23794 & n23797;
  assign n23799 = n1733 & n23798;
  assign n23800 = ~n517 & ~n560;
  assign n23801 = n2654 & n23800;
  assign n23802 = n5090 & n23801;
  assign n23803 = n2444 & n11141;
  assign n23804 = n23802 & n23803;
  assign n23805 = n23799 & n23804;
  assign n23806 = ~n293 & ~n409;
  assign n23807 = ~n567 & ~n592;
  assign n23808 = n23806 & n23807;
  assign n23809 = n1158 & n23808;
  assign n23810 = n3537 & n13380;
  assign n23811 = n23809 & n23810;
  assign n23812 = n23176 & n23811;
  assign n23813 = n23805 & n23812;
  assign n23814 = n3503 & n23813;
  assign n23815 = n4587 & n23814;
  assign n23826 = n23825 ^ n23815;
  assign n23790 = n23644 ^ n23619;
  assign n23791 = ~n23645 & ~n23790;
  assign n23792 = n23791 ^ n23619;
  assign n23827 = n23826 ^ n23792;
  assign n23840 = n23839 ^ n23827;
  assign n23849 = n23848 ^ n23840;
  assign n23787 = n23656 ^ n23613;
  assign n23788 = n23675 & n23787;
  assign n23789 = n23788 ^ n23674;
  assign n23850 = n23849 ^ n23789;
  assign n23779 = n4478 & ~n19696;
  assign n23780 = n4487 & ~n19255;
  assign n23781 = n4484 & n19253;
  assign n23782 = n4480 & ~n19238;
  assign n23783 = ~n23781 & ~n23782;
  assign n23784 = ~n23780 & n23783;
  assign n23785 = ~n23779 & n23784;
  assign n23786 = n23785 ^ x23;
  assign n23851 = n23850 ^ n23786;
  assign n23776 = n23676 ^ n23602;
  assign n23777 = ~n23677 & ~n23776;
  assign n23778 = n23777 ^ n23602;
  assign n23852 = n23851 ^ n23778;
  assign n23773 = n23678 ^ n23591;
  assign n23774 = n23679 & ~n23773;
  assign n23775 = n23774 ^ n23591;
  assign n23853 = n23852 ^ n23775;
  assign n23765 = n4673 & ~n20908;
  assign n23766 = n4688 & ~n19281;
  assign n23767 = n4685 & n19277;
  assign n23768 = ~n4681 & n19260;
  assign n23769 = ~n23767 & ~n23768;
  assign n23770 = ~n23766 & n23769;
  assign n23771 = ~n23765 & n23770;
  assign n23772 = n23771 ^ x20;
  assign n23854 = n23853 ^ n23772;
  assign n23757 = n4963 & n21215;
  assign n23758 = n4972 & n19104;
  assign n23759 = n4970 & n19122;
  assign n23760 = n4976 & ~n19286;
  assign n23761 = ~n23759 & ~n23760;
  assign n23762 = ~n23758 & n23761;
  assign n23763 = ~n23757 & n23762;
  assign n23764 = n23763 ^ x17;
  assign n23855 = n23854 ^ n23764;
  assign n23754 = n23680 ^ n23580;
  assign n23755 = n23681 & ~n23754;
  assign n23756 = n23755 ^ n23580;
  assign n23856 = n23855 ^ n23756;
  assign n23746 = n5749 & n19667;
  assign n23747 = n23746 ^ n19298;
  assign n23748 = n5748 & n23747;
  assign n23749 = ~n5746 & n19096;
  assign n23750 = n5752 & n19292;
  assign n23751 = ~n23749 & ~n23750;
  assign n23752 = ~n23748 & n23751;
  assign n23753 = n23752 ^ x14;
  assign n23857 = n23856 ^ n23753;
  assign n23743 = n23682 ^ n23561;
  assign n23744 = n23683 & ~n23743;
  assign n23745 = n23744 ^ n23561;
  assign n23858 = n23857 ^ n23745;
  assign n23740 = n23684 ^ n23555;
  assign n23741 = ~n23685 & n23740;
  assign n23742 = n23741 ^ n23558;
  assign n23859 = n23858 ^ n23742;
  assign n23732 = n5814 & n22441;
  assign n23733 = n6295 & n19063;
  assign n23734 = n5824 & ~n19078;
  assign n23735 = n5817 & n19303;
  assign n23736 = ~n23734 & ~n23735;
  assign n23737 = ~n23733 & n23736;
  assign n23738 = ~n23732 & n23737;
  assign n23739 = n23738 ^ x11;
  assign n23860 = n23859 ^ n23739;
  assign n23725 = n6306 & ~n23064;
  assign n23726 = n7168 & ~n19512;
  assign n23727 = n6309 & n19439;
  assign n23728 = n6316 & ~n19368;
  assign n23729 = ~n23727 & ~n23728;
  assign n23730 = ~n23726 & n23729;
  assign n23731 = ~n23725 & n23730;
  assign n23861 = n23860 ^ n23731;
  assign n23721 = n23686 ^ x8;
  assign n23722 = n23721 ^ n23543;
  assign n23723 = n23687 & ~n23722;
  assign n23724 = n23723 ^ n23543;
  assign n23862 = n23861 ^ n23724;
  assign n23712 = n23052 ^ n23026;
  assign n23713 = n7515 & n23712;
  assign n23714 = n7518 & n19649;
  assign n23715 = n7520 & ~n19575;
  assign n23716 = ~n23714 & ~n23715;
  assign n23717 = n8029 & n23052;
  assign n23718 = n23716 & ~n23717;
  assign n23719 = ~n23713 & n23718;
  assign n23720 = n23719 ^ x5;
  assign n23863 = n23862 ^ n23720;
  assign n23709 = n23688 ^ n23519;
  assign n23710 = n23689 & ~n23709;
  assign n23711 = n23710 ^ n23519;
  assign n23864 = n23863 ^ n23711;
  assign n23698 = ~x2 & n23052;
  assign n23699 = n33 & n23698;
  assign n23700 = n23699 ^ n33;
  assign n23701 = n23503 & n23700;
  assign n23702 = n8886 & ~n23495;
  assign n23703 = ~n23701 & ~n23702;
  assign n23704 = ~n23491 & ~n23495;
  assign n23705 = n8890 & n23704;
  assign n23706 = n23703 & ~n23705;
  assign n23707 = n8883 & ~n23704;
  assign n23708 = n23706 & ~n23707;
  assign n23865 = n23864 ^ n23708;
  assign n23693 = n23690 ^ n23512;
  assign n23695 = n23693 ^ n23511;
  assign n23696 = n23516 & n23695;
  assign n23694 = ~n23513 & ~n23693;
  assign n23697 = n23696 ^ n23694;
  assign n23866 = n23865 ^ n23697;
  assign n23871 = ~n23516 & n23690;
  assign n24043 = ~n23511 & ~n23871;
  assign n23869 = n23516 & ~n23690;
  assign n24044 = n23708 & ~n23864;
  assign n24045 = ~n23869 & ~n24044;
  assign n24046 = ~n24043 & n24045;
  assign n24047 = ~n23708 & n23864;
  assign n24048 = ~n24046 & ~n24047;
  assign n24041 = n9448 & n23495;
  assign n24042 = x2 & ~n24041;
  assign n24049 = n24048 ^ n24042;
  assign n24025 = n23547 & ~n23686;
  assign n24026 = n23731 ^ n23543;
  assign n24027 = ~n23860 & n24026;
  assign n24028 = ~n23544 & n24027;
  assign n24029 = n24028 ^ n23544;
  assign n24030 = ~n24025 & ~n24029;
  assign n24031 = ~n23547 & n23686;
  assign n24032 = n24031 ^ n23860;
  assign n24033 = n23731 ^ x8;
  assign n24034 = n24033 ^ n23860;
  assign n24035 = n24032 & n24034;
  assign n24036 = n24035 ^ n24031;
  assign n24037 = ~n24030 & ~n24036;
  assign n24014 = n5813 & n22036;
  assign n24015 = n24014 ^ n19368;
  assign n24016 = n5812 & ~n24015;
  assign n24017 = n5817 & n19063;
  assign n24018 = n5824 & n19303;
  assign n24019 = ~n24017 & ~n24018;
  assign n24020 = ~n24016 & n24019;
  assign n24021 = n24020 ^ x11;
  assign n24011 = n23858 ^ n23739;
  assign n24012 = ~n23859 & n24011;
  assign n24013 = n24012 ^ n23742;
  assign n24022 = n24021 ^ n24013;
  assign n23993 = n3285 & ~n20328;
  assign n23994 = n3437 & ~n19238;
  assign n23995 = n3435 & n19233;
  assign n23996 = ~n3440 & n19139;
  assign n23997 = ~n23995 & ~n23996;
  assign n23998 = ~n23994 & n23997;
  assign n23999 = ~n23993 & n23998;
  assign n24000 = n23999 ^ x26;
  assign n23983 = n44 & ~n20045;
  assign n23984 = n3280 & ~n19142;
  assign n23985 = n3275 & ~n19215;
  assign n23986 = ~n23984 & ~n23985;
  assign n23987 = n3277 & ~n19225;
  assign n23988 = n23986 & ~n23987;
  assign n23989 = ~n23983 & n23988;
  assign n23990 = n23989 ^ x29;
  assign n23971 = n41 & ~n19966;
  assign n23972 = n91 & ~n19200;
  assign n23973 = x31 & ~n23822;
  assign n23974 = ~n23972 & n23973;
  assign n23975 = ~n23971 & n23974;
  assign n23976 = ~n54 & ~n19160;
  assign n23977 = n54 & ~n19200;
  assign n23978 = n3640 & ~n23977;
  assign n23979 = ~n23976 & n23978;
  assign n23980 = ~n23975 & ~n23979;
  assign n23957 = n332 & n355;
  assign n23958 = ~n270 & ~n323;
  assign n23959 = ~n527 & n23958;
  assign n23960 = n23957 & n23959;
  assign n23961 = n2233 & n2625;
  assign n23962 = n23960 & n23961;
  assign n23963 = n961 & n2190;
  assign n23964 = n4554 & n23963;
  assign n23965 = n3049 & n23964;
  assign n23966 = n23962 & n23965;
  assign n23967 = n3803 & n3924;
  assign n23968 = n23966 & n23967;
  assign n23969 = n13426 & n23968;
  assign n23970 = n4247 & n23969;
  assign n23981 = n23980 ^ n23970;
  assign n23954 = n23825 ^ n23792;
  assign n23955 = ~n23826 & ~n23954;
  assign n23956 = n23955 ^ n23792;
  assign n23982 = n23981 ^ n23956;
  assign n23991 = n23990 ^ n23982;
  assign n23951 = n23838 ^ n23827;
  assign n23952 = n23839 & n23951;
  assign n23953 = n23952 ^ n23830;
  assign n23992 = n23991 ^ n23953;
  assign n24001 = n24000 ^ n23992;
  assign n23948 = n23848 ^ n23789;
  assign n23949 = n23849 & ~n23948;
  assign n23950 = n23949 ^ n23789;
  assign n24002 = n24001 ^ n23950;
  assign n23940 = n4478 & n20929;
  assign n23941 = n4487 & n19260;
  assign n23942 = n4484 & ~n19255;
  assign n23943 = n4480 & n19253;
  assign n23944 = ~n23942 & ~n23943;
  assign n23945 = ~n23941 & n23944;
  assign n23946 = ~n23940 & n23945;
  assign n23947 = n23946 ^ x23;
  assign n24003 = n24002 ^ n23947;
  assign n23937 = n23850 ^ n23778;
  assign n23938 = ~n23851 & ~n23937;
  assign n23939 = n23938 ^ n23778;
  assign n24004 = n24003 ^ n23939;
  assign n23934 = n23852 ^ n23772;
  assign n23935 = ~n23853 & n23934;
  assign n23936 = n23935 ^ n23775;
  assign n24005 = n24004 ^ n23936;
  assign n23926 = n4673 & n21189;
  assign n23927 = n4688 & n19122;
  assign n23928 = n4685 & ~n19281;
  assign n23929 = ~n4681 & n19277;
  assign n23930 = ~n23928 & ~n23929;
  assign n23931 = ~n23927 & n23930;
  assign n23932 = ~n23926 & n23931;
  assign n23933 = n23932 ^ x20;
  assign n24006 = n24005 ^ n23933;
  assign n23918 = n4963 & n21684;
  assign n23919 = n4972 & n19292;
  assign n23920 = n4976 & n19104;
  assign n23921 = n4970 & ~n19286;
  assign n23922 = ~n23920 & ~n23921;
  assign n23923 = ~n23919 & n23922;
  assign n23924 = ~n23918 & n23923;
  assign n23925 = n23924 ^ x17;
  assign n24007 = n24006 ^ n23925;
  assign n23915 = n23854 ^ n23756;
  assign n23916 = n23855 & ~n23915;
  assign n23917 = n23916 ^ n23756;
  assign n24008 = n24007 ^ n23917;
  assign n23909 = n5749 & ~n21714;
  assign n23910 = n23909 ^ x13;
  assign n23911 = n23910 ^ n19078;
  assign n23902 = x13 & n19298;
  assign n23903 = n13989 & n19096;
  assign n23904 = ~n23902 & ~n23903;
  assign n23899 = n13719 & n19096;
  assign n23900 = ~x13 & n19298;
  assign n23901 = ~n23899 & ~n23900;
  assign n23905 = n23904 ^ n23901;
  assign n23906 = x12 & n23905;
  assign n23907 = n23906 ^ n23904;
  assign n23908 = n23907 ^ x14;
  assign n23912 = n23911 ^ n23908;
  assign n23913 = ~n5748 & n23912;
  assign n23914 = n23913 ^ n23911;
  assign n24009 = n24008 ^ n23914;
  assign n23896 = n23856 ^ n23745;
  assign n23897 = n23857 & ~n23896;
  assign n23898 = n23897 ^ n23745;
  assign n24010 = n24009 ^ n23898;
  assign n24023 = n24022 ^ n24010;
  assign n23888 = n6306 & ~n23468;
  assign n23889 = n6309 & ~n19512;
  assign n23890 = n6316 & n19439;
  assign n23891 = ~n23889 & ~n23890;
  assign n23892 = n7168 & ~n19575;
  assign n23893 = n23891 & ~n23892;
  assign n23894 = ~n23888 & n23893;
  assign n23895 = n23894 ^ x8;
  assign n24024 = n24023 ^ n23895;
  assign n24038 = n24037 ^ n24024;
  assign n23879 = n23292 ^ n23263;
  assign n23880 = n7515 & ~n23879;
  assign n23881 = n8029 & ~n23292;
  assign n23882 = n7518 & n23052;
  assign n23883 = n7520 & n19649;
  assign n23884 = ~n23882 & ~n23883;
  assign n23885 = ~n23881 & n23884;
  assign n23886 = ~n23880 & n23885;
  assign n23887 = n23886 ^ x5;
  assign n24039 = n24038 ^ n23887;
  assign n23876 = n23862 ^ n23711;
  assign n23877 = n23863 & ~n23876;
  assign n23878 = n23877 ^ n23711;
  assign n24040 = n24039 ^ n23878;
  assign n24050 = n24049 ^ n24040;
  assign n23867 = ~n23511 & n23691;
  assign n23868 = n23512 & ~n23867;
  assign n23870 = n23511 & ~n23869;
  assign n23872 = n23871 ^ n23870;
  assign n23873 = ~n23865 & ~n23872;
  assign n23874 = n23873 ^ n23871;
  assign n23875 = n23868 & n23874;
  assign n24051 = n24050 ^ n23875;
  assign n24223 = ~n23887 & n24038;
  assign n24224 = n23878 & ~n24223;
  assign n24225 = n23887 & ~n24038;
  assign n24226 = ~n24224 & ~n24225;
  assign n24200 = n3285 & n20308;
  assign n24201 = n3437 & n19253;
  assign n24202 = n3435 & ~n19238;
  assign n24203 = ~n3440 & n19233;
  assign n24204 = ~n24202 & ~n24203;
  assign n24205 = ~n24201 & n24204;
  assign n24206 = ~n24200 & n24205;
  assign n24207 = n24206 ^ x26;
  assign n24190 = n44 & ~n20031;
  assign n24191 = n3280 & n19139;
  assign n24192 = n3277 & ~n19142;
  assign n24193 = n3275 & ~n19225;
  assign n24194 = ~n24192 & ~n24193;
  assign n24195 = ~n24191 & n24194;
  assign n24196 = ~n24190 & n24195;
  assign n24197 = n24196 ^ x29;
  assign n24168 = n4047 & n12722;
  assign n24169 = n848 & n24168;
  assign n24170 = n1756 & n12893;
  assign n24171 = n551 & n2112;
  assign n24172 = n24170 & n24171;
  assign n24173 = n12232 & n24172;
  assign n24174 = n23625 & n24173;
  assign n24175 = n1210 & n2817;
  assign n24176 = n1530 & n24175;
  assign n24177 = ~n319 & ~n361;
  assign n24178 = n4095 & n24177;
  assign n24179 = n24176 & n24178;
  assign n24180 = n10221 & n21946;
  assign n24181 = ~n126 & ~n163;
  assign n24182 = n2842 & n24181;
  assign n24183 = n2655 & n24182;
  assign n24184 = n24180 & n24183;
  assign n24185 = n24179 & n24184;
  assign n24186 = n24174 & n24185;
  assign n24187 = n24169 & n24186;
  assign n24161 = n41 & ~n20020;
  assign n24162 = n91 & ~n19160;
  assign n24163 = ~n23977 & ~n24162;
  assign n24164 = ~n24161 & n24163;
  assign n24158 = n54 & n19160;
  assign n24159 = n41 & ~n19215;
  assign n24160 = ~n24158 & ~n24159;
  assign n24165 = n24164 ^ n24160;
  assign n24166 = ~x31 & ~n24165;
  assign n24167 = n24166 ^ n24164;
  assign n24188 = n24187 ^ n24167;
  assign n24155 = n23980 ^ n23956;
  assign n24156 = ~n23981 & ~n24155;
  assign n24157 = n24156 ^ n23956;
  assign n24189 = n24188 ^ n24157;
  assign n24198 = n24197 ^ n24189;
  assign n24152 = n23990 ^ n23953;
  assign n24153 = n23991 & n24152;
  assign n24154 = n24153 ^ n23953;
  assign n24199 = n24198 ^ n24154;
  assign n24208 = n24207 ^ n24199;
  assign n24149 = n24000 ^ n23950;
  assign n24150 = n24001 & ~n24149;
  assign n24151 = n24150 ^ n23950;
  assign n24209 = n24208 ^ n24151;
  assign n24133 = n12502 & n20793;
  assign n24134 = n4484 & n19260;
  assign n24135 = n4480 & ~n19255;
  assign n24136 = ~n24134 & ~n24135;
  assign n24137 = x23 & n24136;
  assign n24138 = ~n19277 & n24137;
  assign n24139 = x22 & ~n24138;
  assign n24140 = ~n24133 & n24139;
  assign n24141 = ~n20793 & n24137;
  assign n24142 = n12502 & n19277;
  assign n24143 = ~x22 & ~n24142;
  assign n24144 = ~n24141 & n24143;
  assign n24145 = ~n24140 & ~n24144;
  assign n24146 = ~n12519 & n24136;
  assign n24147 = n24146 ^ x23;
  assign n24148 = ~n24145 & n24147;
  assign n24210 = n24209 ^ n24148;
  assign n24130 = n24002 ^ n23939;
  assign n24131 = ~n24003 & ~n24130;
  assign n24132 = n24131 ^ n23939;
  assign n24211 = n24210 ^ n24132;
  assign n24123 = n4673 & ~n19678;
  assign n24124 = n4685 & n19122;
  assign n24125 = n4688 & ~n19286;
  assign n24126 = ~n4681 & ~n19281;
  assign n24127 = ~n24125 & ~n24126;
  assign n24128 = ~n24124 & n24127;
  assign n24129 = ~n24123 & n24128;
  assign n24212 = n24211 ^ n24129;
  assign n24119 = n24004 ^ x20;
  assign n24120 = n24119 ^ n23932;
  assign n24121 = n24005 & ~n24120;
  assign n24122 = n24121 ^ n23932;
  assign n24213 = n24212 ^ n24122;
  assign n24111 = n4963 & n21699;
  assign n24112 = n4972 & n19096;
  assign n24113 = n4976 & n19292;
  assign n24114 = n4970 & n19104;
  assign n24115 = ~n24113 & ~n24114;
  assign n24116 = ~n24112 & n24115;
  assign n24117 = ~n24111 & n24116;
  assign n24118 = n24117 ^ x17;
  assign n24214 = n24213 ^ n24118;
  assign n24108 = n24006 ^ n23917;
  assign n24109 = n24007 & ~n24108;
  assign n24110 = n24109 ^ n23917;
  assign n24215 = n24214 ^ n24110;
  assign n24102 = n5749 & ~n19657;
  assign n24103 = n24102 ^ x13;
  assign n24104 = n24103 ^ n19303;
  assign n24092 = ~x13 & ~n19078;
  assign n24093 = ~x14 & n23902;
  assign n24094 = x12 & ~n24093;
  assign n24095 = ~n24092 & n24094;
  assign n24096 = x13 & ~n19078;
  assign n24097 = n13989 & n19298;
  assign n24098 = ~x12 & ~n24097;
  assign n24099 = ~n24096 & n24098;
  assign n24100 = ~n24095 & ~n24099;
  assign n24101 = n24100 ^ x14;
  assign n24105 = n24104 ^ n24101;
  assign n24106 = ~n5748 & n24105;
  assign n24107 = n24106 ^ n24104;
  assign n24216 = n24215 ^ n24107;
  assign n24089 = n24008 ^ n23898;
  assign n24090 = n24009 & ~n24089;
  assign n24091 = n24090 ^ n23898;
  assign n24217 = n24216 ^ n24091;
  assign n24081 = n5814 & n22457;
  assign n24082 = n6295 & n19439;
  assign n24083 = n5817 & ~n19368;
  assign n24084 = n5824 & n19063;
  assign n24085 = ~n24083 & ~n24084;
  assign n24086 = ~n24082 & n24085;
  assign n24087 = ~n24081 & n24086;
  assign n24088 = n24087 ^ x11;
  assign n24218 = n24217 ^ n24088;
  assign n24078 = n24021 ^ n24010;
  assign n24079 = n24022 & n24078;
  assign n24080 = n24079 ^ n24013;
  assign n24219 = n24218 ^ n24080;
  assign n24075 = n24037 ^ n24023;
  assign n24076 = n24024 & ~n24075;
  assign n24077 = n24076 ^ n24037;
  assign n24220 = n24219 ^ n24077;
  assign n24067 = n6306 & n23520;
  assign n24068 = n7168 & n19649;
  assign n24069 = n6316 & ~n19512;
  assign n24070 = n6309 & ~n19575;
  assign n24071 = ~n24069 & ~n24070;
  assign n24072 = ~n24068 & n24071;
  assign n24073 = ~n24067 & n24072;
  assign n24074 = n24073 ^ x8;
  assign n24221 = n24220 ^ n24074;
  assign n24059 = n7515 & n23493;
  assign n24060 = n8029 & n23495;
  assign n24061 = n7518 & ~n23292;
  assign n24062 = n7520 & n23052;
  assign n24063 = ~n24061 & ~n24062;
  assign n24064 = ~n24060 & n24063;
  assign n24065 = ~n24059 & n24064;
  assign n24066 = n24065 ^ n4518;
  assign n24222 = n24221 ^ n24066;
  assign n24227 = n24226 ^ n24222;
  assign n24052 = ~n24042 & n24048;
  assign n24053 = n24052 ^ n23875;
  assign n24054 = n24042 & ~n24048;
  assign n24055 = ~n24040 & ~n24054;
  assign n24056 = n24055 ^ n24052;
  assign n24057 = ~n24053 & ~n24056;
  assign n24058 = n24057 ^ n23875;
  assign n24228 = n24227 ^ n24058;
  assign n24411 = n24038 ^ n23878;
  assign n24412 = n24222 ^ n23887;
  assign n24413 = n24039 & n24412;
  assign n24414 = n24411 & n24413;
  assign n24415 = n24414 ^ n24222;
  assign n24416 = ~n24052 & ~n24415;
  assign n24417 = n24226 ^ n24054;
  assign n24418 = n24227 & n24417;
  assign n24419 = n24418 ^ n24054;
  assign n24420 = ~n24416 & ~n24419;
  assign n24396 = n5814 & ~n23064;
  assign n24397 = n6295 & ~n19512;
  assign n24398 = n5817 & n19439;
  assign n24399 = n5824 & ~n19368;
  assign n24400 = ~n24398 & ~n24399;
  assign n24401 = ~n24397 & n24400;
  assign n24402 = ~n24396 & n24401;
  assign n24403 = n24402 ^ x11;
  assign n24378 = n6033 & n22441;
  assign n24379 = n5752 & ~n19078;
  assign n24380 = ~n5746 & n19303;
  assign n24381 = ~n24379 & ~n24380;
  assign n24382 = x14 & n24381;
  assign n24383 = ~n19063 & n24382;
  assign n24384 = x13 & ~n24383;
  assign n24385 = ~n24378 & n24384;
  assign n24386 = ~n22441 & n24382;
  assign n24387 = n6033 & n19063;
  assign n24388 = ~x13 & ~n24387;
  assign n24389 = ~n24386 & n24388;
  assign n24390 = ~n24385 & ~n24389;
  assign n24391 = ~n7589 & n24381;
  assign n24392 = n24391 ^ x14;
  assign n24393 = ~n24390 & n24392;
  assign n24363 = n23936 & ~n24004;
  assign n24364 = n24129 ^ n23932;
  assign n24365 = n24211 & n24364;
  assign n24366 = ~n23933 & n24365;
  assign n24367 = n24366 ^ n23933;
  assign n24368 = ~n24363 & ~n24367;
  assign n24369 = ~n23936 & n24004;
  assign n24370 = n24369 ^ n24211;
  assign n24371 = n24129 ^ x20;
  assign n24372 = n24371 ^ n24211;
  assign n24373 = ~n24370 & ~n24372;
  assign n24374 = n24373 ^ n24369;
  assign n24375 = ~n24368 & ~n24374;
  assign n24344 = ~x22 & ~n20908;
  assign n24345 = x22 & ~n19281;
  assign n24346 = x23 & ~n24345;
  assign n24347 = ~n24344 & n24346;
  assign n24348 = ~n12518 & ~n24347;
  assign n24349 = n4484 & n19277;
  assign n24350 = n4480 & n19260;
  assign n24351 = ~n24349 & ~n24350;
  assign n24352 = ~n24348 & n24351;
  assign n24353 = n14738 & ~n20908;
  assign n24354 = n14740 & ~n19281;
  assign n24355 = n24351 & ~n24354;
  assign n24356 = ~n24353 & n24355;
  assign n24357 = ~x23 & ~n24356;
  assign n24358 = ~n24352 & ~n24357;
  assign n24341 = n24207 ^ n24151;
  assign n24342 = ~n24208 & ~n24341;
  assign n24343 = n24342 ^ n24151;
  assign n24359 = n24358 ^ n24343;
  assign n24330 = n44 & n20294;
  assign n24331 = n3280 & n19233;
  assign n24332 = n3277 & n19139;
  assign n24333 = n3275 & ~n19142;
  assign n24334 = ~n24332 & ~n24333;
  assign n24335 = ~n24331 & n24334;
  assign n24336 = ~n24330 & n24335;
  assign n24337 = n24336 ^ x29;
  assign n24318 = n41 & ~n20210;
  assign n24319 = x31 & ~n24158;
  assign n24320 = n91 & ~n19215;
  assign n24321 = n24319 & ~n24320;
  assign n24322 = ~n24318 & n24321;
  assign n24323 = n41 & ~n19225;
  assign n24324 = n54 & ~n19215;
  assign n24325 = ~x31 & ~n24324;
  assign n24326 = ~n24323 & n24325;
  assign n24327 = ~n24322 & ~n24326;
  assign n24300 = n771 & n3368;
  assign n24301 = n11663 & n24300;
  assign n24302 = n1834 & n4734;
  assign n24303 = n11028 & n24302;
  assign n24304 = ~n456 & ~n709;
  assign n24305 = ~n334 & n24304;
  assign n24306 = ~n656 & n1302;
  assign n24307 = n24305 & n24306;
  assign n24308 = n24303 & n24307;
  assign n24309 = n24301 & n24308;
  assign n24310 = n1897 & n10997;
  assign n24311 = n24309 & n24310;
  assign n24312 = n4225 & n5623;
  assign n24313 = n12161 & n24312;
  assign n24314 = n24311 & n24313;
  assign n24315 = n968 & n24314;
  assign n24316 = n3225 & n24315;
  assign n24317 = n24316 ^ x2;
  assign n24328 = n24327 ^ n24317;
  assign n24297 = n24187 ^ n24157;
  assign n24298 = ~n24188 & n24297;
  assign n24299 = n24298 ^ n24167;
  assign n24329 = n24328 ^ n24299;
  assign n24338 = n24337 ^ n24329;
  assign n24294 = n24197 ^ n24154;
  assign n24295 = ~n24198 & n24294;
  assign n24296 = n24295 ^ n24154;
  assign n24339 = n24338 ^ n24296;
  assign n24286 = n3285 & ~n19696;
  assign n24287 = n3437 & ~n19255;
  assign n24288 = n3435 & n19253;
  assign n24289 = ~n3440 & ~n19238;
  assign n24290 = ~n24288 & ~n24289;
  assign n24291 = ~n24287 & n24290;
  assign n24292 = ~n24286 & n24291;
  assign n24293 = n24292 ^ x26;
  assign n24340 = n24339 ^ n24293;
  assign n24360 = n24359 ^ n24340;
  assign n24278 = n4673 & n21215;
  assign n24279 = n4688 & n19104;
  assign n24280 = ~n4681 & n19122;
  assign n24281 = n4685 & ~n19286;
  assign n24282 = ~n24280 & ~n24281;
  assign n24283 = ~n24279 & n24282;
  assign n24284 = ~n24278 & n24283;
  assign n24285 = n24284 ^ x20;
  assign n24361 = n24360 ^ n24285;
  assign n24275 = n24209 ^ n24132;
  assign n24276 = n24210 & n24275;
  assign n24277 = n24276 ^ n24132;
  assign n24362 = n24361 ^ n24277;
  assign n24376 = n24375 ^ n24362;
  assign n24267 = n4963 & n19668;
  assign n24268 = n4976 & n19096;
  assign n24269 = n4970 & n19292;
  assign n24270 = ~n24268 & ~n24269;
  assign n24271 = n4972 & n19298;
  assign n24272 = n24270 & ~n24271;
  assign n24273 = ~n24267 & n24272;
  assign n24274 = n24273 ^ x17;
  assign n24377 = n24376 ^ n24274;
  assign n24394 = n24393 ^ n24377;
  assign n24264 = n24213 ^ n24110;
  assign n24265 = ~n24214 & n24264;
  assign n24266 = n24265 ^ n24110;
  assign n24395 = n24394 ^ n24266;
  assign n24404 = n24403 ^ n24395;
  assign n24261 = n24215 ^ n24091;
  assign n24262 = n24216 & n24261;
  assign n24263 = n24262 ^ n24091;
  assign n24405 = n24404 ^ n24263;
  assign n24258 = n24217 ^ n24080;
  assign n24259 = n24218 & ~n24258;
  assign n24260 = n24259 ^ n24080;
  assign n24406 = n24405 ^ n24260;
  assign n24250 = n6306 & n23712;
  assign n24251 = n6309 & n19649;
  assign n24252 = n6316 & ~n19575;
  assign n24253 = ~n24251 & ~n24252;
  assign n24254 = n7168 & n23052;
  assign n24255 = n24253 & ~n24254;
  assign n24256 = ~n24250 & n24255;
  assign n24257 = n24256 ^ x8;
  assign n24407 = n24406 ^ n24257;
  assign n24244 = n7515 & ~n23704;
  assign n24245 = n7518 & n23495;
  assign n24246 = n7520 & ~n23292;
  assign n24247 = ~n24245 & ~n24246;
  assign n24248 = ~n24244 & n24247;
  assign n24249 = n24248 ^ x5;
  assign n24408 = n24407 ^ n24249;
  assign n24241 = n24219 ^ n24074;
  assign n24242 = ~n24220 & n24241;
  assign n24243 = n24242 ^ n24077;
  assign n24409 = n24408 ^ n24243;
  assign n24236 = n24221 ^ x2;
  assign n24237 = n24065 ^ x5;
  assign n24238 = n24237 ^ n24221;
  assign n24239 = n24236 & n24238;
  assign n24240 = n24239 ^ x2;
  assign n24410 = n24409 ^ n24240;
  assign n24421 = n24420 ^ n24410;
  assign n24229 = ~n24054 & n24227;
  assign n24230 = n23875 & ~n24229;
  assign n24231 = ~n24052 & ~n24227;
  assign n24232 = n24231 ^ n24049;
  assign n24233 = n24040 & n24232;
  assign n24234 = n24233 ^ n24049;
  assign n24235 = n24230 & ~n24234;
  assign n24422 = n24421 ^ n24235;
  assign n24595 = ~n24240 & ~n24407;
  assign n24596 = n24420 & n24595;
  assign n24597 = ~n24249 & ~n24596;
  assign n24598 = n24420 ^ n24240;
  assign n24599 = n24407 ^ n24240;
  assign n24600 = ~n24598 & ~n24599;
  assign n24601 = n24600 ^ n24420;
  assign n24602 = ~n24597 & n24601;
  assign n24603 = n24243 & ~n24602;
  assign n24604 = ~n24249 & ~n24601;
  assign n24605 = n24240 & n24407;
  assign n24606 = ~n24420 & n24605;
  assign n24607 = ~n24243 & ~n24606;
  assign n24608 = ~n24604 & n24607;
  assign n24609 = ~n24603 & ~n24608;
  assign n24610 = n24606 ^ n24596;
  assign n24611 = ~n24249 & n24610;
  assign n24612 = n24611 ^ n24596;
  assign n24613 = ~n24609 & ~n24612;
  assign n24591 = n7520 & n23495;
  assign n24592 = n24591 ^ x5;
  assign n24588 = n24405 ^ n24257;
  assign n24589 = ~n24406 & n24588;
  assign n24590 = n24589 ^ n24260;
  assign n24593 = n24592 ^ n24590;
  assign n24577 = n16805 & ~n23879;
  assign n24570 = n6316 & n19649;
  assign n24571 = n6309 & n23052;
  assign n24572 = ~n24570 & ~n24571;
  assign n24573 = x8 & n24572;
  assign n24578 = n23292 & n24573;
  assign n24579 = ~n24577 & ~n24578;
  assign n24574 = n23879 & n24573;
  assign n24575 = n16805 & ~n23292;
  assign n24576 = ~n24574 & ~n24575;
  assign n24580 = n24579 ^ n24576;
  assign n24581 = ~x7 & n24580;
  assign n24582 = n24581 ^ n24579;
  assign n24583 = ~n16820 & n24572;
  assign n24584 = n24583 ^ x8;
  assign n24585 = n24582 & n24584;
  assign n24567 = n24403 ^ n24263;
  assign n24568 = n24404 & n24567;
  assign n24569 = n24568 ^ n24263;
  assign n24586 = n24585 ^ n24569;
  assign n24546 = ~x14 & ~n22036;
  assign n24547 = ~n5746 & n19063;
  assign n24548 = n5752 & n19303;
  assign n24549 = ~n24547 & ~n24548;
  assign n24550 = x14 & ~n24549;
  assign n24551 = ~n24546 & ~n24550;
  assign n24552 = ~x13 & n22036;
  assign n24553 = n24551 & ~n24552;
  assign n24554 = ~n6048 & n19368;
  assign n24555 = n24553 & n24554;
  assign n24556 = ~n7589 & n24549;
  assign n24557 = n24556 ^ x14;
  assign n24558 = ~n24555 & n24557;
  assign n24559 = ~n24546 & ~n24552;
  assign n24560 = ~n6048 & ~n19368;
  assign n24561 = ~n24550 & n24560;
  assign n24562 = ~n24559 & n24561;
  assign n24563 = n24558 & ~n24562;
  assign n24536 = n4963 & ~n21715;
  assign n24537 = n4972 & ~n19078;
  assign n24538 = n4976 & n19298;
  assign n24539 = n4970 & n19096;
  assign n24540 = ~n24538 & ~n24539;
  assign n24541 = ~n24537 & n24540;
  assign n24542 = ~n24536 & n24541;
  assign n24543 = n24542 ^ x17;
  assign n24524 = n4478 & n21189;
  assign n24525 = n4487 & n19122;
  assign n24526 = n4484 & ~n19281;
  assign n24527 = n4480 & n19277;
  assign n24528 = ~n24526 & ~n24527;
  assign n24529 = ~n24525 & n24528;
  assign n24530 = ~n24524 & n24529;
  assign n24531 = n24530 ^ x23;
  assign n24506 = n12417 & n20929;
  assign n24507 = n3435 & ~n19255;
  assign n24508 = ~n3440 & n19253;
  assign n24509 = ~n24507 & ~n24508;
  assign n24510 = x26 & n24509;
  assign n24511 = ~n19260 & n24510;
  assign n24512 = x25 & ~n24511;
  assign n24513 = ~n24506 & n24512;
  assign n24514 = ~n20929 & n24510;
  assign n24515 = n12417 & n19260;
  assign n24516 = ~x25 & ~n24515;
  assign n24517 = ~n24514 & n24516;
  assign n24518 = ~n24513 & ~n24517;
  assign n24519 = ~n12432 & n24509;
  assign n24520 = n24519 ^ x26;
  assign n24521 = ~n24518 & n24520;
  assign n24493 = n41 & ~n20045;
  assign n24494 = n91 & ~n19225;
  assign n24495 = x31 & ~n24324;
  assign n24496 = ~n24494 & n24495;
  assign n24497 = ~n24493 & n24496;
  assign n24498 = n41 & ~n19142;
  assign n24499 = n54 & ~n19225;
  assign n24500 = ~n24498 & ~n24499;
  assign n24501 = ~x31 & n24500;
  assign n24502 = ~n24497 & ~n24501;
  assign n24490 = n24337 ^ n24328;
  assign n24491 = n24329 & n24490;
  assign n24492 = n24491 ^ n24337;
  assign n24503 = n24502 ^ n24492;
  assign n24484 = n24316 & ~n24327;
  assign n24485 = x2 & ~n24484;
  assign n24486 = ~n24316 & n24327;
  assign n24487 = ~n24485 & ~n24486;
  assign n24463 = n285 & n4565;
  assign n24464 = ~n234 & ~n362;
  assign n24465 = n1197 & n24464;
  assign n24466 = n24463 & n24465;
  assign n24467 = n2002 & n24466;
  assign n24468 = n58 & n172;
  assign n24469 = n1231 & n2489;
  assign n24470 = n24468 & n24469;
  assign n24471 = n3576 & n3957;
  assign n24472 = n766 & ~n1405;
  assign n24473 = n24471 & n24472;
  assign n24474 = n24470 & n24473;
  assign n24475 = n24467 & n24474;
  assign n24476 = n1685 & n24475;
  assign n24477 = n13515 & n24476;
  assign n24478 = ~n208 & ~n313;
  assign n24479 = n4759 & n24478;
  assign n24480 = n893 & n13488;
  assign n24481 = n24479 & n24480;
  assign n24482 = n1970 & n24481;
  assign n24483 = n24477 & n24482;
  assign n24488 = n24487 ^ n24483;
  assign n24489 = n24488 ^ x2;
  assign n24504 = n24503 ^ n24489;
  assign n24455 = n44 & ~n20328;
  assign n24456 = n3280 & ~n19238;
  assign n24457 = n3277 & n19233;
  assign n24458 = n3275 & n19139;
  assign n24459 = ~n24457 & ~n24458;
  assign n24460 = ~n24456 & n24459;
  assign n24461 = ~n24455 & n24460;
  assign n24462 = n24461 ^ x29;
  assign n24505 = n24504 ^ n24462;
  assign n24522 = n24521 ^ n24505;
  assign n24452 = n24338 ^ n24293;
  assign n24453 = ~n24339 & n24452;
  assign n24454 = n24453 ^ n24296;
  assign n24523 = n24522 ^ n24454;
  assign n24532 = n24531 ^ n24523;
  assign n24449 = n24358 ^ n24340;
  assign n24450 = ~n24359 & n24449;
  assign n24451 = n24450 ^ n24343;
  assign n24533 = n24532 ^ n24451;
  assign n24441 = n4673 & n21684;
  assign n24442 = n4688 & n19292;
  assign n24443 = n4685 & n19104;
  assign n24444 = ~n4681 & ~n19286;
  assign n24445 = ~n24443 & ~n24444;
  assign n24446 = ~n24442 & n24445;
  assign n24447 = ~n24441 & n24446;
  assign n24448 = n24447 ^ x20;
  assign n24534 = n24533 ^ n24448;
  assign n24438 = n24360 ^ n24277;
  assign n24439 = ~n24361 & ~n24438;
  assign n24440 = n24439 ^ n24277;
  assign n24535 = n24534 ^ n24440;
  assign n24544 = n24543 ^ n24535;
  assign n24435 = n24362 ^ n24274;
  assign n24436 = ~n24376 & n24435;
  assign n24437 = n24436 ^ n24375;
  assign n24545 = n24544 ^ n24437;
  assign n24564 = n24563 ^ n24545;
  assign n24432 = n24393 ^ n24266;
  assign n24433 = n24394 & n24432;
  assign n24434 = n24433 ^ n24266;
  assign n24565 = n24564 ^ n24434;
  assign n24424 = n5814 & ~n23468;
  assign n24425 = n5817 & ~n19512;
  assign n24426 = n5824 & n19439;
  assign n24427 = ~n24425 & ~n24426;
  assign n24428 = n6295 & ~n19575;
  assign n24429 = n24427 & ~n24428;
  assign n24430 = ~n24424 & n24429;
  assign n24431 = n24430 ^ x11;
  assign n24566 = n24565 ^ n24431;
  assign n24587 = n24586 ^ n24566;
  assign n24594 = n24593 ^ n24587;
  assign n24614 = n24613 ^ n24594;
  assign n24423 = n24235 & ~n24421;
  assign n24615 = n24614 ^ n24423;
  assign n24792 = n24423 & n24614;
  assign n24777 = ~n24249 & ~n24420;
  assign n24778 = ~n24243 & n24777;
  assign n24779 = ~n24594 & ~n24778;
  assign n24780 = n24249 & n24420;
  assign n24781 = n24243 & n24780;
  assign n24782 = ~n24595 & ~n24781;
  assign n24783 = ~n24779 & n24782;
  assign n24784 = n24243 & ~n24777;
  assign n24785 = ~n24594 & ~n24605;
  assign n24786 = ~n24780 & ~n24785;
  assign n24787 = ~n24784 & n24786;
  assign n24788 = n24594 & n24605;
  assign n24789 = ~n24787 & ~n24788;
  assign n24790 = ~n24783 & n24789;
  assign n24765 = n6306 & n23493;
  assign n24766 = n7168 & n23495;
  assign n24767 = n6309 & ~n23292;
  assign n24768 = n6316 & n23052;
  assign n24769 = ~n24767 & ~n24768;
  assign n24770 = ~n24766 & n24769;
  assign n24771 = ~n24765 & n24770;
  assign n24772 = n24771 ^ x8;
  assign n24755 = n5814 & n23520;
  assign n24756 = n6295 & n19649;
  assign n24757 = n5817 & ~n19575;
  assign n24758 = n5824 & ~n19512;
  assign n24759 = ~n24757 & ~n24758;
  assign n24760 = ~n24756 & n24759;
  assign n24761 = ~n24755 & n24760;
  assign n24762 = n24761 ^ x11;
  assign n24737 = n6033 & n22457;
  assign n24738 = ~n5746 & ~n19368;
  assign n24739 = n5752 & n19063;
  assign n24740 = ~n24738 & ~n24739;
  assign n24741 = x14 & n24740;
  assign n24742 = ~n19439 & n24741;
  assign n24743 = x13 & ~n24742;
  assign n24744 = ~n24737 & n24743;
  assign n24745 = ~n22457 & n24741;
  assign n24746 = n6033 & n19439;
  assign n24747 = ~x13 & ~n24746;
  assign n24748 = ~n24745 & n24747;
  assign n24749 = ~n24744 & ~n24748;
  assign n24750 = ~n7589 & n24740;
  assign n24751 = n24750 ^ x14;
  assign n24752 = ~n24749 & n24751;
  assign n24718 = n5771 & n19658;
  assign n24719 = n4976 & ~n19078;
  assign n24720 = n4970 & n19298;
  assign n24721 = ~n24719 & ~n24720;
  assign n24722 = x17 & n24721;
  assign n24723 = ~n19303 & n24722;
  assign n24724 = ~n24718 & ~n24723;
  assign n24725 = x16 & n24724;
  assign n24726 = ~n19658 & n24722;
  assign n24727 = n5771 & n19303;
  assign n24728 = ~x16 & ~n24727;
  assign n24729 = ~n24726 & n24728;
  assign n24730 = ~n24725 & ~n24729;
  assign n24731 = ~n5786 & n24721;
  assign n24732 = n24731 ^ x17;
  assign n24733 = ~n24730 & n24732;
  assign n24715 = n24532 ^ n24448;
  assign n24716 = ~n24533 & ~n24715;
  assign n24717 = n24716 ^ n24451;
  assign n24734 = n24733 ^ n24717;
  assign n24706 = n4673 & n21699;
  assign n24707 = n4688 & n19096;
  assign n24708 = n4685 & n19292;
  assign n24709 = ~n4681 & n19104;
  assign n24710 = ~n24708 & ~n24709;
  assign n24711 = ~n24707 & n24710;
  assign n24712 = ~n24706 & n24711;
  assign n24713 = n24712 ^ x20;
  assign n24696 = n4478 & ~n19678;
  assign n24697 = n4484 & n19122;
  assign n24698 = n4487 & ~n19286;
  assign n24699 = n4480 & ~n19281;
  assign n24700 = ~n24698 & ~n24699;
  assign n24701 = ~n24697 & n24700;
  assign n24702 = ~n24696 & n24701;
  assign n24703 = n24702 ^ x23;
  assign n24677 = n19230 ^ n19139;
  assign n24678 = n19142 & n24677;
  assign n24679 = n41 & n24678;
  assign n24680 = ~n24499 & ~n24679;
  assign n24681 = x31 & ~n24680;
  assign n24682 = ~n91 & n24677;
  assign n24683 = n12183 & ~n19142;
  assign n24684 = ~n24682 & n24683;
  assign n24685 = ~n54 & ~n19139;
  assign n24686 = n54 & n19142;
  assign n24687 = n3640 & ~n24686;
  assign n24688 = ~n24685 & n24687;
  assign n24689 = ~n24684 & ~n24688;
  assign n24690 = ~n24681 & n24689;
  assign n24674 = n24502 ^ n24489;
  assign n24675 = ~n24503 & ~n24674;
  assign n24676 = n24675 ^ n24492;
  assign n24691 = n24690 ^ n24676;
  assign n24658 = ~n237 & n1075;
  assign n24659 = n2461 & n24658;
  assign n24660 = n3823 & n24659;
  assign n24661 = n12883 & n24660;
  assign n24662 = ~n313 & ~n743;
  assign n24663 = ~n193 & ~n272;
  assign n24664 = n24662 & n24663;
  assign n24665 = n603 & n24664;
  assign n24666 = n813 & n1136;
  assign n24667 = n24665 & n24666;
  assign n24668 = n4121 & n24667;
  assign n24669 = n24661 & n24668;
  assign n24670 = n389 & n24669;
  assign n24671 = n1605 & n24670;
  assign n24672 = n2700 & n24671;
  assign n24653 = n24327 ^ x2;
  assign n24654 = n24327 ^ n24316;
  assign n24655 = n24483 ^ n24316;
  assign n24656 = n24654 & ~n24655;
  assign n24657 = n24653 & n24656;
  assign n24673 = n24672 ^ n24657;
  assign n24692 = n24691 ^ n24673;
  assign n24645 = n3285 & n20793;
  assign n24646 = n3437 & n19277;
  assign n24647 = n3435 & n19260;
  assign n24648 = ~n3440 & ~n19255;
  assign n24649 = ~n24647 & ~n24648;
  assign n24650 = ~n24646 & n24649;
  assign n24651 = ~n24645 & n24650;
  assign n24652 = n24651 ^ x26;
  assign n24693 = n24692 ^ n24652;
  assign n24637 = n44 & n20308;
  assign n24638 = n3280 & n19253;
  assign n24639 = n3277 & ~n19238;
  assign n24640 = n3275 & n19233;
  assign n24641 = ~n24639 & ~n24640;
  assign n24642 = ~n24638 & n24641;
  assign n24643 = ~n24637 & n24642;
  assign n24644 = n24643 ^ x29;
  assign n24694 = n24693 ^ n24644;
  assign n24634 = n24521 ^ n24504;
  assign n24635 = ~n24505 & n24634;
  assign n24636 = n24635 ^ n24521;
  assign n24695 = n24694 ^ n24636;
  assign n24704 = n24703 ^ n24695;
  assign n24631 = n24531 ^ n24454;
  assign n24632 = ~n24523 & n24631;
  assign n24633 = n24632 ^ n24531;
  assign n24705 = n24704 ^ n24633;
  assign n24714 = n24713 ^ n24705;
  assign n24735 = n24734 ^ n24714;
  assign n24628 = n24543 ^ n24440;
  assign n24629 = ~n24535 & ~n24628;
  assign n24630 = n24629 ^ n24543;
  assign n24736 = n24735 ^ n24630;
  assign n24753 = n24752 ^ n24736;
  assign n24625 = n24563 ^ n24437;
  assign n24626 = ~n24545 & n24625;
  assign n24627 = n24626 ^ n24563;
  assign n24754 = n24753 ^ n24627;
  assign n24763 = n24762 ^ n24754;
  assign n24622 = n24564 ^ n24431;
  assign n24623 = n24565 & ~n24622;
  assign n24624 = n24623 ^ n24434;
  assign n24764 = n24763 ^ n24624;
  assign n24773 = n24772 ^ n24764;
  assign n24774 = n24773 ^ x5;
  assign n24619 = n24585 ^ n24566;
  assign n24620 = n24586 & ~n24619;
  assign n24621 = n24620 ^ n24569;
  assign n24775 = n24774 ^ n24621;
  assign n24616 = n24592 ^ n24587;
  assign n24617 = ~n24593 & n24616;
  assign n24618 = n24617 ^ n24590;
  assign n24776 = n24775 ^ n24618;
  assign n24791 = n24790 ^ n24776;
  assign n24793 = n24792 ^ n24791;
  assign n24959 = n24621 & ~n24773;
  assign n24960 = x5 & ~n24959;
  assign n24961 = ~n24621 & n24773;
  assign n24962 = ~n24960 & ~n24961;
  assign n24951 = n6306 & ~n23704;
  assign n24952 = n6309 & n23495;
  assign n24953 = n6316 & ~n23292;
  assign n24954 = ~n24952 & ~n24953;
  assign n24955 = ~n24951 & n24954;
  assign n24956 = n24955 ^ x8;
  assign n24931 = ~x13 & ~n23064;
  assign n24932 = x13 & ~n19512;
  assign n24933 = x14 & ~n24932;
  assign n24934 = ~n24931 & n24933;
  assign n24935 = ~n5746 & n19439;
  assign n24936 = n5752 & ~n19368;
  assign n24937 = ~n24935 & ~n24936;
  assign n24938 = ~n7559 & n24937;
  assign n24939 = ~n24934 & n24938;
  assign n24940 = x14 & ~n24937;
  assign n24941 = ~n24939 & ~n24940;
  assign n24942 = n23064 ^ n19512;
  assign n24943 = x13 & n24942;
  assign n24944 = n24943 ^ n19512;
  assign n24945 = n6033 & ~n24944;
  assign n24946 = ~n24941 & ~n24945;
  assign n24928 = n24752 ^ n24735;
  assign n24929 = n24736 & ~n24928;
  assign n24930 = n24929 ^ n24752;
  assign n24947 = n24946 ^ n24930;
  assign n24918 = n4963 & n22441;
  assign n24919 = n4972 & n19063;
  assign n24920 = n4970 & ~n19078;
  assign n24921 = n4976 & n19303;
  assign n24922 = ~n24920 & ~n24921;
  assign n24923 = ~n24919 & n24922;
  assign n24924 = ~n24918 & n24923;
  assign n24925 = n24924 ^ x17;
  assign n24901 = ~x19 & n19668;
  assign n24902 = x19 & n19298;
  assign n24903 = x20 & ~n24902;
  assign n24904 = ~n24901 & n24903;
  assign n24905 = ~n13667 & ~n24904;
  assign n24906 = n4685 & n19096;
  assign n24907 = ~n4681 & n19292;
  assign n24908 = ~n24906 & ~n24907;
  assign n24909 = ~n24905 & n24908;
  assign n24910 = n15622 & n19668;
  assign n24911 = ~x19 & n4671;
  assign n24912 = n19298 & n24911;
  assign n24913 = n24908 & ~n24912;
  assign n24914 = ~n24910 & n24913;
  assign n24915 = ~x20 & ~n24914;
  assign n24916 = ~n24909 & ~n24915;
  assign n24890 = n4478 & n21215;
  assign n24891 = n4487 & n19104;
  assign n24892 = n4480 & n19122;
  assign n24893 = n4484 & ~n19286;
  assign n24894 = ~n24892 & ~n24893;
  assign n24895 = ~n24891 & n24894;
  assign n24896 = ~n24890 & n24895;
  assign n24897 = n24896 ^ x23;
  assign n24887 = n24703 ^ n24694;
  assign n24888 = ~n24695 & n24887;
  assign n24889 = n24888 ^ n24703;
  assign n24898 = n24897 ^ n24889;
  assign n24869 = n12417 & ~n20908;
  assign n24870 = n3435 & n19277;
  assign n24871 = ~n3440 & n19260;
  assign n24872 = ~n24870 & ~n24871;
  assign n24873 = x26 & n24872;
  assign n24874 = n19281 & n24873;
  assign n24875 = x25 & ~n24874;
  assign n24876 = ~n24869 & n24875;
  assign n24877 = n20908 & n24873;
  assign n24878 = n12417 & ~n19281;
  assign n24879 = ~x25 & ~n24878;
  assign n24880 = ~n24877 & n24879;
  assign n24881 = ~n24876 & ~n24880;
  assign n24882 = ~n12432 & n24872;
  assign n24883 = n24882 ^ x26;
  assign n24884 = ~n24881 & n24883;
  assign n24866 = n24652 ^ n24644;
  assign n24867 = n24693 & ~n24866;
  assign n24868 = n24867 ^ n24692;
  assign n24885 = n24884 ^ n24868;
  assign n24856 = n44 & ~n19696;
  assign n24857 = n3280 & ~n19255;
  assign n24858 = n3277 & n19253;
  assign n24859 = n3275 & ~n19238;
  assign n24860 = ~n24858 & ~n24859;
  assign n24861 = ~n24857 & n24860;
  assign n24862 = ~n24856 & n24861;
  assign n24863 = n24862 ^ x29;
  assign n24839 = n964 & n3087;
  assign n24840 = n4734 & n24839;
  assign n24841 = n11566 & n24840;
  assign n24842 = n4039 & n4723;
  assign n24843 = ~n133 & ~n666;
  assign n24844 = n2771 & n24843;
  assign n24845 = ~n217 & ~n293;
  assign n24846 = ~n115 & n24845;
  assign n24847 = n24844 & n24846;
  assign n24848 = n24842 & n24847;
  assign n24849 = n24841 & n24848;
  assign n24850 = n20715 & n24849;
  assign n24851 = n3605 & n24850;
  assign n24852 = n2064 & n24851;
  assign n24853 = n24852 ^ x5;
  assign n24832 = n41 & ~n20294;
  assign n24833 = n91 & ~n19139;
  assign n24834 = ~n24686 & ~n24833;
  assign n24835 = ~n24832 & n24834;
  assign n24829 = n41 & n19233;
  assign n24830 = n54 & n19139;
  assign n24831 = ~n24829 & ~n24830;
  assign n24836 = n24835 ^ n24831;
  assign n24837 = ~x31 & ~n24836;
  assign n24838 = n24837 ^ n24835;
  assign n24854 = n24853 ^ n24838;
  assign n24824 = ~n24483 & ~n24487;
  assign n24825 = ~n24672 & n24824;
  assign n24822 = n24483 & n24672;
  assign n24823 = n24487 & n24822;
  assign n24826 = n24825 ^ n24823;
  assign n24827 = x2 & n24826;
  assign n24828 = n24827 ^ n24825;
  assign n24855 = n24854 ^ n24828;
  assign n24864 = n24863 ^ n24855;
  assign n24819 = n24690 ^ n24673;
  assign n24820 = n24691 & ~n24819;
  assign n24821 = n24820 ^ n24676;
  assign n24865 = n24864 ^ n24821;
  assign n24886 = n24885 ^ n24865;
  assign n24899 = n24898 ^ n24886;
  assign n24816 = n24713 ^ n24704;
  assign n24817 = ~n24705 & n24816;
  assign n24818 = n24817 ^ n24713;
  assign n24900 = n24899 ^ n24818;
  assign n24917 = n24916 ^ n24900;
  assign n24926 = n24925 ^ n24917;
  assign n24813 = n24717 ^ n24714;
  assign n24814 = ~n24734 & n24813;
  assign n24815 = n24814 ^ n24733;
  assign n24927 = n24926 ^ n24815;
  assign n24948 = n24947 ^ n24927;
  assign n24805 = n5814 & n23712;
  assign n24806 = n5817 & n19649;
  assign n24807 = n5824 & ~n19575;
  assign n24808 = ~n24806 & ~n24807;
  assign n24809 = n6295 & n23052;
  assign n24810 = n24808 & ~n24809;
  assign n24811 = ~n24805 & n24810;
  assign n24812 = n24811 ^ x11;
  assign n24949 = n24948 ^ n24812;
  assign n24802 = n24762 ^ n24627;
  assign n24803 = n24754 & n24802;
  assign n24804 = n24803 ^ n24762;
  assign n24950 = n24949 ^ n24804;
  assign n24957 = n24956 ^ n24950;
  assign n24799 = n24772 ^ n24763;
  assign n24800 = n24764 & ~n24799;
  assign n24801 = n24800 ^ n24772;
  assign n24958 = n24957 ^ n24801;
  assign n24963 = n24962 ^ n24958;
  assign n24794 = n24790 ^ n24618;
  assign n24796 = n24794 ^ n24775;
  assign n24797 = ~n24792 & ~n24796;
  assign n24795 = ~n24776 & ~n24794;
  assign n24798 = n24797 ^ n24795;
  assign n24964 = n24963 ^ n24798;
  assign n25139 = n24776 & n24790;
  assign n25140 = n24963 & n25139;
  assign n25141 = n24963 ^ n24775;
  assign n25142 = ~n24776 & ~n25141;
  assign n25143 = ~n24790 & n25142;
  assign n25144 = ~n25140 & ~n25143;
  assign n25145 = n24792 & ~n25144;
  assign n25136 = n24956 ^ n24801;
  assign n25137 = ~n24957 & n25136;
  assign n25138 = n25137 ^ n24801;
  assign n25146 = n25145 ^ n25138;
  assign n25120 = ~x5 & n24618;
  assign n25121 = n24790 & n25120;
  assign n25122 = ~n24958 & ~n24959;
  assign n25123 = ~n25121 & n25122;
  assign n25124 = ~n24618 & ~n24790;
  assign n25125 = n24960 & n25124;
  assign n25126 = ~n25123 & ~n25125;
  assign n25127 = x5 & ~n24618;
  assign n25128 = n24790 & ~n25127;
  assign n25129 = n24958 & ~n24961;
  assign n25130 = ~n25120 & ~n25129;
  assign n25131 = ~n25128 & n25130;
  assign n25132 = ~n24958 & n24961;
  assign n25133 = ~n25131 & ~n25132;
  assign n25134 = n25126 & n25133;
  assign n25110 = n5814 & ~n23879;
  assign n25111 = n6295 & ~n23292;
  assign n25112 = n5817 & n23052;
  assign n25113 = n5824 & n19649;
  assign n25114 = ~n25112 & ~n25113;
  assign n25115 = ~n25111 & n25114;
  assign n25116 = ~n25110 & n25115;
  assign n25117 = n25116 ^ x11;
  assign n25098 = n4963 & ~n22037;
  assign n25099 = n4972 & ~n19368;
  assign n25100 = n4976 & n19063;
  assign n25101 = n4970 & n19303;
  assign n25102 = ~n25100 & ~n25101;
  assign n25103 = ~n25099 & n25102;
  assign n25104 = ~n25098 & n25103;
  assign n25105 = n25104 ^ x17;
  assign n25088 = n4673 & ~n21715;
  assign n25089 = n4688 & ~n19078;
  assign n25090 = n4685 & n19298;
  assign n25091 = ~n4681 & n19096;
  assign n25092 = ~n25090 & ~n25091;
  assign n25093 = ~n25089 & n25092;
  assign n25094 = ~n25088 & n25093;
  assign n25095 = n25094 ^ x20;
  assign n25078 = n4478 & n21684;
  assign n25079 = n4487 & n19292;
  assign n25080 = n4484 & n19104;
  assign n25081 = n4480 & ~n19286;
  assign n25082 = ~n25080 & ~n25081;
  assign n25083 = ~n25079 & n25082;
  assign n25084 = ~n25078 & n25083;
  assign n25085 = n25084 ^ x23;
  assign n25062 = ~n24838 & n24853;
  assign n25063 = n24825 & ~n25062;
  assign n25064 = n24838 & ~n24853;
  assign n25065 = ~x2 & ~n25064;
  assign n25066 = ~n25063 & n25065;
  assign n25067 = n24838 ^ n24823;
  assign n25068 = x2 & ~n24853;
  assign n25069 = n25068 ^ n24823;
  assign n25070 = ~n25067 & ~n25069;
  assign n25071 = n25070 ^ n24838;
  assign n25072 = ~n25066 & n25071;
  assign n25054 = n44 & n20929;
  assign n25055 = n3280 & n19260;
  assign n25056 = n3277 & ~n19255;
  assign n25057 = n3275 & n19253;
  assign n25058 = ~n25056 & ~n25057;
  assign n25059 = ~n25055 & n25058;
  assign n25060 = ~n25054 & n25059;
  assign n25061 = n25060 ^ x29;
  assign n25073 = n25072 ^ n25061;
  assign n25043 = n41 & ~n20328;
  assign n25044 = n91 & n19233;
  assign n25045 = ~n24830 & ~n25044;
  assign n25046 = ~n25043 & n25045;
  assign n25047 = x31 & ~n25046;
  assign n25048 = ~n54 & n19238;
  assign n25049 = n54 & ~n19233;
  assign n25050 = n3640 & ~n25049;
  assign n25051 = ~n25048 & n25050;
  assign n25052 = ~n25047 & ~n25051;
  assign n25038 = x2 & x5;
  assign n25039 = ~x2 & ~x5;
  assign n25040 = n24852 & ~n25039;
  assign n25041 = ~n25038 & ~n25040;
  assign n25012 = ~n134 & ~n1135;
  assign n25013 = n11807 & n25012;
  assign n25014 = n5651 & n25013;
  assign n25015 = n2822 & n25014;
  assign n25016 = n1496 & n3606;
  assign n25017 = n25015 & n25016;
  assign n25018 = n3840 & n4614;
  assign n25019 = ~n257 & ~n313;
  assign n25020 = n684 & n25019;
  assign n25021 = n1121 & n25020;
  assign n25022 = n25018 & n25021;
  assign n25023 = n2380 & n25022;
  assign n25024 = n25017 & n25023;
  assign n25025 = n756 & n1841;
  assign n25026 = n5616 & n25025;
  assign n25027 = n1288 & n2433;
  assign n25028 = n5113 & n25027;
  assign n25029 = n25026 & n25028;
  assign n25030 = ~n103 & ~n330;
  assign n25031 = ~n263 & n25030;
  assign n25032 = n11069 & n25031;
  assign n25033 = n11080 & n25032;
  assign n25034 = n2920 & n25033;
  assign n25035 = n25029 & n25034;
  assign n25036 = n25024 & n25035;
  assign n25037 = n565 & n25036;
  assign n25042 = n25041 ^ n25037;
  assign n25053 = n25052 ^ n25042;
  assign n25074 = n25073 ^ n25053;
  assign n25009 = n24863 ^ n24821;
  assign n25010 = ~n24864 & n25009;
  assign n25011 = n25010 ^ n24821;
  assign n25075 = n25074 ^ n25011;
  assign n25001 = n3285 & n21189;
  assign n25002 = n3437 & n19122;
  assign n25003 = n3435 & ~n19281;
  assign n25004 = ~n3440 & n19277;
  assign n25005 = ~n25003 & ~n25004;
  assign n25006 = ~n25002 & n25005;
  assign n25007 = ~n25001 & n25006;
  assign n25008 = n25007 ^ x26;
  assign n25076 = n25075 ^ n25008;
  assign n24998 = n24884 ^ n24865;
  assign n24999 = n24885 & ~n24998;
  assign n25000 = n24999 ^ n24868;
  assign n25077 = n25076 ^ n25000;
  assign n25086 = n25085 ^ n25077;
  assign n24995 = n24897 ^ n24886;
  assign n24996 = n24898 & ~n24995;
  assign n24997 = n24996 ^ n24889;
  assign n25087 = n25086 ^ n24997;
  assign n25096 = n25095 ^ n25087;
  assign n24992 = n24916 ^ n24818;
  assign n24993 = ~n24900 & n24992;
  assign n24994 = n24993 ^ n24916;
  assign n25097 = n25096 ^ n24994;
  assign n25106 = n25105 ^ n25097;
  assign n24989 = n24925 ^ n24815;
  assign n24990 = ~n24926 & n24989;
  assign n24991 = n24990 ^ n24815;
  assign n25107 = n25106 ^ n24991;
  assign n24983 = n5749 & ~n22989;
  assign n24984 = n24983 ^ x13;
  assign n24985 = n24984 ^ n19575;
  assign n24974 = ~x13 & ~n19512;
  assign n24975 = n13719 & n19439;
  assign n24976 = x12 & ~n24975;
  assign n24977 = ~n24974 & n24976;
  assign n24978 = n13989 & n19439;
  assign n24979 = ~x12 & ~n24978;
  assign n24980 = ~n24932 & n24979;
  assign n24981 = ~n24977 & ~n24980;
  assign n24982 = n24981 ^ x14;
  assign n24986 = n24985 ^ n24982;
  assign n24987 = ~n5748 & ~n24986;
  assign n24988 = n24987 ^ n24985;
  assign n25108 = n25107 ^ n24988;
  assign n24971 = n24930 ^ n24927;
  assign n24972 = n24947 & ~n24971;
  assign n24973 = n24972 ^ n24946;
  assign n25109 = n25108 ^ n24973;
  assign n25118 = n25117 ^ n25109;
  assign n24968 = n6316 & n23495;
  assign n24969 = n24968 ^ x8;
  assign n24965 = n24812 ^ n24804;
  assign n24966 = n24949 & ~n24965;
  assign n24967 = n24966 ^ n24948;
  assign n24970 = n24969 ^ n24967;
  assign n25119 = n25118 ^ n24970;
  assign n25135 = n25134 ^ n25119;
  assign n25147 = n25146 ^ n25135;
  assign n25303 = n5814 & n23493;
  assign n25304 = n6295 & n23495;
  assign n25305 = n5817 & ~n23292;
  assign n25306 = n5824 & n23052;
  assign n25307 = ~n25305 & ~n25306;
  assign n25308 = ~n25304 & n25307;
  assign n25309 = ~n25303 & n25308;
  assign n25310 = n25309 ^ x11;
  assign n25285 = n6033 & n23520;
  assign n25286 = n5752 & ~n19512;
  assign n25287 = ~n5746 & ~n19575;
  assign n25288 = ~n25286 & ~n25287;
  assign n25289 = x14 & n25288;
  assign n25290 = ~n19649 & n25289;
  assign n25291 = x13 & ~n25290;
  assign n25292 = ~n25285 & n25291;
  assign n25293 = ~n23520 & n25289;
  assign n25294 = n6033 & n19649;
  assign n25295 = ~x13 & ~n25294;
  assign n25296 = ~n25293 & n25295;
  assign n25297 = ~n25292 & ~n25296;
  assign n25298 = ~n7589 & n25288;
  assign n25299 = n25298 ^ x14;
  assign n25300 = ~n25297 & n25299;
  assign n25275 = n4963 & n22457;
  assign n25276 = n4972 & n19439;
  assign n25277 = n4976 & ~n19368;
  assign n25278 = n4970 & n19063;
  assign n25279 = ~n25277 & ~n25278;
  assign n25280 = ~n25276 & n25279;
  assign n25281 = ~n25275 & n25280;
  assign n25282 = n25281 ^ x17;
  assign n25259 = ~x19 & n19657;
  assign n25260 = n25259 ^ n19303;
  assign n25261 = n4671 & n25260;
  assign n25262 = n4685 & ~n19078;
  assign n25263 = ~n4681 & n19298;
  assign n25264 = ~n25262 & ~n25263;
  assign n25265 = x20 & n25264;
  assign n25266 = ~n25261 & n25265;
  assign n25267 = n15622 & n19658;
  assign n25268 = n19303 & n24911;
  assign n25269 = n25264 & ~n25268;
  assign n25270 = ~n25267 & n25269;
  assign n25271 = ~x20 & ~n25270;
  assign n25272 = ~n25266 & ~n25271;
  assign n25249 = n4478 & n21699;
  assign n25250 = n4487 & n19096;
  assign n25251 = n4484 & n19292;
  assign n25252 = n4480 & n19104;
  assign n25253 = ~n25251 & ~n25252;
  assign n25254 = ~n25250 & n25253;
  assign n25255 = ~n25249 & n25254;
  assign n25256 = n25255 ^ x23;
  assign n25231 = n12417 & ~n19678;
  assign n25232 = n3435 & n19122;
  assign n25233 = ~n3440 & ~n19281;
  assign n25234 = ~n25232 & ~n25233;
  assign n25235 = x26 & n25234;
  assign n25236 = n19286 & n25235;
  assign n25237 = ~n25231 & ~n25236;
  assign n25238 = x25 & n25237;
  assign n25239 = n19678 & n25235;
  assign n25240 = n12417 & ~n19286;
  assign n25241 = ~x25 & ~n25240;
  assign n25242 = ~n25239 & n25241;
  assign n25243 = ~n25238 & ~n25242;
  assign n25244 = ~n12432 & n25234;
  assign n25245 = n25244 ^ x26;
  assign n25246 = ~n25243 & n25245;
  assign n25218 = n41 & ~n20308;
  assign n25219 = n91 & n19238;
  assign n25220 = x31 & ~n25049;
  assign n25221 = ~n25219 & n25220;
  assign n25222 = ~n25218 & n25221;
  assign n25223 = ~n54 & ~n19253;
  assign n25224 = n54 & n19238;
  assign n25225 = n3640 & ~n25224;
  assign n25226 = ~n25223 & n25225;
  assign n25227 = ~n25222 & ~n25226;
  assign n25187 = ~n202 & ~n656;
  assign n25188 = ~n51 & ~n283;
  assign n25189 = n25187 & n25188;
  assign n25190 = ~n452 & n1602;
  assign n25191 = n25189 & n25190;
  assign n25192 = n187 & n267;
  assign n25193 = n379 & n1044;
  assign n25194 = n25192 & n25193;
  assign n25195 = n25191 & n25194;
  assign n25196 = ~n192 & ~n227;
  assign n25197 = ~n362 & n25196;
  assign n25198 = n676 & n2753;
  assign n25199 = n25197 & n25198;
  assign n25200 = n3007 & n25199;
  assign n25201 = n3624 & n25200;
  assign n25202 = n25195 & n25201;
  assign n25203 = n3967 & n25202;
  assign n25204 = n2541 & n2765;
  assign n25205 = n2927 & n25204;
  assign n25206 = n10092 & n25205;
  assign n25207 = n768 & n25206;
  assign n25208 = n4397 & n12053;
  assign n25209 = n782 & n10888;
  assign n25210 = ~n138 & ~n319;
  assign n25211 = n2107 & n25210;
  assign n25212 = n25209 & n25211;
  assign n25213 = n25208 & n25212;
  assign n25214 = n25207 & n25213;
  assign n25215 = n25203 & n25214;
  assign n25216 = n11581 & n25215;
  assign n25185 = n25052 ^ n25041;
  assign n25186 = n25042 & n25185;
  assign n25217 = n25216 ^ n25186;
  assign n25228 = n25227 ^ n25217;
  assign n25182 = n25061 ^ n25053;
  assign n25183 = ~n25073 & ~n25182;
  assign n25184 = n25183 ^ n25072;
  assign n25229 = n25228 ^ n25184;
  assign n25174 = n44 & n20793;
  assign n25175 = n3280 & n19277;
  assign n25176 = n3277 & n19260;
  assign n25177 = n3275 & ~n19255;
  assign n25178 = ~n25176 & ~n25177;
  assign n25179 = ~n25175 & n25178;
  assign n25180 = ~n25174 & n25179;
  assign n25181 = n25180 ^ x29;
  assign n25230 = n25229 ^ n25181;
  assign n25247 = n25246 ^ n25230;
  assign n25171 = n25074 ^ n25008;
  assign n25172 = ~n25075 & n25171;
  assign n25173 = n25172 ^ n25011;
  assign n25248 = n25247 ^ n25173;
  assign n25257 = n25256 ^ n25248;
  assign n25168 = n25085 ^ n25000;
  assign n25169 = n25077 & n25168;
  assign n25170 = n25169 ^ n25085;
  assign n25258 = n25257 ^ n25170;
  assign n25273 = n25272 ^ n25258;
  assign n25165 = n25095 ^ n24997;
  assign n25166 = n25087 & n25165;
  assign n25167 = n25166 ^ n25095;
  assign n25274 = n25273 ^ n25167;
  assign n25283 = n25282 ^ n25274;
  assign n25162 = n25105 ^ n24994;
  assign n25163 = n25097 & n25162;
  assign n25164 = n25163 ^ n25105;
  assign n25284 = n25283 ^ n25164;
  assign n25301 = n25300 ^ n25284;
  assign n25159 = n24991 ^ n24988;
  assign n25160 = n25107 & n25159;
  assign n25161 = n25160 ^ n24988;
  assign n25302 = n25301 ^ n25161;
  assign n25311 = n25310 ^ n25302;
  assign n25312 = n25311 ^ x8;
  assign n25156 = n25117 ^ n24973;
  assign n25157 = n25109 & n25156;
  assign n25158 = n25157 ^ n25117;
  assign n25313 = n25312 ^ n25158;
  assign n25153 = n25118 ^ n24967;
  assign n25154 = n24970 & ~n25153;
  assign n25155 = n25154 ^ n25118;
  assign n25314 = n25313 ^ n25155;
  assign n25148 = n25138 ^ n25134;
  assign n25150 = n25148 ^ n25119;
  assign n25151 = ~n25145 & ~n25150;
  assign n25149 = ~n25135 & ~n25148;
  assign n25152 = n25151 ^ n25149;
  assign n25315 = n25314 ^ n25152;
  assign n25472 = ~n25119 & ~n25134;
  assign n25473 = ~n25138 & ~n25314;
  assign n25474 = ~n25472 & ~n25473;
  assign n25475 = ~n25138 & ~n25474;
  assign n25476 = n25119 & n25134;
  assign n25477 = ~n25314 & ~n25476;
  assign n25478 = ~n25475 & ~n25477;
  assign n25479 = ~n25474 & n25477;
  assign n25480 = n25145 & ~n25479;
  assign n25481 = ~n25478 & n25480;
  assign n25452 = n24969 & n25118;
  assign n25453 = n24967 & n25138;
  assign n25454 = ~n25313 & ~n25453;
  assign n25455 = ~n25452 & ~n25454;
  assign n25456 = ~n24967 & ~n25138;
  assign n25457 = ~n24969 & ~n25118;
  assign n25458 = ~n25313 & ~n25457;
  assign n25459 = ~n25456 & ~n25458;
  assign n25460 = ~n25455 & ~n25459;
  assign n25461 = ~n25132 & ~n25460;
  assign n25462 = ~n25131 & n25461;
  assign n25463 = n25126 & n25462;
  assign n25464 = n25138 & ~n25452;
  assign n25465 = n25155 & ~n25464;
  assign n25466 = n25313 & ~n25465;
  assign n25467 = n25453 & ~n25458;
  assign n25468 = ~n25466 & ~n25467;
  assign n25469 = ~n25463 & n25468;
  assign n25446 = n5814 & ~n23704;
  assign n25447 = n5817 & n23495;
  assign n25448 = n5824 & ~n23292;
  assign n25449 = ~n25447 & ~n25448;
  assign n25450 = ~n25446 & n25449;
  assign n25451 = n25450 ^ x11;
  assign n25470 = n25469 ^ n25451;
  assign n25441 = n25311 ^ n25158;
  assign n25442 = n25312 & n25441;
  assign n25443 = n25442 ^ x8;
  assign n25438 = n25310 ^ n25161;
  assign n25439 = n25302 & n25438;
  assign n25440 = n25439 ^ n25310;
  assign n25444 = n25443 ^ n25440;
  assign n25420 = n6033 & n23712;
  assign n25421 = ~n5746 & n19649;
  assign n25422 = n5752 & ~n19575;
  assign n25423 = ~n25421 & ~n25422;
  assign n25424 = x14 & n25423;
  assign n25425 = ~n23052 & n25424;
  assign n25426 = ~n25420 & ~n25425;
  assign n25427 = x13 & n25426;
  assign n25428 = ~n23712 & n25424;
  assign n25429 = n6033 & n23052;
  assign n25430 = ~x13 & ~n25429;
  assign n25431 = ~n25428 & n25430;
  assign n25432 = ~n25427 & ~n25431;
  assign n25433 = ~n7589 & n25423;
  assign n25434 = n25433 ^ x14;
  assign n25435 = ~n25432 & n25434;
  assign n25417 = n25300 ^ n25283;
  assign n25418 = n25284 & ~n25417;
  assign n25419 = n25418 ^ n25300;
  assign n25436 = n25435 ^ n25419;
  assign n25407 = n4963 & ~n23064;
  assign n25408 = n4972 & ~n19512;
  assign n25409 = n4976 & n19439;
  assign n25410 = n4970 & ~n19368;
  assign n25411 = ~n25409 & ~n25410;
  assign n25412 = ~n25408 & n25411;
  assign n25413 = ~n25407 & n25412;
  assign n25414 = n25413 ^ x17;
  assign n25397 = n4673 & n22441;
  assign n25398 = n4688 & n19063;
  assign n25399 = ~n4681 & ~n19078;
  assign n25400 = n4685 & n19303;
  assign n25401 = ~n25399 & ~n25400;
  assign n25402 = ~n25398 & n25401;
  assign n25403 = ~n25397 & n25402;
  assign n25404 = n25403 ^ x20;
  assign n25385 = n3285 & n21215;
  assign n25386 = n3437 & n19104;
  assign n25387 = ~n3440 & n19122;
  assign n25388 = n3435 & ~n19286;
  assign n25389 = ~n25387 & ~n25388;
  assign n25390 = ~n25386 & n25389;
  assign n25391 = ~n25385 & n25390;
  assign n25392 = n25391 ^ x26;
  assign n25369 = n20745 & ~n20908;
  assign n25370 = ~n19281 & n20747;
  assign n25371 = n3277 & n19277;
  assign n25372 = n3275 & n19260;
  assign n25373 = ~n25371 & ~n25372;
  assign n25374 = ~n25370 & n25373;
  assign n25375 = ~n25369 & n25374;
  assign n25376 = ~x29 & ~n25375;
  assign n25377 = n20747 & ~n20908;
  assign n25378 = ~n19281 & n20745;
  assign n25379 = x29 & n25373;
  assign n25380 = ~n25378 & n25379;
  assign n25381 = ~n25377 & n25380;
  assign n25382 = ~n25376 & ~n25381;
  assign n25357 = n41 & n19696;
  assign n25358 = n91 & ~n19253;
  assign n25359 = ~n25224 & ~n25358;
  assign n25360 = ~n25357 & n25359;
  assign n25361 = x31 & ~n25360;
  assign n25362 = n41 & ~n19255;
  assign n25363 = n54 & n19253;
  assign n25364 = ~x31 & ~n25363;
  assign n25365 = ~n25362 & n25364;
  assign n25366 = ~n25361 & ~n25365;
  assign n25353 = n25216 ^ n25037;
  assign n25354 = n25042 & ~n25353;
  assign n25355 = n25185 & n25354;
  assign n25356 = n25355 ^ n25037;
  assign n25367 = n25366 ^ n25356;
  assign n25339 = n1767 & n4562;
  assign n25340 = n3035 & n25339;
  assign n25341 = n999 & n3149;
  assign n25342 = n2398 & n25341;
  assign n25343 = n11530 & n11545;
  assign n25344 = n25342 & n25343;
  assign n25345 = n769 & n12872;
  assign n25346 = n247 & n2912;
  assign n25347 = n25345 & n25346;
  assign n25348 = n25344 & n25347;
  assign n25349 = n1204 & n25348;
  assign n25350 = n25340 & n25349;
  assign n25351 = n25350 ^ n25037;
  assign n25352 = n25351 ^ x8;
  assign n25368 = n25367 ^ n25352;
  assign n25383 = n25382 ^ n25368;
  assign n25336 = n25217 ^ n25184;
  assign n25337 = ~n25228 & ~n25336;
  assign n25338 = n25337 ^ n25184;
  assign n25384 = n25383 ^ n25338;
  assign n25393 = n25392 ^ n25384;
  assign n25333 = n25246 ^ n25229;
  assign n25334 = n25230 & ~n25333;
  assign n25335 = n25334 ^ n25246;
  assign n25394 = n25393 ^ n25335;
  assign n25330 = n25256 ^ n25247;
  assign n25331 = n25248 & ~n25330;
  assign n25332 = n25331 ^ n25256;
  assign n25395 = n25394 ^ n25332;
  assign n25322 = n4478 & n19668;
  assign n25323 = n4484 & n19096;
  assign n25324 = n4480 & n19292;
  assign n25325 = ~n25323 & ~n25324;
  assign n25326 = n4487 & n19298;
  assign n25327 = n25325 & ~n25326;
  assign n25328 = ~n25322 & n25327;
  assign n25329 = n25328 ^ x23;
  assign n25396 = n25395 ^ n25329;
  assign n25405 = n25404 ^ n25396;
  assign n25319 = n25272 ^ n25257;
  assign n25320 = n25258 & ~n25319;
  assign n25321 = n25320 ^ n25272;
  assign n25406 = n25405 ^ n25321;
  assign n25415 = n25414 ^ n25406;
  assign n25316 = n25282 ^ n25273;
  assign n25317 = n25274 & ~n25316;
  assign n25318 = n25317 ^ n25282;
  assign n25416 = n25415 ^ n25318;
  assign n25437 = n25436 ^ n25416;
  assign n25445 = n25444 ^ n25437;
  assign n25471 = n25470 ^ n25445;
  assign n25482 = n25481 ^ n25471;
  assign n25614 = n25440 & ~n25443;
  assign n25615 = n25469 & ~n25614;
  assign n25616 = ~n25440 & n25443;
  assign n25617 = ~n25615 & ~n25616;
  assign n25618 = n25451 & n25617;
  assign n25619 = ~n25469 & n25614;
  assign n25620 = ~n25618 & ~n25619;
  assign n25621 = ~n25437 & ~n25620;
  assign n25622 = n25437 & ~n25617;
  assign n25623 = n25469 & n25616;
  assign n25624 = n25451 & ~n25623;
  assign n25625 = n25622 & ~n25624;
  assign n25626 = n25451 & ~n25469;
  assign n25627 = n25614 & n25626;
  assign n25628 = ~n25451 & n25623;
  assign n25629 = ~n25627 & ~n25628;
  assign n25630 = ~n25625 & n25629;
  assign n25631 = ~n25621 & n25630;
  assign n25603 = n6033 & ~n23879;
  assign n25596 = n5752 & n19649;
  assign n25597 = ~n5746 & n23052;
  assign n25598 = ~n25596 & ~n25597;
  assign n25599 = x14 & n25598;
  assign n25604 = n23292 & n25599;
  assign n25605 = ~n25603 & ~n25604;
  assign n25600 = n23879 & n25599;
  assign n25601 = n6033 & ~n23292;
  assign n25602 = ~n25600 & ~n25601;
  assign n25606 = n25605 ^ n25602;
  assign n25607 = ~x13 & n25606;
  assign n25608 = n25607 ^ n25605;
  assign n25609 = ~n7589 & n25598;
  assign n25610 = n25609 ^ x14;
  assign n25611 = n25608 & n25610;
  assign n25586 = n4963 & ~n23468;
  assign n25587 = n4976 & ~n19512;
  assign n25588 = n4970 & n19439;
  assign n25589 = ~n25587 & ~n25588;
  assign n25590 = n4972 & ~n19575;
  assign n25591 = n25589 & ~n25590;
  assign n25592 = ~n25586 & n25591;
  assign n25593 = n25592 ^ x17;
  assign n25576 = n4673 & ~n22037;
  assign n25577 = n4688 & ~n19368;
  assign n25578 = n4685 & n19063;
  assign n25579 = ~n4681 & n19303;
  assign n25580 = ~n25578 & ~n25579;
  assign n25581 = ~n25577 & n25580;
  assign n25582 = ~n25576 & n25581;
  assign n25583 = n25582 ^ x20;
  assign n25566 = n4478 & ~n21715;
  assign n25567 = n4487 & ~n19078;
  assign n25568 = n4480 & n19096;
  assign n25569 = n4484 & n19298;
  assign n25570 = ~n25568 & ~n25569;
  assign n25571 = ~n25567 & n25570;
  assign n25572 = ~n25566 & n25571;
  assign n25573 = n25572 ^ x23;
  assign n25548 = n12417 & n21684;
  assign n25549 = n3435 & n19104;
  assign n25550 = ~n3440 & ~n19286;
  assign n25551 = ~n25549 & ~n25550;
  assign n25552 = x26 & n25551;
  assign n25553 = ~n19292 & n25552;
  assign n25554 = ~n25548 & ~n25553;
  assign n25555 = x25 & n25554;
  assign n25556 = ~n21684 & n25552;
  assign n25557 = n12417 & n19292;
  assign n25558 = ~x25 & ~n25557;
  assign n25559 = ~n25556 & n25558;
  assign n25560 = ~n25555 & ~n25559;
  assign n25561 = ~n12432 & n25551;
  assign n25562 = n25561 ^ x26;
  assign n25563 = ~n25560 & n25562;
  assign n25538 = n44 & n21189;
  assign n25539 = n3280 & n19122;
  assign n25540 = n3277 & ~n19281;
  assign n25541 = n3275 & n19277;
  assign n25542 = ~n25540 & ~n25541;
  assign n25543 = ~n25539 & n25542;
  assign n25544 = ~n25538 & n25543;
  assign n25545 = n25544 ^ x29;
  assign n25525 = n41 & ~n20929;
  assign n25526 = n91 & n19255;
  assign n25527 = n54 & ~n19253;
  assign n25528 = x31 & ~n25527;
  assign n25529 = ~n25526 & n25528;
  assign n25530 = ~n25525 & n25529;
  assign n25531 = ~n54 & ~n19260;
  assign n25532 = n54 & n19255;
  assign n25533 = n3640 & ~n25532;
  assign n25534 = ~n25531 & n25533;
  assign n25535 = ~n25530 & ~n25534;
  assign n25511 = n1001 & n2595;
  assign n25512 = n12225 & n25012;
  assign n25513 = n25511 & n25512;
  assign n25514 = ~n238 & ~n919;
  assign n25515 = ~n174 & ~n929;
  assign n25516 = n25514 & n25515;
  assign n25517 = n4740 & n25516;
  assign n25518 = n25513 & n25517;
  assign n25519 = n4799 & n12136;
  assign n25520 = n25518 & n25519;
  assign n25521 = n10105 & n25520;
  assign n25522 = n3079 & n25521;
  assign n25523 = n2111 & n25522;
  assign n25508 = n25037 ^ x8;
  assign n25509 = ~n25351 & n25508;
  assign n25510 = n25509 ^ x8;
  assign n25524 = n25523 ^ n25510;
  assign n25536 = n25535 ^ n25524;
  assign n25505 = n25356 ^ n25352;
  assign n25506 = n25367 & n25505;
  assign n25507 = n25506 ^ n25366;
  assign n25537 = n25536 ^ n25507;
  assign n25546 = n25545 ^ n25537;
  assign n25502 = n25382 ^ n25338;
  assign n25503 = ~n25383 & ~n25502;
  assign n25504 = n25503 ^ n25338;
  assign n25547 = n25546 ^ n25504;
  assign n25564 = n25563 ^ n25547;
  assign n25499 = n25392 ^ n25335;
  assign n25500 = n25393 & n25499;
  assign n25501 = n25500 ^ n25335;
  assign n25565 = n25564 ^ n25501;
  assign n25574 = n25573 ^ n25565;
  assign n25496 = n25394 ^ n25329;
  assign n25497 = ~n25395 & n25496;
  assign n25498 = n25497 ^ n25332;
  assign n25575 = n25574 ^ n25498;
  assign n25584 = n25583 ^ n25575;
  assign n25493 = n25404 ^ n25321;
  assign n25494 = n25405 & n25493;
  assign n25495 = n25494 ^ n25321;
  assign n25585 = n25584 ^ n25495;
  assign n25594 = n25593 ^ n25585;
  assign n25490 = n25406 ^ n25318;
  assign n25491 = ~n25415 & n25490;
  assign n25492 = n25491 ^ n25414;
  assign n25595 = n25594 ^ n25492;
  assign n25612 = n25611 ^ n25595;
  assign n25487 = n5824 & n23495;
  assign n25488 = n25487 ^ x11;
  assign n25484 = n25419 ^ n25416;
  assign n25485 = n25436 & n25484;
  assign n25486 = n25485 ^ n25435;
  assign n25489 = n25488 ^ n25486;
  assign n25613 = n25612 ^ n25489;
  assign n25632 = n25631 ^ n25613;
  assign n25483 = n25471 & n25481;
  assign n25633 = n25632 ^ n25483;
  assign n25780 = n25483 & ~n25632;
  assign n25764 = n25440 ^ n25437;
  assign n25765 = n25613 ^ n25437;
  assign n25766 = n25764 & ~n25765;
  assign n25767 = n25444 & n25766;
  assign n25768 = n25767 ^ n25613;
  assign n25769 = ~n25626 & ~n25768;
  assign n25770 = n25437 & ~n25614;
  assign n25771 = ~n25616 & ~n25770;
  assign n25772 = ~n25613 & ~n25771;
  assign n25773 = ~n25769 & ~n25772;
  assign n25774 = ~n25451 & n25469;
  assign n25775 = n25613 & ~n25770;
  assign n25776 = n25774 & ~n25775;
  assign n25777 = ~n25628 & ~n25776;
  assign n25778 = n25773 & n25777;
  assign n25759 = n25612 ^ n25486;
  assign n25760 = n25489 & ~n25759;
  assign n25761 = n25760 ^ n25612;
  assign n25756 = n25611 ^ n25492;
  assign n25757 = n25595 & n25756;
  assign n25758 = n25757 ^ n25611;
  assign n25762 = n25761 ^ n25758;
  assign n25739 = n5796 & n23493;
  assign n25740 = ~n5746 & ~n23292;
  assign n25741 = n5752 & n23052;
  assign n25742 = ~n25740 & ~n25741;
  assign n25743 = ~n25739 & n25742;
  assign n25744 = ~x13 & n23495;
  assign n25745 = n5748 & n25744;
  assign n25746 = n25743 & ~n25745;
  assign n25747 = ~x14 & ~n25746;
  assign n25748 = n13989 & ~n23493;
  assign n25749 = n14928 & ~n23495;
  assign n25750 = ~n7559 & ~n25749;
  assign n25751 = ~n25748 & n25750;
  assign n25752 = n25742 & ~n25751;
  assign n25753 = ~n25747 & ~n25752;
  assign n25721 = n5771 & n23520;
  assign n25722 = n4970 & ~n19512;
  assign n25723 = n4976 & ~n19575;
  assign n25724 = ~n25722 & ~n25723;
  assign n25725 = x17 & n25724;
  assign n25726 = ~n19649 & n25725;
  assign n25727 = x16 & ~n25726;
  assign n25728 = ~n25721 & n25727;
  assign n25729 = ~n23520 & n25725;
  assign n25730 = n5771 & n19649;
  assign n25731 = ~x16 & ~n25730;
  assign n25732 = ~n25729 & n25731;
  assign n25733 = ~n25728 & ~n25732;
  assign n25734 = ~n5786 & n25724;
  assign n25735 = n25734 ^ x17;
  assign n25736 = ~n25733 & n25735;
  assign n25711 = n4673 & n22457;
  assign n25712 = n4688 & n19439;
  assign n25713 = n4685 & ~n19368;
  assign n25714 = ~n4681 & n19063;
  assign n25715 = ~n25713 & ~n25714;
  assign n25716 = ~n25712 & n25715;
  assign n25717 = ~n25711 & n25716;
  assign n25718 = n25717 ^ x20;
  assign n25701 = n4478 & n19658;
  assign n25702 = n4484 & ~n19078;
  assign n25703 = n4487 & n19303;
  assign n25704 = n4480 & n19298;
  assign n25705 = ~n25703 & ~n25704;
  assign n25706 = ~n25702 & n25705;
  assign n25707 = ~n25701 & n25706;
  assign n25708 = n25707 ^ x23;
  assign n25691 = n3285 & n21699;
  assign n25692 = n3437 & n19096;
  assign n25693 = n3435 & n19292;
  assign n25694 = ~n3440 & n19104;
  assign n25695 = ~n25693 & ~n25694;
  assign n25696 = ~n25692 & n25695;
  assign n25697 = ~n25691 & n25696;
  assign n25698 = n25697 ^ x26;
  assign n25681 = n44 & ~n19678;
  assign n25682 = n3277 & n19122;
  assign n25683 = n3280 & ~n19286;
  assign n25684 = n3275 & ~n19281;
  assign n25685 = ~n25683 & ~n25684;
  assign n25686 = ~n25682 & n25685;
  assign n25687 = ~n25681 & n25686;
  assign n25688 = n25687 ^ x29;
  assign n25664 = n676 & n1787;
  assign n25665 = n2435 & n25664;
  assign n25666 = ~n110 & ~n216;
  assign n25667 = n1124 & n25666;
  assign n25668 = n25665 & n25667;
  assign n25669 = n223 & n12301;
  assign n25670 = n25668 & n25669;
  assign n25671 = n1586 & n2466;
  assign n25672 = n4774 & n10208;
  assign n25673 = n25671 & n25672;
  assign n25674 = n25670 & n25673;
  assign n25675 = n11541 & n12854;
  assign n25676 = n25674 & n25675;
  assign n25677 = n25035 & n25676;
  assign n25678 = n4247 & n25677;
  assign n25660 = n25510 & n25535;
  assign n25659 = ~n25510 & ~n25535;
  assign n25661 = n25660 ^ n25659;
  assign n25662 = ~n25523 & n25661;
  assign n25663 = n25662 ^ n25660;
  assign n25679 = n25678 ^ n25663;
  assign n25652 = n41 & ~n20793;
  assign n25653 = n91 & ~n19260;
  assign n25654 = ~n25532 & ~n25653;
  assign n25655 = ~n25652 & n25654;
  assign n25649 = n41 & n19277;
  assign n25650 = n54 & n19260;
  assign n25651 = ~n25649 & ~n25650;
  assign n25656 = n25655 ^ n25651;
  assign n25657 = ~x31 & ~n25656;
  assign n25658 = n25657 ^ n25655;
  assign n25680 = n25679 ^ n25658;
  assign n25689 = n25688 ^ n25680;
  assign n25646 = n25545 ^ n25507;
  assign n25647 = ~n25537 & ~n25646;
  assign n25648 = n25647 ^ n25545;
  assign n25690 = n25689 ^ n25648;
  assign n25699 = n25698 ^ n25690;
  assign n25643 = n25563 ^ n25504;
  assign n25644 = n25547 & ~n25643;
  assign n25645 = n25644 ^ n25563;
  assign n25700 = n25699 ^ n25645;
  assign n25709 = n25708 ^ n25700;
  assign n25640 = n25573 ^ n25501;
  assign n25641 = n25565 & n25640;
  assign n25642 = n25641 ^ n25573;
  assign n25710 = n25709 ^ n25642;
  assign n25719 = n25718 ^ n25710;
  assign n25637 = n25583 ^ n25574;
  assign n25638 = n25575 & ~n25637;
  assign n25639 = n25638 ^ n25583;
  assign n25720 = n25719 ^ n25639;
  assign n25737 = n25736 ^ n25720;
  assign n25634 = n25593 ^ n25495;
  assign n25635 = n25585 & n25634;
  assign n25636 = n25635 ^ n25593;
  assign n25738 = n25737 ^ n25636;
  assign n25754 = n25753 ^ n25738;
  assign n25755 = n25754 ^ x11;
  assign n25763 = n25762 ^ n25755;
  assign n25779 = n25778 ^ n25763;
  assign n25781 = n25780 ^ n25779;
  assign n25907 = ~n25754 & n25778;
  assign n25908 = n25758 & n25907;
  assign n25909 = n25761 & ~n25908;
  assign n25910 = n25778 ^ n25758;
  assign n25911 = n25758 ^ n25754;
  assign n25912 = n25910 & n25911;
  assign n25913 = n25912 ^ n25778;
  assign n25914 = ~n25909 & n25913;
  assign n25915 = ~x11 & ~n25914;
  assign n25916 = n25761 & ~n25913;
  assign n25917 = n25754 & ~n25778;
  assign n25918 = ~n25758 & n25917;
  assign n25919 = x11 & ~n25918;
  assign n25920 = ~n25916 & n25919;
  assign n25921 = ~n25915 & ~n25920;
  assign n25922 = ~n25908 & ~n25918;
  assign n25923 = n25762 & ~n25922;
  assign n25924 = ~n25921 & ~n25923;
  assign n25890 = n5796 & ~n23704;
  assign n25891 = n13719 & ~n23292;
  assign n25892 = ~n25744 & ~n25891;
  assign n25893 = n5742 & ~n25892;
  assign n25894 = ~n13989 & ~n23495;
  assign n25895 = ~x13 & n23292;
  assign n25896 = n5744 & ~n25895;
  assign n25897 = ~n25894 & n25896;
  assign n25898 = ~n25893 & ~n25897;
  assign n25899 = n25898 ^ x14;
  assign n25900 = n5748 & ~n23704;
  assign n25901 = n25898 & n25900;
  assign n25902 = ~n25899 & n25901;
  assign n25903 = n25902 ^ n25899;
  assign n25904 = ~n25890 & n25903;
  assign n25880 = n4963 & n23712;
  assign n25881 = n4976 & n19649;
  assign n25882 = n4970 & ~n19575;
  assign n25883 = ~n25881 & ~n25882;
  assign n25884 = n4972 & n23052;
  assign n25885 = n25883 & ~n25884;
  assign n25886 = ~n25880 & n25885;
  assign n25887 = n25886 ^ x17;
  assign n25870 = n4673 & ~n23064;
  assign n25871 = n4688 & ~n19512;
  assign n25872 = n4685 & n19439;
  assign n25873 = ~n4681 & ~n19368;
  assign n25874 = ~n25872 & ~n25873;
  assign n25875 = ~n25871 & n25874;
  assign n25876 = ~n25870 & n25875;
  assign n25877 = n25876 ^ x20;
  assign n25867 = n25718 ^ n25709;
  assign n25868 = n25710 & ~n25867;
  assign n25869 = n25868 ^ n25718;
  assign n25878 = n25877 ^ n25869;
  assign n25857 = n4478 & n22441;
  assign n25858 = n4487 & n19063;
  assign n25859 = n4480 & ~n19078;
  assign n25860 = n4484 & n19303;
  assign n25861 = ~n25859 & ~n25860;
  assign n25862 = ~n25858 & n25861;
  assign n25863 = ~n25857 & n25862;
  assign n25864 = n25863 ^ x23;
  assign n25847 = n3285 & n19668;
  assign n25848 = n3435 & n19096;
  assign n25849 = ~n3440 & n19292;
  assign n25850 = ~n25848 & ~n25849;
  assign n25851 = n3437 & n19298;
  assign n25852 = n25850 & ~n25851;
  assign n25853 = ~n25847 & n25852;
  assign n25854 = n25853 ^ x26;
  assign n25831 = ~x28 & n21214;
  assign n25832 = n25831 ^ n19104;
  assign n25833 = n42 & n25832;
  assign n25834 = n3275 & n19122;
  assign n25835 = n3277 & ~n19286;
  assign n25836 = ~n25834 & ~n25835;
  assign n25837 = x29 & n25836;
  assign n25838 = ~n25833 & n25837;
  assign n25839 = x28 & ~n21215;
  assign n25840 = ~x28 & ~n19104;
  assign n25841 = n12466 & ~n25840;
  assign n25842 = ~n25839 & n25841;
  assign n25843 = ~x29 & ~n25836;
  assign n25844 = ~n25842 & ~n25843;
  assign n25845 = ~n25838 & n25844;
  assign n25818 = n41 & ~n20908;
  assign n25819 = n91 & n19277;
  assign n25820 = x31 & ~n25650;
  assign n25821 = ~n25819 & n25820;
  assign n25822 = ~n25818 & n25821;
  assign n25823 = n41 & ~n19281;
  assign n25824 = n54 & n19277;
  assign n25825 = ~x31 & ~n25824;
  assign n25826 = ~n25823 & n25825;
  assign n25827 = ~n25822 & ~n25826;
  assign n25803 = n1785 & n11293;
  assign n25804 = n4066 & n25803;
  assign n25805 = n3290 & n25804;
  assign n25806 = n2894 & n25805;
  assign n25807 = ~n256 & ~n298;
  assign n25808 = n11388 & n25807;
  assign n25809 = n25190 & n25808;
  assign n25810 = n252 & n2022;
  assign n25811 = n25809 & n25810;
  assign n25812 = n1618 & n4097;
  assign n25813 = n25811 & n25812;
  assign n25814 = n1559 & n25813;
  assign n25815 = n2421 & n25814;
  assign n25816 = n25806 & n25815;
  assign n25817 = n25816 ^ x11;
  assign n25828 = n25827 ^ n25817;
  assign n25799 = n25659 & ~n25678;
  assign n25798 = n25660 & n25678;
  assign n25800 = n25799 ^ n25798;
  assign n25801 = n25523 & n25800;
  assign n25802 = n25801 ^ n25799;
  assign n25829 = n25828 ^ n25802;
  assign n25795 = n25688 ^ n25679;
  assign n25796 = n25680 & n25795;
  assign n25797 = n25796 ^ n25688;
  assign n25830 = n25829 ^ n25797;
  assign n25846 = n25845 ^ n25830;
  assign n25855 = n25854 ^ n25846;
  assign n25792 = n25698 ^ n25689;
  assign n25793 = n25690 & ~n25792;
  assign n25794 = n25793 ^ n25698;
  assign n25856 = n25855 ^ n25794;
  assign n25865 = n25864 ^ n25856;
  assign n25789 = n25708 ^ n25699;
  assign n25790 = n25700 & ~n25789;
  assign n25791 = n25790 ^ n25708;
  assign n25866 = n25865 ^ n25791;
  assign n25879 = n25878 ^ n25866;
  assign n25888 = n25887 ^ n25879;
  assign n25786 = n25736 ^ n25719;
  assign n25787 = n25720 & ~n25786;
  assign n25788 = n25787 ^ n25736;
  assign n25889 = n25888 ^ n25788;
  assign n25905 = n25904 ^ n25889;
  assign n25783 = n25753 ^ n25737;
  assign n25784 = n25738 & ~n25783;
  assign n25785 = n25784 ^ n25753;
  assign n25906 = n25905 ^ n25785;
  assign n25925 = n25924 ^ n25906;
  assign n25782 = n25779 & n25780;
  assign n25926 = n25925 ^ n25782;
  assign n26055 = n25782 & ~n25925;
  assign n26039 = n25761 ^ x11;
  assign n26040 = n25906 ^ n25758;
  assign n26041 = n25762 & n26040;
  assign n26042 = ~n26039 & n26041;
  assign n26043 = n26042 ^ n25906;
  assign n26044 = ~n25917 & n26043;
  assign n26045 = n25907 ^ n25906;
  assign n26046 = n25758 & ~n25761;
  assign n26047 = x11 & ~n26046;
  assign n26048 = ~n25758 & n25761;
  assign n26049 = ~n26047 & ~n26048;
  assign n26050 = n26049 ^ n25906;
  assign n26051 = n26045 & ~n26050;
  assign n26052 = n26051 ^ n25907;
  assign n26053 = ~n26044 & ~n26052;
  assign n26027 = n4963 & ~n23879;
  assign n26028 = n4972 & ~n23292;
  assign n26029 = n4976 & n23052;
  assign n26030 = n4970 & n19649;
  assign n26031 = ~n26029 & ~n26030;
  assign n26032 = ~n26028 & n26031;
  assign n26033 = ~n26027 & n26032;
  assign n26034 = n26033 ^ x17;
  assign n26017 = n4673 & ~n23468;
  assign n26018 = n4685 & ~n19512;
  assign n26019 = ~n4681 & n19439;
  assign n26020 = ~n26018 & ~n26019;
  assign n26021 = n4688 & ~n19575;
  assign n26022 = n26020 & ~n26021;
  assign n26023 = ~n26017 & n26022;
  assign n26024 = n26023 ^ x20;
  assign n26007 = n4478 & ~n22037;
  assign n26008 = n4487 & ~n19368;
  assign n26009 = n4484 & n19063;
  assign n26010 = n4480 & n19303;
  assign n26011 = ~n26009 & ~n26010;
  assign n26012 = ~n26008 & n26011;
  assign n26013 = ~n26007 & n26012;
  assign n26014 = n26013 ^ x23;
  assign n25997 = n3285 & ~n21715;
  assign n25998 = n3437 & ~n19078;
  assign n25999 = n3435 & n19298;
  assign n26000 = ~n3440 & n19096;
  assign n26001 = ~n25999 & ~n26000;
  assign n26002 = ~n25998 & n26001;
  assign n26003 = ~n25997 & n26002;
  assign n26004 = n26003 ^ x26;
  assign n25987 = n44 & n21684;
  assign n25988 = n3280 & n19292;
  assign n25989 = n3277 & n19104;
  assign n25990 = n3275 & ~n19286;
  assign n25991 = ~n25989 & ~n25990;
  assign n25992 = ~n25988 & n25991;
  assign n25993 = ~n25987 & n25992;
  assign n25994 = n25993 ^ x29;
  assign n25976 = n41 & n21189;
  assign n25977 = n91 & ~n19281;
  assign n25978 = ~n25824 & ~n25977;
  assign n25979 = ~n25976 & n25978;
  assign n25980 = x31 & ~n25979;
  assign n25981 = n3676 & n19122;
  assign n25982 = n3671 & ~n19281;
  assign n25983 = ~n25981 & ~n25982;
  assign n25984 = ~n25980 & n25983;
  assign n25962 = ~n659 & n806;
  assign n25963 = n1021 & n4424;
  assign n25964 = n25962 & n25963;
  assign n25965 = n11039 & n25964;
  assign n25966 = n12856 & n25965;
  assign n25967 = ~n527 & n834;
  assign n25968 = n786 & n1825;
  assign n25969 = n25967 & n25968;
  assign n25970 = n3362 & n25969;
  assign n25971 = n24179 & n25970;
  assign n25972 = n23812 & n25971;
  assign n25973 = n11076 & n25972;
  assign n25974 = n25966 & n25973;
  assign n25958 = n25523 ^ x11;
  assign n25959 = n25816 ^ n25523;
  assign n25960 = n25958 & ~n25959;
  assign n25961 = n25960 ^ x11;
  assign n25975 = n25974 ^ n25961;
  assign n25985 = n25984 ^ n25975;
  assign n25947 = n25817 & n25827;
  assign n25948 = n25798 & ~n25947;
  assign n25949 = ~n25817 & ~n25827;
  assign n25950 = n25523 & ~n25949;
  assign n25951 = ~n25948 & n25950;
  assign n25952 = n25827 ^ n25799;
  assign n25953 = ~n25523 & ~n25817;
  assign n25954 = n25953 ^ n25827;
  assign n25955 = n25952 & ~n25954;
  assign n25956 = n25955 ^ n25799;
  assign n25957 = ~n25951 & ~n25956;
  assign n25986 = n25985 ^ n25957;
  assign n25995 = n25994 ^ n25986;
  assign n25944 = n25845 ^ n25797;
  assign n25945 = ~n25830 & n25944;
  assign n25946 = n25945 ^ n25845;
  assign n25996 = n25995 ^ n25946;
  assign n26005 = n26004 ^ n25996;
  assign n25941 = n25846 ^ n25794;
  assign n25942 = n25855 & ~n25941;
  assign n25943 = n25942 ^ n25854;
  assign n26006 = n26005 ^ n25943;
  assign n26015 = n26014 ^ n26006;
  assign n25938 = n25864 ^ n25791;
  assign n25939 = ~n25865 & n25938;
  assign n25940 = n25939 ^ n25791;
  assign n26016 = n26015 ^ n25940;
  assign n26025 = n26024 ^ n26016;
  assign n25935 = n25869 ^ n25866;
  assign n25936 = n25878 & ~n25935;
  assign n25937 = n25936 ^ n25877;
  assign n26026 = n26025 ^ n25937;
  assign n26035 = n26034 ^ n26026;
  assign n25933 = n5752 & n23495;
  assign n25934 = n25933 ^ x14;
  assign n26036 = n26035 ^ n25934;
  assign n25930 = n25887 ^ n25788;
  assign n25931 = ~n25888 & n25930;
  assign n25932 = n25931 ^ n25788;
  assign n26037 = n26036 ^ n25932;
  assign n25927 = n25904 ^ n25785;
  assign n25928 = ~n25905 & n25927;
  assign n25929 = n25928 ^ n25785;
  assign n26038 = n26037 ^ n25929;
  assign n26054 = n26053 ^ n26038;
  assign n26056 = n26055 ^ n26054;
  assign n26187 = n26054 & n26055;
  assign n26184 = n26035 ^ n25932;
  assign n26185 = ~n26036 & ~n26184;
  assign n26186 = n26185 ^ n25932;
  assign n26188 = n26187 ^ n26186;
  assign n26172 = n4963 & n23493;
  assign n26173 = n4972 & n23495;
  assign n26174 = n4976 & ~n23292;
  assign n26175 = n4970 & n23052;
  assign n26176 = ~n26174 & ~n26175;
  assign n26177 = ~n26173 & n26176;
  assign n26178 = ~n26172 & n26177;
  assign n26179 = n26178 ^ x17;
  assign n26154 = n13653 & n23520;
  assign n26155 = ~n4681 & ~n19512;
  assign n26156 = n4685 & ~n19575;
  assign n26157 = ~n26155 & ~n26156;
  assign n26158 = x20 & n26157;
  assign n26159 = ~n19649 & n26158;
  assign n26160 = x19 & ~n26159;
  assign n26161 = ~n26154 & n26160;
  assign n26162 = ~n23520 & n26158;
  assign n26163 = n13653 & n19649;
  assign n26164 = ~x19 & ~n26163;
  assign n26165 = ~n26162 & n26164;
  assign n26166 = ~n26161 & ~n26165;
  assign n26167 = ~n13668 & n26157;
  assign n26168 = n26167 ^ x20;
  assign n26169 = ~n26166 & n26168;
  assign n26136 = n12502 & n22457;
  assign n26137 = n4484 & ~n19368;
  assign n26138 = n4480 & n19063;
  assign n26139 = ~n26137 & ~n26138;
  assign n26140 = x23 & n26139;
  assign n26141 = ~n19439 & n26140;
  assign n26142 = x22 & ~n26141;
  assign n26143 = ~n26136 & n26142;
  assign n26144 = ~n22457 & n26140;
  assign n26145 = n12502 & n19439;
  assign n26146 = ~x22 & ~n26145;
  assign n26147 = ~n26144 & n26146;
  assign n26148 = ~n26143 & ~n26147;
  assign n26149 = ~n12519 & n26139;
  assign n26150 = n26149 ^ x23;
  assign n26151 = ~n26148 & n26150;
  assign n26126 = n3285 & n19658;
  assign n26127 = n3435 & ~n19078;
  assign n26128 = n3437 & n19303;
  assign n26129 = ~n3440 & n19298;
  assign n26130 = ~n26128 & ~n26129;
  assign n26131 = ~n26127 & n26130;
  assign n26132 = ~n26126 & n26131;
  assign n26133 = n26132 ^ x26;
  assign n26106 = n25994 ^ n25961;
  assign n26107 = n25961 ^ n25957;
  assign n26108 = n26106 & ~n26107;
  assign n26109 = n26108 ^ n25994;
  assign n26110 = n25974 & ~n26109;
  assign n26111 = ~n25957 & ~n25994;
  assign n26112 = ~n25961 & n26111;
  assign n26113 = ~n25984 & ~n26112;
  assign n26114 = ~n26110 & n26113;
  assign n26115 = ~n25974 & n26109;
  assign n26116 = n25957 & n25994;
  assign n26117 = n25961 & n26116;
  assign n26118 = n25984 & ~n26117;
  assign n26119 = ~n26115 & n26118;
  assign n26120 = ~n26114 & ~n26119;
  assign n26121 = ~n26112 & ~n26117;
  assign n26122 = n25975 & ~n26121;
  assign n26123 = ~n26120 & ~n26122;
  assign n26093 = n41 & n19678;
  assign n26094 = n91 & ~n19122;
  assign n26095 = n54 & n19281;
  assign n26096 = x31 & ~n26095;
  assign n26097 = ~n26094 & n26096;
  assign n26098 = ~n26093 & n26097;
  assign n26099 = n54 & ~n19122;
  assign n26100 = ~x31 & ~n26099;
  assign n26101 = ~n91 & ~n19286;
  assign n26102 = ~n54 & ~n26101;
  assign n26103 = n26100 & ~n26102;
  assign n26104 = ~n26098 & ~n26103;
  assign n26080 = n3133 & n11386;
  assign n26081 = n4129 & n26080;
  assign n26082 = n2771 & n2936;
  assign n26083 = n1377 & n2292;
  assign n26084 = n26082 & n26083;
  assign n26085 = n2240 & n11276;
  assign n26086 = n26084 & n26085;
  assign n26087 = n1612 & n10900;
  assign n26088 = n26086 & n26087;
  assign n26089 = n941 & n26088;
  assign n26090 = n26081 & n26089;
  assign n26091 = n11638 & n26090;
  assign n26092 = n26091 ^ n25974;
  assign n26105 = n26104 ^ n26092;
  assign n26124 = n26123 ^ n26105;
  assign n26072 = n44 & n21699;
  assign n26073 = n3280 & n19096;
  assign n26074 = n3277 & n19292;
  assign n26075 = n3275 & n19104;
  assign n26076 = ~n26074 & ~n26075;
  assign n26077 = ~n26073 & n26076;
  assign n26078 = ~n26072 & n26077;
  assign n26079 = n26078 ^ x29;
  assign n26125 = n26124 ^ n26079;
  assign n26134 = n26133 ^ n26125;
  assign n26069 = n26004 ^ n25946;
  assign n26070 = n25996 & n26069;
  assign n26071 = n26070 ^ n26004;
  assign n26135 = n26134 ^ n26071;
  assign n26152 = n26151 ^ n26135;
  assign n26066 = n26014 ^ n26005;
  assign n26067 = n26006 & ~n26066;
  assign n26068 = n26067 ^ n26014;
  assign n26153 = n26152 ^ n26068;
  assign n26170 = n26169 ^ n26153;
  assign n26063 = n26024 ^ n25940;
  assign n26064 = n26016 & n26063;
  assign n26065 = n26064 ^ n26024;
  assign n26171 = n26170 ^ n26065;
  assign n26180 = n26179 ^ n26171;
  assign n26060 = n26034 ^ n25937;
  assign n26061 = n26026 & n26060;
  assign n26062 = n26061 ^ n26034;
  assign n26181 = n26180 ^ n26062;
  assign n26182 = n26181 ^ x14;
  assign n26057 = n26053 ^ n25929;
  assign n26058 = ~n26038 & ~n26057;
  assign n26059 = n26058 ^ n26053;
  assign n26183 = n26182 ^ n26059;
  assign n26189 = n26188 ^ n26183;
  assign n26292 = n4963 & ~n23704;
  assign n26293 = n4976 & n23495;
  assign n26294 = n4970 & ~n23292;
  assign n26295 = ~n26293 & ~n26294;
  assign n26296 = ~n26292 & n26295;
  assign n26297 = n26296 ^ x17;
  assign n26282 = n4673 & n23712;
  assign n26283 = n4685 & n19649;
  assign n26284 = ~n4681 & ~n19575;
  assign n26285 = ~n26283 & ~n26284;
  assign n26286 = n4688 & n23052;
  assign n26287 = n26285 & ~n26286;
  assign n26288 = ~n26282 & n26287;
  assign n26289 = n26288 ^ x20;
  assign n26273 = n4478 & ~n23064;
  assign n26274 = n4487 & ~n19512;
  assign n26275 = n4484 & n19439;
  assign n26276 = n4480 & ~n19368;
  assign n26277 = ~n26275 & ~n26276;
  assign n26278 = ~n26274 & n26277;
  assign n26279 = ~n26273 & n26278;
  assign n26280 = n26279 ^ x23;
  assign n26261 = n44 & n19668;
  assign n26262 = n3277 & n19096;
  assign n26263 = n3275 & n19292;
  assign n26264 = ~n26262 & ~n26263;
  assign n26265 = n3280 & n19298;
  assign n26266 = n26264 & ~n26265;
  assign n26267 = ~n26261 & n26266;
  assign n26268 = n26267 ^ x29;
  assign n26245 = n25961 & ~n25974;
  assign n26246 = n25984 & n26245;
  assign n26247 = ~n26116 & ~n26246;
  assign n26248 = n25984 ^ n25961;
  assign n26249 = n25975 & n26248;
  assign n26250 = n26249 ^ n25984;
  assign n26251 = ~n26247 & n26250;
  assign n26252 = n26105 & ~n26251;
  assign n26253 = ~n26105 & n26250;
  assign n26254 = n26111 & ~n26253;
  assign n26255 = ~n25961 & n25974;
  assign n26256 = ~n25984 & n26255;
  assign n26257 = ~n26116 & n26256;
  assign n26258 = ~n26254 & ~n26257;
  assign n26259 = ~n26252 & n26258;
  assign n26234 = n41 & ~n21215;
  assign n26235 = x31 & ~n19286;
  assign n26236 = ~n11234 & ~n26235;
  assign n26237 = ~n26099 & ~n26236;
  assign n26238 = ~n26234 & n26237;
  assign n26239 = n3676 & n19104;
  assign n26240 = n3671 & ~n19286;
  assign n26241 = ~n26239 & ~n26240;
  assign n26242 = ~n26238 & n26241;
  assign n26221 = ~n83 & ~n134;
  assign n26222 = ~n518 & n26221;
  assign n26223 = n1567 & n3594;
  assign n26224 = n26222 & n26223;
  assign n26225 = n2180 & n26224;
  assign n26226 = n980 & n12294;
  assign n26227 = n26225 & n26226;
  assign n26228 = n2642 & n4727;
  assign n26229 = n26227 & n26228;
  assign n26230 = n5607 & n26229;
  assign n26231 = n12080 & n26230;
  assign n26232 = n2481 & n26231;
  assign n26233 = n26232 ^ x14;
  assign n26243 = n26242 ^ n26233;
  assign n26218 = n26104 ^ n25974;
  assign n26219 = n26104 ^ n26091;
  assign n26220 = ~n26218 & ~n26219;
  assign n26244 = n26243 ^ n26220;
  assign n26260 = n26259 ^ n26244;
  assign n26269 = n26268 ^ n26260;
  assign n26215 = n26133 ^ n26124;
  assign n26216 = n26125 & ~n26215;
  assign n26217 = n26216 ^ n26133;
  assign n26270 = n26269 ^ n26217;
  assign n26207 = n3285 & n22441;
  assign n26208 = n3437 & n19063;
  assign n26209 = ~n3440 & ~n19078;
  assign n26210 = n3435 & n19303;
  assign n26211 = ~n26209 & ~n26210;
  assign n26212 = ~n26208 & n26211;
  assign n26213 = ~n26207 & n26212;
  assign n26214 = n26213 ^ x26;
  assign n26271 = n26270 ^ n26214;
  assign n26204 = n26151 ^ n26134;
  assign n26205 = n26135 & ~n26204;
  assign n26206 = n26205 ^ n26151;
  assign n26272 = n26271 ^ n26206;
  assign n26281 = n26280 ^ n26272;
  assign n26290 = n26289 ^ n26281;
  assign n26201 = n26169 ^ n26152;
  assign n26202 = n26153 & ~n26201;
  assign n26203 = n26202 ^ n26169;
  assign n26291 = n26290 ^ n26203;
  assign n26298 = n26297 ^ n26291;
  assign n26198 = n26179 ^ n26170;
  assign n26199 = n26171 & ~n26198;
  assign n26200 = n26199 ^ n26179;
  assign n26299 = n26298 ^ n26200;
  assign n26195 = n26180 ^ x14;
  assign n26196 = n26181 & n26195;
  assign n26197 = n26196 ^ x14;
  assign n26300 = n26299 ^ n26197;
  assign n26190 = n26186 ^ n26059;
  assign n26192 = n26190 ^ n26182;
  assign n26193 = ~n26187 & n26192;
  assign n26191 = n26183 & n26190;
  assign n26194 = n26193 ^ n26191;
  assign n26301 = n26300 ^ n26194;
  assign n26427 = n26059 & ~n26182;
  assign n26428 = ~n26300 & ~n26427;
  assign n26429 = ~n26059 & n26182;
  assign n26430 = ~n26186 & n26300;
  assign n26431 = ~n26429 & n26430;
  assign n26432 = ~n26428 & ~n26431;
  assign n26433 = n26183 & n26186;
  assign n26434 = n26432 & ~n26433;
  assign n26435 = n26187 & n26434;
  assign n26407 = ~n26180 & n26186;
  assign n26408 = x14 & ~n26407;
  assign n26409 = n26180 & ~n26186;
  assign n26410 = ~n26408 & ~n26409;
  assign n26411 = n26299 & ~n26410;
  assign n26412 = n26062 & ~n26411;
  assign n26413 = n26186 ^ x14;
  assign n26414 = n26186 ^ n26180;
  assign n26415 = n26299 ^ n26180;
  assign n26416 = n26414 & n26415;
  assign n26417 = n26413 & n26416;
  assign n26418 = n26417 ^ n26299;
  assign n26419 = ~n26412 & n26418;
  assign n26420 = ~n26059 & ~n26419;
  assign n26421 = n26062 & ~n26418;
  assign n26422 = ~n26299 & n26410;
  assign n26423 = ~n26421 & ~n26422;
  assign n26424 = ~n26420 & n26423;
  assign n26396 = n4673 & ~n23879;
  assign n26397 = n4688 & ~n23292;
  assign n26398 = n4685 & n23052;
  assign n26399 = ~n4681 & n19649;
  assign n26400 = ~n26398 & ~n26399;
  assign n26401 = ~n26397 & n26400;
  assign n26402 = ~n26396 & n26401;
  assign n26403 = n26402 ^ x20;
  assign n26386 = n4478 & ~n23468;
  assign n26387 = n4484 & ~n19512;
  assign n26388 = n4480 & n19439;
  assign n26389 = ~n26387 & ~n26388;
  assign n26390 = n4487 & ~n19575;
  assign n26391 = n26389 & ~n26390;
  assign n26392 = ~n26386 & n26391;
  assign n26393 = n26392 ^ x23;
  assign n26376 = n3285 & ~n22037;
  assign n26377 = n3437 & ~n19368;
  assign n26378 = n3435 & n19063;
  assign n26379 = ~n3440 & n19303;
  assign n26380 = ~n26378 & ~n26379;
  assign n26381 = ~n26377 & n26380;
  assign n26382 = ~n26376 & n26381;
  assign n26383 = n26382 ^ x26;
  assign n26358 = ~x28 & ~n21715;
  assign n26359 = x28 & ~n19078;
  assign n26360 = x29 & ~n26359;
  assign n26361 = ~n26358 & n26360;
  assign n26362 = ~n12475 & ~n26361;
  assign n26363 = n3275 & n19096;
  assign n26364 = n3277 & n19298;
  assign n26365 = ~n26363 & ~n26364;
  assign n26366 = ~n26362 & n26365;
  assign n26367 = x28 & n21715;
  assign n26368 = ~x28 & n19078;
  assign n26369 = n12466 & ~n26368;
  assign n26370 = ~n26367 & n26369;
  assign n26371 = ~x29 & ~n26365;
  assign n26372 = ~n26370 & ~n26371;
  assign n26373 = ~n26366 & n26372;
  assign n26344 = n26091 & n26104;
  assign n26345 = n26233 & ~n26242;
  assign n26346 = n26344 & ~n26345;
  assign n26347 = ~n26233 & n26242;
  assign n26348 = n25974 & ~n26347;
  assign n26349 = ~n26346 & n26348;
  assign n26350 = ~n26091 & ~n26104;
  assign n26351 = n26350 ^ n26242;
  assign n26352 = ~n25974 & ~n26233;
  assign n26353 = n26352 ^ n26242;
  assign n26354 = ~n26351 & n26353;
  assign n26355 = n26354 ^ n26350;
  assign n26356 = ~n26349 & ~n26355;
  assign n26336 = n3667 & n21684;
  assign n26337 = ~n3673 & n19104;
  assign n26338 = n3669 & ~n19286;
  assign n26339 = ~n26337 & ~n26338;
  assign n26340 = n3676 & n19292;
  assign n26341 = n26339 & ~n26340;
  assign n26342 = ~n26336 & n26341;
  assign n26323 = ~n133 & ~n284;
  assign n26324 = n1324 & n26323;
  assign n26325 = n2378 & n26324;
  assign n26326 = n21265 & n26325;
  assign n26327 = n12743 & n13507;
  assign n26328 = n411 & n26327;
  assign n26329 = n3109 & n26328;
  assign n26330 = n26326 & n26329;
  assign n26331 = n4548 & n26330;
  assign n26332 = n12254 & n26331;
  assign n26333 = n4104 & n26332;
  assign n26334 = n1207 & n26333;
  assign n26319 = n25974 ^ x14;
  assign n26320 = n26232 ^ n25974;
  assign n26321 = n26319 & ~n26320;
  assign n26322 = n26321 ^ x14;
  assign n26335 = n26334 ^ n26322;
  assign n26343 = n26342 ^ n26335;
  assign n26357 = n26356 ^ n26343;
  assign n26374 = n26373 ^ n26357;
  assign n26316 = n26268 ^ n26259;
  assign n26317 = n26260 & n26316;
  assign n26318 = n26317 ^ n26268;
  assign n26375 = n26374 ^ n26318;
  assign n26384 = n26383 ^ n26375;
  assign n26313 = n26269 ^ n26214;
  assign n26314 = ~n26270 & n26313;
  assign n26315 = n26314 ^ n26217;
  assign n26385 = n26384 ^ n26315;
  assign n26394 = n26393 ^ n26385;
  assign n26310 = n26280 ^ n26206;
  assign n26311 = n26272 & n26310;
  assign n26312 = n26311 ^ n26280;
  assign n26395 = n26394 ^ n26312;
  assign n26404 = n26403 ^ n26395;
  assign n26308 = n4970 & n23495;
  assign n26309 = n26308 ^ x17;
  assign n26405 = n26404 ^ n26309;
  assign n26305 = n26289 ^ n26203;
  assign n26306 = n26290 & n26305;
  assign n26307 = n26306 ^ n26203;
  assign n26406 = n26405 ^ n26307;
  assign n26425 = n26424 ^ n26406;
  assign n26302 = n26297 ^ n26200;
  assign n26303 = n26298 & n26302;
  assign n26304 = n26303 ^ n26200;
  assign n26426 = n26425 ^ n26304;
  assign n26436 = n26435 ^ n26426;
  assign n26531 = n26426 & n26435;
  assign n26532 = n26406 ^ n26304;
  assign n26533 = ~n26425 & ~n26532;
  assign n26534 = n26533 ^ n26424;
  assign n26535 = ~n26531 & ~n26534;
  assign n26536 = ~n26406 & n26424;
  assign n26537 = ~n26304 & n26536;
  assign n26538 = n26435 & n26537;
  assign n26539 = ~n26535 & ~n26538;
  assign n26519 = n4673 & n23493;
  assign n26520 = n4688 & n23495;
  assign n26521 = n4685 & ~n23292;
  assign n26522 = ~n4681 & n23052;
  assign n26523 = ~n26521 & ~n26522;
  assign n26524 = ~n26520 & n26523;
  assign n26525 = ~n26519 & n26524;
  assign n26526 = n26525 ^ x20;
  assign n26501 = n12502 & n23520;
  assign n26502 = n4480 & ~n19512;
  assign n26503 = n4484 & ~n19575;
  assign n26504 = ~n26502 & ~n26503;
  assign n26505 = x23 & n26504;
  assign n26506 = ~n19649 & n26505;
  assign n26507 = x22 & ~n26506;
  assign n26508 = ~n26501 & n26507;
  assign n26509 = ~n23520 & n26505;
  assign n26510 = n12502 & n19649;
  assign n26511 = ~x22 & ~n26510;
  assign n26512 = ~n26509 & n26511;
  assign n26513 = ~n26508 & ~n26512;
  assign n26514 = ~n12519 & n26504;
  assign n26515 = n26514 ^ x23;
  assign n26516 = ~n26513 & n26515;
  assign n26491 = n3285 & n22457;
  assign n26492 = n3437 & n19439;
  assign n26493 = n3435 & ~n19368;
  assign n26494 = ~n3440 & n19063;
  assign n26495 = ~n26493 & ~n26494;
  assign n26496 = ~n26492 & n26495;
  assign n26497 = ~n26491 & n26496;
  assign n26498 = n26497 ^ x26;
  assign n26481 = n44 & n19658;
  assign n26482 = n3277 & ~n19078;
  assign n26483 = n3280 & n19303;
  assign n26484 = n3275 & n19298;
  assign n26485 = ~n26483 & ~n26484;
  assign n26486 = ~n26482 & n26485;
  assign n26487 = ~n26481 & n26486;
  assign n26488 = n26487 ^ x29;
  assign n26469 = ~n54 & n21699;
  assign n26470 = n54 & n19104;
  assign n26471 = n11234 & ~n26470;
  assign n26472 = ~n26469 & n26471;
  assign n26473 = n41 & n19096;
  assign n26474 = ~x31 & ~n19292;
  assign n26475 = ~n5358 & ~n26474;
  assign n26476 = ~n26473 & ~n26475;
  assign n26477 = n91 & ~n19292;
  assign n26478 = ~n26476 & ~n26477;
  assign n26479 = ~n26472 & n26478;
  assign n26463 = n26322 & n26342;
  assign n26464 = n26334 & n26463;
  assign n26465 = ~n26322 & ~n26342;
  assign n26466 = ~n26334 & n26465;
  assign n26467 = ~n26464 & ~n26466;
  assign n26452 = n3215 & n12155;
  assign n26453 = n4554 & n11393;
  assign n26454 = n13405 & n26453;
  assign n26455 = n834 & n4906;
  assign n26456 = n1497 & n26455;
  assign n26457 = n26454 & n26456;
  assign n26458 = n26452 & n26457;
  assign n26459 = n917 & n11264;
  assign n26460 = n26458 & n26459;
  assign n26461 = n2568 & n4186;
  assign n26462 = n26460 & n26461;
  assign n26468 = n26467 ^ n26462;
  assign n26480 = n26479 ^ n26468;
  assign n26489 = n26488 ^ n26480;
  assign n26449 = n26373 ^ n26356;
  assign n26450 = n26357 & n26449;
  assign n26451 = n26450 ^ n26373;
  assign n26490 = n26489 ^ n26451;
  assign n26499 = n26498 ^ n26490;
  assign n26446 = n26383 ^ n26374;
  assign n26447 = n26375 & ~n26446;
  assign n26448 = n26447 ^ n26383;
  assign n26500 = n26499 ^ n26448;
  assign n26517 = n26516 ^ n26500;
  assign n26443 = n26393 ^ n26315;
  assign n26444 = n26385 & n26443;
  assign n26445 = n26444 ^ n26393;
  assign n26518 = n26517 ^ n26445;
  assign n26527 = n26526 ^ n26518;
  assign n26528 = n26527 ^ x17;
  assign n26440 = n26403 ^ n26312;
  assign n26441 = n26395 & n26440;
  assign n26442 = n26441 ^ n26403;
  assign n26529 = n26528 ^ n26442;
  assign n26437 = n26404 ^ n26307;
  assign n26438 = ~n26405 & ~n26437;
  assign n26439 = n26438 ^ n26307;
  assign n26530 = n26529 ^ n26439;
  assign n26540 = n26539 ^ n26530;
  assign n26631 = ~n26442 & ~n26527;
  assign n26632 = ~x17 & ~n26631;
  assign n26633 = n26442 & n26527;
  assign n26634 = ~n26632 & ~n26633;
  assign n26623 = n4673 & ~n23704;
  assign n26624 = n4685 & n23495;
  assign n26625 = ~n4681 & ~n23292;
  assign n26626 = ~n26624 & ~n26625;
  assign n26627 = ~n26623 & n26626;
  assign n26628 = n26627 ^ x20;
  assign n26613 = n4478 & n23712;
  assign n26614 = n4484 & n19649;
  assign n26615 = n4480 & ~n19575;
  assign n26616 = ~n26614 & ~n26615;
  assign n26617 = n4487 & n23052;
  assign n26618 = n26616 & ~n26617;
  assign n26619 = ~n26613 & n26618;
  assign n26620 = n26619 ^ x23;
  assign n26603 = n3285 & ~n23064;
  assign n26604 = n3437 & ~n19512;
  assign n26605 = n3435 & n19439;
  assign n26606 = ~n3440 & ~n19368;
  assign n26607 = ~n26605 & ~n26606;
  assign n26608 = ~n26604 & n26607;
  assign n26609 = ~n26603 & n26608;
  assign n26610 = n26609 ^ x26;
  assign n26600 = n26498 ^ n26451;
  assign n26601 = ~n26490 & n26600;
  assign n26602 = n26601 ^ n26498;
  assign n26611 = n26610 ^ n26602;
  assign n26590 = n44 & n22441;
  assign n26591 = n3280 & n19063;
  assign n26592 = n3275 & ~n19078;
  assign n26593 = n3277 & n19303;
  assign n26594 = ~n26592 & ~n26593;
  assign n26595 = ~n26591 & n26594;
  assign n26596 = ~n26590 & n26595;
  assign n26597 = n26596 ^ x29;
  assign n26576 = x31 & n19667;
  assign n26577 = n26576 ^ n19298;
  assign n26578 = x30 & ~n26577;
  assign n26579 = ~x29 & x31;
  assign n26580 = n19096 & n26579;
  assign n26581 = ~n60 & ~n26580;
  assign n26582 = ~n26578 & ~n26581;
  assign n26583 = n45 & n26577;
  assign n26584 = n3671 & n19096;
  assign n26585 = n3669 & n19292;
  assign n26586 = ~n26584 & ~n26585;
  assign n26587 = ~n26583 & n26586;
  assign n26588 = ~n26582 & n26587;
  assign n26573 = ~n26462 & ~n26466;
  assign n26574 = ~n26464 & ~n26573;
  assign n26558 = n3376 & n11242;
  assign n26559 = ~n185 & ~n262;
  assign n26560 = ~n99 & n26559;
  assign n26561 = n11069 & n26560;
  assign n26562 = n26558 & n26561;
  assign n26563 = n294 & n1866;
  assign n26564 = n1205 & n21261;
  assign n26565 = n26563 & n26564;
  assign n26566 = n2782 & n26565;
  assign n26567 = n11018 & n26566;
  assign n26568 = n26562 & n26567;
  assign n26569 = n564 & n26568;
  assign n26570 = n4769 & n26569;
  assign n26571 = n3706 & n26570;
  assign n26557 = n26462 ^ x17;
  assign n26572 = n26571 ^ n26557;
  assign n26575 = n26574 ^ n26572;
  assign n26589 = n26588 ^ n26575;
  assign n26598 = n26597 ^ n26589;
  assign n26554 = n26488 ^ n26479;
  assign n26555 = ~n26480 & ~n26554;
  assign n26556 = n26555 ^ n26488;
  assign n26599 = n26598 ^ n26556;
  assign n26612 = n26611 ^ n26599;
  assign n26621 = n26620 ^ n26612;
  assign n26551 = n26516 ^ n26499;
  assign n26552 = ~n26500 & n26551;
  assign n26553 = n26552 ^ n26516;
  assign n26622 = n26621 ^ n26553;
  assign n26629 = n26628 ^ n26622;
  assign n26548 = n26526 ^ n26517;
  assign n26549 = ~n26518 & n26548;
  assign n26550 = n26549 ^ n26526;
  assign n26630 = n26629 ^ n26550;
  assign n26635 = n26634 ^ n26630;
  assign n26541 = ~n26439 & n26529;
  assign n26542 = n26541 ^ n26538;
  assign n26543 = n26439 & ~n26529;
  assign n26544 = ~n26535 & ~n26543;
  assign n26545 = ~n26541 & n26544;
  assign n26546 = ~n26542 & n26545;
  assign n26547 = n26546 ^ n26542;
  assign n26636 = n26635 ^ n26547;
  assign n26723 = ~n26439 & n26534;
  assign n26724 = n26442 ^ x17;
  assign n26725 = n26527 ^ n26442;
  assign n26726 = n26630 ^ n26527;
  assign n26727 = ~n26725 & ~n26726;
  assign n26728 = n26724 & n26727;
  assign n26729 = n26728 ^ n26630;
  assign n26730 = ~n26723 & ~n26729;
  assign n26731 = n26439 & ~n26534;
  assign n26732 = n26731 ^ n26630;
  assign n26733 = n26635 & n26732;
  assign n26734 = n26733 ^ n26634;
  assign n26735 = ~n26730 & n26734;
  assign n26711 = n4478 & ~n23879;
  assign n26712 = n4487 & ~n23292;
  assign n26713 = n4484 & n23052;
  assign n26714 = n4480 & n19649;
  assign n26715 = ~n26713 & ~n26714;
  assign n26716 = ~n26712 & n26715;
  assign n26717 = ~n26711 & n26716;
  assign n26718 = n26717 ^ x23;
  assign n26701 = n3285 & ~n23468;
  assign n26702 = n3435 & ~n19512;
  assign n26703 = ~n3440 & n19439;
  assign n26704 = ~n26702 & ~n26703;
  assign n26705 = n3437 & ~n19575;
  assign n26706 = n26704 & ~n26705;
  assign n26707 = ~n26701 & n26706;
  assign n26708 = n26707 ^ x26;
  assign n26691 = n44 & ~n22037;
  assign n26692 = n3280 & ~n19368;
  assign n26693 = n3277 & n19063;
  assign n26694 = n3275 & n19303;
  assign n26695 = ~n26693 & ~n26694;
  assign n26696 = ~n26692 & n26695;
  assign n26697 = ~n26691 & n26696;
  assign n26698 = n26697 ^ x29;
  assign n26677 = n41 & ~n21715;
  assign n26678 = n54 & n19096;
  assign n26679 = n91 & n19298;
  assign n26680 = ~n26678 & ~n26679;
  assign n26681 = x31 & n26680;
  assign n26682 = ~n26677 & n26681;
  assign n26683 = n41 & ~n19078;
  assign n26684 = ~x31 & ~n19298;
  assign n26685 = ~n5358 & ~n26684;
  assign n26686 = ~n26683 & ~n26685;
  assign n26687 = ~n26682 & ~n26686;
  assign n26664 = n4750 & n5659;
  assign n26665 = n11809 & n26664;
  assign n26666 = ~n683 & ~n850;
  assign n26667 = ~n217 & n26666;
  assign n26668 = n2040 & n13416;
  assign n26669 = n26667 & n26668;
  assign n26670 = n533 & n728;
  assign n26671 = n26669 & n26670;
  assign n26672 = n26665 & n26671;
  assign n26673 = n2887 & n26672;
  assign n26674 = n981 & n26673;
  assign n26675 = n5412 & n25214;
  assign n26676 = n26674 & n26675;
  assign n26688 = n26687 ^ n26676;
  assign n26661 = n26588 ^ n26574;
  assign n26662 = n26575 & ~n26661;
  assign n26663 = n26662 ^ n26588;
  assign n26689 = n26688 ^ n26663;
  assign n26658 = n26571 ^ n26462;
  assign n26659 = n26557 & ~n26658;
  assign n26660 = n26659 ^ x17;
  assign n26690 = n26689 ^ n26660;
  assign n26699 = n26698 ^ n26690;
  assign n26655 = n26589 ^ n26556;
  assign n26656 = ~n26598 & n26655;
  assign n26657 = n26656 ^ n26597;
  assign n26700 = n26699 ^ n26657;
  assign n26709 = n26708 ^ n26700;
  assign n26652 = n26602 ^ n26599;
  assign n26653 = n26611 & n26652;
  assign n26654 = n26653 ^ n26610;
  assign n26710 = n26709 ^ n26654;
  assign n26719 = n26718 ^ n26710;
  assign n26650 = ~n4681 & n23495;
  assign n26651 = n26650 ^ x20;
  assign n26720 = n26719 ^ n26651;
  assign n26647 = n26620 ^ n26553;
  assign n26648 = n26621 & n26647;
  assign n26649 = n26648 ^ n26553;
  assign n26721 = n26720 ^ n26649;
  assign n26644 = n26628 ^ n26550;
  assign n26645 = n26629 & n26644;
  assign n26646 = n26645 ^ n26550;
  assign n26722 = n26721 ^ n26646;
  assign n26736 = n26735 ^ n26722;
  assign n26637 = ~n26541 & ~n26635;
  assign n26638 = ~n26543 & n26635;
  assign n26639 = n26638 ^ n26530;
  assign n26640 = n26534 & n26639;
  assign n26641 = n26640 ^ n26530;
  assign n26642 = ~n26637 & ~n26641;
  assign n26643 = n26531 & n26642;
  assign n26737 = n26736 ^ n26643;
  assign n26826 = n4478 & n23493;
  assign n26827 = n4487 & n23495;
  assign n26828 = n4484 & ~n23292;
  assign n26829 = n4480 & n23052;
  assign n26830 = ~n26828 & ~n26829;
  assign n26831 = ~n26827 & n26830;
  assign n26832 = ~n26826 & n26831;
  assign n26833 = n26832 ^ x23;
  assign n26808 = n12417 & n23520;
  assign n26809 = ~n3440 & ~n19512;
  assign n26810 = n3435 & ~n19575;
  assign n26811 = ~n26809 & ~n26810;
  assign n26812 = x26 & n26811;
  assign n26813 = ~n19649 & n26812;
  assign n26814 = x25 & ~n26813;
  assign n26815 = ~n26808 & n26814;
  assign n26816 = ~n23520 & n26812;
  assign n26817 = n12417 & n19649;
  assign n26818 = ~x25 & ~n26817;
  assign n26819 = ~n26816 & n26818;
  assign n26820 = ~n26815 & ~n26819;
  assign n26821 = ~n12432 & n26811;
  assign n26822 = n26821 ^ x26;
  assign n26823 = ~n26820 & n26822;
  assign n26785 = n26663 & n26698;
  assign n26786 = ~n26676 & n26785;
  assign n26787 = n26687 & ~n26786;
  assign n26788 = n26676 ^ n26663;
  assign n26789 = n26698 ^ n26663;
  assign n26790 = n26788 & n26789;
  assign n26791 = n26790 ^ n26698;
  assign n26792 = ~n26787 & n26791;
  assign n26793 = n26660 & ~n26792;
  assign n26794 = ~n26663 & ~n26698;
  assign n26795 = ~n26676 & ~n26687;
  assign n26796 = n26794 & ~n26795;
  assign n26797 = ~n26660 & ~n26796;
  assign n26798 = n26676 & n26687;
  assign n26799 = ~n26785 & n26798;
  assign n26800 = n26797 & ~n26799;
  assign n26801 = ~n26793 & ~n26800;
  assign n26802 = n26794 & n26798;
  assign n26803 = n26785 & n26795;
  assign n26804 = ~n26802 & ~n26803;
  assign n26805 = ~n26801 & n26804;
  assign n26775 = n3667 & n19658;
  assign n26776 = ~n12591 & ~n19078;
  assign n26777 = ~n5354 & ~n26776;
  assign n26778 = n3669 & ~n19298;
  assign n26779 = ~n26777 & ~n26778;
  assign n26780 = ~x31 & n19303;
  assign n26781 = n41 & ~n26780;
  assign n26782 = n26779 & ~n26781;
  assign n26783 = ~n26775 & ~n26782;
  assign n26760 = n1575 & n11583;
  assign n26761 = ~n141 & ~n248;
  assign n26762 = n1180 & n26761;
  assign n26763 = n26760 & n26762;
  assign n26764 = n24481 & n26763;
  assign n26765 = ~n593 & ~n1166;
  assign n26766 = ~n353 & n26765;
  assign n26767 = n12728 & n26766;
  assign n26768 = n13405 & n26767;
  assign n26769 = n26764 & n26768;
  assign n26770 = n3692 & n26769;
  assign n26771 = n4919 & n5460;
  assign n26772 = n26770 & n26771;
  assign n26773 = n565 & n26772;
  assign n26774 = n26773 ^ n26676;
  assign n26784 = n26783 ^ n26774;
  assign n26806 = n26805 ^ n26784;
  assign n26752 = n44 & n22457;
  assign n26753 = n3280 & n19439;
  assign n26754 = n3277 & ~n19368;
  assign n26755 = n3275 & n19063;
  assign n26756 = ~n26754 & ~n26755;
  assign n26757 = ~n26753 & n26756;
  assign n26758 = ~n26752 & n26757;
  assign n26759 = n26758 ^ x29;
  assign n26807 = n26806 ^ n26759;
  assign n26824 = n26823 ^ n26807;
  assign n26749 = n26708 ^ n26699;
  assign n26750 = ~n26700 & n26749;
  assign n26751 = n26750 ^ n26708;
  assign n26825 = n26824 ^ n26751;
  assign n26834 = n26833 ^ n26825;
  assign n26835 = n26834 ^ x20;
  assign n26746 = n26718 ^ n26654;
  assign n26747 = ~n26710 & n26746;
  assign n26748 = n26747 ^ n26718;
  assign n26836 = n26835 ^ n26748;
  assign n26743 = n26719 ^ n26649;
  assign n26744 = n26720 & n26743;
  assign n26745 = n26744 ^ n26649;
  assign n26837 = n26836 ^ n26745;
  assign n26740 = n26722 ^ n26643;
  assign n26741 = ~n26735 & ~n26740;
  assign n26738 = n26721 ^ n26643;
  assign n26739 = n26722 & ~n26738;
  assign n26742 = n26741 ^ n26739;
  assign n26838 = n26837 ^ n26742;
  assign n26932 = n12417 & n23712;
  assign n26933 = n3435 & n19649;
  assign n26934 = ~n3440 & ~n19575;
  assign n26935 = ~n26933 & ~n26934;
  assign n26936 = x26 & n26935;
  assign n26937 = ~n23052 & n26936;
  assign n26938 = ~n26932 & ~n26937;
  assign n26939 = x25 & n26938;
  assign n26940 = ~n23712 & n26936;
  assign n26941 = n12417 & n23052;
  assign n26942 = ~x25 & ~n26941;
  assign n26943 = ~n26940 & n26942;
  assign n26944 = ~n26939 & ~n26943;
  assign n26945 = ~n12432 & n26935;
  assign n26946 = n26945 ^ x26;
  assign n26947 = ~n26944 & n26946;
  assign n26929 = n26823 ^ n26806;
  assign n26930 = n26807 & ~n26929;
  assign n26931 = n26930 ^ n26823;
  assign n26948 = n26947 ^ n26931;
  assign n26912 = ~x28 & ~n23064;
  assign n26913 = x28 & ~n19512;
  assign n26914 = x29 & ~n26913;
  assign n26915 = ~n26912 & n26914;
  assign n26916 = ~n12475 & ~n26915;
  assign n26917 = n3277 & n19439;
  assign n26918 = n3275 & ~n19368;
  assign n26919 = ~n26917 & ~n26918;
  assign n26920 = ~n26916 & n26919;
  assign n26921 = x28 & n23064;
  assign n26922 = ~x28 & n19512;
  assign n26923 = n12466 & ~n26922;
  assign n26924 = ~n26921 & n26923;
  assign n26925 = ~x29 & ~n26919;
  assign n26926 = ~n26924 & ~n26925;
  assign n26927 = ~n26920 & n26926;
  assign n26898 = n26784 & ~n26785;
  assign n26899 = ~n26660 & ~n26795;
  assign n26900 = ~n26798 & ~n26899;
  assign n26901 = ~n26898 & n26900;
  assign n26902 = n26676 ^ n26660;
  assign n26903 = n26784 ^ n26660;
  assign n26904 = n26902 & ~n26903;
  assign n26905 = ~n26688 & n26904;
  assign n26906 = n26905 ^ n26784;
  assign n26907 = ~n26794 & ~n26906;
  assign n26908 = ~n26784 & n26785;
  assign n26909 = ~n26907 & ~n26908;
  assign n26910 = ~n26901 & n26909;
  assign n26891 = n26773 & n26783;
  assign n26892 = n26676 & n26891;
  assign n26893 = ~n26773 & ~n26783;
  assign n26894 = ~n26676 & n26893;
  assign n26895 = ~n26892 & ~n26894;
  assign n26875 = ~n385 & n3183;
  assign n26876 = n1834 & n11642;
  assign n26877 = n26875 & n26876;
  assign n26878 = ~n518 & ~n525;
  assign n26879 = n441 & n26878;
  assign n26880 = n2521 & n26879;
  assign n26881 = n26877 & n26880;
  assign n26882 = n916 & n26881;
  assign n26883 = n13414 & n26882;
  assign n26884 = n474 & n1036;
  assign n26885 = n4194 & n26884;
  assign n26886 = n12729 & n26885;
  assign n26887 = n26883 & n26886;
  assign n26888 = n2668 & n26887;
  assign n26889 = n4379 & n26888;
  assign n26890 = n26889 ^ x20;
  assign n26896 = n26895 ^ n26890;
  assign n26864 = n41 & ~n22441;
  assign n26865 = x31 & ~n19078;
  assign n26866 = ~n12183 & ~n26865;
  assign n26867 = ~n26864 & ~n26866;
  assign n26868 = n91 & ~n19303;
  assign n26869 = n26867 & ~n26868;
  assign n26870 = n41 & n19063;
  assign n26871 = n54 & n19303;
  assign n26872 = ~n26870 & ~n26871;
  assign n26873 = ~x31 & ~n26872;
  assign n26874 = ~n26869 & ~n26873;
  assign n26897 = n26896 ^ n26874;
  assign n26911 = n26910 ^ n26897;
  assign n26928 = n26927 ^ n26911;
  assign n26949 = n26948 ^ n26928;
  assign n26858 = n4478 & ~n23704;
  assign n26859 = n4484 & n23495;
  assign n26860 = n4480 & ~n23292;
  assign n26861 = ~n26859 & ~n26860;
  assign n26862 = ~n26858 & n26861;
  assign n26863 = n26862 ^ x23;
  assign n26950 = n26949 ^ n26863;
  assign n26855 = n26833 ^ n26824;
  assign n26856 = n26825 & ~n26855;
  assign n26857 = n26856 ^ n26833;
  assign n26951 = n26950 ^ n26857;
  assign n26852 = n26834 ^ n26748;
  assign n26853 = n26835 & n26852;
  assign n26854 = n26853 ^ x20;
  assign n26952 = n26951 ^ n26854;
  assign n26839 = n26646 & ~n26721;
  assign n26840 = n26735 & ~n26839;
  assign n26843 = ~n26646 & n26721;
  assign n26848 = ~n26840 & ~n26843;
  assign n26849 = n26848 ^ n26745;
  assign n26850 = ~n26837 & n26849;
  assign n26851 = n26850 ^ n26848;
  assign n26953 = n26952 ^ n26851;
  assign n26841 = n26837 & n26840;
  assign n26842 = n26722 & ~n26735;
  assign n26844 = ~n26837 & ~n26843;
  assign n26845 = n26643 & ~n26844;
  assign n26846 = ~n26842 & n26845;
  assign n26847 = ~n26841 & n26846;
  assign n26954 = n26953 ^ n26847;
  assign n27034 = n26847 & ~n26953;
  assign n27031 = n26949 ^ n26857;
  assign n27032 = n26950 & ~n27031;
  assign n27033 = n27032 ^ n26857;
  assign n27035 = n27034 ^ n27033;
  assign n27019 = n3285 & ~n23879;
  assign n27020 = n3437 & ~n23292;
  assign n27021 = n3435 & n23052;
  assign n27022 = ~n3440 & n19649;
  assign n27023 = ~n27021 & ~n27022;
  assign n27024 = ~n27020 & n27023;
  assign n27025 = ~n27019 & n27024;
  assign n27026 = n27025 ^ x26;
  assign n27008 = n44 & ~n23468;
  assign n27009 = n3277 & ~n19512;
  assign n27010 = n3275 & n19439;
  assign n27011 = ~n27009 & ~n27010;
  assign n27012 = n3280 & ~n19575;
  assign n27013 = n27011 & ~n27012;
  assign n27014 = ~n27008 & n27013;
  assign n27015 = n27014 ^ x29;
  assign n26997 = ~n26874 & ~n26892;
  assign n26998 = ~n26894 & ~n26997;
  assign n26999 = ~n26890 & ~n26998;
  assign n27000 = n26783 ^ n26773;
  assign n27001 = n26874 ^ n26773;
  assign n27002 = n26676 & n26890;
  assign n27003 = n27002 ^ n26874;
  assign n27004 = ~n27001 & ~n27003;
  assign n27005 = ~n27000 & n27004;
  assign n27006 = n27005 ^ n27002;
  assign n27007 = ~n26999 & ~n27006;
  assign n27016 = n27015 ^ n27007;
  assign n26981 = n2102 & n13510;
  assign n26982 = n3706 & n26981;
  assign n26983 = ~n228 & ~n1060;
  assign n26984 = ~n115 & ~n336;
  assign n26985 = n26983 & n26984;
  assign n26986 = n1934 & n26985;
  assign n26987 = n2182 & n3893;
  assign n26988 = n430 & n584;
  assign n26989 = n26987 & n26988;
  assign n26990 = n26986 & n26989;
  assign n26991 = n2226 & n26990;
  assign n26992 = n3604 & n26991;
  assign n26993 = n12276 & n26992;
  assign n26994 = n26982 & n26993;
  assign n26977 = n26676 ^ x20;
  assign n26978 = n26889 ^ n26676;
  assign n26979 = n26977 & ~n26978;
  assign n26980 = n26979 ^ x20;
  assign n26995 = n26994 ^ n26980;
  assign n26969 = n41 & n22037;
  assign n26970 = n91 & ~n19063;
  assign n26971 = n54 & ~n19303;
  assign n26972 = ~n26970 & ~n26971;
  assign n26973 = ~n26969 & n26972;
  assign n26966 = n41 & ~n19368;
  assign n26967 = n54 & n19063;
  assign n26968 = ~n26966 & ~n26967;
  assign n26974 = n26973 ^ n26968;
  assign n26975 = ~x31 & ~n26974;
  assign n26976 = n26975 ^ n26973;
  assign n26996 = n26995 ^ n26976;
  assign n27017 = n27016 ^ n26996;
  assign n26963 = n26927 ^ n26910;
  assign n26964 = n26911 & ~n26963;
  assign n26965 = n26964 ^ n26927;
  assign n27018 = n27017 ^ n26965;
  assign n27027 = n27026 ^ n27018;
  assign n26961 = n4480 & n23495;
  assign n26962 = n26961 ^ x23;
  assign n27028 = n27027 ^ n26962;
  assign n26958 = n26931 ^ n26928;
  assign n26959 = n26948 & n26958;
  assign n26960 = n26959 ^ n26947;
  assign n27029 = n27028 ^ n26960;
  assign n26955 = n26854 ^ n26851;
  assign n26956 = ~n26952 & ~n26955;
  assign n26957 = n26956 ^ n26851;
  assign n27030 = n27029 ^ n26957;
  assign n27036 = n27035 ^ n27030;
  assign n27099 = n3285 & n23493;
  assign n27100 = n3437 & n23495;
  assign n27101 = n3435 & ~n23292;
  assign n27102 = ~n3440 & n23052;
  assign n27103 = ~n27101 & ~n27102;
  assign n27104 = ~n27100 & n27103;
  assign n27105 = ~n27099 & n27104;
  assign n27106 = n27105 ^ x26;
  assign n27090 = n26980 & n26994;
  assign n27091 = ~n26976 & n27090;
  assign n27092 = ~n26980 & ~n26994;
  assign n27093 = n26976 & n27092;
  assign n27094 = ~n27091 & ~n27093;
  assign n27077 = ~n209 & ~n524;
  assign n27078 = n893 & n27077;
  assign n27079 = n236 & n27078;
  assign n27080 = n962 & n13311;
  assign n27081 = n27079 & n27080;
  assign n27082 = n1046 & n1225;
  assign n27083 = n584 & n3075;
  assign n27084 = n27082 & n27083;
  assign n27085 = n27081 & n27084;
  assign n27086 = n25200 & n27085;
  assign n27087 = n19399 & n27086;
  assign n27088 = n20728 & n27087;
  assign n27089 = n10104 & n27088;
  assign n27095 = n27094 ^ n27089;
  assign n27067 = n41 & n22457;
  assign n27068 = n91 & ~n19368;
  assign n27069 = x31 & ~n26967;
  assign n27070 = ~n27068 & n27069;
  assign n27071 = ~n27067 & n27070;
  assign n27072 = n41 & n19439;
  assign n27073 = n54 & ~n19368;
  assign n27074 = ~x31 & ~n27073;
  assign n27075 = ~n27072 & n27074;
  assign n27076 = ~n27071 & ~n27075;
  assign n27096 = n27095 ^ n27076;
  assign n27064 = n27007 ^ n26996;
  assign n27065 = n27016 & ~n27064;
  assign n27066 = n27065 ^ n27015;
  assign n27097 = n27096 ^ n27066;
  assign n27048 = n12466 & n23520;
  assign n27049 = n3275 & ~n19512;
  assign n27050 = n3277 & ~n19575;
  assign n27051 = ~n27049 & ~n27050;
  assign n27052 = x29 & n27051;
  assign n27053 = ~n19649 & n27052;
  assign n27054 = x28 & ~n27053;
  assign n27055 = ~n27048 & n27054;
  assign n27056 = ~n23520 & n27052;
  assign n27057 = n12466 & n19649;
  assign n27058 = ~x28 & ~n27057;
  assign n27059 = ~n27056 & n27058;
  assign n27060 = ~n27055 & ~n27059;
  assign n27061 = ~n12476 & n27051;
  assign n27062 = n27061 ^ x29;
  assign n27063 = ~n27060 & n27062;
  assign n27098 = n27097 ^ n27063;
  assign n27107 = n27106 ^ n27098;
  assign n27045 = n27026 ^ n26965;
  assign n27046 = ~n27018 & n27045;
  assign n27047 = n27046 ^ n27026;
  assign n27108 = n27107 ^ n27047;
  assign n27109 = n27108 ^ x23;
  assign n27042 = n27027 ^ n26960;
  assign n27043 = n27028 & n27042;
  assign n27044 = n27043 ^ n26960;
  assign n27110 = n27109 ^ n27044;
  assign n27037 = n27033 ^ n26957;
  assign n27039 = n27037 ^ n27029;
  assign n27040 = ~n27034 & n27039;
  assign n27038 = n27030 & ~n27037;
  assign n27041 = n27040 ^ n27038;
  assign n27111 = n27110 ^ n27041;
  assign n27181 = ~n26957 & n27029;
  assign n27182 = n27110 & ~n27181;
  assign n27183 = n27034 & ~n27182;
  assign n27184 = n26957 & ~n27029;
  assign n27185 = ~n27033 & ~n27110;
  assign n27186 = ~n27184 & n27185;
  assign n27187 = n27183 & ~n27186;
  assign n27188 = n27030 & n27033;
  assign n27189 = n27187 & ~n27188;
  assign n27164 = ~n26960 & ~n27027;
  assign n27165 = ~n27109 & ~n27164;
  assign n27166 = ~n27033 & ~n27165;
  assign n27167 = n26960 & n27027;
  assign n27168 = n27109 & ~n27167;
  assign n27169 = ~n27166 & ~n27168;
  assign n27170 = n26962 & ~n27169;
  assign n27171 = n27033 & ~n27164;
  assign n27172 = n27168 & ~n27171;
  assign n27173 = ~n27170 & ~n27172;
  assign n27174 = n26957 & n27173;
  assign n27175 = ~n27167 & ~n27171;
  assign n27176 = ~n27109 & ~n27175;
  assign n27177 = ~n26962 & n27169;
  assign n27178 = ~n27176 & ~n27177;
  assign n27179 = ~n27174 & n27178;
  assign n27155 = n3285 & ~n23704;
  assign n27156 = n3435 & n23495;
  assign n27157 = ~n3440 & ~n23292;
  assign n27158 = ~n27156 & ~n27157;
  assign n27159 = ~n27155 & n27158;
  assign n27160 = n27159 ^ x26;
  assign n27145 = n44 & n23712;
  assign n27146 = n3277 & n19649;
  assign n27147 = n3275 & ~n19575;
  assign n27148 = ~n27146 & ~n27147;
  assign n27149 = n3280 & n23052;
  assign n27150 = n27148 & ~n27149;
  assign n27151 = ~n27145 & n27150;
  assign n27152 = n27151 ^ x29;
  assign n27136 = x31 & n23064;
  assign n27137 = ~x31 & n19512;
  assign n27138 = n41 & ~n27137;
  assign n27139 = ~n27136 & n27138;
  assign n27140 = ~n3673 & n19439;
  assign n27141 = x31 & n27073;
  assign n27142 = ~n27140 & ~n27141;
  assign n27143 = ~n27139 & n27142;
  assign n27133 = n27089 & ~n27091;
  assign n27134 = ~n27093 & ~n27133;
  assign n27131 = n27089 ^ x23;
  assign n27121 = ~n61 & ~n449;
  assign n27122 = n2314 & n27121;
  assign n27123 = n184 & n321;
  assign n27124 = n27122 & n27123;
  assign n27125 = n1576 & n4087;
  assign n27126 = n27124 & n27125;
  assign n27127 = n1070 & n4725;
  assign n27128 = n27126 & n27127;
  assign n27129 = n3373 & n27128;
  assign n27130 = n11742 & n27129;
  assign n27132 = n27131 ^ n27130;
  assign n27135 = n27134 ^ n27132;
  assign n27144 = n27143 ^ n27135;
  assign n27153 = n27152 ^ n27144;
  assign n27118 = n27095 ^ n27066;
  assign n27119 = ~n27096 & ~n27118;
  assign n27120 = n27119 ^ n27066;
  assign n27154 = n27153 ^ n27120;
  assign n27161 = n27160 ^ n27154;
  assign n27115 = n27106 ^ n27097;
  assign n27116 = ~n27098 & n27115;
  assign n27117 = n27116 ^ n27106;
  assign n27162 = n27161 ^ n27117;
  assign n27112 = n27047 ^ x23;
  assign n27113 = ~n27108 & ~n27112;
  assign n27114 = n27113 ^ x23;
  assign n27163 = n27162 ^ n27114;
  assign n27180 = n27179 ^ n27163;
  assign n27190 = n27189 ^ n27180;
  assign n27269 = ~n27180 & n27189;
  assign n27249 = n27114 & ~n27117;
  assign n27250 = n27154 & n27160;
  assign n27251 = ~n27249 & n27250;
  assign n27252 = ~n27179 & n27251;
  assign n27253 = n27117 ^ n27114;
  assign n27254 = n27160 ^ n27117;
  assign n27255 = ~n27161 & ~n27254;
  assign n27256 = n27253 & n27255;
  assign n27257 = ~n27252 & ~n27256;
  assign n27258 = ~n27154 & ~n27160;
  assign n27259 = ~n27114 & n27117;
  assign n27261 = n27258 & ~n27259;
  assign n27262 = n27249 & ~n27250;
  assign n27263 = ~n27261 & ~n27262;
  assign n27260 = ~n27258 & n27259;
  assign n27264 = n27263 ^ n27260;
  assign n27265 = ~n27179 & ~n27264;
  assign n27266 = n27265 ^ n27263;
  assign n27267 = n27257 & n27266;
  assign n27238 = n12466 & ~n23879;
  assign n27231 = n3275 & n19649;
  assign n27232 = n3277 & n23052;
  assign n27233 = ~n27231 & ~n27232;
  assign n27234 = x29 & n27233;
  assign n27239 = n23292 & n27234;
  assign n27240 = ~n27238 & ~n27239;
  assign n27235 = n23879 & n27234;
  assign n27236 = n12466 & ~n23292;
  assign n27237 = ~n27235 & ~n27236;
  assign n27241 = n27240 ^ n27237;
  assign n27242 = ~x28 & n27241;
  assign n27243 = n27242 ^ n27240;
  assign n27244 = ~n12476 & n27233;
  assign n27245 = n27244 ^ x29;
  assign n27246 = n27243 & n27245;
  assign n27214 = n1172 & n4906;
  assign n27215 = n4071 & n5091;
  assign n27216 = n27214 & n27215;
  assign n27217 = n2038 & n3122;
  assign n27218 = n2311 & n3372;
  assign n27219 = n27217 & n27218;
  assign n27220 = n27216 & n27219;
  assign n27221 = n12886 & n19519;
  assign n27222 = n27220 & n27221;
  assign n27223 = n2094 & n11518;
  assign n27224 = n12765 & n27223;
  assign n27225 = n3349 & n27224;
  assign n27226 = n27222 & n27225;
  assign n27227 = n13337 & n27226;
  assign n27211 = n27130 ^ n27089;
  assign n27212 = n27131 & ~n27211;
  assign n27213 = n27212 ^ x23;
  assign n27228 = n27227 ^ n27213;
  assign n27203 = n41 & n23468;
  assign n27204 = n91 & n19512;
  assign n27205 = n54 & ~n19439;
  assign n27206 = ~n27204 & ~n27205;
  assign n27207 = ~n27203 & n27206;
  assign n27200 = n41 & ~n19575;
  assign n27201 = n54 & ~n19512;
  assign n27202 = ~n27200 & ~n27201;
  assign n27208 = n27207 ^ n27202;
  assign n27209 = ~x31 & ~n27208;
  assign n27210 = n27209 ^ n27207;
  assign n27229 = n27228 ^ n27210;
  assign n27197 = n27143 ^ n27134;
  assign n27198 = ~n27135 & n27197;
  assign n27199 = n27198 ^ n27143;
  assign n27230 = n27229 ^ n27199;
  assign n27247 = n27246 ^ n27230;
  assign n27194 = ~n3440 & n23495;
  assign n27195 = n27194 ^ x26;
  assign n27191 = n27152 ^ n27120;
  assign n27192 = ~n27153 & n27191;
  assign n27193 = n27192 ^ n27120;
  assign n27196 = n27195 ^ n27193;
  assign n27248 = n27247 ^ n27196;
  assign n27268 = n27267 ^ n27248;
  assign n27270 = n27269 ^ n27268;
  assign n27322 = n27268 & n27269;
  assign n27311 = n44 & n23493;
  assign n27312 = n3280 & n23495;
  assign n27313 = n3277 & ~n23292;
  assign n27314 = n3275 & n23052;
  assign n27315 = ~n27313 & ~n27314;
  assign n27316 = ~n27312 & n27315;
  assign n27317 = ~n27311 & n27316;
  assign n27318 = n27317 ^ x29;
  assign n27301 = ~n54 & n23520;
  assign n27302 = n11234 & ~n27201;
  assign n27303 = ~n27301 & n27302;
  assign n27304 = ~x31 & ~n19649;
  assign n27305 = ~n5354 & n19575;
  assign n27306 = ~n12591 & ~n27305;
  assign n27307 = ~n27304 & n27306;
  assign n27308 = ~n27303 & n27307;
  assign n27293 = n1481 & n3083;
  assign n27294 = n19519 & n27293;
  assign n27295 = ~n755 & ~n3381;
  assign n27296 = n3428 & n27295;
  assign n27297 = n3368 & n27296;
  assign n27298 = n27294 & n27297;
  assign n27299 = n11841 & n27298;
  assign n27291 = n27213 ^ n27210;
  assign n27292 = ~n27228 & n27291;
  assign n27300 = n27299 ^ n27292;
  assign n27309 = n27308 ^ n27300;
  assign n27310 = n27309 ^ x26;
  assign n27319 = n27318 ^ n27310;
  assign n27288 = n27246 ^ n27199;
  assign n27289 = ~n27230 & n27288;
  assign n27290 = n27289 ^ n27246;
  assign n27320 = n27319 ^ n27290;
  assign n27274 = ~n27154 & ~n27259;
  assign n27275 = ~n27248 & ~n27249;
  assign n27276 = ~n27274 & n27275;
  assign n27277 = ~n27252 & ~n27276;
  assign n27278 = ~n27154 & ~n27275;
  assign n27279 = n27248 & ~n27259;
  assign n27280 = n27160 & ~n27279;
  assign n27281 = ~n27278 & n27280;
  assign n27282 = n27179 & ~n27281;
  assign n27283 = ~n27160 & n27278;
  assign n27284 = ~n27279 & ~n27283;
  assign n27285 = ~n27282 & n27284;
  assign n27286 = n27277 & ~n27285;
  assign n27271 = n27247 ^ n27193;
  assign n27272 = n27196 & n27271;
  assign n27273 = n27272 ^ n27247;
  assign n27287 = n27286 ^ n27273;
  assign n27321 = n27320 ^ n27287;
  assign n27323 = n27322 ^ n27321;
  assign n27366 = n27273 & n27320;
  assign n27367 = n27286 & ~n27366;
  assign n27368 = ~n27273 & ~n27320;
  assign n27369 = ~n27367 & ~n27368;
  assign n27370 = ~n27286 & n27366;
  assign n27371 = n27322 & ~n27370;
  assign n27372 = n27369 & ~n27371;
  assign n27373 = n27286 & n27368;
  assign n27374 = n27322 & n27373;
  assign n27375 = ~n27372 & ~n27374;
  assign n27346 = n27318 ^ n27290;
  assign n27347 = n27318 ^ n27308;
  assign n27348 = n27346 & n27347;
  assign n27349 = n27348 ^ n27290;
  assign n27350 = x26 & ~n27349;
  assign n27351 = ~n27290 & n27308;
  assign n27352 = ~n27318 & n27351;
  assign n27353 = n27300 & ~n27352;
  assign n27354 = n27350 & ~n27353;
  assign n27355 = ~x26 & n27300;
  assign n27356 = n27349 & n27355;
  assign n27357 = ~n27300 & n27352;
  assign n27358 = n27290 & ~n27308;
  assign n27359 = x26 & ~n27300;
  assign n27360 = n27318 & ~n27359;
  assign n27361 = n27358 & n27360;
  assign n27362 = ~n27357 & ~n27361;
  assign n27363 = ~n27356 & n27362;
  assign n27364 = ~n27354 & n27363;
  assign n27342 = n44 & ~n23704;
  assign n27343 = n3275 & ~n23292;
  assign n27344 = ~n27342 & ~n27343;
  assign n27337 = n3425 & n3872;
  assign n27336 = x29 ^ x26;
  assign n27338 = n27337 ^ n27336;
  assign n27339 = n27338 ^ n27227;
  assign n27332 = n27299 ^ n27227;
  assign n27333 = ~n27228 & ~n27332;
  assign n27334 = n27291 & n27333;
  assign n27335 = n27334 ^ n27227;
  assign n27340 = n27339 ^ n27335;
  assign n27324 = x31 & n23026;
  assign n27325 = n27324 ^ n23052;
  assign n27326 = n41 & ~n27325;
  assign n27327 = n91 & ~n19649;
  assign n27328 = n3669 & n19575;
  assign n27329 = ~n12591 & ~n27328;
  assign n27330 = ~n27327 & n27329;
  assign n27331 = ~n27326 & n27330;
  assign n27341 = n27340 ^ n27331;
  assign n27345 = n27344 ^ n27341;
  assign n27365 = n27364 ^ n27345;
  assign n27376 = n27375 ^ n27365;
  assign y0 = n23014;
  assign y1 = n23259;
  assign y2 = ~n23489;
  assign y3 = ~n23692;
  assign y4 = n23866;
  assign y5 = ~n24051;
  assign y6 = ~n24228;
  assign y7 = ~n24422;
  assign y8 = n24615;
  assign y9 = ~n24793;
  assign y10 = ~n24964;
  assign y11 = ~n25147;
  assign y12 = n25315;
  assign y13 = n25482;
  assign y14 = ~n25633;
  assign y15 = n25781;
  assign y16 = ~n25926;
  assign y17 = n26056;
  assign y18 = n26189;
  assign y19 = ~n26301;
  assign y20 = n26436;
  assign y21 = ~n26540;
  assign y22 = n26636;
  assign y23 = ~n26737;
  assign y24 = ~n26838;
  assign y25 = ~n26954;
  assign y26 = n27036;
  assign y27 = n27111;
  assign y28 = ~n27190;
  assign y29 = n27270;
  assign y30 = n27323;
  assign y31 = n27376;
endmodule
