module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127;
  wire n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285;
  assign n129 = ~x126 & ~x127;
  assign n130 = ~x125 & n129;
  assign n131 = ~x124 & n130;
  assign n132 = ~x123 & n131;
  assign n133 = x122 & n132;
  assign n134 = ~x122 & n132;
  assign n135 = ~x121 & n134;
  assign n9801 = ~x120 & n135;
  assign n9802 = ~x119 & n9801;
  assign n9803 = ~x118 & n9802;
  assign n136 = ~x118 & ~x119;
  assign n137 = ~x117 & n136;
  assign n138 = ~x116 & ~x120;
  assign n139 = n137 & n138;
  assign n140 = n135 & n139;
  assign n141 = ~x115 & n140;
  assign n9087 = ~x114 & n141;
  assign n142 = ~x111 & ~x112;
  assign n143 = ~x113 & ~x114;
  assign n144 = n142 & n143;
  assign n145 = n141 & n144;
  assign n146 = ~x110 & n145;
  assign n147 = ~x109 & n146;
  assign n148 = ~x104 & ~x105;
  assign n149 = ~x108 & n148;
  assign n150 = ~x106 & ~x107;
  assign n151 = n149 & n150;
  assign n152 = n147 & n151;
  assign n153 = ~x103 & n152;
  assign n154 = ~x102 & n153;
  assign n155 = ~x101 & n154;
  assign n156 = ~x97 & ~x98;
  assign n157 = ~x99 & ~x100;
  assign n158 = n156 & n157;
  assign n159 = ~x96 & n158;
  assign n160 = n155 & n159;
  assign n161 = ~x95 & n160;
  assign n162 = ~x94 & n161;
  assign n163 = ~x93 & n162;
  assign n164 = ~x92 & n163;
  assign n165 = ~x91 & n164;
  assign n166 = ~x90 & n165;
  assign n167 = ~x89 & n166;
  assign n168 = ~x88 & n167;
  assign n169 = ~x85 & ~x86;
  assign n170 = ~x84 & ~x87;
  assign n171 = n169 & n170;
  assign n172 = n168 & n171;
  assign n173 = ~x83 & n172;
  assign n174 = ~x82 & n173;
  assign n175 = ~x81 & n174;
  assign n176 = ~x79 & ~x80;
  assign n177 = n175 & n176;
  assign n178 = ~x78 & n177;
  assign n179 = ~x77 & n178;
  assign n180 = ~x76 & n179;
  assign n181 = ~x75 & n180;
  assign n182 = ~x74 & n181;
  assign n183 = ~x73 & n182;
  assign n184 = ~x71 & ~x72;
  assign n185 = n183 & n184;
  assign n186 = ~x70 & n185;
  assign n187 = ~x69 & n186;
  assign n188 = ~x68 & n187;
  assign n189 = ~x67 & n188;
  assign n190 = ~x63 & x65;
  assign n191 = ~x66 & ~n190;
  assign n192 = n189 & n191;
  assign n193 = ~x61 & x65;
  assign n194 = x62 & ~n193;
  assign n195 = ~n192 & n194;
  assign n196 = x61 & ~x65;
  assign n197 = x64 & ~n196;
  assign n198 = ~x62 & x65;
  assign n199 = ~n197 & ~n198;
  assign n200 = ~n195 & ~n199;
  assign n201 = x64 & ~n198;
  assign n202 = ~x64 & x65;
  assign n203 = ~x66 & ~n202;
  assign n204 = ~n201 & n203;
  assign n205 = n204 ^ x66;
  assign n206 = ~n200 & n205;
  assign n207 = n206 ^ x66;
  assign n208 = n189 & ~n207;
  assign n209 = x63 & ~n208;
  assign n210 = n189 & n209;
  assign n211 = x63 & n204;
  assign n212 = n200 & ~n211;
  assign n213 = ~x63 & x66;
  assign n214 = n189 & ~n213;
  assign n215 = ~n212 & n214;
  assign n216 = x64 & n215;
  assign n217 = n193 & ~n216;
  assign n218 = x65 ^ x60;
  assign n219 = n215 ^ x61;
  assign n220 = n219 ^ x60;
  assign n221 = ~n218 & n220;
  assign n222 = n221 ^ x60;
  assign n223 = x64 & ~n222;
  assign n224 = ~n217 & ~n223;
  assign n225 = n224 ^ x66;
  assign n226 = x65 & n215;
  assign n227 = x64 & n192;
  assign n228 = x62 & ~n227;
  assign n229 = ~n226 & ~n228;
  assign n230 = x64 & ~n192;
  assign n231 = ~n202 & ~n230;
  assign n232 = ~n196 & ~n231;
  assign n233 = n215 & n232;
  assign n234 = n192 & n193;
  assign n235 = ~n233 & ~n234;
  assign n236 = ~n229 & n235;
  assign n237 = n236 ^ n224;
  assign n238 = ~n225 & ~n237;
  assign n239 = n238 ^ x66;
  assign n240 = n210 & ~n239;
  assign n242 = n239 ^ x67;
  assign n243 = n188 & n242;
  assign n244 = n209 & ~n243;
  assign n247 = ~x63 & x67;
  assign n248 = n188 & ~n247;
  assign n249 = ~n239 & n248;
  assign n250 = ~n210 & ~n249;
  assign n251 = x65 & ~n250;
  assign n252 = n216 & ~n251;
  assign n253 = n215 ^ x60;
  assign n254 = n253 ^ x60;
  assign n255 = n218 ^ x60;
  assign n256 = n254 & n255;
  assign n257 = n256 ^ x60;
  assign n258 = x64 & ~n257;
  assign n259 = n258 ^ x65;
  assign n260 = ~n250 & n259;
  assign n261 = ~n252 & ~n260;
  assign n262 = n261 ^ x61;
  assign n263 = n262 ^ x66;
  assign n264 = n250 ^ x60;
  assign n265 = ~x59 & x65;
  assign n266 = ~n264 & ~n265;
  assign n267 = x59 & ~x65;
  assign n268 = x64 & ~n267;
  assign n269 = ~n266 & n268;
  assign n270 = ~x60 & x65;
  assign n271 = x64 & ~n250;
  assign n272 = n270 & ~n271;
  assign n273 = ~n269 & ~n272;
  assign n274 = n273 ^ n262;
  assign n275 = n263 & n274;
  assign n276 = n275 ^ x66;
  assign n277 = n276 ^ x67;
  assign n278 = ~n225 & ~n250;
  assign n279 = n278 ^ n236;
  assign n280 = n279 ^ n276;
  assign n281 = n277 & n280;
  assign n282 = n281 ^ x67;
  assign n283 = n282 ^ x68;
  assign n284 = n244 & n283;
  assign n285 = n187 & n284;
  assign n286 = n285 ^ n244;
  assign n245 = x69 & ~n244;
  assign n246 = n186 & ~n245;
  assign n287 = ~x69 & n286;
  assign n288 = x64 & ~x65;
  assign n289 = n288 ^ x65;
  assign n290 = n250 & n289;
  assign n291 = n290 ^ x65;
  assign n292 = ~x59 & n291;
  assign n293 = ~n202 & ~n292;
  assign n294 = x59 & ~n251;
  assign n295 = x65 & n294;
  assign n296 = n293 & ~n295;
  assign n297 = n296 ^ n271;
  assign n298 = n296 ^ n294;
  assign n299 = n282 ^ n244;
  assign n300 = n283 & n299;
  assign n301 = n300 ^ x68;
  assign n302 = n187 & ~n301;
  assign n303 = n302 ^ n296;
  assign n304 = n296 & n303;
  assign n305 = n304 ^ n296;
  assign n306 = n298 & n305;
  assign n307 = n306 ^ n304;
  assign n308 = n307 ^ n296;
  assign n309 = n308 ^ n302;
  assign n310 = ~n297 & n309;
  assign n311 = n310 ^ n271;
  assign n312 = n311 ^ x60;
  assign n313 = n312 ^ x66;
  assign n314 = x65 ^ x59;
  assign n315 = n314 ^ n302;
  assign n316 = n302 ^ x65;
  assign n317 = x65 ^ x58;
  assign n318 = n317 ^ n302;
  assign n319 = ~n302 & n318;
  assign n320 = n319 ^ n302;
  assign n321 = ~n316 & ~n320;
  assign n322 = n321 ^ n319;
  assign n323 = n322 ^ n302;
  assign n324 = n323 ^ n317;
  assign n325 = n315 & n324;
  assign n326 = n325 ^ x58;
  assign n327 = x64 & ~n326;
  assign n328 = x64 & n302;
  assign n329 = n265 & ~n328;
  assign n330 = ~n327 & ~n329;
  assign n331 = n330 ^ n312;
  assign n332 = ~n313 & ~n331;
  assign n333 = n332 ^ x66;
  assign n334 = n333 ^ x67;
  assign n335 = n273 ^ x66;
  assign n336 = n302 & ~n335;
  assign n337 = n336 ^ n262;
  assign n338 = n337 ^ n333;
  assign n339 = n334 & ~n338;
  assign n340 = n339 ^ x67;
  assign n341 = n340 ^ x68;
  assign n342 = n277 & n302;
  assign n343 = n342 ^ n279;
  assign n344 = n343 ^ n340;
  assign n345 = n341 & ~n344;
  assign n346 = n345 ^ n340;
  assign n347 = ~n287 & n346;
  assign n348 = n246 & ~n347;
  assign n349 = n286 & ~n348;
  assign n350 = ~n240 & ~n349;
  assign n351 = ~x72 & n183;
  assign n352 = ~n350 & ~n351;
  assign n353 = x65 & n348;
  assign n354 = ~n328 & ~n353;
  assign n355 = x65 & n302;
  assign n356 = x58 & ~n355;
  assign n357 = ~n354 & n356;
  assign n358 = n289 & ~n302;
  assign n359 = n358 ^ x65;
  assign n360 = ~x58 & n359;
  assign n361 = ~n202 & ~n360;
  assign n362 = n361 ^ n328;
  assign n363 = n348 & ~n362;
  assign n364 = n363 ^ n328;
  assign n365 = ~n357 & ~n364;
  assign n366 = n365 ^ x59;
  assign n367 = n366 ^ x66;
  assign n370 = x58 & ~x65;
  assign n371 = ~x57 & ~n370;
  assign n368 = x57 & ~x65;
  assign n369 = x58 & ~n368;
  assign n372 = n371 ^ n369;
  assign n373 = n369 ^ x65;
  assign n374 = n369 ^ n348;
  assign n375 = ~n369 & ~n374;
  assign n376 = n375 ^ n369;
  assign n377 = ~n373 & ~n376;
  assign n378 = n377 ^ n375;
  assign n379 = n378 ^ n369;
  assign n380 = n379 ^ n348;
  assign n381 = n372 & ~n380;
  assign n382 = n381 ^ n371;
  assign n383 = x64 & n382;
  assign n384 = x64 & n348;
  assign n385 = ~x58 & x65;
  assign n386 = ~n384 & n385;
  assign n387 = ~n383 & ~n386;
  assign n388 = n387 ^ n366;
  assign n389 = n367 & n388;
  assign n390 = n389 ^ x66;
  assign n391 = n390 ^ x67;
  assign n392 = n330 ^ x66;
  assign n393 = n348 & ~n392;
  assign n394 = n393 ^ n312;
  assign n395 = n394 ^ n390;
  assign n396 = n391 & n395;
  assign n397 = n396 ^ x67;
  assign n398 = n397 ^ x68;
  assign n399 = n334 & n348;
  assign n400 = n399 ^ n337;
  assign n401 = n400 ^ n397;
  assign n402 = n398 & ~n401;
  assign n403 = n402 ^ x68;
  assign n404 = n403 ^ x69;
  assign n405 = n341 & n348;
  assign n406 = n405 ^ n343;
  assign n407 = n406 ^ n403;
  assign n408 = n404 & n407;
  assign n409 = n408 ^ x69;
  assign n410 = n409 ^ x70;
  assign n411 = n409 ^ n350;
  assign n412 = n410 & n411;
  assign n413 = n412 ^ n409;
  assign n414 = n185 & ~n413;
  assign n415 = ~n350 & ~n414;
  assign n416 = n415 ^ x72;
  assign n417 = n416 ^ n415;
  assign n418 = x70 & ~x71;
  assign n419 = ~n350 & n418;
  assign n420 = n409 & n419;
  assign n421 = x71 & n350;
  assign n424 = ~x56 & ~n368;
  assign n422 = x56 & ~x65;
  assign n423 = x57 & ~n422;
  assign n425 = n424 ^ n423;
  assign n426 = n423 ^ x65;
  assign n427 = n423 ^ n414;
  assign n428 = ~n423 & ~n427;
  assign n429 = n428 ^ n423;
  assign n430 = ~n426 & ~n429;
  assign n431 = n430 ^ n428;
  assign n432 = n431 ^ n423;
  assign n433 = n432 ^ n414;
  assign n434 = n425 & ~n433;
  assign n435 = n434 ^ n424;
  assign n436 = x64 & n435;
  assign n437 = x64 & n414;
  assign n438 = ~x57 & x65;
  assign n439 = ~n437 & n438;
  assign n440 = ~n436 & ~n439;
  assign n441 = n440 ^ x66;
  assign n442 = x65 & n414;
  assign n443 = x57 & ~n353;
  assign n444 = n442 & n443;
  assign n445 = n289 & ~n348;
  assign n446 = n445 ^ x65;
  assign n447 = ~x57 & n446;
  assign n448 = ~n202 & ~n447;
  assign n449 = n414 & ~n448;
  assign n450 = ~n444 & ~n449;
  assign n451 = n414 & ~n443;
  assign n452 = n384 & ~n451;
  assign n453 = n450 & ~n452;
  assign n454 = n453 ^ x58;
  assign n455 = n454 ^ n440;
  assign n456 = ~n441 & n455;
  assign n457 = n456 ^ x66;
  assign n458 = n457 ^ x67;
  assign n459 = n387 ^ x66;
  assign n460 = n414 & ~n459;
  assign n461 = n460 ^ n366;
  assign n462 = n461 ^ n457;
  assign n463 = n458 & ~n462;
  assign n464 = n463 ^ x67;
  assign n465 = n464 ^ x68;
  assign n466 = n391 & n414;
  assign n467 = n466 ^ n394;
  assign n468 = n467 ^ n464;
  assign n469 = n465 & n468;
  assign n470 = n469 ^ x68;
  assign n471 = n470 ^ x69;
  assign n472 = n398 & n414;
  assign n473 = n472 ^ n400;
  assign n474 = n473 ^ n470;
  assign n475 = n471 & ~n474;
  assign n476 = n475 ^ x69;
  assign n477 = n476 ^ x70;
  assign n478 = n404 & n414;
  assign n479 = n478 ^ n406;
  assign n480 = n479 ^ n476;
  assign n481 = n477 & ~n480;
  assign n482 = n481 ^ n476;
  assign n483 = ~n421 & ~n482;
  assign n484 = ~n420 & ~n483;
  assign n485 = n351 & ~n484;
  assign n486 = n415 & ~n485;
  assign n487 = ~n240 & ~n486;
  assign n488 = n487 ^ n415;
  assign n489 = ~n417 & n488;
  assign n490 = n489 ^ n415;
  assign n491 = n183 & n490;
  assign n492 = x65 ^ x56;
  assign n493 = n492 ^ n485;
  assign n494 = n485 ^ x65;
  assign n495 = x65 ^ x55;
  assign n496 = n495 ^ n485;
  assign n497 = ~n485 & n496;
  assign n498 = n497 ^ n485;
  assign n499 = ~n494 & ~n498;
  assign n500 = n499 ^ n497;
  assign n501 = n500 ^ n485;
  assign n502 = n501 ^ n495;
  assign n503 = n493 & n502;
  assign n504 = n503 ^ x55;
  assign n505 = x64 & ~n504;
  assign n506 = x64 & n485;
  assign n507 = ~x56 & x65;
  assign n508 = ~n506 & n507;
  assign n509 = ~n505 & ~n508;
  assign n510 = n509 ^ x66;
  assign n511 = x65 & n485;
  assign n512 = x56 & ~n442;
  assign n513 = n511 & n512;
  assign n514 = n289 & ~n414;
  assign n515 = n514 ^ x65;
  assign n516 = ~x56 & n515;
  assign n517 = ~n202 & ~n516;
  assign n518 = n485 & ~n517;
  assign n519 = ~n513 & ~n518;
  assign n520 = n485 & ~n512;
  assign n521 = n437 & ~n520;
  assign n522 = n519 & ~n521;
  assign n523 = n522 ^ x57;
  assign n524 = n523 ^ n509;
  assign n525 = ~n510 & n524;
  assign n526 = n525 ^ x66;
  assign n527 = n526 ^ x67;
  assign n528 = ~n441 & n485;
  assign n529 = n528 ^ n454;
  assign n530 = n529 ^ n526;
  assign n531 = n527 & ~n530;
  assign n532 = n531 ^ x67;
  assign n533 = n532 ^ x68;
  assign n534 = n458 & n485;
  assign n535 = n534 ^ n461;
  assign n536 = n535 ^ n532;
  assign n537 = n533 & ~n536;
  assign n538 = n537 ^ x68;
  assign n539 = n538 ^ x69;
  assign n540 = n465 & n485;
  assign n541 = n540 ^ n467;
  assign n542 = n541 ^ n538;
  assign n543 = n539 & n542;
  assign n544 = n543 ^ x69;
  assign n545 = n544 ^ x70;
  assign n546 = n471 & n485;
  assign n547 = n546 ^ n473;
  assign n548 = n547 ^ n544;
  assign n549 = n545 & ~n548;
  assign n550 = n549 ^ x70;
  assign n551 = n550 ^ x71;
  assign n552 = n477 & n485;
  assign n553 = n552 ^ n479;
  assign n554 = n553 ^ n550;
  assign n555 = n551 & ~n554;
  assign n556 = n555 ^ n550;
  assign n557 = n491 & ~n556;
  assign n558 = n352 & ~n557;
  assign n559 = n415 & n484;
  assign n560 = ~n240 & ~n559;
  assign n561 = n351 & ~n560;
  assign n562 = ~n557 & ~n561;
  assign n563 = n539 & ~n562;
  assign n564 = n563 ^ n541;
  assign n565 = ~x70 & n564;
  assign n566 = x65 & ~n562;
  assign n567 = x55 & ~n511;
  assign n568 = n566 & n567;
  assign n569 = n289 & ~n485;
  assign n570 = n569 ^ x65;
  assign n571 = ~x55 & n570;
  assign n572 = ~n202 & ~n571;
  assign n573 = ~n562 & ~n572;
  assign n574 = ~n568 & ~n573;
  assign n575 = ~n562 & ~n567;
  assign n576 = n506 & ~n575;
  assign n577 = n574 & ~n576;
  assign n578 = n577 ^ x56;
  assign n579 = n578 ^ x66;
  assign n580 = ~x65 & ~n562;
  assign n581 = x55 & ~x65;
  assign n582 = ~x54 & x64;
  assign n583 = ~n581 & n582;
  assign n584 = ~n580 & n583;
  assign n586 = x64 & ~n562;
  assign n585 = ~x55 & x65;
  assign n587 = n586 ^ n585;
  assign n588 = n587 ^ n585;
  assign n589 = x54 & n581;
  assign n590 = n589 ^ x55;
  assign n591 = n590 ^ n585;
  assign n592 = n588 & n591;
  assign n593 = n592 ^ n585;
  assign n594 = ~n584 & ~n593;
  assign n595 = n594 ^ n578;
  assign n596 = n579 & n595;
  assign n597 = n596 ^ x66;
  assign n598 = n597 ^ x67;
  assign n599 = ~n510 & ~n562;
  assign n600 = n599 ^ n523;
  assign n601 = n600 ^ n597;
  assign n602 = n598 & ~n601;
  assign n603 = n602 ^ x67;
  assign n604 = n603 ^ x68;
  assign n605 = n527 & ~n562;
  assign n606 = n605 ^ n529;
  assign n607 = n606 ^ n603;
  assign n608 = n604 & ~n607;
  assign n609 = n608 ^ x68;
  assign n610 = n609 ^ x69;
  assign n611 = n533 & ~n562;
  assign n612 = n611 ^ n535;
  assign n613 = n612 ^ n609;
  assign n614 = n610 & ~n613;
  assign n615 = n614 ^ x69;
  assign n616 = ~n565 & n615;
  assign n617 = n545 & ~n562;
  assign n618 = n617 ^ n547;
  assign n619 = x70 & x71;
  assign n620 = ~n618 & ~n619;
  assign n621 = n616 & ~n620;
  assign n622 = x71 & ~n564;
  assign n623 = n615 & n622;
  assign n624 = n618 ^ x71;
  assign n625 = x70 & ~n564;
  assign n626 = n625 ^ n618;
  assign n627 = n624 & ~n626;
  assign n628 = n627 ^ x71;
  assign n629 = ~n623 & ~n628;
  assign n630 = ~n621 & n629;
  assign n631 = n551 & ~n562;
  assign n632 = n631 ^ n553;
  assign n633 = ~x72 & n632;
  assign n634 = ~x73 & n558;
  assign n635 = ~n633 & ~n634;
  assign n636 = ~n630 & n635;
  assign n637 = x72 & ~n634;
  assign n638 = ~n632 & n637;
  assign n639 = x73 & ~n558;
  assign n640 = n182 & ~n639;
  assign n641 = ~n638 & n640;
  assign n642 = ~n636 & n641;
  assign n643 = n558 & ~n642;
  assign n644 = ~n240 & ~n643;
  assign n645 = n182 & ~n644;
  assign n646 = x74 & n644;
  assign n647 = n181 & ~n646;
  assign n648 = x65 & n642;
  assign n649 = x54 & ~n566;
  assign n650 = n648 & n649;
  assign n651 = n289 & n562;
  assign n652 = n651 ^ x65;
  assign n653 = ~x54 & n652;
  assign n654 = ~n202 & ~n653;
  assign n655 = n642 & ~n654;
  assign n656 = ~n650 & ~n655;
  assign n657 = n642 & ~n649;
  assign n658 = n586 & ~n657;
  assign n659 = n656 & ~n658;
  assign n660 = n659 ^ x55;
  assign n661 = n660 ^ x66;
  assign n662 = ~x53 & ~x54;
  assign n663 = ~n642 & n662;
  assign n664 = ~x53 & x65;
  assign n665 = ~n663 & ~n664;
  assign n666 = x64 & ~n665;
  assign n667 = x64 & n642;
  assign n668 = n667 ^ x54;
  assign n669 = n667 ^ x65;
  assign n670 = n669 ^ x65;
  assign n671 = x53 & ~x65;
  assign n672 = n671 ^ x65;
  assign n673 = n670 & ~n672;
  assign n674 = n673 ^ x65;
  assign n675 = ~n668 & n674;
  assign n676 = ~n666 & ~n675;
  assign n677 = n676 ^ n660;
  assign n678 = n661 & n677;
  assign n679 = n678 ^ x66;
  assign n680 = n679 ^ x67;
  assign n681 = n594 ^ x66;
  assign n682 = n642 & ~n681;
  assign n683 = n682 ^ n578;
  assign n684 = n683 ^ n679;
  assign n685 = n680 & ~n684;
  assign n686 = n685 ^ x67;
  assign n687 = n686 ^ x68;
  assign n688 = n598 & n642;
  assign n689 = n688 ^ n600;
  assign n690 = n689 ^ n686;
  assign n691 = n687 & ~n690;
  assign n692 = n691 ^ x68;
  assign n693 = n692 ^ x69;
  assign n694 = n604 & n642;
  assign n695 = n694 ^ n606;
  assign n696 = n695 ^ n692;
  assign n697 = n693 & ~n696;
  assign n698 = n697 ^ x69;
  assign n699 = n698 ^ x70;
  assign n700 = n610 & n642;
  assign n701 = n700 ^ n612;
  assign n702 = n701 ^ n698;
  assign n703 = n699 & ~n702;
  assign n704 = n703 ^ x70;
  assign n705 = n704 ^ x71;
  assign n706 = n615 ^ x70;
  assign n707 = n642 & n706;
  assign n708 = n707 ^ n564;
  assign n709 = n708 ^ n704;
  assign n710 = n705 & n709;
  assign n711 = n710 ^ x71;
  assign n712 = n711 ^ x72;
  assign n713 = ~n616 & ~n625;
  assign n714 = n713 ^ x71;
  assign n715 = n642 & ~n714;
  assign n716 = n715 ^ n618;
  assign n717 = n716 ^ n711;
  assign n718 = n712 & ~n717;
  assign n719 = n718 ^ x72;
  assign n720 = n719 ^ x73;
  assign n721 = n630 ^ x72;
  assign n722 = n642 & ~n721;
  assign n723 = n722 ^ n632;
  assign n724 = n723 ^ n719;
  assign n725 = n720 & ~n724;
  assign n726 = n725 ^ n719;
  assign n727 = n647 & ~n726;
  assign n728 = ~n645 & ~n727;
  assign n729 = ~x65 & ~n728;
  assign n730 = ~x52 & x64;
  assign n731 = ~n671 & n730;
  assign n732 = ~n729 & n731;
  assign n733 = x64 & ~n728;
  assign n734 = x52 & ~x65;
  assign n735 = x53 & ~n734;
  assign n736 = n735 ^ n664;
  assign n737 = n733 & n736;
  assign n738 = n737 ^ n664;
  assign n739 = ~n732 & ~n738;
  assign n740 = n739 ^ x66;
  assign n741 = n289 & ~n642;
  assign n742 = n741 ^ x65;
  assign n743 = ~x53 & n742;
  assign n744 = x53 & x65;
  assign n745 = ~n642 & n744;
  assign n746 = ~n202 & ~n745;
  assign n747 = ~n743 & n746;
  assign n748 = n747 ^ n667;
  assign n749 = n747 ^ n671;
  assign n750 = n747 ^ n728;
  assign n751 = n747 & ~n750;
  assign n752 = n751 ^ n747;
  assign n753 = n749 & n752;
  assign n754 = n753 ^ n751;
  assign n755 = n754 ^ n747;
  assign n756 = n755 ^ n728;
  assign n757 = ~n748 & ~n756;
  assign n758 = n757 ^ n667;
  assign n759 = n758 ^ x54;
  assign n760 = n759 ^ n739;
  assign n761 = ~n740 & ~n760;
  assign n762 = n761 ^ x66;
  assign n763 = n762 ^ x67;
  assign n764 = n676 ^ x66;
  assign n765 = ~n728 & ~n764;
  assign n766 = n765 ^ n660;
  assign n767 = n766 ^ n762;
  assign n768 = n763 & ~n767;
  assign n769 = n768 ^ x67;
  assign n770 = n769 ^ x68;
  assign n771 = n680 & ~n728;
  assign n772 = n771 ^ n683;
  assign n773 = n772 ^ n769;
  assign n774 = n770 & ~n773;
  assign n775 = n774 ^ x68;
  assign n776 = n775 ^ x69;
  assign n777 = n687 & ~n728;
  assign n778 = n777 ^ n689;
  assign n779 = n778 ^ n775;
  assign n780 = n776 & ~n779;
  assign n781 = n780 ^ x69;
  assign n782 = n781 ^ x70;
  assign n783 = n693 & ~n728;
  assign n784 = n783 ^ n695;
  assign n785 = n784 ^ n781;
  assign n786 = n782 & ~n785;
  assign n787 = n786 ^ x70;
  assign n788 = n787 ^ x71;
  assign n789 = n699 & ~n728;
  assign n790 = n789 ^ n701;
  assign n791 = n790 ^ n787;
  assign n792 = n788 & ~n791;
  assign n793 = n792 ^ x71;
  assign n794 = n793 ^ x72;
  assign n795 = n705 & ~n728;
  assign n796 = n795 ^ n708;
  assign n797 = n796 ^ n793;
  assign n798 = n794 & n797;
  assign n799 = n798 ^ x72;
  assign n800 = n799 ^ x73;
  assign n801 = n712 & ~n728;
  assign n802 = n801 ^ n716;
  assign n803 = n802 ^ n799;
  assign n804 = n800 & ~n803;
  assign n805 = n804 ^ x73;
  assign n806 = n805 ^ x74;
  assign n807 = n720 & ~n728;
  assign n808 = n807 ^ n723;
  assign n809 = n808 ^ n805;
  assign n810 = n806 & n809;
  assign n811 = n810 ^ x74;
  assign n812 = x75 & n811;
  assign n813 = n180 & ~n812;
  assign n814 = ~n240 & ~n728;
  assign n815 = ~n644 & ~n814;
  assign n816 = ~n813 & n815;
  assign n817 = n811 ^ x75;
  assign n818 = n815 ^ x75;
  assign n819 = n817 & ~n818;
  assign n820 = n819 ^ x75;
  assign n821 = n180 & ~n820;
  assign n822 = n806 & n821;
  assign n823 = n822 ^ n808;
  assign n824 = ~x75 & n823;
  assign n825 = ~x76 & n816;
  assign n826 = ~n824 & ~n825;
  assign n827 = ~x51 & x64;
  assign n828 = n827 ^ x65;
  assign n829 = n821 ^ x52;
  assign n830 = n829 ^ n827;
  assign n833 = n830 ^ n821;
  assign n834 = n833 ^ n830;
  assign n831 = n830 ^ x64;
  assign n832 = n831 ^ n830;
  assign n835 = n834 ^ n832;
  assign n836 = n830 ^ n827;
  assign n837 = n836 ^ n830;
  assign n838 = n837 ^ n834;
  assign n839 = n834 & ~n838;
  assign n840 = n839 ^ n834;
  assign n841 = ~n835 & n840;
  assign n842 = n841 ^ n839;
  assign n843 = n842 ^ n830;
  assign n844 = n843 ^ n834;
  assign n845 = n828 & n844;
  assign n846 = n845 ^ x65;
  assign n847 = n846 ^ x66;
  assign n848 = x52 & n733;
  assign n849 = n728 & n730;
  assign n850 = n849 ^ x65;
  assign n851 = ~n848 & n850;
  assign n852 = n851 ^ n733;
  assign n853 = n851 ^ n734;
  assign n854 = n851 ^ n821;
  assign n855 = ~n851 & ~n854;
  assign n856 = n855 ^ n851;
  assign n857 = ~n853 & ~n856;
  assign n858 = n857 ^ n855;
  assign n859 = n858 ^ n851;
  assign n860 = n859 ^ n821;
  assign n861 = n852 & ~n860;
  assign n862 = n861 ^ n733;
  assign n863 = n862 ^ x53;
  assign n864 = n863 ^ n846;
  assign n865 = n847 & n864;
  assign n866 = n865 ^ x66;
  assign n867 = n866 ^ x67;
  assign n868 = ~n740 & n821;
  assign n869 = n868 ^ n759;
  assign n870 = n869 ^ n866;
  assign n871 = n867 & n870;
  assign n872 = n871 ^ x67;
  assign n873 = n872 ^ x68;
  assign n874 = n763 & n821;
  assign n875 = n874 ^ n766;
  assign n876 = n875 ^ n872;
  assign n877 = n873 & ~n876;
  assign n878 = n877 ^ x68;
  assign n879 = n878 ^ x69;
  assign n880 = n770 & n821;
  assign n881 = n880 ^ n772;
  assign n882 = n881 ^ n878;
  assign n883 = n879 & ~n882;
  assign n884 = n883 ^ x69;
  assign n885 = n884 ^ x70;
  assign n886 = n776 & n821;
  assign n887 = n886 ^ n778;
  assign n888 = n887 ^ n884;
  assign n889 = n885 & ~n888;
  assign n890 = n889 ^ x70;
  assign n891 = n890 ^ x71;
  assign n892 = n782 & n821;
  assign n893 = n892 ^ n784;
  assign n894 = n893 ^ n890;
  assign n895 = n891 & ~n894;
  assign n896 = n895 ^ x71;
  assign n897 = n896 ^ x72;
  assign n898 = n788 & n821;
  assign n899 = n898 ^ n790;
  assign n900 = n899 ^ n896;
  assign n901 = n897 & ~n900;
  assign n902 = n901 ^ x72;
  assign n903 = n902 ^ x73;
  assign n904 = n794 & n821;
  assign n905 = n904 ^ n796;
  assign n906 = n905 ^ n902;
  assign n907 = n903 & n906;
  assign n908 = n907 ^ x73;
  assign n909 = n908 ^ x74;
  assign n910 = n800 & n821;
  assign n911 = n910 ^ n802;
  assign n912 = n911 ^ n908;
  assign n913 = n909 & ~n912;
  assign n914 = n913 ^ x74;
  assign n915 = n826 & n914;
  assign n916 = x75 & ~n825;
  assign n917 = ~n823 & n916;
  assign n918 = x76 & ~n815;
  assign n919 = n179 & ~n918;
  assign n920 = ~n917 & n919;
  assign n921 = ~n915 & n920;
  assign n922 = n816 & ~n921;
  assign n923 = ~n178 & n922;
  assign n924 = ~n240 & ~n922;
  assign n925 = ~x77 & ~n924;
  assign n926 = x77 & n924;
  assign n927 = ~x50 & n827;
  assign n928 = ~n921 & n927;
  assign n929 = ~x50 & x65;
  assign n930 = x64 & n929;
  assign n931 = ~n928 & ~n930;
  assign n934 = x64 & n921;
  assign n932 = x50 & ~x65;
  assign n933 = x51 & ~n932;
  assign n935 = n934 ^ n933;
  assign n936 = n935 ^ n933;
  assign n937 = ~x51 & x65;
  assign n938 = n937 ^ n933;
  assign n939 = ~n936 & n938;
  assign n940 = n939 ^ n933;
  assign n941 = n931 & ~n940;
  assign n942 = n941 ^ x66;
  assign n950 = x64 & n821;
  assign n943 = n821 ^ x65;
  assign n944 = n827 & ~n943;
  assign n945 = ~n202 & ~n944;
  assign n946 = x65 & n821;
  assign n947 = x51 & ~n946;
  assign n948 = x65 & n947;
  assign n949 = n945 & ~n948;
  assign n951 = n950 ^ n949;
  assign n952 = n949 ^ n947;
  assign n953 = n949 ^ n921;
  assign n954 = n949 & n953;
  assign n955 = n954 ^ n949;
  assign n956 = n952 & n955;
  assign n957 = n956 ^ n954;
  assign n958 = n957 ^ n949;
  assign n959 = n958 ^ n921;
  assign n960 = ~n951 & n959;
  assign n961 = n960 ^ n950;
  assign n962 = n961 ^ x52;
  assign n963 = n962 ^ n941;
  assign n964 = ~n942 & ~n963;
  assign n965 = n964 ^ x66;
  assign n966 = n965 ^ x67;
  assign n967 = n847 & n921;
  assign n968 = n967 ^ n863;
  assign n969 = n968 ^ n965;
  assign n970 = n966 & n969;
  assign n971 = n970 ^ x67;
  assign n972 = n971 ^ x68;
  assign n973 = n867 & n921;
  assign n974 = n973 ^ n869;
  assign n975 = n974 ^ n971;
  assign n976 = n972 & n975;
  assign n977 = n976 ^ x68;
  assign n978 = n977 ^ x69;
  assign n979 = n873 & n921;
  assign n980 = n979 ^ n875;
  assign n981 = n980 ^ n977;
  assign n982 = n978 & ~n981;
  assign n983 = n982 ^ x69;
  assign n984 = n983 ^ x70;
  assign n985 = n879 & n921;
  assign n986 = n985 ^ n881;
  assign n987 = n986 ^ n983;
  assign n988 = n984 & ~n987;
  assign n989 = n988 ^ x70;
  assign n990 = n989 ^ x71;
  assign n991 = n885 & n921;
  assign n992 = n991 ^ n887;
  assign n993 = n992 ^ n989;
  assign n994 = n990 & ~n993;
  assign n995 = n994 ^ x71;
  assign n996 = n995 ^ x72;
  assign n997 = n891 & n921;
  assign n998 = n997 ^ n893;
  assign n999 = n998 ^ n995;
  assign n1000 = n996 & ~n999;
  assign n1001 = n1000 ^ x72;
  assign n1002 = n1001 ^ x73;
  assign n1003 = n897 & n921;
  assign n1004 = n1003 ^ n899;
  assign n1005 = n1004 ^ n1001;
  assign n1006 = n1002 & ~n1005;
  assign n1007 = n1006 ^ x73;
  assign n1008 = n1007 ^ x74;
  assign n1009 = n903 & n921;
  assign n1010 = n1009 ^ n905;
  assign n1011 = n1010 ^ n1007;
  assign n1012 = n1008 & n1011;
  assign n1013 = n1012 ^ x74;
  assign n1014 = n1013 ^ x75;
  assign n1015 = n909 & n921;
  assign n1016 = n1015 ^ n911;
  assign n1017 = n1016 ^ n1013;
  assign n1018 = n1014 & ~n1017;
  assign n1019 = n1018 ^ x75;
  assign n1020 = n1019 ^ x76;
  assign n1021 = n914 ^ x75;
  assign n1022 = n921 & n1021;
  assign n1023 = n1022 ^ n823;
  assign n1024 = n1023 ^ n1019;
  assign n1025 = n1020 & ~n1024;
  assign n1026 = n1025 ^ n1019;
  assign n1027 = ~n926 & ~n1026;
  assign n1028 = ~n925 & ~n1027;
  assign n1029 = n178 & ~n1028;
  assign n1030 = n922 & ~n1029;
  assign n1031 = ~n240 & ~n1030;
  assign n1032 = n1031 ^ x78;
  assign n1033 = n177 & n1032;
  assign n1034 = ~x49 & x64;
  assign n1035 = n1029 ^ x50;
  assign n1036 = n1034 & ~n1035;
  assign n1037 = x64 & x65;
  assign n1038 = x50 & n1037;
  assign n1039 = n1038 ^ n929;
  assign n1040 = n1029 & n1039;
  assign n1041 = n1040 ^ n929;
  assign n1042 = ~n1036 & ~n1041;
  assign n1043 = x65 & n1034;
  assign n1044 = ~x50 & n202;
  assign n1045 = ~n1043 & ~n1044;
  assign n1046 = n1042 & n1045;
  assign n1047 = n1046 ^ x66;
  assign n1048 = x65 & n178;
  assign n1049 = n1048 ^ n288;
  assign n1050 = n1049 ^ n288;
  assign n1051 = n1028 ^ n288;
  assign n1052 = n1051 ^ n288;
  assign n1053 = n1050 & ~n1052;
  assign n1054 = n1053 ^ n288;
  assign n1055 = ~n921 & n1054;
  assign n1056 = n1055 ^ n288;
  assign n1057 = x50 & n1056;
  assign n1058 = ~n288 & ~n921;
  assign n1059 = ~x50 & ~n1058;
  assign n1060 = ~n202 & ~n1059;
  assign n1061 = ~x65 & n921;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = n1062 ^ n934;
  assign n1064 = n1029 & n1063;
  assign n1065 = n1064 ^ n934;
  assign n1066 = ~n1057 & ~n1065;
  assign n1067 = n1066 ^ x51;
  assign n1068 = n1067 ^ n1046;
  assign n1069 = ~n1047 & n1068;
  assign n1070 = n1069 ^ x66;
  assign n1071 = n1070 ^ x67;
  assign n1072 = ~n942 & n1029;
  assign n1073 = n1072 ^ n962;
  assign n1074 = n1073 ^ n1070;
  assign n1075 = n1071 & n1074;
  assign n1076 = n1075 ^ x67;
  assign n1077 = n1076 ^ x68;
  assign n1078 = n966 & n1029;
  assign n1079 = n1078 ^ n968;
  assign n1080 = n1079 ^ n1076;
  assign n1081 = n1077 & n1080;
  assign n1082 = n1081 ^ x68;
  assign n1083 = n1082 ^ x69;
  assign n1084 = n972 & n1029;
  assign n1085 = n1084 ^ n974;
  assign n1086 = n1085 ^ n1082;
  assign n1087 = n1083 & n1086;
  assign n1088 = n1087 ^ x69;
  assign n1089 = n1088 ^ x70;
  assign n1090 = n978 & n1029;
  assign n1091 = n1090 ^ n980;
  assign n1092 = n1091 ^ n1088;
  assign n1093 = n1089 & ~n1092;
  assign n1094 = n1093 ^ x70;
  assign n1095 = n1094 ^ x71;
  assign n1096 = n984 & n1029;
  assign n1097 = n1096 ^ n986;
  assign n1098 = n1097 ^ n1094;
  assign n1099 = n1095 & ~n1098;
  assign n1100 = n1099 ^ x71;
  assign n1101 = n1100 ^ x72;
  assign n1102 = n990 & n1029;
  assign n1103 = n1102 ^ n992;
  assign n1104 = n1103 ^ n1100;
  assign n1105 = n1101 & ~n1104;
  assign n1106 = n1105 ^ x72;
  assign n1107 = n1106 ^ x73;
  assign n1108 = n996 & n1029;
  assign n1109 = n1108 ^ n998;
  assign n1110 = n1109 ^ n1106;
  assign n1111 = n1107 & ~n1110;
  assign n1112 = n1111 ^ x73;
  assign n1113 = n1112 ^ x74;
  assign n1114 = n1002 & n1029;
  assign n1115 = n1114 ^ n1004;
  assign n1116 = n1115 ^ n1112;
  assign n1117 = n1113 & ~n1116;
  assign n1118 = n1117 ^ x74;
  assign n1119 = n1118 ^ x75;
  assign n1120 = n1008 & n1029;
  assign n1121 = n1120 ^ n1010;
  assign n1122 = n1121 ^ n1118;
  assign n1123 = n1119 & n1122;
  assign n1124 = n1123 ^ x75;
  assign n1125 = n1124 ^ x76;
  assign n1126 = n1014 & n1029;
  assign n1127 = n1126 ^ n1016;
  assign n1128 = n1127 ^ n1124;
  assign n1129 = n1125 & ~n1128;
  assign n1130 = n1129 ^ x76;
  assign n1131 = n1130 ^ x77;
  assign n1132 = n1020 & n1029;
  assign n1133 = n1132 ^ n1023;
  assign n1134 = n1133 ^ n1130;
  assign n1135 = n1131 & ~n1134;
  assign n1136 = n1135 ^ n1130;
  assign n1137 = n1033 & ~n1136;
  assign n1138 = n923 & ~n1137;
  assign n1139 = n178 & ~n1031;
  assign n1140 = ~n1137 & ~n1139;
  assign n1141 = n1131 & ~n1140;
  assign n1142 = n1141 ^ n1133;
  assign n1143 = ~x78 & n1142;
  assign n1144 = ~n240 & ~n1138;
  assign n1145 = ~x79 & ~n1144;
  assign n1146 = ~n1143 & ~n1145;
  assign n1147 = ~x48 & x64;
  assign n1148 = x64 & ~n1140;
  assign n1149 = n1148 ^ x49;
  assign n1150 = ~n1147 & n1149;
  assign n1151 = x65 & n1150;
  assign n1152 = n1151 ^ x65;
  assign n1153 = n1140 ^ x49;
  assign n1154 = n1147 & n1153;
  assign n1155 = ~n1152 & ~n1154;
  assign n1156 = n1155 ^ x66;
  assign n1157 = ~x49 & ~n1140;
  assign n1158 = x64 & n1029;
  assign n1159 = ~n1157 & n1158;
  assign n1160 = x65 & ~n1140;
  assign n1161 = n1159 & ~n1160;
  assign n1162 = n289 & ~n1029;
  assign n1163 = n1162 ^ x65;
  assign n1164 = n1157 & n1163;
  assign n1165 = x65 & ~n1034;
  assign n1166 = ~n1158 & n1165;
  assign n1167 = ~n1140 & n1166;
  assign n1168 = ~n1164 & ~n1167;
  assign n1169 = ~n1161 & n1168;
  assign n1170 = n1169 ^ x50;
  assign n1171 = n1170 ^ n1155;
  assign n1172 = ~n1156 & n1171;
  assign n1173 = n1172 ^ x66;
  assign n1174 = n1173 ^ x67;
  assign n1175 = ~n1047 & ~n1140;
  assign n1176 = n1175 ^ n1067;
  assign n1177 = n1176 ^ n1173;
  assign n1178 = n1174 & ~n1177;
  assign n1179 = n1178 ^ x67;
  assign n1180 = n1179 ^ x68;
  assign n1181 = n1071 & ~n1140;
  assign n1182 = n1181 ^ n1073;
  assign n1183 = n1182 ^ n1179;
  assign n1184 = n1180 & n1183;
  assign n1185 = n1184 ^ x68;
  assign n1186 = n1185 ^ x69;
  assign n1187 = n1077 & ~n1140;
  assign n1188 = n1187 ^ n1079;
  assign n1189 = n1188 ^ n1185;
  assign n1190 = n1186 & n1189;
  assign n1191 = n1190 ^ x69;
  assign n1192 = n1191 ^ x70;
  assign n1193 = n1083 & ~n1140;
  assign n1194 = n1193 ^ n1085;
  assign n1195 = n1194 ^ n1191;
  assign n1196 = n1192 & n1195;
  assign n1197 = n1196 ^ x70;
  assign n1198 = n1197 ^ x71;
  assign n1199 = n1089 & ~n1140;
  assign n1200 = n1199 ^ n1091;
  assign n1201 = n1200 ^ n1197;
  assign n1202 = n1198 & ~n1201;
  assign n1203 = n1202 ^ x71;
  assign n1204 = n1203 ^ x72;
  assign n1205 = n1095 & ~n1140;
  assign n1206 = n1205 ^ n1097;
  assign n1207 = n1206 ^ n1203;
  assign n1208 = n1204 & ~n1207;
  assign n1209 = n1208 ^ x72;
  assign n1210 = n1209 ^ x73;
  assign n1211 = n1101 & ~n1140;
  assign n1212 = n1211 ^ n1103;
  assign n1213 = n1212 ^ n1209;
  assign n1214 = n1210 & ~n1213;
  assign n1215 = n1214 ^ x73;
  assign n1216 = n1215 ^ x74;
  assign n1217 = n1107 & ~n1140;
  assign n1218 = n1217 ^ n1109;
  assign n1219 = n1218 ^ n1215;
  assign n1220 = n1216 & ~n1219;
  assign n1221 = n1220 ^ x74;
  assign n1222 = n1221 ^ x75;
  assign n1223 = n1113 & ~n1140;
  assign n1224 = n1223 ^ n1115;
  assign n1225 = n1224 ^ n1221;
  assign n1226 = n1222 & ~n1225;
  assign n1227 = n1226 ^ x75;
  assign n1228 = n1227 ^ x76;
  assign n1229 = n1119 & ~n1140;
  assign n1230 = n1229 ^ n1121;
  assign n1231 = n1230 ^ n1227;
  assign n1232 = n1228 & n1231;
  assign n1233 = n1232 ^ x76;
  assign n1234 = n1233 ^ x77;
  assign n1235 = n1125 & ~n1140;
  assign n1236 = n1235 ^ n1127;
  assign n1237 = n1236 ^ n1233;
  assign n1238 = n1234 & ~n1237;
  assign n1239 = n1238 ^ x77;
  assign n1240 = n1146 & n1239;
  assign n1241 = x78 & ~n1145;
  assign n1242 = ~n1142 & n1241;
  assign n1243 = ~x80 & n175;
  assign n1244 = ~n1144 & n1243;
  assign n1245 = ~n177 & ~n1244;
  assign n1246 = ~n1242 & ~n1245;
  assign n1247 = ~n1240 & n1246;
  assign n1248 = n1138 & ~n1247;
  assign n1249 = ~n240 & ~n1248;
  assign n1250 = n1249 ^ x80;
  assign n1251 = n1239 ^ x78;
  assign n1252 = n1247 & n1251;
  assign n1253 = n1252 ^ n1142;
  assign n1254 = n1253 ^ n1249;
  assign n1255 = n1254 ^ n1249;
  assign n1256 = n1249 ^ x79;
  assign n1257 = n1256 ^ n1249;
  assign n1258 = ~n1255 & n1257;
  assign n1259 = n1258 ^ n1249;
  assign n1260 = n1250 & ~n1259;
  assign n1261 = n1260 ^ x80;
  assign n1263 = ~x80 & ~n1249;
  assign n1264 = ~n1253 & ~n1263;
  assign n1265 = x79 & x80;
  assign n1266 = ~n1264 & ~n1265;
  assign n1262 = x79 & n1249;
  assign n1267 = n1266 ^ n1262;
  assign n1268 = ~n1156 & n1247;
  assign n1269 = n1268 ^ n1170;
  assign n1270 = n1269 ^ x67;
  assign n1271 = ~x47 & n1147;
  assign n1272 = ~n1247 & n1271;
  assign n1273 = ~x47 & x65;
  assign n1274 = x64 & n1273;
  assign n1275 = ~n1272 & ~n1274;
  assign n1276 = x64 & n1247;
  assign n1277 = n1276 ^ x47;
  assign n1278 = n1276 ^ x48;
  assign n1279 = n1278 ^ n1276;
  assign n1280 = n1276 & ~n1279;
  assign n1281 = n1280 ^ n1276;
  assign n1282 = ~n1277 & n1281;
  assign n1283 = n1282 ^ n1280;
  assign n1284 = n1283 ^ n1276;
  assign n1285 = n1284 ^ n1278;
  assign n1286 = ~x65 & ~n1285;
  assign n1287 = n1286 ^ n1278;
  assign n1288 = n1275 & n1287;
  assign n1289 = ~x66 & n1288;
  assign n1290 = n1140 ^ x65;
  assign n1291 = n1147 & n1290;
  assign n1292 = ~n202 & ~n1291;
  assign n1293 = x48 & ~n1160;
  assign n1294 = x65 & n1293;
  assign n1295 = n1292 & ~n1294;
  assign n1296 = n1295 ^ n1148;
  assign n1297 = n1295 ^ n1293;
  assign n1298 = n1295 ^ n1247;
  assign n1299 = n1295 & n1298;
  assign n1300 = n1299 ^ n1295;
  assign n1301 = n1297 & n1300;
  assign n1302 = n1301 ^ n1299;
  assign n1303 = n1302 ^ n1295;
  assign n1304 = n1303 ^ n1247;
  assign n1305 = ~n1296 & n1304;
  assign n1306 = n1305 ^ n1148;
  assign n1307 = n1306 ^ x49;
  assign n1308 = ~n1289 & ~n1307;
  assign n1309 = n1308 ^ n1269;
  assign n1310 = n1309 ^ n1269;
  assign n1311 = x66 & ~n1288;
  assign n1312 = n1311 ^ n1269;
  assign n1313 = n1312 ^ n1269;
  assign n1314 = ~n1310 & ~n1313;
  assign n1315 = n1314 ^ n1269;
  assign n1316 = n1270 & n1315;
  assign n1317 = n1316 ^ x67;
  assign n1318 = n1317 ^ x68;
  assign n1319 = n1174 & n1247;
  assign n1320 = n1319 ^ n1176;
  assign n1321 = n1320 ^ n1317;
  assign n1322 = n1318 & ~n1321;
  assign n1323 = n1322 ^ x68;
  assign n1324 = n1323 ^ x69;
  assign n1325 = n1180 & n1247;
  assign n1326 = n1325 ^ n1182;
  assign n1327 = n1326 ^ n1323;
  assign n1328 = n1324 & n1327;
  assign n1329 = n1328 ^ x69;
  assign n1330 = n1329 ^ x70;
  assign n1331 = n1186 & n1247;
  assign n1332 = n1331 ^ n1188;
  assign n1333 = n1332 ^ n1329;
  assign n1334 = n1330 & n1333;
  assign n1335 = n1334 ^ x70;
  assign n1336 = n1335 ^ x71;
  assign n1337 = n1192 & n1247;
  assign n1338 = n1337 ^ n1194;
  assign n1339 = n1338 ^ n1335;
  assign n1340 = n1336 & n1339;
  assign n1341 = n1340 ^ x71;
  assign n1342 = n1341 ^ x72;
  assign n1343 = n1198 & n1247;
  assign n1344 = n1343 ^ n1200;
  assign n1345 = n1344 ^ n1341;
  assign n1346 = n1342 & ~n1345;
  assign n1347 = n1346 ^ x72;
  assign n1348 = n1347 ^ x73;
  assign n1349 = n1204 & n1247;
  assign n1350 = n1349 ^ n1206;
  assign n1351 = n1350 ^ n1347;
  assign n1352 = n1348 & ~n1351;
  assign n1353 = n1352 ^ x73;
  assign n1354 = n1353 ^ x74;
  assign n1355 = n1210 & n1247;
  assign n1356 = n1355 ^ n1212;
  assign n1357 = n1356 ^ n1353;
  assign n1358 = n1354 & ~n1357;
  assign n1359 = n1358 ^ x74;
  assign n1360 = n1359 ^ x75;
  assign n1361 = n1216 & n1247;
  assign n1362 = n1361 ^ n1218;
  assign n1363 = n1362 ^ n1359;
  assign n1364 = n1360 & ~n1363;
  assign n1365 = n1364 ^ x75;
  assign n1366 = n1365 ^ x76;
  assign n1367 = n1222 & n1247;
  assign n1368 = n1367 ^ n1224;
  assign n1369 = n1368 ^ n1365;
  assign n1370 = n1366 & ~n1369;
  assign n1371 = n1370 ^ x76;
  assign n1372 = n1371 ^ x77;
  assign n1373 = n1228 & n1247;
  assign n1374 = n1373 ^ n1230;
  assign n1375 = n1374 ^ n1371;
  assign n1376 = n1372 & n1375;
  assign n1377 = n1376 ^ x77;
  assign n1378 = n1377 ^ x78;
  assign n1379 = n1234 & n1247;
  assign n1380 = n1379 ^ n1236;
  assign n1381 = n1380 ^ n1377;
  assign n1382 = n1378 & ~n1381;
  assign n1383 = n1382 ^ x78;
  assign n1384 = n1383 ^ n1262;
  assign n1385 = ~n1262 & ~n1384;
  assign n1386 = n1385 ^ n1262;
  assign n1387 = ~n1267 & ~n1386;
  assign n1388 = n1387 ^ n1385;
  assign n1389 = n1388 ^ n1262;
  assign n1390 = n1389 ^ n1383;
  assign n1391 = ~n1261 & ~n1390;
  assign n1392 = n1391 ^ n1261;
  assign n1393 = n175 & ~n1392;
  assign n1394 = ~n240 & n1393;
  assign n1395 = ~n1249 & ~n1394;
  assign n1396 = n1395 ^ x81;
  assign n1397 = n174 & ~n1396;
  assign n1398 = ~x46 & ~x47;
  assign n1399 = ~n1393 & n1398;
  assign n1400 = ~x46 & x65;
  assign n1401 = ~n1399 & ~n1400;
  assign n1402 = x64 & ~n1401;
  assign n1403 = x64 & n1393;
  assign n1404 = x46 & ~x65;
  assign n1405 = x47 & ~n1404;
  assign n1406 = n1405 ^ n1273;
  assign n1407 = n1403 & n1406;
  assign n1408 = n1407 ^ n1273;
  assign n1409 = ~n1402 & ~n1408;
  assign n1410 = n1409 ^ x66;
  assign n1411 = x65 & n175;
  assign n1412 = n1411 ^ n288;
  assign n1413 = n1412 ^ n288;
  assign n1414 = n1392 ^ n288;
  assign n1415 = n1414 ^ n288;
  assign n1416 = n1413 & ~n1415;
  assign n1417 = n1416 ^ n288;
  assign n1418 = ~n1247 & n1417;
  assign n1419 = n1418 ^ n288;
  assign n1420 = x47 & n1419;
  assign n1421 = ~n288 & ~n1247;
  assign n1422 = ~x47 & ~n1421;
  assign n1423 = ~n202 & ~n1422;
  assign n1424 = ~x65 & n1247;
  assign n1425 = ~n1423 & ~n1424;
  assign n1426 = n1425 ^ n1276;
  assign n1427 = n1393 & n1426;
  assign n1428 = n1427 ^ n1276;
  assign n1429 = ~n1420 & ~n1428;
  assign n1430 = n1429 ^ x48;
  assign n1431 = n1430 ^ n1409;
  assign n1432 = ~n1410 & n1431;
  assign n1433 = n1432 ^ x66;
  assign n1434 = n1433 ^ x67;
  assign n1435 = n1288 ^ x66;
  assign n1436 = n1393 & ~n1435;
  assign n1437 = n1436 ^ n1307;
  assign n1438 = n1437 ^ n1433;
  assign n1439 = n1434 & n1438;
  assign n1440 = n1439 ^ x67;
  assign n1441 = n1440 ^ x68;
  assign n1442 = ~n1308 & ~n1311;
  assign n1443 = n1442 ^ x67;
  assign n1444 = n1393 & ~n1443;
  assign n1445 = n1444 ^ n1269;
  assign n1446 = n1445 ^ n1440;
  assign n1447 = n1441 & ~n1446;
  assign n1448 = n1447 ^ x68;
  assign n1449 = n1448 ^ x69;
  assign n1450 = n1318 & n1393;
  assign n1451 = n1450 ^ n1320;
  assign n1452 = n1451 ^ n1448;
  assign n1453 = n1449 & ~n1452;
  assign n1454 = n1453 ^ x69;
  assign n1455 = n1454 ^ x70;
  assign n1456 = n1324 & n1393;
  assign n1457 = n1456 ^ n1326;
  assign n1458 = n1457 ^ n1454;
  assign n1459 = n1455 & n1458;
  assign n1460 = n1459 ^ x70;
  assign n1461 = n1460 ^ x71;
  assign n1462 = n1330 & n1393;
  assign n1463 = n1462 ^ n1332;
  assign n1464 = n1463 ^ n1460;
  assign n1465 = n1461 & n1464;
  assign n1466 = n1465 ^ x71;
  assign n1467 = n1466 ^ x72;
  assign n1468 = n1336 & n1393;
  assign n1469 = n1468 ^ n1338;
  assign n1470 = n1469 ^ n1466;
  assign n1471 = n1467 & n1470;
  assign n1472 = n1471 ^ x72;
  assign n1473 = n1472 ^ x73;
  assign n1474 = n1342 & n1393;
  assign n1475 = n1474 ^ n1344;
  assign n1476 = n1475 ^ n1472;
  assign n1477 = n1473 & ~n1476;
  assign n1478 = n1477 ^ x73;
  assign n1479 = n1478 ^ x74;
  assign n1480 = n1348 & n1393;
  assign n1481 = n1480 ^ n1350;
  assign n1482 = n1481 ^ n1478;
  assign n1483 = n1479 & ~n1482;
  assign n1484 = n1483 ^ x74;
  assign n1485 = n1484 ^ x75;
  assign n1486 = n1354 & n1393;
  assign n1487 = n1486 ^ n1356;
  assign n1488 = n1487 ^ n1484;
  assign n1489 = n1485 & ~n1488;
  assign n1490 = n1489 ^ x75;
  assign n1491 = n1490 ^ x76;
  assign n1492 = n1360 & n1393;
  assign n1493 = n1492 ^ n1362;
  assign n1494 = n1493 ^ n1490;
  assign n1495 = n1491 & ~n1494;
  assign n1496 = n1495 ^ x76;
  assign n1497 = n1496 ^ x77;
  assign n1498 = n1366 & n1393;
  assign n1499 = n1498 ^ n1368;
  assign n1500 = n1499 ^ n1496;
  assign n1501 = n1497 & ~n1500;
  assign n1502 = n1501 ^ x77;
  assign n1503 = n1502 ^ x78;
  assign n1504 = n1372 & n1393;
  assign n1505 = n1504 ^ n1374;
  assign n1506 = n1505 ^ n1502;
  assign n1507 = n1503 & n1506;
  assign n1508 = n1507 ^ x78;
  assign n1509 = n1508 ^ x79;
  assign n1510 = n1378 & n1393;
  assign n1511 = n1510 ^ n1380;
  assign n1512 = n1511 ^ n1508;
  assign n1513 = n1509 & ~n1512;
  assign n1514 = n1513 ^ x79;
  assign n1515 = n1514 ^ x80;
  assign n1516 = n1383 ^ x79;
  assign n1517 = n1393 & n1516;
  assign n1518 = n1517 ^ n1253;
  assign n1519 = n1518 ^ n1514;
  assign n1520 = n1515 & n1519;
  assign n1521 = n1520 ^ x80;
  assign n1522 = n1397 & ~n1521;
  assign n1523 = ~n175 & n1248;
  assign n1524 = ~n1522 & n1523;
  assign n1525 = ~n240 & ~n1524;
  assign n1526 = x82 & n1525;
  assign n1527 = ~x82 & ~n1525;
  assign n1528 = n175 & n1395;
  assign n1529 = ~n1522 & ~n1528;
  assign n1530 = n1434 & ~n1529;
  assign n1531 = n1530 ^ n1437;
  assign n1532 = ~x68 & n1531;
  assign n1533 = n1441 & ~n1529;
  assign n1534 = n1533 ^ n1445;
  assign n1535 = ~x69 & ~n1534;
  assign n1536 = ~n1532 & ~n1535;
  assign n1537 = ~x45 & x64;
  assign n1538 = n1537 ^ x65;
  assign n1539 = n1529 ^ x46;
  assign n1540 = n1539 ^ n1537;
  assign n1543 = n1540 ^ n1529;
  assign n1544 = n1543 ^ n1540;
  assign n1541 = n1540 ^ x64;
  assign n1542 = n1541 ^ n1540;
  assign n1545 = n1544 ^ n1542;
  assign n1546 = n1540 ^ n1537;
  assign n1547 = n1546 ^ n1540;
  assign n1548 = n1547 ^ n1544;
  assign n1549 = ~n1544 & n1548;
  assign n1550 = n1549 ^ n1544;
  assign n1551 = n1545 & ~n1550;
  assign n1552 = n1551 ^ n1549;
  assign n1553 = n1552 ^ n1540;
  assign n1554 = n1553 ^ n1544;
  assign n1555 = n1538 & n1554;
  assign n1556 = n1555 ^ x65;
  assign n1557 = n1556 ^ x66;
  assign n1558 = n1400 ^ n1393;
  assign n1559 = n1558 ^ n1400;
  assign n1560 = ~x46 & ~x64;
  assign n1561 = x65 ^ x46;
  assign n1562 = ~n1560 & ~n1561;
  assign n1563 = n1562 ^ n1400;
  assign n1564 = ~n1559 & n1563;
  assign n1565 = n1564 ^ n1400;
  assign n1566 = ~n202 & ~n1565;
  assign n1567 = n1566 ^ n1403;
  assign n1568 = n1566 ^ n1404;
  assign n1569 = n1566 ^ n1529;
  assign n1570 = n1566 & ~n1569;
  assign n1571 = n1570 ^ n1566;
  assign n1572 = n1568 & n1571;
  assign n1573 = n1572 ^ n1570;
  assign n1574 = n1573 ^ n1566;
  assign n1575 = n1574 ^ n1529;
  assign n1576 = ~n1567 & ~n1575;
  assign n1577 = n1576 ^ n1403;
  assign n1578 = n1577 ^ x47;
  assign n1579 = n1578 ^ n1556;
  assign n1580 = n1557 & n1579;
  assign n1581 = n1580 ^ x66;
  assign n1582 = n1581 ^ x67;
  assign n1583 = ~n1410 & ~n1529;
  assign n1584 = n1583 ^ n1430;
  assign n1585 = n1584 ^ n1581;
  assign n1586 = n1582 & ~n1585;
  assign n1587 = n1586 ^ x67;
  assign n1588 = n1536 & n1587;
  assign n1589 = n1534 ^ x69;
  assign n1590 = x68 & ~n1531;
  assign n1591 = n1590 ^ n1534;
  assign n1592 = n1589 & ~n1591;
  assign n1593 = n1592 ^ x69;
  assign n1594 = ~n1588 & ~n1593;
  assign n1595 = n1594 ^ x70;
  assign n1596 = n1449 & ~n1529;
  assign n1597 = n1596 ^ n1451;
  assign n1598 = n1597 ^ n1594;
  assign n1599 = ~n1595 & n1598;
  assign n1600 = n1599 ^ x70;
  assign n1601 = n1600 ^ x71;
  assign n1602 = n1455 & ~n1529;
  assign n1603 = n1602 ^ n1457;
  assign n1604 = n1603 ^ n1600;
  assign n1605 = n1601 & n1604;
  assign n1606 = n1605 ^ x71;
  assign n1607 = n1606 ^ x72;
  assign n1608 = n1461 & ~n1529;
  assign n1609 = n1608 ^ n1463;
  assign n1610 = n1609 ^ n1606;
  assign n1611 = n1607 & n1610;
  assign n1612 = n1611 ^ x72;
  assign n1613 = n1612 ^ x73;
  assign n1614 = n1467 & ~n1529;
  assign n1615 = n1614 ^ n1469;
  assign n1616 = n1615 ^ n1612;
  assign n1617 = n1613 & n1616;
  assign n1618 = n1617 ^ x73;
  assign n1619 = n1618 ^ x74;
  assign n1620 = n1473 & ~n1529;
  assign n1621 = n1620 ^ n1475;
  assign n1622 = n1621 ^ n1618;
  assign n1623 = n1619 & ~n1622;
  assign n1624 = n1623 ^ x74;
  assign n1625 = n1624 ^ x75;
  assign n1626 = n1479 & ~n1529;
  assign n1627 = n1626 ^ n1481;
  assign n1628 = n1627 ^ n1624;
  assign n1629 = n1625 & ~n1628;
  assign n1630 = n1629 ^ x75;
  assign n1631 = n1630 ^ x76;
  assign n1632 = n1485 & ~n1529;
  assign n1633 = n1632 ^ n1487;
  assign n1634 = n1633 ^ n1630;
  assign n1635 = n1631 & ~n1634;
  assign n1636 = n1635 ^ x76;
  assign n1637 = n1636 ^ x77;
  assign n1638 = n1491 & ~n1529;
  assign n1639 = n1638 ^ n1493;
  assign n1640 = n1639 ^ n1636;
  assign n1641 = n1637 & ~n1640;
  assign n1642 = n1641 ^ x77;
  assign n1643 = n1642 ^ x78;
  assign n1644 = n1497 & ~n1529;
  assign n1645 = n1644 ^ n1499;
  assign n1646 = n1645 ^ n1642;
  assign n1647 = n1643 & ~n1646;
  assign n1648 = n1647 ^ x78;
  assign n1649 = n1648 ^ x79;
  assign n1650 = n1503 & ~n1529;
  assign n1651 = n1650 ^ n1505;
  assign n1652 = n1651 ^ n1648;
  assign n1653 = n1649 & n1652;
  assign n1654 = n1653 ^ x79;
  assign n1655 = n1654 ^ x80;
  assign n1656 = n1509 & ~n1529;
  assign n1657 = n1656 ^ n1511;
  assign n1658 = n1657 ^ n1654;
  assign n1659 = n1655 & ~n1658;
  assign n1660 = n1659 ^ x80;
  assign n1661 = n1660 ^ x81;
  assign n1662 = n1515 & ~n1529;
  assign n1663 = n1662 ^ n1518;
  assign n1664 = n1663 ^ n1660;
  assign n1665 = n1661 & ~n1664;
  assign n1666 = n1665 ^ n1660;
  assign n1667 = ~n1527 & n1666;
  assign n1668 = ~n1526 & ~n1667;
  assign n1669 = n173 & n1668;
  assign n1821 = n1669 ^ x65;
  assign n1822 = n1669 ^ x64;
  assign n1823 = n1822 ^ x64;
  assign n1670 = n1524 & ~n1669;
  assign n1671 = ~n240 & ~n1670;
  assign n1672 = ~x83 & ~n1671;
  assign n1673 = x83 & n1671;
  assign n1674 = x65 & n1529;
  assign n1675 = n173 & n1674;
  assign n1676 = n1668 & n1675;
  assign n1677 = n288 & ~n1529;
  assign n1678 = ~n1676 & ~n1677;
  assign n1679 = x45 & ~n1678;
  assign n1689 = x64 & ~n1529;
  assign n1680 = n202 ^ x65;
  assign n1681 = n1680 ^ n1529;
  assign n1682 = n1537 ^ n1529;
  assign n1683 = n1529 ^ n202;
  assign n1684 = n1683 ^ n1529;
  assign n1685 = ~n1682 & ~n1684;
  assign n1686 = n1685 ^ n1529;
  assign n1687 = n1681 & ~n1686;
  assign n1688 = n1687 ^ n202;
  assign n1690 = n1689 ^ n1688;
  assign n1691 = n1669 & n1690;
  assign n1692 = n1691 ^ n1689;
  assign n1693 = ~n1679 & ~n1692;
  assign n1694 = n1693 ^ x46;
  assign n1695 = n1694 ^ x66;
  assign n1696 = x64 & n1669;
  assign n1697 = x44 & ~x65;
  assign n1698 = x45 & ~n1697;
  assign n1699 = n1696 & n1698;
  assign n1700 = ~x44 & n1537;
  assign n1701 = ~x45 & x65;
  assign n1702 = ~n1700 & ~n1701;
  assign n1703 = ~n1669 & ~n1702;
  assign n1704 = ~x44 & x65;
  assign n1705 = n1704 ^ n1701;
  assign n1706 = x64 & n1705;
  assign n1707 = n1706 ^ n1701;
  assign n1708 = ~n1703 & ~n1707;
  assign n1709 = ~n1699 & n1708;
  assign n1710 = n1709 ^ n1694;
  assign n1711 = n1695 & n1710;
  assign n1712 = n1711 ^ x66;
  assign n1713 = n1712 ^ x67;
  assign n1714 = n1557 & n1669;
  assign n1715 = n1714 ^ n1578;
  assign n1716 = n1715 ^ n1712;
  assign n1717 = n1713 & n1716;
  assign n1718 = n1717 ^ x67;
  assign n1719 = n1718 ^ x68;
  assign n1720 = n1582 & n1669;
  assign n1721 = n1720 ^ n1584;
  assign n1722 = n1721 ^ n1718;
  assign n1723 = n1719 & ~n1722;
  assign n1724 = n1723 ^ x68;
  assign n1725 = n1724 ^ x69;
  assign n1726 = n1587 ^ x68;
  assign n1727 = n1669 & n1726;
  assign n1728 = n1727 ^ n1531;
  assign n1729 = n1728 ^ n1724;
  assign n1730 = n1725 & n1729;
  assign n1731 = n1730 ^ x69;
  assign n1732 = n1731 ^ x70;
  assign n1733 = n1587 ^ n1531;
  assign n1734 = n1726 & n1733;
  assign n1735 = n1734 ^ x68;
  assign n1736 = n1735 ^ x69;
  assign n1737 = n1669 & n1736;
  assign n1738 = n1737 ^ n1534;
  assign n1739 = n1738 ^ n1731;
  assign n1740 = n1732 & ~n1739;
  assign n1741 = n1740 ^ x70;
  assign n1742 = n1741 ^ x71;
  assign n1743 = ~n1595 & n1669;
  assign n1744 = n1743 ^ n1597;
  assign n1745 = n1744 ^ n1741;
  assign n1746 = n1742 & ~n1745;
  assign n1747 = n1746 ^ x71;
  assign n1748 = n1747 ^ x72;
  assign n1749 = n1601 & n1669;
  assign n1750 = n1749 ^ n1603;
  assign n1751 = n1750 ^ n1747;
  assign n1752 = n1748 & n1751;
  assign n1753 = n1752 ^ x72;
  assign n1754 = n1753 ^ x73;
  assign n1755 = n1607 & n1669;
  assign n1756 = n1755 ^ n1609;
  assign n1757 = n1756 ^ n1753;
  assign n1758 = n1754 & n1757;
  assign n1759 = n1758 ^ x73;
  assign n1760 = n1759 ^ x74;
  assign n1761 = n1613 & n1669;
  assign n1762 = n1761 ^ n1615;
  assign n1763 = n1762 ^ n1759;
  assign n1764 = n1760 & n1763;
  assign n1765 = n1764 ^ x74;
  assign n1766 = n1765 ^ x75;
  assign n1767 = n1619 & n1669;
  assign n1768 = n1767 ^ n1621;
  assign n1769 = n1768 ^ n1765;
  assign n1770 = n1766 & ~n1769;
  assign n1771 = n1770 ^ x75;
  assign n1772 = n1771 ^ x76;
  assign n1773 = n1625 & n1669;
  assign n1774 = n1773 ^ n1627;
  assign n1775 = n1774 ^ n1771;
  assign n1776 = n1772 & ~n1775;
  assign n1777 = n1776 ^ x76;
  assign n1778 = n1777 ^ x77;
  assign n1779 = n1631 & n1669;
  assign n1780 = n1779 ^ n1633;
  assign n1781 = n1780 ^ n1777;
  assign n1782 = n1778 & ~n1781;
  assign n1783 = n1782 ^ x77;
  assign n1784 = n1783 ^ x78;
  assign n1785 = n1637 & n1669;
  assign n1786 = n1785 ^ n1639;
  assign n1787 = n1786 ^ n1783;
  assign n1788 = n1784 & ~n1787;
  assign n1789 = n1788 ^ x78;
  assign n1790 = n1789 ^ x79;
  assign n1791 = n1643 & n1669;
  assign n1792 = n1791 ^ n1645;
  assign n1793 = n1792 ^ n1789;
  assign n1794 = n1790 & ~n1793;
  assign n1795 = n1794 ^ x79;
  assign n1796 = n1795 ^ x80;
  assign n1797 = n1649 & n1669;
  assign n1798 = n1797 ^ n1651;
  assign n1799 = n1798 ^ n1795;
  assign n1800 = n1796 & n1799;
  assign n1801 = n1800 ^ x80;
  assign n1802 = n1801 ^ x81;
  assign n1803 = n1655 & n1669;
  assign n1804 = n1803 ^ n1657;
  assign n1805 = n1804 ^ n1801;
  assign n1806 = n1802 & ~n1805;
  assign n1807 = n1806 ^ x81;
  assign n1808 = n1807 ^ x82;
  assign n1809 = n1661 & n1669;
  assign n1810 = n1809 ^ n1663;
  assign n1811 = n1810 ^ n1807;
  assign n1812 = n1808 & ~n1811;
  assign n1813 = n1812 ^ n1807;
  assign n1814 = ~n1673 & ~n1813;
  assign n1815 = ~n1672 & ~n1814;
  assign n1816 = n172 & ~n1815;
  assign n1824 = n1816 ^ x64;
  assign n1825 = ~n1823 & n1824;
  assign n1826 = n1825 ^ x64;
  assign n1827 = n1821 & n1826;
  assign n1828 = x44 & n1827;
  assign n1829 = ~x65 & n1669;
  assign n1830 = ~x44 & ~n1829;
  assign n1831 = ~n288 & ~n1669;
  assign n1832 = n1830 & ~n1831;
  assign n1833 = ~n202 & ~n1832;
  assign n1834 = n1833 ^ n1696;
  assign n1835 = n1816 & ~n1834;
  assign n1836 = n1835 ^ n1696;
  assign n1837 = ~n1828 & ~n1836;
  assign n1838 = n1837 ^ x45;
  assign n1839 = ~x43 & ~x44;
  assign n1840 = ~n1816 & n1839;
  assign n1841 = ~x43 & x65;
  assign n1842 = ~n1840 & ~n1841;
  assign n1843 = x64 & ~n1842;
  assign n1844 = x64 & n1816;
  assign n1845 = x43 & n1697;
  assign n1846 = n1845 ^ x44;
  assign n1847 = n1846 ^ n1704;
  assign n1848 = n1844 & n1847;
  assign n1849 = n1848 ^ n1704;
  assign n1850 = ~n1843 & ~n1849;
  assign n1851 = ~x66 & n1850;
  assign n1852 = n1838 & ~n1851;
  assign n1853 = n1709 ^ x66;
  assign n1854 = n1816 & ~n1853;
  assign n1855 = n1854 ^ n1694;
  assign n1856 = n1852 & n1855;
  assign n1857 = x67 & ~n1850;
  assign n1858 = n1838 & n1857;
  assign n1859 = x66 & ~n1850;
  assign n1860 = ~x67 & ~n1855;
  assign n1861 = n1859 & ~n1860;
  assign n1862 = ~n1858 & ~n1861;
  assign n1863 = ~n1856 & n1862;
  assign n1864 = x66 & x67;
  assign n1865 = n1838 & n1864;
  assign n1866 = x67 & n1855;
  assign n1867 = ~n1865 & ~n1866;
  assign n1868 = n1863 & n1867;
  assign n1869 = n1868 ^ x68;
  assign n1870 = n1713 & n1816;
  assign n1871 = n1870 ^ n1715;
  assign n1872 = n1871 ^ n1868;
  assign n1873 = ~n1869 & ~n1872;
  assign n1874 = n1873 ^ x68;
  assign n1875 = n1874 ^ x69;
  assign n1876 = n1719 & n1816;
  assign n1877 = n1876 ^ n1721;
  assign n1878 = n1877 ^ n1874;
  assign n1879 = n1875 & ~n1878;
  assign n1880 = n1879 ^ x69;
  assign n1881 = n1880 ^ x70;
  assign n1882 = n1725 & n1816;
  assign n1883 = n1882 ^ n1728;
  assign n1884 = n1883 ^ n1880;
  assign n1885 = n1881 & n1884;
  assign n1886 = n1885 ^ x70;
  assign n1887 = n1886 ^ x71;
  assign n1888 = n1732 & n1816;
  assign n1889 = n1888 ^ n1738;
  assign n1890 = n1889 ^ n1886;
  assign n1891 = n1887 & ~n1890;
  assign n1892 = n1891 ^ x71;
  assign n1893 = n1892 ^ x72;
  assign n1894 = n1742 & n1816;
  assign n1895 = n1894 ^ n1744;
  assign n1896 = n1895 ^ n1892;
  assign n1897 = n1893 & ~n1896;
  assign n1898 = n1897 ^ x72;
  assign n1899 = n1898 ^ x73;
  assign n1900 = n1748 & n1816;
  assign n1901 = n1900 ^ n1750;
  assign n1902 = n1901 ^ n1898;
  assign n1903 = n1899 & n1902;
  assign n1904 = n1903 ^ x73;
  assign n1905 = n1904 ^ x74;
  assign n1906 = n1754 & n1816;
  assign n1907 = n1906 ^ n1756;
  assign n1908 = n1907 ^ n1904;
  assign n1909 = n1905 & n1908;
  assign n1910 = n1909 ^ x74;
  assign n1911 = n1910 ^ x75;
  assign n1819 = ~x87 & n168;
  assign n1820 = n169 & n1819;
  assign n1912 = n1760 & n1816;
  assign n1913 = n1912 ^ n1762;
  assign n1914 = n1913 ^ n1910;
  assign n1915 = n1911 & n1914;
  assign n1916 = n1915 ^ x75;
  assign n1917 = n1916 ^ x76;
  assign n1918 = n1766 & n1816;
  assign n1919 = n1918 ^ n1768;
  assign n1920 = n1919 ^ n1916;
  assign n1921 = n1917 & ~n1920;
  assign n1922 = n1921 ^ x76;
  assign n1923 = n1922 ^ x77;
  assign n1924 = n1772 & n1816;
  assign n1925 = n1924 ^ n1774;
  assign n1926 = n1925 ^ n1922;
  assign n1927 = n1923 & ~n1926;
  assign n1928 = n1927 ^ x77;
  assign n1929 = n1928 ^ x78;
  assign n1930 = n1778 & n1816;
  assign n1931 = n1930 ^ n1780;
  assign n1932 = n1931 ^ n1928;
  assign n1933 = n1929 & ~n1932;
  assign n1934 = n1933 ^ x78;
  assign n1935 = n1934 ^ x79;
  assign n1936 = n1784 & n1816;
  assign n1937 = n1936 ^ n1786;
  assign n1938 = n1937 ^ n1934;
  assign n1939 = n1935 & ~n1938;
  assign n1940 = n1939 ^ x79;
  assign n1941 = n1940 ^ x80;
  assign n1942 = n1790 & n1816;
  assign n1943 = n1942 ^ n1792;
  assign n1944 = n1943 ^ n1940;
  assign n1945 = n1941 & ~n1944;
  assign n1946 = n1945 ^ x80;
  assign n1947 = n1946 ^ x81;
  assign n1948 = n1796 & n1816;
  assign n1949 = n1948 ^ n1798;
  assign n1950 = n1949 ^ n1946;
  assign n1951 = n1947 & n1950;
  assign n1952 = n1951 ^ x81;
  assign n1953 = n1952 ^ x82;
  assign n1954 = n1802 & n1816;
  assign n1955 = n1954 ^ n1804;
  assign n1956 = n1955 ^ n1952;
  assign n1957 = n1953 & ~n1956;
  assign n1958 = n1957 ^ x82;
  assign n1959 = n1958 ^ x83;
  assign n1960 = n1808 & n1816;
  assign n1961 = n1960 ^ n1810;
  assign n1962 = n1961 ^ n1958;
  assign n1963 = n1959 & n1962;
  assign n1964 = n1963 ^ x83;
  assign n1969 = n1964 ^ x84;
  assign n1817 = ~n240 & n1816;
  assign n1818 = ~n1671 & ~n1817;
  assign n1970 = n1964 ^ n1818;
  assign n1971 = n1969 & n1970;
  assign n1972 = n1971 ^ x84;
  assign n1973 = n1820 & ~n1972;
  assign n1974 = n1911 & n1973;
  assign n1975 = n1974 ^ n1913;
  assign n1976 = n1975 ^ x76;
  assign n1977 = n1905 & n1973;
  assign n1978 = n1977 ^ n1907;
  assign n1979 = ~x75 & n1978;
  assign n1980 = x65 & n1820;
  assign n1981 = n1980 ^ n288;
  assign n1982 = n1981 ^ n288;
  assign n1983 = n1972 ^ n288;
  assign n1984 = n1983 ^ n288;
  assign n1985 = n1982 & ~n1984;
  assign n1986 = n1985 ^ n288;
  assign n1987 = ~n1816 & n1986;
  assign n1988 = n1987 ^ n288;
  assign n1989 = x43 & n1988;
  assign n1990 = n1841 ^ n1816;
  assign n1991 = n1990 ^ n1841;
  assign n1992 = ~x43 & n288;
  assign n1993 = n1992 ^ n1841;
  assign n1994 = ~n1991 & n1993;
  assign n1995 = n1994 ^ n1841;
  assign n1996 = ~n202 & ~n1995;
  assign n1997 = n1996 ^ n1844;
  assign n1998 = n1973 & ~n1997;
  assign n1999 = n1998 ^ n1844;
  assign n2000 = ~n1989 & ~n1999;
  assign n2001 = n2000 ^ x44;
  assign n2002 = n2001 ^ x66;
  assign n2003 = x64 & n1973;
  assign n2004 = x42 & ~x65;
  assign n2005 = x43 & ~n2004;
  assign n2006 = n2003 & n2005;
  assign n2008 = x65 ^ x43;
  assign n2015 = n2008 ^ x65;
  assign n2007 = x65 ^ x42;
  assign n2009 = n2008 ^ n2007;
  assign n2010 = n2009 ^ x65;
  assign n2011 = n2007 ^ x64;
  assign n2012 = n2011 ^ n2007;
  assign n2013 = n2012 ^ n2010;
  assign n2014 = ~n2010 & ~n2013;
  assign n2016 = n2015 ^ n2014;
  assign n2017 = n2016 ^ n2010;
  assign n2018 = n1973 ^ x65;
  assign n2019 = n2018 ^ x65;
  assign n2020 = n2014 ^ n2010;
  assign n2021 = ~n2019 & ~n2020;
  assign n2022 = n2021 ^ x65;
  assign n2023 = ~n2017 & n2022;
  assign n2024 = n2023 ^ x65;
  assign n2025 = n2024 ^ x65;
  assign n2026 = n2025 ^ x65;
  assign n2027 = ~n2006 & ~n2026;
  assign n2028 = n2027 ^ n2001;
  assign n2029 = n2002 & n2028;
  assign n2030 = n2029 ^ x66;
  assign n2031 = n2030 ^ x67;
  assign n2032 = n1850 ^ x66;
  assign n2033 = n1973 & ~n2032;
  assign n2034 = n2033 ^ n1838;
  assign n2035 = n2034 ^ n2030;
  assign n2036 = n2031 & ~n2035;
  assign n2037 = n2036 ^ x67;
  assign n2038 = n2037 ^ x68;
  assign n2039 = ~n1852 & ~n1859;
  assign n2040 = n2039 ^ x67;
  assign n2041 = n1973 & ~n2040;
  assign n2042 = n2041 ^ n1855;
  assign n2043 = n2042 ^ n2037;
  assign n2044 = n2038 & ~n2043;
  assign n2045 = n2044 ^ x68;
  assign n2046 = n2045 ^ x69;
  assign n2047 = ~n1869 & n1973;
  assign n2048 = n2047 ^ n1871;
  assign n2049 = n2048 ^ n2045;
  assign n2050 = n2046 & n2049;
  assign n2051 = n2050 ^ x69;
  assign n2052 = n2051 ^ x70;
  assign n2053 = n1875 & n1973;
  assign n2054 = n2053 ^ n1877;
  assign n2055 = n2054 ^ n2051;
  assign n2056 = n2052 & ~n2055;
  assign n2057 = n2056 ^ x70;
  assign n2058 = n2057 ^ x71;
  assign n2059 = n1881 & n1973;
  assign n2060 = n2059 ^ n1883;
  assign n2061 = n2060 ^ n2057;
  assign n2062 = n2058 & n2061;
  assign n2063 = n2062 ^ x71;
  assign n2064 = n2063 ^ x72;
  assign n2065 = n1887 & n1973;
  assign n2066 = n2065 ^ n1889;
  assign n2067 = n2066 ^ n2063;
  assign n2068 = n2064 & ~n2067;
  assign n2069 = n2068 ^ x72;
  assign n2070 = n2069 ^ x73;
  assign n2071 = n1893 & n1973;
  assign n2072 = n2071 ^ n1895;
  assign n2073 = n2072 ^ n2069;
  assign n2074 = n2070 & ~n2073;
  assign n2075 = n2074 ^ x73;
  assign n2076 = n2075 ^ x74;
  assign n2077 = n1899 & n1973;
  assign n2078 = n2077 ^ n1901;
  assign n2079 = n2078 ^ n2075;
  assign n2080 = n2076 & n2079;
  assign n2081 = n2080 ^ x74;
  assign n2082 = ~n1979 & n2081;
  assign n2083 = n2082 ^ n1975;
  assign n2084 = n2083 ^ n1975;
  assign n2085 = x75 & ~n1978;
  assign n2086 = n2085 ^ n1975;
  assign n2087 = n2086 ^ n1975;
  assign n2088 = ~n2084 & ~n2087;
  assign n2089 = n2088 ^ n1975;
  assign n2090 = ~n1976 & ~n2089;
  assign n2091 = n2090 ^ x76;
  assign n2092 = n2091 ^ x77;
  assign n2093 = n1917 & n1973;
  assign n2094 = n2093 ^ n1919;
  assign n2095 = n2094 ^ n2091;
  assign n2096 = n2092 & ~n2095;
  assign n2097 = n2096 ^ x77;
  assign n2098 = n2097 ^ x78;
  assign n2099 = n1923 & n1973;
  assign n2100 = n2099 ^ n1925;
  assign n2101 = n2100 ^ n2097;
  assign n2102 = n2098 & ~n2101;
  assign n2103 = n2102 ^ x78;
  assign n2104 = n2103 ^ x79;
  assign n2105 = n1929 & n1973;
  assign n2106 = n2105 ^ n1931;
  assign n2107 = n2106 ^ n2103;
  assign n2108 = n2104 & ~n2107;
  assign n2109 = n2108 ^ x79;
  assign n2110 = n2109 ^ x80;
  assign n2111 = n1935 & n1973;
  assign n2112 = n2111 ^ n1937;
  assign n2113 = n2112 ^ n2109;
  assign n2114 = n2110 & ~n2113;
  assign n2115 = n2114 ^ x80;
  assign n2116 = n2115 ^ x81;
  assign n2117 = n1941 & n1973;
  assign n2118 = n2117 ^ n1943;
  assign n2119 = n2118 ^ n2115;
  assign n2120 = n2116 & ~n2119;
  assign n2121 = n2120 ^ x81;
  assign n2122 = n2121 ^ x82;
  assign n2123 = n1947 & n1973;
  assign n2124 = n2123 ^ n1949;
  assign n2125 = n2124 ^ n2121;
  assign n2126 = n2122 & n2125;
  assign n2127 = n2126 ^ x82;
  assign n2128 = n2127 ^ x83;
  assign n2129 = n1953 & n1973;
  assign n2130 = n2129 ^ n1955;
  assign n2131 = n2130 ^ n2127;
  assign n2132 = n2128 & ~n2131;
  assign n2133 = n2132 ^ x83;
  assign n2134 = n2133 ^ x84;
  assign n2135 = n1959 & n1973;
  assign n2136 = n2135 ^ n1961;
  assign n2137 = n2136 ^ n2133;
  assign n2138 = n2134 & n2137;
  assign n2139 = n2138 ^ x84;
  assign n2140 = n2139 ^ x85;
  assign n2141 = n2139 ^ n1818;
  assign n2142 = n2141 ^ n1818;
  assign n1965 = x84 & n1964;
  assign n1966 = n1820 & ~n1965;
  assign n1967 = n1818 & ~n1966;
  assign n2143 = n1967 ^ n1818;
  assign n2144 = n2142 & ~n2143;
  assign n2145 = n2144 ^ n1818;
  assign n2146 = n2140 & n2145;
  assign n2147 = n2146 ^ x85;
  assign n1968 = ~x86 & n1819;
  assign n2160 = x42 & x65;
  assign n2161 = n1968 & n2160;
  assign n2162 = ~n1973 & n2161;
  assign n2163 = ~n2147 & n2162;
  assign n2164 = n2003 & n2004;
  assign n2165 = ~n2163 & ~n2164;
  assign n2148 = n1968 & ~n2147;
  assign n2166 = ~x42 & x64;
  assign n2167 = ~n2018 & n2166;
  assign n2168 = ~n202 & ~n2167;
  assign n2169 = n2168 ^ n2003;
  assign n2170 = n2148 & ~n2169;
  assign n2171 = n2170 ^ n2003;
  assign n2172 = n2165 & ~n2171;
  assign n2173 = n2172 ^ x43;
  assign n2174 = n2173 ^ x66;
  assign n2175 = x64 & n2148;
  assign n2176 = x41 & n2004;
  assign n2177 = n2176 ^ x42;
  assign n2178 = n2175 & n2177;
  assign n2179 = ~x41 & n2166;
  assign n2180 = ~x42 & x65;
  assign n2181 = ~n2179 & ~n2180;
  assign n2182 = ~n2148 & ~n2181;
  assign n2183 = ~x41 & x65;
  assign n2184 = n2183 ^ n2180;
  assign n2185 = x64 & n2184;
  assign n2186 = n2185 ^ n2180;
  assign n2187 = ~n2182 & ~n2186;
  assign n2188 = ~n2178 & n2187;
  assign n2189 = n2188 ^ n2173;
  assign n2190 = n2174 & n2189;
  assign n2191 = n2190 ^ x66;
  assign n2192 = n2191 ^ x67;
  assign n2193 = n2027 ^ x66;
  assign n2194 = n2148 & ~n2193;
  assign n2195 = n2194 ^ n2001;
  assign n2196 = n2195 ^ n2191;
  assign n2197 = n2192 & ~n2196;
  assign n2198 = n2197 ^ x67;
  assign n2199 = n2198 ^ x68;
  assign n2151 = n2128 & n2148;
  assign n2152 = n2151 ^ n2130;
  assign n2153 = x84 & n2152;
  assign n2154 = n2110 & n2148;
  assign n2155 = n2154 ^ n2112;
  assign n2156 = n2155 ^ x81;
  assign n2157 = n2104 & n2148;
  assign n2158 = n2157 ^ n2106;
  assign n2159 = x80 & n2158;
  assign n2200 = n2031 & n2148;
  assign n2201 = n2200 ^ n2034;
  assign n2202 = n2201 ^ n2198;
  assign n2203 = n2199 & ~n2202;
  assign n2204 = n2203 ^ x68;
  assign n2205 = n2204 ^ x69;
  assign n2206 = n2038 & n2148;
  assign n2207 = n2206 ^ n2042;
  assign n2208 = n2207 ^ n2204;
  assign n2209 = n2205 & ~n2208;
  assign n2210 = n2209 ^ x69;
  assign n2211 = n2210 ^ x70;
  assign n2212 = n2046 & n2148;
  assign n2213 = n2212 ^ n2048;
  assign n2214 = n2213 ^ n2210;
  assign n2215 = n2211 & n2214;
  assign n2216 = n2215 ^ x70;
  assign n2217 = n2216 ^ x71;
  assign n2218 = n2052 & n2148;
  assign n2219 = n2218 ^ n2054;
  assign n2220 = n2219 ^ n2216;
  assign n2221 = n2217 & ~n2220;
  assign n2222 = n2221 ^ x71;
  assign n2223 = n2222 ^ x72;
  assign n2224 = n2058 & n2148;
  assign n2225 = n2224 ^ n2060;
  assign n2226 = n2225 ^ n2222;
  assign n2227 = n2223 & n2226;
  assign n2228 = n2227 ^ x72;
  assign n2229 = n2228 ^ x73;
  assign n2230 = n2064 & n2148;
  assign n2231 = n2230 ^ n2066;
  assign n2232 = n2231 ^ n2228;
  assign n2233 = n2229 & ~n2232;
  assign n2234 = n2233 ^ x73;
  assign n2235 = n2234 ^ x74;
  assign n2236 = n2070 & n2148;
  assign n2237 = n2236 ^ n2072;
  assign n2238 = n2237 ^ n2234;
  assign n2239 = n2235 & ~n2238;
  assign n2240 = n2239 ^ x74;
  assign n2241 = n2240 ^ x75;
  assign n2242 = n2076 & n2148;
  assign n2243 = n2242 ^ n2078;
  assign n2244 = n2243 ^ n2240;
  assign n2245 = n2241 & n2244;
  assign n2246 = n2245 ^ x75;
  assign n2247 = n2246 ^ x76;
  assign n2248 = n2081 ^ x75;
  assign n2249 = n2148 & n2248;
  assign n2250 = n2249 ^ n1978;
  assign n2251 = n2250 ^ n2246;
  assign n2252 = n2247 & n2251;
  assign n2253 = n2252 ^ x76;
  assign n2254 = n2253 ^ x77;
  assign n2255 = ~n2082 & ~n2085;
  assign n2256 = n2255 ^ x76;
  assign n2257 = n2148 & ~n2256;
  assign n2258 = n2257 ^ n1975;
  assign n2259 = n2258 ^ n2253;
  assign n2260 = n2254 & n2259;
  assign n2261 = n2260 ^ x77;
  assign n2262 = n2261 ^ x78;
  assign n2263 = n2092 & n2148;
  assign n2264 = n2263 ^ n2094;
  assign n2265 = n2264 ^ n2261;
  assign n2266 = n2262 & ~n2265;
  assign n2267 = n2266 ^ x78;
  assign n2268 = n2267 ^ x79;
  assign n2269 = n2098 & n2148;
  assign n2270 = n2269 ^ n2100;
  assign n2271 = n2270 ^ n2267;
  assign n2272 = n2268 & ~n2271;
  assign n2273 = n2272 ^ x79;
  assign n2274 = ~n2159 & ~n2273;
  assign n2275 = n2274 ^ n2155;
  assign n2276 = n2275 ^ n2155;
  assign n2277 = ~x80 & ~n2158;
  assign n2278 = n2277 ^ n2155;
  assign n2279 = n2278 ^ n2155;
  assign n2280 = ~n2276 & ~n2279;
  assign n2281 = n2280 ^ n2155;
  assign n2282 = n2156 & ~n2281;
  assign n2283 = n2282 ^ x81;
  assign n2284 = n2283 ^ x82;
  assign n2285 = n2116 & n2148;
  assign n2286 = n2285 ^ n2118;
  assign n2287 = n2286 ^ n2283;
  assign n2288 = n2284 & ~n2287;
  assign n2289 = n2288 ^ x82;
  assign n2290 = n2289 ^ x83;
  assign n2291 = n2122 & n2148;
  assign n2292 = n2291 ^ n2124;
  assign n2293 = n2292 ^ n2289;
  assign n2294 = n2290 & n2293;
  assign n2295 = n2294 ^ x83;
  assign n2296 = ~n2153 & ~n2295;
  assign n2297 = ~x84 & ~n2152;
  assign n2298 = n2134 & n2148;
  assign n2299 = n2298 ^ n2136;
  assign n2300 = ~x85 & n2299;
  assign n2301 = ~n2297 & ~n2300;
  assign n2302 = ~n2296 & n2301;
  assign n2149 = n1967 & ~n2148;
  assign n2150 = ~n240 & ~n2149;
  assign n2303 = x86 & n2150;
  assign n2304 = n1819 & ~n2303;
  assign n2305 = x85 & ~n2299;
  assign n2306 = n2304 & ~n2305;
  assign n2307 = ~n2302 & n2306;
  assign n2308 = n1968 & ~n2150;
  assign n2309 = ~n2307 & ~n2308;
  assign n2314 = n2199 & ~n2309;
  assign n2315 = n2314 ^ n2201;
  assign n2316 = n2315 ^ x69;
  assign n2317 = n2192 & ~n2309;
  assign n2318 = n2317 ^ n2195;
  assign n2319 = x68 & n2318;
  assign n2320 = n2309 ^ n288;
  assign n2321 = n2320 ^ n288;
  assign n2322 = n289 ^ n288;
  assign n2323 = ~n2321 & n2322;
  assign n2324 = n2323 ^ n288;
  assign n2325 = ~n2148 & n2324;
  assign n2326 = n2325 ^ n288;
  assign n2327 = x41 & n2326;
  assign n2328 = n2183 ^ n2148;
  assign n2329 = n2328 ^ n2183;
  assign n2330 = ~x41 & n288;
  assign n2331 = n2330 ^ n2183;
  assign n2332 = ~n2329 & n2331;
  assign n2333 = n2332 ^ n2183;
  assign n2334 = ~n202 & ~n2333;
  assign n2335 = n2334 ^ n2175;
  assign n2336 = ~n2309 & ~n2335;
  assign n2337 = n2336 ^ n2175;
  assign n2338 = ~n2327 & ~n2337;
  assign n2339 = n2338 ^ x42;
  assign n2340 = n2339 ^ x66;
  assign n2341 = x64 & ~n2309;
  assign n2342 = x41 & ~x65;
  assign n2343 = x40 & n2342;
  assign n2344 = n2343 ^ x41;
  assign n2345 = n2341 & n2344;
  assign n2346 = ~x40 & x64;
  assign n2347 = ~x65 & ~n2346;
  assign n2348 = ~x41 & ~n2347;
  assign n2349 = n2309 & n2348;
  assign n2350 = ~x40 & x65;
  assign n2351 = x64 & n2350;
  assign n2352 = ~x41 & n202;
  assign n2353 = ~n2351 & ~n2352;
  assign n2354 = ~n2349 & n2353;
  assign n2355 = ~n2345 & n2354;
  assign n2356 = n2355 ^ n2339;
  assign n2357 = n2340 & n2356;
  assign n2358 = n2357 ^ x66;
  assign n2359 = n2358 ^ x67;
  assign n2360 = n2188 ^ x66;
  assign n2361 = ~n2309 & ~n2360;
  assign n2362 = n2361 ^ n2173;
  assign n2363 = n2362 ^ n2358;
  assign n2364 = n2359 & ~n2363;
  assign n2365 = n2364 ^ x67;
  assign n2366 = ~n2319 & ~n2365;
  assign n2367 = n2366 ^ n2315;
  assign n2368 = n2367 ^ n2315;
  assign n2369 = ~x68 & ~n2318;
  assign n2370 = n2369 ^ n2315;
  assign n2371 = n2370 ^ n2315;
  assign n2372 = ~n2368 & ~n2371;
  assign n2373 = n2372 ^ n2315;
  assign n2374 = n2316 & ~n2373;
  assign n2375 = n2374 ^ x69;
  assign n2376 = n2375 ^ x70;
  assign n2377 = n2205 & ~n2309;
  assign n2378 = n2377 ^ n2207;
  assign n2379 = n2378 ^ n2375;
  assign n2380 = n2376 & ~n2379;
  assign n2381 = n2380 ^ x70;
  assign n2382 = n2381 ^ x71;
  assign n2383 = n2211 & ~n2309;
  assign n2384 = n2383 ^ n2213;
  assign n2385 = n2384 ^ n2381;
  assign n2386 = n2382 & n2385;
  assign n2387 = n2386 ^ x71;
  assign n2388 = n2387 ^ x72;
  assign n2389 = n2217 & ~n2309;
  assign n2390 = n2389 ^ n2219;
  assign n2391 = n2390 ^ n2387;
  assign n2392 = n2388 & ~n2391;
  assign n2393 = n2392 ^ x72;
  assign n2394 = n2393 ^ x73;
  assign n2395 = n2223 & ~n2309;
  assign n2396 = n2395 ^ n2225;
  assign n2397 = n2396 ^ n2393;
  assign n2398 = n2394 & n2397;
  assign n2399 = n2398 ^ x73;
  assign n2400 = n2399 ^ x74;
  assign n2401 = n2229 & ~n2309;
  assign n2402 = n2401 ^ n2231;
  assign n2403 = n2402 ^ n2399;
  assign n2404 = n2400 & ~n2403;
  assign n2405 = n2404 ^ x74;
  assign n2406 = n2405 ^ x75;
  assign n2407 = n2235 & ~n2309;
  assign n2408 = n2407 ^ n2237;
  assign n2409 = n2408 ^ n2405;
  assign n2410 = n2406 & ~n2409;
  assign n2411 = n2410 ^ x75;
  assign n2412 = n2411 ^ x76;
  assign n2413 = n2241 & ~n2309;
  assign n2414 = n2413 ^ n2243;
  assign n2415 = n2414 ^ n2411;
  assign n2416 = n2412 & n2415;
  assign n2417 = n2416 ^ x76;
  assign n2418 = n2417 ^ x77;
  assign n2419 = n2247 & ~n2309;
  assign n2420 = n2419 ^ n2250;
  assign n2421 = n2420 ^ n2417;
  assign n2422 = n2418 & n2421;
  assign n2423 = n2422 ^ x77;
  assign n2424 = n2423 ^ x78;
  assign n2425 = n2254 & ~n2309;
  assign n2426 = n2425 ^ n2258;
  assign n2427 = n2426 ^ n2423;
  assign n2428 = n2424 & n2427;
  assign n2429 = n2428 ^ x78;
  assign n2430 = n2429 ^ x79;
  assign n2431 = n2262 & ~n2309;
  assign n2432 = n2431 ^ n2264;
  assign n2433 = n2432 ^ n2429;
  assign n2434 = n2430 & ~n2433;
  assign n2435 = n2434 ^ x79;
  assign n2436 = n2435 ^ x80;
  assign n2437 = n2268 & ~n2309;
  assign n2438 = n2437 ^ n2270;
  assign n2439 = n2438 ^ n2435;
  assign n2440 = n2436 & ~n2439;
  assign n2441 = n2440 ^ x80;
  assign n2442 = n2441 ^ x81;
  assign n2443 = n2273 ^ x80;
  assign n2444 = ~n2309 & n2443;
  assign n2445 = n2444 ^ n2158;
  assign n2446 = n2445 ^ n2441;
  assign n2447 = n2442 & ~n2446;
  assign n2448 = n2447 ^ x81;
  assign n2449 = n2448 ^ x82;
  assign n2450 = ~n2274 & ~n2277;
  assign n2451 = n2450 ^ x81;
  assign n2452 = ~n2309 & n2451;
  assign n2453 = n2452 ^ n2155;
  assign n2454 = n2453 ^ n2448;
  assign n2455 = n2449 & ~n2454;
  assign n2456 = n2455 ^ x82;
  assign n2457 = n2456 ^ x83;
  assign n2458 = n2284 & ~n2309;
  assign n2459 = n2458 ^ n2286;
  assign n2460 = n2459 ^ n2456;
  assign n2461 = n2457 & ~n2460;
  assign n2462 = n2461 ^ x83;
  assign n2463 = n2462 ^ x84;
  assign n2464 = n2290 & ~n2309;
  assign n2465 = n2464 ^ n2292;
  assign n2466 = n2465 ^ n2462;
  assign n2467 = n2463 & n2466;
  assign n2468 = n2467 ^ x84;
  assign n2469 = n2468 ^ x85;
  assign n2470 = n2295 ^ x84;
  assign n2471 = ~n2309 & n2470;
  assign n2472 = n2471 ^ n2152;
  assign n2473 = n2472 ^ n2468;
  assign n2474 = n2469 & ~n2473;
  assign n2475 = n2474 ^ x85;
  assign n2476 = n2475 ^ x86;
  assign n2477 = ~n2296 & ~n2297;
  assign n2478 = n2477 ^ x85;
  assign n2479 = ~n2309 & n2478;
  assign n2480 = n2479 ^ n2299;
  assign n2481 = n2480 ^ n2475;
  assign n2482 = n2476 & n2481;
  assign n2483 = n2482 ^ x86;
  assign n2488 = n2483 ^ x87;
  assign n2310 = ~n240 & ~n2309;
  assign n2311 = ~n2150 & ~n2310;
  assign n2489 = n2483 ^ n2311;
  assign n2490 = n2488 & n2489;
  assign n2491 = n2490 ^ x87;
  assign n2492 = n168 & ~n2491;
  assign n2680 = n2492 ^ x65;
  assign n2681 = n2492 ^ x64;
  assign n2682 = n2681 ^ x64;
  assign n2312 = x88 & ~n2311;
  assign n2313 = n167 & ~n2312;
  assign n2484 = n168 & ~n2483;
  assign n2485 = ~n1819 & n2311;
  assign n2486 = ~n2484 & n2485;
  assign n2487 = ~x88 & n2486;
  assign n2493 = n2394 & n2492;
  assign n2494 = n2493 ^ n2396;
  assign n2495 = n2494 ^ x74;
  assign n2496 = n2388 & n2492;
  assign n2497 = n2496 ^ n2390;
  assign n2498 = x73 & n2497;
  assign n2499 = x65 & n168;
  assign n2500 = n2499 ^ n288;
  assign n2501 = n2500 ^ n288;
  assign n2502 = n2491 ^ n288;
  assign n2503 = n2502 ^ n288;
  assign n2504 = n2501 & ~n2503;
  assign n2505 = n2504 ^ n288;
  assign n2506 = n2309 & n2505;
  assign n2507 = n2506 ^ n288;
  assign n2508 = x40 & n2507;
  assign n2509 = n2351 ^ n2309;
  assign n2510 = n2509 ^ n2351;
  assign n2511 = ~x65 & n2346;
  assign n2512 = n2511 ^ n2351;
  assign n2513 = n2510 & n2512;
  assign n2514 = n2513 ^ n2351;
  assign n2515 = ~n202 & ~n2514;
  assign n2516 = n2515 ^ n2341;
  assign n2517 = n2492 & ~n2516;
  assign n2518 = n2517 ^ n2341;
  assign n2519 = ~n2508 & ~n2518;
  assign n2520 = n2519 ^ x41;
  assign n2521 = n2520 ^ x66;
  assign n2522 = x64 & n2492;
  assign n2523 = x39 & ~x65;
  assign n2524 = x40 & ~n2523;
  assign n2525 = n2522 & n2524;
  assign n2526 = ~x39 & n2346;
  assign n2527 = ~n2350 & ~n2526;
  assign n2528 = ~n2492 & ~n2527;
  assign n2529 = ~x39 & x65;
  assign n2530 = n2529 ^ n2350;
  assign n2531 = x64 & n2530;
  assign n2532 = n2531 ^ n2350;
  assign n2533 = ~n2528 & ~n2532;
  assign n2534 = ~n2525 & n2533;
  assign n2535 = n2534 ^ n2520;
  assign n2536 = n2521 & n2535;
  assign n2537 = n2536 ^ x66;
  assign n2538 = n2537 ^ x67;
  assign n2539 = n2355 ^ x66;
  assign n2540 = n2492 & ~n2539;
  assign n2541 = n2540 ^ n2339;
  assign n2542 = n2541 ^ n2537;
  assign n2543 = n2538 & ~n2542;
  assign n2544 = n2543 ^ x67;
  assign n2545 = n2544 ^ x68;
  assign n2546 = n2359 & n2492;
  assign n2547 = n2546 ^ n2362;
  assign n2548 = n2547 ^ n2544;
  assign n2549 = n2545 & ~n2548;
  assign n2550 = n2549 ^ x68;
  assign n2551 = n2550 ^ x69;
  assign n2552 = n2365 ^ x68;
  assign n2553 = n2492 & n2552;
  assign n2554 = n2553 ^ n2318;
  assign n2555 = n2554 ^ n2550;
  assign n2556 = n2551 & ~n2555;
  assign n2557 = n2556 ^ x69;
  assign n2558 = n2557 ^ x70;
  assign n2559 = ~n2366 & ~n2369;
  assign n2560 = n2559 ^ n2316;
  assign n2561 = n2560 ^ n2315;
  assign n2562 = n2492 & n2561;
  assign n2563 = n2562 ^ n2315;
  assign n2564 = n2563 ^ n2557;
  assign n2565 = n2558 & ~n2564;
  assign n2566 = n2565 ^ x70;
  assign n2567 = n2566 ^ x71;
  assign n2568 = n2376 & n2492;
  assign n2569 = n2568 ^ n2378;
  assign n2570 = n2569 ^ n2566;
  assign n2571 = n2567 & ~n2570;
  assign n2572 = n2571 ^ x71;
  assign n2573 = n2572 ^ x72;
  assign n2574 = n2382 & n2492;
  assign n2575 = n2574 ^ n2384;
  assign n2576 = n2575 ^ n2572;
  assign n2577 = n2573 & n2576;
  assign n2578 = n2577 ^ x72;
  assign n2579 = ~n2498 & ~n2578;
  assign n2580 = n2579 ^ n2494;
  assign n2581 = n2580 ^ n2494;
  assign n2582 = ~x73 & ~n2497;
  assign n2583 = n2582 ^ n2494;
  assign n2584 = n2583 ^ n2494;
  assign n2585 = ~n2581 & ~n2584;
  assign n2586 = n2585 ^ n2494;
  assign n2587 = ~n2495 & n2586;
  assign n2588 = n2587 ^ x74;
  assign n2589 = n2588 ^ x75;
  assign n2590 = n2400 & n2492;
  assign n2591 = n2590 ^ n2402;
  assign n2592 = n2591 ^ n2588;
  assign n2593 = n2589 & ~n2592;
  assign n2594 = n2593 ^ x75;
  assign n2595 = n2594 ^ x76;
  assign n2596 = n2406 & n2492;
  assign n2597 = n2596 ^ n2408;
  assign n2598 = n2597 ^ n2594;
  assign n2599 = n2595 & ~n2598;
  assign n2600 = n2599 ^ x76;
  assign n2601 = n2600 ^ x77;
  assign n2602 = n2412 & n2492;
  assign n2603 = n2602 ^ n2414;
  assign n2604 = n2603 ^ n2600;
  assign n2605 = n2601 & n2604;
  assign n2606 = n2605 ^ x77;
  assign n2607 = n2606 ^ x78;
  assign n2608 = n2418 & n2492;
  assign n2609 = n2608 ^ n2420;
  assign n2610 = n2609 ^ n2606;
  assign n2611 = n2607 & n2610;
  assign n2612 = n2611 ^ x78;
  assign n2613 = n2612 ^ x79;
  assign n2614 = n2424 & n2492;
  assign n2615 = n2614 ^ n2426;
  assign n2616 = n2615 ^ n2612;
  assign n2617 = n2613 & n2616;
  assign n2618 = n2617 ^ x79;
  assign n2619 = n2618 ^ x80;
  assign n2620 = n2430 & n2492;
  assign n2621 = n2620 ^ n2432;
  assign n2622 = n2621 ^ n2618;
  assign n2623 = n2619 & ~n2622;
  assign n2624 = n2623 ^ x80;
  assign n2625 = n2624 ^ x81;
  assign n2626 = n2436 & n2492;
  assign n2627 = n2626 ^ n2438;
  assign n2628 = n2627 ^ n2624;
  assign n2629 = n2625 & ~n2628;
  assign n2630 = n2629 ^ x81;
  assign n2631 = n2630 ^ x82;
  assign n2632 = n2442 & n2492;
  assign n2633 = n2632 ^ n2445;
  assign n2634 = n2633 ^ n2630;
  assign n2635 = n2631 & ~n2634;
  assign n2636 = n2635 ^ x82;
  assign n2637 = n2636 ^ x83;
  assign n2638 = n2449 & n2492;
  assign n2639 = n2638 ^ n2453;
  assign n2640 = n2639 ^ n2636;
  assign n2641 = n2637 & ~n2640;
  assign n2642 = n2641 ^ x83;
  assign n2643 = n2642 ^ x84;
  assign n2644 = n2457 & n2492;
  assign n2645 = n2644 ^ n2459;
  assign n2646 = n2645 ^ n2642;
  assign n2647 = n2643 & ~n2646;
  assign n2648 = n2647 ^ x84;
  assign n2649 = n2648 ^ x85;
  assign n2650 = n2463 & n2492;
  assign n2651 = n2650 ^ n2465;
  assign n2652 = n2651 ^ n2648;
  assign n2653 = n2649 & n2652;
  assign n2654 = n2653 ^ x85;
  assign n2655 = n2654 ^ x86;
  assign n2656 = n2469 & n2492;
  assign n2657 = n2656 ^ n2472;
  assign n2658 = n2657 ^ n2654;
  assign n2659 = n2655 & ~n2658;
  assign n2660 = n2659 ^ x86;
  assign n2661 = n2660 ^ x87;
  assign n2662 = n2476 & n2492;
  assign n2663 = n2662 ^ n2480;
  assign n2664 = n2663 ^ n2660;
  assign n2665 = n2661 & ~n2664;
  assign n2666 = n2665 ^ n2660;
  assign n2667 = ~n2487 & n2666;
  assign n2668 = n2313 & ~n2667;
  assign n2683 = n2668 ^ x64;
  assign n2684 = ~n2682 & n2683;
  assign n2685 = n2684 ^ x64;
  assign n2686 = n2680 & n2685;
  assign n2687 = x39 & n2686;
  assign n2688 = ~x65 & n2492;
  assign n2689 = ~n288 & ~n2492;
  assign n2690 = ~x39 & ~n2689;
  assign n2691 = ~n202 & ~n2690;
  assign n2692 = ~n2688 & ~n2691;
  assign n2693 = n2692 ^ n2522;
  assign n2694 = n2668 & n2693;
  assign n2695 = n2694 ^ n2522;
  assign n2696 = ~n2687 & ~n2695;
  assign n2697 = n2696 ^ x40;
  assign n2698 = n2697 ^ x66;
  assign n2699 = ~x38 & ~n2668;
  assign n2700 = ~x38 & x65;
  assign n2701 = ~n2699 & ~n2700;
  assign n2702 = x64 & ~n2523;
  assign n2703 = ~n2701 & n2702;
  assign n2704 = x64 & n2668;
  assign n2705 = x38 & n2523;
  assign n2706 = n2705 ^ x39;
  assign n2707 = n2706 ^ n2529;
  assign n2708 = n2704 & n2707;
  assign n2709 = n2708 ^ n2529;
  assign n2710 = ~n2703 & ~n2709;
  assign n2711 = n2710 ^ n2697;
  assign n2712 = n2698 & n2711;
  assign n2713 = n2712 ^ x66;
  assign n2714 = n2713 ^ x67;
  assign n2715 = n2534 ^ x66;
  assign n2716 = n2668 & ~n2715;
  assign n2717 = n2716 ^ n2520;
  assign n2718 = n2717 ^ n2713;
  assign n2719 = n2714 & ~n2718;
  assign n2720 = n2719 ^ x67;
  assign n2721 = n2720 ^ x68;
  assign n2722 = n2538 & n2668;
  assign n2723 = n2722 ^ n2541;
  assign n2724 = n2723 ^ n2720;
  assign n2725 = n2721 & ~n2724;
  assign n2726 = n2725 ^ x68;
  assign n2727 = n2726 ^ x69;
  assign n2728 = n2545 & n2668;
  assign n2729 = n2728 ^ n2547;
  assign n2730 = n2729 ^ n2726;
  assign n2731 = n2727 & ~n2730;
  assign n2732 = n2731 ^ x69;
  assign n2733 = n2732 ^ x70;
  assign n2674 = n2661 & n2668;
  assign n2675 = n2674 ^ n2663;
  assign n2676 = n2675 ^ x88;
  assign n2677 = n2655 & n2668;
  assign n2678 = n2677 ^ n2657;
  assign n2679 = x87 & n2678;
  assign n2669 = n2554 ^ x69;
  assign n2670 = n2669 ^ n2550;
  assign n2671 = n2670 ^ n2554;
  assign n2672 = n2668 & n2671;
  assign n2673 = n2672 ^ n2554;
  assign n2734 = n2732 ^ n2673;
  assign n2735 = n2733 & ~n2734;
  assign n2736 = n2735 ^ x70;
  assign n2737 = n2736 ^ x71;
  assign n2738 = n2558 & n2668;
  assign n2739 = n2738 ^ n2563;
  assign n2740 = n2739 ^ n2736;
  assign n2741 = n2737 & ~n2740;
  assign n2742 = n2741 ^ x71;
  assign n2743 = n2742 ^ x72;
  assign n2744 = n2567 & n2668;
  assign n2745 = n2744 ^ n2569;
  assign n2746 = n2745 ^ n2742;
  assign n2747 = n2743 & ~n2746;
  assign n2748 = n2747 ^ x72;
  assign n2749 = n2748 ^ x73;
  assign n2750 = n2573 & n2668;
  assign n2751 = n2750 ^ n2575;
  assign n2752 = n2751 ^ n2748;
  assign n2753 = n2749 & n2752;
  assign n2754 = n2753 ^ x73;
  assign n2755 = n2754 ^ x74;
  assign n2756 = n2578 ^ x73;
  assign n2757 = n2668 & n2756;
  assign n2758 = n2757 ^ n2497;
  assign n2759 = n2758 ^ n2754;
  assign n2760 = n2755 & ~n2759;
  assign n2761 = n2760 ^ x74;
  assign n2762 = n2761 ^ x75;
  assign n2763 = ~n2579 & ~n2582;
  assign n2764 = n2763 ^ x74;
  assign n2765 = n2668 & n2764;
  assign n2766 = n2765 ^ n2494;
  assign n2767 = n2766 ^ n2761;
  assign n2768 = n2762 & n2767;
  assign n2769 = n2768 ^ x75;
  assign n2770 = n2769 ^ x76;
  assign n2771 = n2589 & n2668;
  assign n2772 = n2771 ^ n2591;
  assign n2773 = n2772 ^ n2769;
  assign n2774 = n2770 & ~n2773;
  assign n2775 = n2774 ^ x76;
  assign n2776 = n2775 ^ x77;
  assign n2777 = n2595 & n2668;
  assign n2778 = n2777 ^ n2597;
  assign n2779 = n2778 ^ n2775;
  assign n2780 = n2776 & ~n2779;
  assign n2781 = n2780 ^ x77;
  assign n2782 = n2781 ^ x78;
  assign n2783 = n2601 & n2668;
  assign n2784 = n2783 ^ n2603;
  assign n2785 = n2784 ^ n2781;
  assign n2786 = n2782 & n2785;
  assign n2787 = n2786 ^ x78;
  assign n2788 = n2787 ^ x79;
  assign n2789 = n2607 & n2668;
  assign n2790 = n2789 ^ n2609;
  assign n2791 = n2790 ^ n2787;
  assign n2792 = n2788 & n2791;
  assign n2793 = n2792 ^ x79;
  assign n2794 = n2793 ^ x80;
  assign n2795 = n2613 & n2668;
  assign n2796 = n2795 ^ n2615;
  assign n2797 = n2796 ^ n2793;
  assign n2798 = n2794 & n2797;
  assign n2799 = n2798 ^ x80;
  assign n2800 = n2799 ^ x81;
  assign n2801 = n2619 & n2668;
  assign n2802 = n2801 ^ n2621;
  assign n2803 = n2802 ^ n2799;
  assign n2804 = n2800 & ~n2803;
  assign n2805 = n2804 ^ x81;
  assign n2806 = n2805 ^ x82;
  assign n2807 = n2625 & n2668;
  assign n2808 = n2807 ^ n2627;
  assign n2809 = n2808 ^ n2805;
  assign n2810 = n2806 & ~n2809;
  assign n2811 = n2810 ^ x82;
  assign n2812 = n2811 ^ x83;
  assign n2813 = n2631 & n2668;
  assign n2814 = n2813 ^ n2633;
  assign n2815 = n2814 ^ n2811;
  assign n2816 = n2812 & ~n2815;
  assign n2817 = n2816 ^ x83;
  assign n2818 = n2817 ^ x84;
  assign n2819 = n2637 & n2668;
  assign n2820 = n2819 ^ n2639;
  assign n2821 = n2820 ^ n2817;
  assign n2822 = n2818 & ~n2821;
  assign n2823 = n2822 ^ x84;
  assign n2824 = n2823 ^ x85;
  assign n2825 = n2643 & n2668;
  assign n2826 = n2825 ^ n2645;
  assign n2827 = n2826 ^ n2823;
  assign n2828 = n2824 & ~n2827;
  assign n2829 = n2828 ^ x85;
  assign n2830 = n2829 ^ x86;
  assign n2831 = n2649 & n2668;
  assign n2832 = n2831 ^ n2651;
  assign n2833 = n2832 ^ n2829;
  assign n2834 = n2830 & n2833;
  assign n2835 = n2834 ^ x86;
  assign n2836 = ~n2679 & ~n2835;
  assign n2837 = n2836 ^ n2675;
  assign n2838 = n2837 ^ n2675;
  assign n2839 = ~x87 & ~n2678;
  assign n2840 = n2839 ^ n2675;
  assign n2841 = n2840 ^ n2675;
  assign n2842 = ~n2838 & ~n2841;
  assign n2843 = n2842 ^ n2675;
  assign n2844 = ~n2676 & n2843;
  assign n2845 = n2844 ^ x88;
  assign n2846 = n2845 ^ x89;
  assign n2847 = n2486 & ~n2668;
  assign n2848 = ~n240 & ~n2847;
  assign n2849 = n2848 ^ n2845;
  assign n2850 = n2846 & ~n2849;
  assign n2851 = n2850 ^ x89;
  assign n2852 = n166 & ~n2851;
  assign n2853 = n2733 & n2852;
  assign n2854 = n2853 ^ n2673;
  assign n2855 = ~x71 & ~n2854;
  assign n2856 = n2737 & n2852;
  assign n2857 = n2856 ^ n2739;
  assign n2858 = ~x72 & ~n2857;
  assign n2859 = ~n2855 & ~n2858;
  assign n2860 = n2668 ^ x65;
  assign n2861 = n2860 ^ x38;
  assign n2862 = n2683 ^ x64;
  assign n2863 = n2852 ^ x64;
  assign n2864 = ~n2862 & n2863;
  assign n2865 = n2864 ^ x64;
  assign n2866 = n2865 ^ n2860;
  assign n2867 = n2861 & n2866;
  assign n2868 = n2867 ^ n2864;
  assign n2869 = n2868 ^ x64;
  assign n2870 = n2869 ^ x38;
  assign n2871 = n2860 & n2870;
  assign n2872 = n2871 ^ n2860;
  assign n2873 = ~n288 & ~n2668;
  assign n2874 = ~n2701 & ~n2873;
  assign n2875 = ~n202 & ~n2874;
  assign n2876 = n2875 ^ n2704;
  assign n2877 = n2852 & ~n2876;
  assign n2878 = n2877 ^ n2704;
  assign n2879 = ~n2872 & ~n2878;
  assign n2880 = n2879 ^ x39;
  assign n2881 = n2880 ^ x66;
  assign n2882 = ~x38 & ~n2852;
  assign n2883 = ~x65 & ~n2882;
  assign n2884 = ~x37 & x64;
  assign n2885 = ~n2883 & n2884;
  assign n2886 = x64 & n2852;
  assign n2887 = x38 & ~x65;
  assign n2888 = x37 & n2887;
  assign n2889 = n2888 ^ x38;
  assign n2890 = n2889 ^ n2700;
  assign n2891 = n2886 & n2890;
  assign n2892 = n2891 ^ n2700;
  assign n2893 = ~n2885 & ~n2892;
  assign n2894 = n2893 ^ n2880;
  assign n2895 = n2881 & n2894;
  assign n2896 = n2895 ^ x66;
  assign n2897 = n2896 ^ x67;
  assign n2898 = n2710 ^ x66;
  assign n2899 = n2852 & ~n2898;
  assign n2900 = n2899 ^ n2697;
  assign n2901 = n2900 ^ n2896;
  assign n2902 = n2897 & ~n2901;
  assign n2903 = n2902 ^ x67;
  assign n2904 = n2903 ^ x68;
  assign n2905 = n2714 & n2852;
  assign n2906 = n2905 ^ n2717;
  assign n2907 = n2906 ^ n2903;
  assign n2908 = n2904 & ~n2907;
  assign n2909 = n2908 ^ x68;
  assign n2910 = n2909 ^ x69;
  assign n2911 = n2721 & n2852;
  assign n2912 = n2911 ^ n2723;
  assign n2913 = n2912 ^ n2909;
  assign n2914 = n2910 & ~n2913;
  assign n2915 = n2914 ^ x69;
  assign n2916 = n2915 ^ x70;
  assign n2917 = n2727 & n2852;
  assign n2918 = n2917 ^ n2729;
  assign n2919 = n2918 ^ n2915;
  assign n2920 = n2916 & ~n2919;
  assign n2921 = n2920 ^ x70;
  assign n2922 = n2859 & n2921;
  assign n2923 = n2857 ^ x72;
  assign n2924 = x71 & n2854;
  assign n2925 = n2924 ^ n2857;
  assign n2926 = n2923 & ~n2925;
  assign n2927 = n2926 ^ x72;
  assign n2928 = ~n2922 & ~n2927;
  assign n2929 = n2928 ^ x73;
  assign n2930 = n2743 & n2852;
  assign n2931 = n2930 ^ n2745;
  assign n2932 = n2931 ^ n2928;
  assign n2933 = ~n2929 & n2932;
  assign n2934 = n2933 ^ x73;
  assign n2935 = n2934 ^ x74;
  assign n2936 = n2749 & n2852;
  assign n2937 = n2936 ^ n2751;
  assign n2938 = n2937 ^ n2934;
  assign n2939 = n2935 & n2938;
  assign n2940 = n2939 ^ x74;
  assign n2941 = n2940 ^ x75;
  assign n2942 = n2755 & n2852;
  assign n2943 = n2942 ^ n2758;
  assign n2944 = n2943 ^ n2940;
  assign n2945 = n2941 & ~n2944;
  assign n2946 = n2945 ^ x75;
  assign n2947 = n2946 ^ x76;
  assign n2948 = n2762 & n2852;
  assign n2949 = n2948 ^ n2766;
  assign n2950 = n2949 ^ n2946;
  assign n2951 = n2947 & n2950;
  assign n2952 = n2951 ^ x76;
  assign n2953 = n2952 ^ x77;
  assign n2954 = n2770 & n2852;
  assign n2955 = n2954 ^ n2772;
  assign n2956 = n2955 ^ n2952;
  assign n2957 = n2953 & ~n2956;
  assign n2958 = n2957 ^ x77;
  assign n2959 = n2958 ^ x78;
  assign n2960 = n2776 & n2852;
  assign n2961 = n2960 ^ n2778;
  assign n2962 = n2961 ^ n2958;
  assign n2963 = n2959 & ~n2962;
  assign n2964 = n2963 ^ x78;
  assign n2965 = n2964 ^ x79;
  assign n2966 = n2782 & n2852;
  assign n2967 = n2966 ^ n2784;
  assign n2968 = n2967 ^ n2964;
  assign n2969 = n2965 & n2968;
  assign n2970 = n2969 ^ x79;
  assign n2971 = n2970 ^ x80;
  assign n2972 = n2788 & n2852;
  assign n2973 = n2972 ^ n2790;
  assign n2974 = n2973 ^ n2970;
  assign n2975 = n2971 & n2974;
  assign n2976 = n2975 ^ x80;
  assign n2977 = n2976 ^ x81;
  assign n2978 = n2794 & n2852;
  assign n2979 = n2978 ^ n2796;
  assign n2980 = n2979 ^ n2976;
  assign n2981 = n2977 & n2980;
  assign n2982 = n2981 ^ x81;
  assign n2983 = n2982 ^ x82;
  assign n2984 = n2800 & n2852;
  assign n2985 = n2984 ^ n2802;
  assign n2986 = n2985 ^ n2982;
  assign n2987 = n2983 & ~n2986;
  assign n2988 = n2987 ^ x82;
  assign n2989 = n2988 ^ x83;
  assign n2990 = n2806 & n2852;
  assign n2991 = n2990 ^ n2808;
  assign n2992 = n2991 ^ n2988;
  assign n2993 = n2989 & ~n2992;
  assign n2994 = n2993 ^ x83;
  assign n2995 = n2994 ^ x84;
  assign n2996 = n2812 & n2852;
  assign n2997 = n2996 ^ n2814;
  assign n2998 = n2997 ^ n2994;
  assign n2999 = n2995 & ~n2998;
  assign n3000 = n2999 ^ x84;
  assign n3001 = n3000 ^ x85;
  assign n3002 = n2818 & n2852;
  assign n3003 = n3002 ^ n2820;
  assign n3004 = n3003 ^ n3000;
  assign n3005 = n3001 & ~n3004;
  assign n3006 = n3005 ^ x85;
  assign n3007 = n3006 ^ x86;
  assign n3008 = n2824 & n2852;
  assign n3009 = n3008 ^ n2826;
  assign n3010 = n3009 ^ n3006;
  assign n3011 = n3007 & ~n3010;
  assign n3012 = n3011 ^ x86;
  assign n3013 = n3012 ^ x87;
  assign n3014 = n2830 & n2852;
  assign n3015 = n3014 ^ n2832;
  assign n3016 = n3015 ^ n3012;
  assign n3017 = n3013 & n3016;
  assign n3018 = n3017 ^ x87;
  assign n3019 = n3018 ^ x88;
  assign n3020 = n2835 ^ x87;
  assign n3021 = n2852 & n3020;
  assign n3022 = n3021 ^ n2678;
  assign n3023 = n3022 ^ n3018;
  assign n3024 = n3019 & ~n3023;
  assign n3025 = n3024 ^ x88;
  assign n3026 = n3025 ^ x89;
  assign n3027 = ~n2836 & ~n2839;
  assign n3028 = n3027 ^ x88;
  assign n3029 = n2852 & n3028;
  assign n3030 = n3029 ^ n2675;
  assign n3031 = n3030 ^ n3025;
  assign n3032 = n3026 & n3031;
  assign n3033 = n3032 ^ x89;
  assign n3034 = n3033 ^ x90;
  assign n3035 = ~x90 & ~n2851;
  assign n3036 = ~n2848 & ~n3035;
  assign n3037 = ~n240 & ~n3036;
  assign n3038 = n3037 ^ n3033;
  assign n3039 = n3034 & ~n3038;
  assign n3040 = n3039 ^ x90;
  assign n3041 = n165 & ~n3040;
  assign n3042 = n3026 & n3041;
  assign n3043 = n3042 ^ n3030;
  assign n3044 = n3043 ^ x90;
  assign n3045 = n3019 & n3041;
  assign n3046 = n3045 ^ n3022;
  assign n3047 = x89 & n3046;
  assign n3048 = n2971 & n3041;
  assign n3049 = n3048 ^ n2973;
  assign n3050 = n3049 ^ x81;
  assign n3051 = n2965 & n3041;
  assign n3052 = n3051 ^ n2967;
  assign n3053 = x80 & ~n3052;
  assign n3054 = n2852 ^ x65;
  assign n3055 = n2884 & ~n3054;
  assign n3056 = ~n202 & ~n3055;
  assign n3057 = x65 & n2852;
  assign n3058 = x37 & ~n3057;
  assign n3059 = x65 & n3058;
  assign n3060 = n3056 & ~n3059;
  assign n3061 = n3060 ^ n2886;
  assign n3062 = n3060 ^ n3058;
  assign n3063 = n3060 ^ n3041;
  assign n3064 = n3060 & n3063;
  assign n3065 = n3064 ^ n3060;
  assign n3066 = n3062 & n3065;
  assign n3067 = n3066 ^ n3064;
  assign n3068 = n3067 ^ n3060;
  assign n3069 = n3068 ^ n3041;
  assign n3070 = ~n3061 & n3069;
  assign n3071 = n3070 ^ n2886;
  assign n3072 = n3071 ^ x38;
  assign n3073 = n3072 ^ x66;
  assign n3074 = x64 & n3041;
  assign n3075 = x37 & ~x65;
  assign n3076 = x36 & n3075;
  assign n3077 = n3076 ^ x37;
  assign n3078 = n3074 & n3077;
  assign n3080 = x65 ^ x37;
  assign n3087 = n3080 ^ x65;
  assign n3079 = x65 ^ x36;
  assign n3081 = n3080 ^ n3079;
  assign n3082 = n3081 ^ x65;
  assign n3083 = n3079 ^ x64;
  assign n3084 = n3083 ^ n3079;
  assign n3085 = n3084 ^ n3082;
  assign n3086 = ~n3082 & ~n3085;
  assign n3088 = n3087 ^ n3086;
  assign n3089 = n3088 ^ n3082;
  assign n3090 = n3041 ^ x65;
  assign n3091 = n3090 ^ x65;
  assign n3092 = n3086 ^ n3082;
  assign n3093 = ~n3091 & ~n3092;
  assign n3094 = n3093 ^ x65;
  assign n3095 = ~n3089 & n3094;
  assign n3096 = n3095 ^ x65;
  assign n3097 = n3096 ^ x65;
  assign n3098 = n3097 ^ x65;
  assign n3099 = ~n3078 & ~n3098;
  assign n3100 = n3099 ^ n3072;
  assign n3101 = ~n3073 & ~n3100;
  assign n3102 = n3101 ^ x66;
  assign n3103 = n3102 ^ x67;
  assign n3104 = n2893 ^ x66;
  assign n3105 = n3041 & ~n3104;
  assign n3106 = n3105 ^ n2880;
  assign n3107 = n3106 ^ n3102;
  assign n3108 = n3103 & ~n3107;
  assign n3109 = n3108 ^ x67;
  assign n3110 = n3109 ^ x68;
  assign n3111 = n2897 & n3041;
  assign n3112 = n3111 ^ n2900;
  assign n3113 = n3112 ^ n3109;
  assign n3114 = n3110 & ~n3113;
  assign n3115 = n3114 ^ x68;
  assign n3116 = n3115 ^ x69;
  assign n3117 = n2904 & n3041;
  assign n3118 = n3117 ^ n2906;
  assign n3119 = n3118 ^ n3115;
  assign n3120 = n3116 & ~n3119;
  assign n3121 = n3120 ^ x69;
  assign n3122 = n3121 ^ x70;
  assign n3123 = n2910 & n3041;
  assign n3124 = n3123 ^ n2912;
  assign n3125 = n3124 ^ n3121;
  assign n3126 = n3122 & ~n3125;
  assign n3127 = n3126 ^ x70;
  assign n3128 = n3127 ^ x71;
  assign n3129 = n2916 & n3041;
  assign n3130 = n3129 ^ n2918;
  assign n3131 = n3130 ^ n3127;
  assign n3132 = n3128 & ~n3131;
  assign n3133 = n3132 ^ x71;
  assign n3134 = n3133 ^ x72;
  assign n3135 = n2921 ^ x71;
  assign n3136 = n3041 & n3135;
  assign n3137 = n3136 ^ n2854;
  assign n3138 = n3137 ^ n3133;
  assign n3139 = n3134 & ~n3138;
  assign n3140 = n3139 ^ x72;
  assign n3141 = n3140 ^ x73;
  assign n3142 = n2921 ^ n2854;
  assign n3143 = n3135 & ~n3142;
  assign n3144 = n3143 ^ x71;
  assign n3145 = n3144 ^ x72;
  assign n3146 = n3041 & n3145;
  assign n3147 = n3146 ^ n2857;
  assign n3148 = n3147 ^ n3140;
  assign n3149 = n3141 & ~n3148;
  assign n3150 = n3149 ^ x73;
  assign n3151 = n3150 ^ x74;
  assign n3152 = ~n2929 & n3041;
  assign n3153 = n3152 ^ n2931;
  assign n3154 = n3153 ^ n3150;
  assign n3155 = n3151 & ~n3154;
  assign n3156 = n3155 ^ x74;
  assign n3157 = n3156 ^ x75;
  assign n3158 = n2935 & n3041;
  assign n3159 = n3158 ^ n2937;
  assign n3160 = n3159 ^ n3156;
  assign n3161 = n3157 & n3160;
  assign n3162 = n3161 ^ x75;
  assign n3163 = n3162 ^ x76;
  assign n3164 = n2941 & n3041;
  assign n3165 = n3164 ^ n2943;
  assign n3166 = n3165 ^ n3162;
  assign n3167 = n3163 & ~n3166;
  assign n3168 = n3167 ^ x76;
  assign n3169 = n3168 ^ x77;
  assign n3170 = n2947 & n3041;
  assign n3171 = n3170 ^ n2949;
  assign n3172 = n3171 ^ n3168;
  assign n3173 = n3169 & n3172;
  assign n3174 = n3173 ^ x77;
  assign n3175 = n3174 ^ x78;
  assign n3176 = n2953 & n3041;
  assign n3177 = n3176 ^ n2955;
  assign n3178 = n3177 ^ n3174;
  assign n3179 = n3175 & ~n3178;
  assign n3180 = n3179 ^ x78;
  assign n3181 = n3180 ^ x79;
  assign n3182 = n2959 & n3041;
  assign n3183 = n3182 ^ n2961;
  assign n3184 = n3183 ^ n3180;
  assign n3185 = n3181 & ~n3184;
  assign n3186 = n3185 ^ x79;
  assign n3187 = ~n3053 & ~n3186;
  assign n3188 = n3187 ^ n3049;
  assign n3189 = n3188 ^ n3049;
  assign n3190 = ~x80 & n3052;
  assign n3191 = n3190 ^ n3049;
  assign n3192 = n3191 ^ n3049;
  assign n3193 = ~n3189 & ~n3192;
  assign n3194 = n3193 ^ n3049;
  assign n3195 = ~n3050 & n3194;
  assign n3196 = n3195 ^ x81;
  assign n3197 = n3196 ^ x82;
  assign n3198 = n2977 & n3041;
  assign n3199 = n3198 ^ n2979;
  assign n3200 = n3199 ^ n3196;
  assign n3201 = n3197 & n3200;
  assign n3202 = n3201 ^ x82;
  assign n3203 = n3202 ^ x83;
  assign n3204 = n2983 & n3041;
  assign n3205 = n3204 ^ n2985;
  assign n3206 = n3205 ^ n3202;
  assign n3207 = n3203 & ~n3206;
  assign n3208 = n3207 ^ x83;
  assign n3209 = n3208 ^ x84;
  assign n3210 = n2989 & n3041;
  assign n3211 = n3210 ^ n2991;
  assign n3212 = n3211 ^ n3208;
  assign n3213 = n3209 & ~n3212;
  assign n3214 = n3213 ^ x84;
  assign n3215 = n3214 ^ x85;
  assign n3216 = n2995 & n3041;
  assign n3217 = n3216 ^ n2997;
  assign n3218 = n3217 ^ n3214;
  assign n3219 = n3215 & ~n3218;
  assign n3220 = n3219 ^ x85;
  assign n3221 = n3220 ^ x86;
  assign n3222 = n3001 & n3041;
  assign n3223 = n3222 ^ n3003;
  assign n3224 = n3223 ^ n3220;
  assign n3225 = n3221 & ~n3224;
  assign n3226 = n3225 ^ x86;
  assign n3227 = n3226 ^ x87;
  assign n3228 = n3007 & n3041;
  assign n3229 = n3228 ^ n3009;
  assign n3230 = n3229 ^ n3226;
  assign n3231 = n3227 & ~n3230;
  assign n3232 = n3231 ^ x87;
  assign n3233 = n3232 ^ x88;
  assign n3234 = n3013 & n3041;
  assign n3235 = n3234 ^ n3015;
  assign n3236 = n3235 ^ n3232;
  assign n3237 = n3233 & n3236;
  assign n3238 = n3237 ^ x88;
  assign n3239 = ~n3047 & ~n3238;
  assign n3240 = n3239 ^ n3043;
  assign n3241 = n3240 ^ n3043;
  assign n3242 = ~x89 & ~n3046;
  assign n3243 = n3242 ^ n3043;
  assign n3244 = n3243 ^ n3043;
  assign n3245 = ~n3241 & ~n3244;
  assign n3246 = n3245 ^ n3043;
  assign n3247 = ~n3044 & n3246;
  assign n3248 = n3247 ^ x90;
  assign n3249 = n3248 ^ x91;
  assign n3250 = x90 & n3033;
  assign n3251 = n165 & ~n240;
  assign n3252 = ~n3250 & n3251;
  assign n3253 = ~n2848 & ~n3252;
  assign n3254 = n3253 ^ n3248;
  assign n3255 = n3249 & n3254;
  assign n3256 = n3255 ^ x91;
  assign n3257 = n164 & ~n3256;
  assign n3258 = ~n3239 & ~n3242;
  assign n3259 = n3258 ^ x90;
  assign n3260 = n3257 & n3259;
  assign n3261 = n3260 ^ n3043;
  assign n3262 = ~x91 & n3261;
  assign n3263 = n3253 & ~n3257;
  assign n3264 = ~n240 & ~n3263;
  assign n3265 = ~x92 & ~n3264;
  assign n3266 = ~n3262 & ~n3265;
  assign n3267 = n3238 ^ x89;
  assign n3268 = n3257 & n3267;
  assign n3269 = n3268 ^ n3046;
  assign n3270 = n3269 ^ x90;
  assign n3271 = n3233 & n3257;
  assign n3272 = n3271 ^ n3235;
  assign n3273 = ~x89 & n3272;
  assign n3274 = n3273 ^ n3269;
  assign n3275 = n3274 ^ n3269;
  assign n3276 = n3221 & n3257;
  assign n3277 = n3276 ^ n3223;
  assign n3278 = ~x87 & ~n3277;
  assign n3279 = n3227 & n3257;
  assign n3280 = n3279 ^ n3229;
  assign n3281 = ~x88 & ~n3280;
  assign n3282 = ~n3278 & ~n3281;
  assign n3283 = n3103 & n3257;
  assign n3284 = n3283 ^ n3106;
  assign n3285 = ~x68 & ~n3284;
  assign n3286 = n3110 & n3257;
  assign n3287 = n3286 ^ n3112;
  assign n3288 = ~x69 & ~n3287;
  assign n3289 = ~n3285 & ~n3288;
  assign n3290 = ~x36 & x64;
  assign n3291 = ~x35 & n3290;
  assign n3292 = ~n3257 & n3291;
  assign n3293 = ~x35 & x65;
  assign n3294 = x64 & n3293;
  assign n3295 = ~n3292 & ~n3294;
  assign n3296 = x64 & n3257;
  assign n3297 = n3296 ^ x35;
  assign n3298 = n3296 ^ x36;
  assign n3299 = n3298 ^ n3296;
  assign n3300 = n3296 & ~n3299;
  assign n3301 = n3300 ^ n3296;
  assign n3302 = ~n3297 & n3301;
  assign n3303 = n3302 ^ n3300;
  assign n3304 = n3303 ^ n3296;
  assign n3305 = n3304 ^ n3298;
  assign n3306 = ~x65 & ~n3305;
  assign n3307 = n3306 ^ n3298;
  assign n3308 = n3295 & n3307;
  assign n3309 = n3308 ^ x66;
  assign n3310 = x65 & n164;
  assign n3311 = n3310 ^ n288;
  assign n3312 = n3311 ^ n288;
  assign n3313 = n3256 ^ n288;
  assign n3314 = n3313 ^ n288;
  assign n3315 = n3312 & ~n3314;
  assign n3316 = n3315 ^ n288;
  assign n3317 = ~n3041 & n3316;
  assign n3318 = n3317 ^ n288;
  assign n3319 = x36 & n3318;
  assign n3320 = ~n3090 & n3290;
  assign n3321 = ~n202 & ~n3320;
  assign n3322 = n3321 ^ n3074;
  assign n3323 = n3257 & ~n3322;
  assign n3324 = n3323 ^ n3074;
  assign n3325 = ~n3319 & ~n3324;
  assign n3326 = n3325 ^ x37;
  assign n3327 = n3326 ^ n3308;
  assign n3328 = ~n3309 & n3327;
  assign n3329 = n3328 ^ x66;
  assign n3330 = n3329 ^ x67;
  assign n3331 = n3099 ^ x66;
  assign n3332 = n3257 & ~n3331;
  assign n3333 = n3332 ^ n3072;
  assign n3334 = n3333 ^ n3329;
  assign n3335 = n3330 & n3334;
  assign n3336 = n3335 ^ x67;
  assign n3337 = n3289 & n3336;
  assign n3338 = n3287 ^ x69;
  assign n3339 = x68 & n3284;
  assign n3340 = n3339 ^ n3287;
  assign n3341 = n3338 & ~n3340;
  assign n3342 = n3341 ^ x69;
  assign n3343 = ~n3337 & ~n3342;
  assign n3344 = n3343 ^ x70;
  assign n3345 = n3116 & n3257;
  assign n3346 = n3345 ^ n3118;
  assign n3347 = n3346 ^ n3343;
  assign n3348 = ~n3344 & n3347;
  assign n3349 = n3348 ^ x70;
  assign n3350 = n3349 ^ x71;
  assign n3351 = n3122 & n3257;
  assign n3352 = n3351 ^ n3124;
  assign n3353 = n3352 ^ n3349;
  assign n3354 = n3350 & ~n3353;
  assign n3355 = n3354 ^ x71;
  assign n3356 = n3355 ^ x72;
  assign n3357 = n3128 & n3257;
  assign n3358 = n3357 ^ n3130;
  assign n3359 = n3358 ^ n3355;
  assign n3360 = n3356 & ~n3359;
  assign n3361 = n3360 ^ x72;
  assign n3362 = n3361 ^ x73;
  assign n3363 = n3134 & n3257;
  assign n3364 = n3363 ^ n3137;
  assign n3365 = n3364 ^ n3361;
  assign n3366 = n3362 & ~n3365;
  assign n3367 = n3366 ^ x73;
  assign n3368 = n3367 ^ x74;
  assign n3369 = n3141 & n3257;
  assign n3370 = n3369 ^ n3147;
  assign n3371 = n3370 ^ n3367;
  assign n3372 = n3368 & ~n3371;
  assign n3373 = n3372 ^ x74;
  assign n3374 = n3373 ^ x75;
  assign n3375 = n3151 & n3257;
  assign n3376 = n3375 ^ n3153;
  assign n3377 = n3376 ^ n3373;
  assign n3378 = n3374 & ~n3377;
  assign n3379 = n3378 ^ x75;
  assign n3380 = n3379 ^ x76;
  assign n3381 = n3157 & n3257;
  assign n3382 = n3381 ^ n3159;
  assign n3383 = n3382 ^ n3379;
  assign n3384 = n3380 & n3383;
  assign n3385 = n3384 ^ x76;
  assign n3386 = n3385 ^ x77;
  assign n3387 = n3163 & n3257;
  assign n3388 = n3387 ^ n3165;
  assign n3389 = n3388 ^ n3385;
  assign n3390 = n3386 & ~n3389;
  assign n3391 = n3390 ^ x77;
  assign n3392 = n3391 ^ x78;
  assign n3393 = n3169 & n3257;
  assign n3394 = n3393 ^ n3171;
  assign n3395 = n3394 ^ n3391;
  assign n3396 = n3392 & n3395;
  assign n3397 = n3396 ^ x78;
  assign n3398 = n3397 ^ x79;
  assign n3399 = n3175 & n3257;
  assign n3400 = n3399 ^ n3177;
  assign n3401 = n3400 ^ n3397;
  assign n3402 = n3398 & ~n3401;
  assign n3403 = n3402 ^ x79;
  assign n3404 = n3403 ^ x80;
  assign n3405 = n3181 & n3257;
  assign n3406 = n3405 ^ n3183;
  assign n3407 = n3406 ^ n3403;
  assign n3408 = n3404 & ~n3407;
  assign n3409 = n3408 ^ x80;
  assign n3410 = n3409 ^ x81;
  assign n3411 = n3186 ^ x80;
  assign n3412 = n3257 & n3411;
  assign n3413 = n3412 ^ n3052;
  assign n3414 = n3413 ^ n3409;
  assign n3415 = n3410 & n3414;
  assign n3416 = n3415 ^ x81;
  assign n3417 = n3416 ^ x82;
  assign n3418 = ~n3187 & ~n3190;
  assign n3419 = n3418 ^ x81;
  assign n3420 = n3257 & n3419;
  assign n3421 = n3420 ^ n3049;
  assign n3422 = n3421 ^ n3416;
  assign n3423 = n3417 & n3422;
  assign n3424 = n3423 ^ x82;
  assign n3425 = n3424 ^ x83;
  assign n3426 = n3197 & n3257;
  assign n3427 = n3426 ^ n3199;
  assign n3428 = n3427 ^ n3424;
  assign n3429 = n3425 & n3428;
  assign n3430 = n3429 ^ x83;
  assign n3431 = n3430 ^ x84;
  assign n3432 = n3203 & n3257;
  assign n3433 = n3432 ^ n3205;
  assign n3434 = n3433 ^ n3430;
  assign n3435 = n3431 & ~n3434;
  assign n3436 = n3435 ^ x84;
  assign n3437 = n3436 ^ x85;
  assign n3438 = n3209 & n3257;
  assign n3439 = n3438 ^ n3211;
  assign n3440 = n3439 ^ n3436;
  assign n3441 = n3437 & ~n3440;
  assign n3442 = n3441 ^ x85;
  assign n3443 = n3442 ^ x86;
  assign n3444 = n3215 & n3257;
  assign n3445 = n3444 ^ n3217;
  assign n3446 = n3445 ^ n3442;
  assign n3447 = n3443 & ~n3446;
  assign n3448 = n3447 ^ x86;
  assign n3449 = n3282 & n3448;
  assign n3450 = n3280 ^ x88;
  assign n3451 = x87 & n3277;
  assign n3452 = n3451 ^ n3280;
  assign n3453 = n3450 & ~n3452;
  assign n3454 = n3453 ^ x88;
  assign n3455 = ~n3449 & ~n3454;
  assign n3456 = x89 & ~n3272;
  assign n3457 = n3455 & ~n3456;
  assign n3458 = n3457 ^ n3269;
  assign n3459 = n3458 ^ n3269;
  assign n3460 = ~n3275 & ~n3459;
  assign n3461 = n3460 ^ n3269;
  assign n3462 = n3270 & ~n3461;
  assign n3463 = n3462 ^ x90;
  assign n3464 = n3266 & n3463;
  assign n3465 = n3264 ^ x92;
  assign n3466 = x91 & ~n3261;
  assign n3467 = n3466 ^ x92;
  assign n3468 = n3465 & n3467;
  assign n3469 = n3468 ^ x92;
  assign n3470 = n163 & ~n3469;
  assign n3471 = ~n3464 & n3470;
  assign n3472 = n3455 ^ x89;
  assign n3473 = n3471 & ~n3472;
  assign n3474 = n3473 ^ n3272;
  assign n3475 = ~x90 & n3474;
  assign n3476 = ~n3273 & ~n3457;
  assign n3477 = n3476 ^ x90;
  assign n3478 = n3471 & n3477;
  assign n3479 = n3478 ^ n3269;
  assign n3480 = ~x91 & ~n3479;
  assign n3481 = ~n3475 & ~n3480;
  assign n3482 = n3374 & n3471;
  assign n3483 = n3482 ^ n3376;
  assign n3484 = ~x76 & ~n3483;
  assign n3485 = n3380 & n3471;
  assign n3486 = n3485 ^ n3382;
  assign n3487 = ~x77 & n3486;
  assign n3488 = ~n3484 & ~n3487;
  assign n3489 = ~x34 & ~x35;
  assign n3490 = ~n3471 & n3489;
  assign n3491 = ~x34 & x65;
  assign n3492 = ~n3490 & ~n3491;
  assign n3493 = x64 & ~n3492;
  assign n3494 = x64 & n3471;
  assign n3495 = x34 & ~x65;
  assign n3496 = x35 & ~n3495;
  assign n3497 = n3496 ^ n3293;
  assign n3498 = n3494 & n3497;
  assign n3499 = n3498 ^ n3293;
  assign n3500 = ~n3493 & ~n3499;
  assign n3501 = n3500 ^ x66;
  assign n3502 = n289 & ~n3257;
  assign n3503 = n3502 ^ x65;
  assign n3504 = ~x35 & n3503;
  assign n3505 = ~n202 & ~n3504;
  assign n3506 = x65 & n3257;
  assign n3507 = x35 & ~n3506;
  assign n3508 = x65 & n3507;
  assign n3509 = n3505 & ~n3508;
  assign n3510 = n3509 ^ n3296;
  assign n3511 = n3509 ^ n3507;
  assign n3512 = n3509 ^ n3471;
  assign n3513 = n3509 & n3512;
  assign n3514 = n3513 ^ n3509;
  assign n3515 = n3511 & n3514;
  assign n3516 = n3515 ^ n3513;
  assign n3517 = n3516 ^ n3509;
  assign n3518 = n3517 ^ n3471;
  assign n3519 = ~n3510 & n3518;
  assign n3520 = n3519 ^ n3296;
  assign n3521 = n3520 ^ x36;
  assign n3522 = n3521 ^ n3500;
  assign n3523 = ~n3501 & ~n3522;
  assign n3524 = n3523 ^ x66;
  assign n3525 = n3524 ^ x67;
  assign n3526 = ~n3309 & n3471;
  assign n3527 = n3526 ^ n3326;
  assign n3528 = n3527 ^ n3524;
  assign n3529 = n3525 & ~n3528;
  assign n3530 = n3529 ^ x67;
  assign n3531 = n3530 ^ x68;
  assign n3532 = n3330 & n3471;
  assign n3533 = n3532 ^ n3333;
  assign n3534 = n3533 ^ n3530;
  assign n3535 = n3531 & n3534;
  assign n3536 = n3535 ^ x68;
  assign n3537 = n3536 ^ x69;
  assign n3538 = n3336 ^ x68;
  assign n3539 = n3471 & n3538;
  assign n3540 = n3539 ^ n3284;
  assign n3541 = n3540 ^ n3536;
  assign n3542 = n3537 & ~n3541;
  assign n3543 = n3542 ^ x69;
  assign n3544 = n3543 ^ x70;
  assign n3545 = n3336 ^ n3284;
  assign n3546 = n3538 & ~n3545;
  assign n3547 = n3546 ^ x68;
  assign n3548 = n3547 ^ x69;
  assign n3549 = n3471 & n3548;
  assign n3550 = n3549 ^ n3287;
  assign n3551 = n3550 ^ n3543;
  assign n3552 = n3544 & ~n3551;
  assign n3553 = n3552 ^ x70;
  assign n3554 = n3553 ^ x71;
  assign n3555 = ~n3344 & n3471;
  assign n3556 = n3555 ^ n3346;
  assign n3557 = n3556 ^ n3553;
  assign n3558 = n3554 & ~n3557;
  assign n3559 = n3558 ^ x71;
  assign n3560 = n3559 ^ x72;
  assign n3561 = n3350 & n3471;
  assign n3562 = n3561 ^ n3352;
  assign n3563 = n3562 ^ n3559;
  assign n3564 = n3560 & ~n3563;
  assign n3565 = n3564 ^ x72;
  assign n3566 = n3565 ^ x73;
  assign n3567 = n3356 & n3471;
  assign n3568 = n3567 ^ n3358;
  assign n3569 = n3568 ^ n3565;
  assign n3570 = n3566 & ~n3569;
  assign n3571 = n3570 ^ x73;
  assign n3572 = n3571 ^ x74;
  assign n3573 = n3362 & n3471;
  assign n3574 = n3573 ^ n3364;
  assign n3575 = n3574 ^ n3571;
  assign n3576 = n3572 & ~n3575;
  assign n3577 = n3576 ^ x74;
  assign n3578 = n3577 ^ x75;
  assign n3579 = n3368 & n3471;
  assign n3580 = n3579 ^ n3370;
  assign n3581 = n3580 ^ n3577;
  assign n3582 = n3578 & ~n3581;
  assign n3583 = n3582 ^ x75;
  assign n3584 = n3488 & n3583;
  assign n3585 = n3486 ^ x77;
  assign n3586 = x76 & n3483;
  assign n3587 = n3586 ^ n3486;
  assign n3588 = ~n3585 & n3587;
  assign n3589 = n3588 ^ x77;
  assign n3590 = ~n3584 & ~n3589;
  assign n3591 = n3590 ^ x78;
  assign n3592 = n3386 & n3471;
  assign n3593 = n3592 ^ n3388;
  assign n3594 = n3593 ^ n3590;
  assign n3595 = ~n3591 & n3594;
  assign n3596 = n3595 ^ x78;
  assign n3597 = n3596 ^ x79;
  assign n3598 = n3392 & n3471;
  assign n3599 = n3598 ^ n3394;
  assign n3600 = n3599 ^ n3596;
  assign n3601 = n3597 & n3600;
  assign n3602 = n3601 ^ x79;
  assign n3603 = n3602 ^ x80;
  assign n3604 = n3398 & n3471;
  assign n3605 = n3604 ^ n3400;
  assign n3606 = n3605 ^ n3602;
  assign n3607 = n3603 & ~n3606;
  assign n3608 = n3607 ^ x80;
  assign n3609 = n3608 ^ x81;
  assign n3610 = n3404 & n3471;
  assign n3611 = n3610 ^ n3406;
  assign n3612 = n3611 ^ n3608;
  assign n3613 = n3609 & ~n3612;
  assign n3614 = n3613 ^ x81;
  assign n3615 = n3614 ^ x82;
  assign n3616 = n3410 & n3471;
  assign n3617 = n3616 ^ n3413;
  assign n3618 = n3617 ^ n3614;
  assign n3619 = n3615 & n3618;
  assign n3620 = n3619 ^ x82;
  assign n3621 = n3620 ^ x83;
  assign n3622 = n3417 & n3471;
  assign n3623 = n3622 ^ n3421;
  assign n3624 = n3623 ^ n3620;
  assign n3625 = n3621 & n3624;
  assign n3626 = n3625 ^ x83;
  assign n3627 = n3626 ^ x84;
  assign n3628 = n3425 & n3471;
  assign n3629 = n3628 ^ n3427;
  assign n3630 = n3629 ^ n3626;
  assign n3631 = n3627 & n3630;
  assign n3632 = n3631 ^ x84;
  assign n3633 = n3632 ^ x85;
  assign n3634 = n3431 & n3471;
  assign n3635 = n3634 ^ n3433;
  assign n3636 = n3635 ^ n3632;
  assign n3637 = n3633 & ~n3636;
  assign n3638 = n3637 ^ x85;
  assign n3639 = n3638 ^ x86;
  assign n3640 = n3437 & n3471;
  assign n3641 = n3640 ^ n3439;
  assign n3642 = n3641 ^ n3638;
  assign n3643 = n3639 & ~n3642;
  assign n3644 = n3643 ^ x86;
  assign n3645 = n3644 ^ x87;
  assign n3646 = n3443 & n3471;
  assign n3647 = n3646 ^ n3445;
  assign n3648 = n3647 ^ n3644;
  assign n3649 = n3645 & ~n3648;
  assign n3650 = n3649 ^ x87;
  assign n3651 = n3650 ^ x88;
  assign n3652 = n3448 ^ x87;
  assign n3653 = n3471 & n3652;
  assign n3654 = n3653 ^ n3277;
  assign n3655 = n3654 ^ n3650;
  assign n3656 = n3651 & ~n3655;
  assign n3657 = n3656 ^ x88;
  assign n3658 = n3657 ^ x89;
  assign n3659 = n3448 ^ n3277;
  assign n3660 = n3652 & ~n3659;
  assign n3661 = n3660 ^ x87;
  assign n3662 = n3661 ^ x88;
  assign n3663 = n3471 & n3662;
  assign n3664 = n3663 ^ n3280;
  assign n3665 = n3664 ^ n3657;
  assign n3666 = n3658 & ~n3665;
  assign n3667 = n3666 ^ x89;
  assign n3668 = n3481 & n3667;
  assign n3669 = n3479 ^ x91;
  assign n3670 = x90 & ~n3474;
  assign n3671 = n3670 ^ n3479;
  assign n3672 = n3669 & ~n3671;
  assign n3673 = n3672 ^ x91;
  assign n3674 = ~n3668 & ~n3673;
  assign n3675 = n3674 ^ x92;
  assign n3676 = n3463 ^ x91;
  assign n3677 = n3471 & n3676;
  assign n3678 = n3677 ^ n3261;
  assign n3679 = n3678 ^ n3674;
  assign n3680 = ~n3675 & ~n3679;
  assign n3681 = n3680 ^ x92;
  assign n3682 = n162 & ~n3681;
  assign n3683 = ~n3264 & ~n3471;
  assign n3684 = ~n240 & ~n3683;
  assign n3685 = ~n163 & ~n3684;
  assign n3686 = ~n3682 & n3685;
  assign n3687 = n3684 ^ x93;
  assign n3688 = n3681 ^ x93;
  assign n3689 = n3687 & n3688;
  assign n3690 = n3689 ^ x93;
  assign n3691 = n162 & ~n3690;
  assign n3692 = ~n3675 & n3691;
  assign n3693 = n3692 ^ n3678;
  assign n3694 = ~x93 & n3693;
  assign n3695 = ~x94 & n3686;
  assign n3696 = ~n3694 & ~n3695;
  assign n3697 = n3615 & n3691;
  assign n3698 = n3697 ^ n3617;
  assign n3699 = ~x83 & n3698;
  assign n3700 = n3621 & n3691;
  assign n3701 = n3700 ^ n3623;
  assign n3702 = ~x84 & n3701;
  assign n3703 = ~n3699 & ~n3702;
  assign n3704 = ~x65 & n3691;
  assign n3705 = ~x33 & x64;
  assign n3706 = ~n3495 & n3705;
  assign n3707 = ~n3704 & n3706;
  assign n3708 = x64 & n3691;
  assign n3709 = n3708 ^ x33;
  assign n3710 = n3708 ^ x34;
  assign n3711 = n3710 ^ n3708;
  assign n3712 = n3708 & ~n3711;
  assign n3713 = n3712 ^ n3708;
  assign n3714 = ~n3709 & n3713;
  assign n3715 = n3714 ^ n3712;
  assign n3716 = n3715 ^ n3708;
  assign n3717 = n3716 ^ n3710;
  assign n3718 = ~x65 & ~n3717;
  assign n3719 = n3718 ^ n3710;
  assign n3720 = ~n3707 & n3719;
  assign n3721 = n3720 ^ x66;
  assign n3722 = n289 & ~n3471;
  assign n3723 = n3722 ^ x65;
  assign n3724 = ~x34 & n3723;
  assign n3725 = ~n202 & ~n3724;
  assign n3726 = x65 & n3471;
  assign n3727 = x34 & ~n3726;
  assign n3728 = x65 & n3727;
  assign n3729 = n3725 & ~n3728;
  assign n3730 = n3729 ^ n3494;
  assign n3731 = n3729 ^ n3727;
  assign n3732 = n3729 ^ n3691;
  assign n3733 = n3729 & n3732;
  assign n3734 = n3733 ^ n3729;
  assign n3735 = n3731 & n3734;
  assign n3736 = n3735 ^ n3733;
  assign n3737 = n3736 ^ n3729;
  assign n3738 = n3737 ^ n3691;
  assign n3739 = ~n3730 & n3738;
  assign n3740 = n3739 ^ n3494;
  assign n3741 = n3740 ^ x35;
  assign n3742 = n3741 ^ n3720;
  assign n3743 = ~n3721 & ~n3742;
  assign n3744 = n3743 ^ x66;
  assign n3745 = n3744 ^ x67;
  assign n3746 = ~n3501 & n3691;
  assign n3747 = n3746 ^ n3521;
  assign n3748 = n3747 ^ n3744;
  assign n3749 = n3745 & n3748;
  assign n3750 = n3749 ^ x67;
  assign n3751 = n3750 ^ x68;
  assign n3752 = n3525 & n3691;
  assign n3753 = n3752 ^ n3527;
  assign n3754 = n3753 ^ n3750;
  assign n3755 = n3751 & ~n3754;
  assign n3756 = n3755 ^ x68;
  assign n3757 = n3756 ^ x69;
  assign n3758 = n3531 & n3691;
  assign n3759 = n3758 ^ n3533;
  assign n3760 = n3759 ^ n3756;
  assign n3761 = n3757 & n3760;
  assign n3762 = n3761 ^ x69;
  assign n3763 = n3762 ^ x70;
  assign n3764 = n3537 & n3691;
  assign n3765 = n3764 ^ n3540;
  assign n3766 = n3765 ^ n3762;
  assign n3767 = n3763 & ~n3766;
  assign n3768 = n3767 ^ x70;
  assign n3769 = n3768 ^ x71;
  assign n3770 = n3544 & n3691;
  assign n3771 = n3770 ^ n3550;
  assign n3772 = n3771 ^ n3768;
  assign n3773 = n3769 & ~n3772;
  assign n3774 = n3773 ^ x71;
  assign n3775 = n3774 ^ x72;
  assign n3776 = n3554 & n3691;
  assign n3777 = n3776 ^ n3556;
  assign n3778 = n3777 ^ n3774;
  assign n3779 = n3775 & ~n3778;
  assign n3780 = n3779 ^ x72;
  assign n3781 = n3780 ^ x73;
  assign n3782 = n3560 & n3691;
  assign n3783 = n3782 ^ n3562;
  assign n3784 = n3783 ^ n3780;
  assign n3785 = n3781 & ~n3784;
  assign n3786 = n3785 ^ x73;
  assign n3787 = n3786 ^ x74;
  assign n3788 = n3566 & n3691;
  assign n3789 = n3788 ^ n3568;
  assign n3790 = n3789 ^ n3786;
  assign n3791 = n3787 & ~n3790;
  assign n3792 = n3791 ^ x74;
  assign n3793 = n3792 ^ x75;
  assign n3794 = n3572 & n3691;
  assign n3795 = n3794 ^ n3574;
  assign n3796 = n3795 ^ n3792;
  assign n3797 = n3793 & ~n3796;
  assign n3798 = n3797 ^ x75;
  assign n3799 = n3798 ^ x76;
  assign n3800 = n3578 & n3691;
  assign n3801 = n3800 ^ n3580;
  assign n3802 = n3801 ^ n3798;
  assign n3803 = n3799 & ~n3802;
  assign n3804 = n3803 ^ x76;
  assign n3805 = n3804 ^ x77;
  assign n3806 = n3583 ^ x76;
  assign n3807 = n3691 & n3806;
  assign n3808 = n3807 ^ n3483;
  assign n3809 = n3808 ^ n3804;
  assign n3810 = n3805 & ~n3809;
  assign n3811 = n3810 ^ x77;
  assign n3812 = n3811 ^ x78;
  assign n3813 = n3583 ^ n3483;
  assign n3814 = n3806 & ~n3813;
  assign n3815 = n3814 ^ x76;
  assign n3816 = n3815 ^ x77;
  assign n3817 = n3691 & n3816;
  assign n3818 = n3817 ^ n3486;
  assign n3819 = n3818 ^ n3811;
  assign n3820 = n3812 & n3819;
  assign n3821 = n3820 ^ x78;
  assign n3822 = n3821 ^ x79;
  assign n3823 = ~n3591 & n3691;
  assign n3824 = n3823 ^ n3593;
  assign n3825 = n3824 ^ n3821;
  assign n3826 = n3822 & ~n3825;
  assign n3827 = n3826 ^ x79;
  assign n3828 = n3827 ^ x80;
  assign n3829 = n3597 & n3691;
  assign n3830 = n3829 ^ n3599;
  assign n3831 = n3830 ^ n3827;
  assign n3832 = n3828 & n3831;
  assign n3833 = n3832 ^ x80;
  assign n3834 = n3833 ^ x81;
  assign n3835 = n3603 & n3691;
  assign n3836 = n3835 ^ n3605;
  assign n3837 = n3836 ^ n3833;
  assign n3838 = n3834 & ~n3837;
  assign n3839 = n3838 ^ x81;
  assign n3840 = n3839 ^ x82;
  assign n3841 = n3609 & n3691;
  assign n3842 = n3841 ^ n3611;
  assign n3843 = n3842 ^ n3839;
  assign n3844 = n3840 & ~n3843;
  assign n3845 = n3844 ^ x82;
  assign n3846 = n3703 & n3845;
  assign n3847 = n3701 ^ x84;
  assign n3848 = x83 & ~n3698;
  assign n3849 = n3848 ^ n3701;
  assign n3850 = ~n3847 & n3849;
  assign n3851 = n3850 ^ x84;
  assign n3852 = ~n3846 & ~n3851;
  assign n3853 = n3852 ^ x85;
  assign n3854 = n3627 & n3691;
  assign n3855 = n3854 ^ n3629;
  assign n3856 = n3855 ^ n3852;
  assign n3857 = ~n3853 & ~n3856;
  assign n3858 = n3857 ^ x85;
  assign n3859 = n3858 ^ x86;
  assign n3860 = n3633 & n3691;
  assign n3861 = n3860 ^ n3635;
  assign n3862 = n3861 ^ n3858;
  assign n3863 = n3859 & ~n3862;
  assign n3864 = n3863 ^ x86;
  assign n3865 = n3864 ^ x87;
  assign n3866 = n3639 & n3691;
  assign n3867 = n3866 ^ n3641;
  assign n3868 = n3867 ^ n3864;
  assign n3869 = n3865 & ~n3868;
  assign n3870 = n3869 ^ x87;
  assign n3871 = n3870 ^ x88;
  assign n3872 = n3645 & n3691;
  assign n3873 = n3872 ^ n3647;
  assign n3874 = n3873 ^ n3870;
  assign n3875 = n3871 & ~n3874;
  assign n3876 = n3875 ^ x88;
  assign n3877 = n3876 ^ x89;
  assign n3878 = n3651 & n3691;
  assign n3879 = n3878 ^ n3654;
  assign n3880 = n3879 ^ n3876;
  assign n3881 = n3877 & ~n3880;
  assign n3882 = n3881 ^ x89;
  assign n3883 = n3882 ^ x90;
  assign n3884 = n3658 & n3691;
  assign n3885 = n3884 ^ n3664;
  assign n3886 = n3885 ^ n3882;
  assign n3887 = n3883 & ~n3886;
  assign n3888 = n3887 ^ x90;
  assign n3889 = n3888 ^ x91;
  assign n3890 = n3667 ^ x90;
  assign n3891 = n3691 & n3890;
  assign n3892 = n3891 ^ n3474;
  assign n3893 = n3892 ^ n3888;
  assign n3894 = n3889 & n3893;
  assign n3895 = n3894 ^ x91;
  assign n3896 = n3895 ^ x92;
  assign n3897 = n3667 ^ n3474;
  assign n3898 = n3890 & n3897;
  assign n3899 = n3898 ^ x90;
  assign n3900 = n3899 ^ x91;
  assign n3901 = n3691 & n3900;
  assign n3902 = n3901 ^ n3479;
  assign n3903 = n3902 ^ n3895;
  assign n3904 = n3896 & ~n3903;
  assign n3905 = n3904 ^ x92;
  assign n3906 = n3696 & n3905;
  assign n3907 = x93 & ~n3695;
  assign n3908 = ~n3693 & n3907;
  assign n3909 = n161 & ~n3684;
  assign n3910 = ~n162 & ~n3909;
  assign n3911 = ~n3908 & ~n3910;
  assign n3912 = ~n3906 & n3911;
  assign n3913 = n3686 & ~n3912;
  assign n3914 = ~n240 & ~n3913;
  assign n3915 = n161 & ~n3914;
  assign n3916 = x95 & n3914;
  assign n3917 = n160 & ~n3916;
  assign n3918 = n3845 ^ x83;
  assign n3919 = n3845 ^ n3698;
  assign n3920 = n3918 & n3919;
  assign n3921 = n3920 ^ x83;
  assign n3922 = n3921 ^ x84;
  assign n3923 = n3912 & n3922;
  assign n3924 = n3923 ^ n3701;
  assign n3925 = ~x85 & n3924;
  assign n3926 = ~n3853 & n3912;
  assign n3927 = n3926 ^ n3855;
  assign n3928 = ~x86 & n3927;
  assign n3929 = ~n3925 & ~n3928;
  assign n3930 = n3691 ^ x65;
  assign n3931 = n3705 & ~n3930;
  assign n3932 = ~n202 & ~n3931;
  assign n3933 = x65 & n3691;
  assign n3934 = x33 & ~n3933;
  assign n3935 = x65 & n3934;
  assign n3936 = n3932 & ~n3935;
  assign n3937 = n3936 ^ n3708;
  assign n3938 = n3936 ^ n3934;
  assign n3939 = n3936 ^ n3912;
  assign n3940 = n3936 & n3939;
  assign n3941 = n3940 ^ n3936;
  assign n3942 = n3938 & n3941;
  assign n3943 = n3942 ^ n3940;
  assign n3944 = n3943 ^ n3936;
  assign n3945 = n3944 ^ n3912;
  assign n3946 = ~n3937 & n3945;
  assign n3947 = n3946 ^ n3708;
  assign n3948 = n3947 ^ x34;
  assign n3949 = n3948 ^ x66;
  assign n3950 = x64 & n3912;
  assign n3951 = x33 & ~x65;
  assign n3952 = x32 & n3951;
  assign n3953 = n3952 ^ x33;
  assign n3954 = n3950 & n3953;
  assign n3955 = ~x32 & n288;
  assign n3956 = n3955 ^ x65;
  assign n3957 = ~x33 & n3956;
  assign n3958 = ~n3912 & n3957;
  assign n3959 = x33 ^ x32;
  assign n3960 = x64 ^ x33;
  assign n3961 = n3960 ^ x33;
  assign n3962 = n3959 & n3961;
  assign n3963 = n3962 ^ x33;
  assign n3964 = x65 & ~n3963;
  assign n3965 = ~n3958 & ~n3964;
  assign n3966 = ~n3954 & n3965;
  assign n3967 = n3966 ^ n3948;
  assign n3968 = ~n3949 & ~n3967;
  assign n3969 = n3968 ^ x66;
  assign n3970 = n3969 ^ x67;
  assign n3971 = ~n3721 & n3912;
  assign n3972 = n3971 ^ n3741;
  assign n3973 = n3972 ^ n3969;
  assign n3974 = n3970 & n3973;
  assign n3975 = n3974 ^ x67;
  assign n3976 = n3975 ^ x68;
  assign n3977 = n3745 & n3912;
  assign n3978 = n3977 ^ n3747;
  assign n3979 = n3978 ^ n3975;
  assign n3980 = n3976 & n3979;
  assign n3981 = n3980 ^ x68;
  assign n3982 = n3981 ^ x69;
  assign n3983 = n3751 & n3912;
  assign n3984 = n3983 ^ n3753;
  assign n3985 = n3984 ^ n3981;
  assign n3986 = n3982 & ~n3985;
  assign n3987 = n3986 ^ x69;
  assign n3988 = n3987 ^ x70;
  assign n3989 = n3757 & n3912;
  assign n3990 = n3989 ^ n3759;
  assign n3991 = n3990 ^ n3987;
  assign n3992 = n3988 & n3991;
  assign n3993 = n3992 ^ x70;
  assign n3994 = n3993 ^ x71;
  assign n3995 = n3763 & n3912;
  assign n3996 = n3995 ^ n3765;
  assign n3997 = n3996 ^ n3993;
  assign n3998 = n3994 & ~n3997;
  assign n3999 = n3998 ^ x71;
  assign n4000 = n3999 ^ x72;
  assign n4001 = n3771 ^ x71;
  assign n4002 = n4001 ^ n3768;
  assign n4003 = n4002 ^ n3771;
  assign n4004 = n3912 & n4003;
  assign n4005 = n4004 ^ n3771;
  assign n4006 = n4005 ^ n3999;
  assign n4007 = n4000 & ~n4006;
  assign n4008 = n4007 ^ x72;
  assign n4009 = n4008 ^ x73;
  assign n4010 = n3775 & n3912;
  assign n4011 = n4010 ^ n3777;
  assign n4012 = n4011 ^ n4008;
  assign n4013 = n4009 & ~n4012;
  assign n4014 = n4013 ^ x73;
  assign n4015 = n4014 ^ x74;
  assign n4016 = n3781 & n3912;
  assign n4017 = n4016 ^ n3783;
  assign n4018 = n4017 ^ n4014;
  assign n4019 = n4015 & ~n4018;
  assign n4020 = n4019 ^ x74;
  assign n4021 = n4020 ^ x75;
  assign n4022 = n3787 & n3912;
  assign n4023 = n4022 ^ n3789;
  assign n4024 = n4023 ^ n4020;
  assign n4025 = n4021 & ~n4024;
  assign n4026 = n4025 ^ x75;
  assign n4027 = n4026 ^ x76;
  assign n4028 = n3793 & n3912;
  assign n4029 = n4028 ^ n3795;
  assign n4030 = n4029 ^ n4026;
  assign n4031 = n4027 & ~n4030;
  assign n4032 = n4031 ^ x76;
  assign n4033 = n4032 ^ x77;
  assign n4034 = n3799 & n3912;
  assign n4035 = n4034 ^ n3801;
  assign n4036 = n4035 ^ n4032;
  assign n4037 = n4033 & ~n4036;
  assign n4038 = n4037 ^ x77;
  assign n4039 = n4038 ^ x78;
  assign n4040 = n3805 & n3912;
  assign n4041 = n4040 ^ n3808;
  assign n4042 = n4041 ^ n4038;
  assign n4043 = n4039 & ~n4042;
  assign n4044 = n4043 ^ x78;
  assign n4045 = n4044 ^ x79;
  assign n4046 = n3812 & n3912;
  assign n4047 = n4046 ^ n3818;
  assign n4048 = n4047 ^ n4044;
  assign n4049 = n4045 & n4048;
  assign n4050 = n4049 ^ x79;
  assign n4051 = n4050 ^ x80;
  assign n4052 = n3822 & n3912;
  assign n4053 = n4052 ^ n3824;
  assign n4054 = n4053 ^ n4050;
  assign n4055 = n4051 & ~n4054;
  assign n4056 = n4055 ^ x80;
  assign n4057 = n4056 ^ x81;
  assign n4058 = n3828 & n3912;
  assign n4059 = n4058 ^ n3830;
  assign n4060 = n4059 ^ n4056;
  assign n4061 = n4057 & n4060;
  assign n4062 = n4061 ^ x81;
  assign n4063 = n4062 ^ x82;
  assign n4064 = n3834 & n3912;
  assign n4065 = n4064 ^ n3836;
  assign n4066 = n4065 ^ n4062;
  assign n4067 = n4063 & ~n4066;
  assign n4068 = n4067 ^ x82;
  assign n4069 = n4068 ^ x83;
  assign n4070 = n3840 & n3912;
  assign n4071 = n4070 ^ n3842;
  assign n4072 = n4071 ^ n4068;
  assign n4073 = n4069 & ~n4072;
  assign n4074 = n4073 ^ x83;
  assign n4075 = n4074 ^ x84;
  assign n4076 = n3912 & n3918;
  assign n4077 = n4076 ^ n3698;
  assign n4078 = n4077 ^ n4074;
  assign n4079 = n4075 & n4078;
  assign n4080 = n4079 ^ x84;
  assign n4081 = n3929 & n4080;
  assign n4082 = n3927 ^ x86;
  assign n4083 = x85 & ~n3924;
  assign n4084 = n4083 ^ n3927;
  assign n4085 = ~n4082 & n4084;
  assign n4086 = n4085 ^ x86;
  assign n4087 = ~n4081 & ~n4086;
  assign n4088 = n4087 ^ x87;
  assign n4089 = n3859 & n3912;
  assign n4090 = n4089 ^ n3861;
  assign n4091 = n4090 ^ n4087;
  assign n4092 = ~n4088 & n4091;
  assign n4093 = n4092 ^ x87;
  assign n4094 = n4093 ^ x88;
  assign n4095 = n3865 & n3912;
  assign n4096 = n4095 ^ n3867;
  assign n4097 = n4096 ^ n4093;
  assign n4098 = n4094 & ~n4097;
  assign n4099 = n4098 ^ x88;
  assign n4100 = n4099 ^ x89;
  assign n4101 = n3871 & n3912;
  assign n4102 = n4101 ^ n3873;
  assign n4103 = n4102 ^ n4099;
  assign n4104 = n4100 & ~n4103;
  assign n4105 = n4104 ^ x89;
  assign n4106 = n4105 ^ x90;
  assign n4107 = n3877 & n3912;
  assign n4108 = n4107 ^ n3879;
  assign n4109 = n4108 ^ n4105;
  assign n4110 = n4106 & ~n4109;
  assign n4111 = n4110 ^ x90;
  assign n4112 = n4111 ^ x91;
  assign n4113 = n3883 & n3912;
  assign n4114 = n4113 ^ n3885;
  assign n4115 = n4114 ^ n4111;
  assign n4116 = n4112 & ~n4115;
  assign n4117 = n4116 ^ x91;
  assign n4118 = n4117 ^ x92;
  assign n4119 = n3889 & n3912;
  assign n4120 = n4119 ^ n3892;
  assign n4121 = n4120 ^ n4117;
  assign n4122 = n4118 & n4121;
  assign n4123 = n4122 ^ x92;
  assign n4124 = n4123 ^ x93;
  assign n4125 = n3896 & n3912;
  assign n4126 = n4125 ^ n3902;
  assign n4127 = n4126 ^ n4123;
  assign n4128 = n4124 & ~n4127;
  assign n4129 = n4128 ^ x93;
  assign n4130 = n4129 ^ x94;
  assign n4131 = n3905 ^ x93;
  assign n4132 = n3912 & n4131;
  assign n4133 = n4132 ^ n3693;
  assign n4134 = n4133 ^ n4129;
  assign n4135 = n4130 & ~n4134;
  assign n4136 = n4135 ^ n4129;
  assign n4137 = n3917 & ~n4136;
  assign n4138 = ~n3915 & ~n4137;
  assign n4375 = x64 & ~n4138;
  assign n4171 = ~x31 & x64;
  assign n4368 = n4138 ^ x65;
  assign n4369 = n4171 & n4368;
  assign n4370 = ~n202 & ~n4369;
  assign n4371 = x65 & ~n4138;
  assign n4372 = x31 & ~n4371;
  assign n4373 = x65 & n4372;
  assign n4374 = n4370 & ~n4373;
  assign n4376 = n4375 ^ n4374;
  assign n4377 = n4374 ^ n4372;
  assign n4145 = n4039 & ~n4138;
  assign n4146 = n4145 ^ n4041;
  assign n4147 = ~x79 & ~n4146;
  assign n4148 = n4045 & ~n4138;
  assign n4149 = n4148 ^ n4047;
  assign n4150 = ~x80 & n4149;
  assign n4151 = ~n4147 & ~n4150;
  assign n4152 = n4138 ^ n288;
  assign n4153 = n4152 ^ n288;
  assign n4154 = n2322 & ~n4153;
  assign n4155 = n4154 ^ n288;
  assign n4156 = ~n3912 & n4155;
  assign n4157 = n4156 ^ n288;
  assign n4158 = x32 & n4157;
  assign n4159 = ~n288 & ~n3912;
  assign n4160 = ~x32 & ~n4159;
  assign n4161 = ~n202 & ~n4160;
  assign n4162 = ~x65 & n3912;
  assign n4163 = ~n4161 & ~n4162;
  assign n4164 = n4163 ^ n3950;
  assign n4165 = ~n4138 & n4164;
  assign n4166 = n4165 ^ n3950;
  assign n4167 = ~n4158 & ~n4166;
  assign n4168 = n4167 ^ x33;
  assign n4169 = n4168 ^ x66;
  assign n4170 = ~x65 & n4138;
  assign n4172 = n4170 & ~n4171;
  assign n4173 = x32 & x64;
  assign n4174 = x31 & ~x65;
  assign n4175 = n4173 & ~n4174;
  assign n4176 = n4175 ^ x32;
  assign n4177 = ~n4138 & ~n4176;
  assign n4178 = n4177 ^ x32;
  assign n4179 = ~n4172 & ~n4178;
  assign n4180 = x32 ^ x31;
  assign n4181 = ~x64 & n4180;
  assign n4182 = n4181 ^ x31;
  assign n4183 = x65 & ~n4182;
  assign n4184 = ~n4179 & ~n4183;
  assign n4185 = n4184 ^ n4168;
  assign n4186 = n4169 & n4185;
  assign n4187 = n4186 ^ x66;
  assign n4188 = n4187 ^ x67;
  assign n4189 = n3966 ^ x66;
  assign n4190 = ~n4138 & ~n4189;
  assign n4191 = n4190 ^ n3948;
  assign n4192 = n4191 ^ n4187;
  assign n4193 = n4188 & n4192;
  assign n4194 = n4193 ^ x67;
  assign n4195 = n4194 ^ x68;
  assign n4196 = n3970 & ~n4138;
  assign n4197 = n4196 ^ n3972;
  assign n4198 = n4197 ^ n4194;
  assign n4199 = n4195 & n4198;
  assign n4200 = n4199 ^ x68;
  assign n4201 = n4200 ^ x69;
  assign n4202 = n3976 & ~n4138;
  assign n4203 = n4202 ^ n3978;
  assign n4204 = n4203 ^ n4200;
  assign n4205 = n4201 & n4204;
  assign n4206 = n4205 ^ x69;
  assign n4207 = n4206 ^ x70;
  assign n4208 = n3982 & ~n4138;
  assign n4209 = n4208 ^ n3984;
  assign n4210 = n4209 ^ n4206;
  assign n4211 = n4207 & ~n4210;
  assign n4212 = n4211 ^ x70;
  assign n4213 = n4212 ^ x71;
  assign n4214 = n3988 & ~n4138;
  assign n4215 = n4214 ^ n3990;
  assign n4216 = n4215 ^ n4212;
  assign n4217 = n4213 & n4216;
  assign n4218 = n4217 ^ x71;
  assign n4219 = n4218 ^ x72;
  assign n4220 = n3994 & ~n4138;
  assign n4221 = n4220 ^ n3996;
  assign n4222 = n4221 ^ n4218;
  assign n4223 = n4219 & ~n4222;
  assign n4224 = n4223 ^ x72;
  assign n4225 = n4224 ^ x73;
  assign n4226 = n4000 & ~n4138;
  assign n4227 = n4226 ^ n4005;
  assign n4228 = n4227 ^ n4224;
  assign n4229 = n4225 & ~n4228;
  assign n4230 = n4229 ^ x73;
  assign n4231 = n4230 ^ x74;
  assign n4232 = n4009 & ~n4138;
  assign n4233 = n4232 ^ n4011;
  assign n4234 = n4233 ^ n4230;
  assign n4235 = n4231 & ~n4234;
  assign n4236 = n4235 ^ x74;
  assign n4237 = n4236 ^ x75;
  assign n4238 = n4015 & ~n4138;
  assign n4239 = n4238 ^ n4017;
  assign n4240 = n4239 ^ n4236;
  assign n4241 = n4237 & ~n4240;
  assign n4242 = n4241 ^ x75;
  assign n4243 = n4242 ^ x76;
  assign n4244 = n4021 & ~n4138;
  assign n4245 = n4244 ^ n4023;
  assign n4246 = n4245 ^ n4242;
  assign n4247 = n4243 & ~n4246;
  assign n4248 = n4247 ^ x76;
  assign n4249 = n4248 ^ x77;
  assign n4250 = n4027 & ~n4138;
  assign n4251 = n4250 ^ n4029;
  assign n4252 = n4251 ^ n4248;
  assign n4253 = n4249 & ~n4252;
  assign n4254 = n4253 ^ x77;
  assign n4255 = n4254 ^ x78;
  assign n4256 = n4033 & ~n4138;
  assign n4257 = n4256 ^ n4035;
  assign n4258 = n4257 ^ n4254;
  assign n4259 = n4255 & ~n4258;
  assign n4260 = n4259 ^ x78;
  assign n4261 = n4151 & n4260;
  assign n4262 = n4149 ^ x80;
  assign n4263 = x79 & n4146;
  assign n4264 = n4263 ^ n4149;
  assign n4265 = ~n4262 & n4264;
  assign n4266 = n4265 ^ x80;
  assign n4267 = ~n4261 & ~n4266;
  assign n4268 = n4267 ^ x81;
  assign n4269 = n4051 & ~n4138;
  assign n4270 = n4269 ^ n4053;
  assign n4271 = n4270 ^ n4267;
  assign n4272 = ~n4268 & n4271;
  assign n4273 = n4272 ^ x81;
  assign n4274 = n4273 ^ x82;
  assign n4275 = n4057 & ~n4138;
  assign n4276 = n4275 ^ n4059;
  assign n4277 = n4276 ^ n4273;
  assign n4278 = n4274 & n4277;
  assign n4279 = n4278 ^ x82;
  assign n4280 = n4279 ^ x83;
  assign n4281 = n4063 & ~n4138;
  assign n4282 = n4281 ^ n4065;
  assign n4283 = n4282 ^ n4279;
  assign n4284 = n4280 & ~n4283;
  assign n4285 = n4284 ^ x83;
  assign n4286 = n4285 ^ x84;
  assign n4287 = n4069 & ~n4138;
  assign n4288 = n4287 ^ n4071;
  assign n4289 = n4288 ^ n4285;
  assign n4290 = n4286 & ~n4289;
  assign n4291 = n4290 ^ x84;
  assign n4292 = n4291 ^ x85;
  assign n4293 = n4075 & ~n4138;
  assign n4294 = n4293 ^ n4077;
  assign n4295 = n4294 ^ n4291;
  assign n4296 = n4292 & n4295;
  assign n4297 = n4296 ^ x85;
  assign n4298 = n4297 ^ x86;
  assign n4299 = n4080 ^ x85;
  assign n4300 = ~n4138 & n4299;
  assign n4301 = n4300 ^ n3924;
  assign n4302 = n4301 ^ n4297;
  assign n4303 = n4298 & n4302;
  assign n4304 = n4303 ^ x86;
  assign n4305 = n4304 ^ x87;
  assign n4306 = n4080 ^ n3924;
  assign n4307 = n4299 & n4306;
  assign n4308 = n4307 ^ x85;
  assign n4309 = n4308 ^ x86;
  assign n4310 = ~n4138 & n4309;
  assign n4311 = n4310 ^ n3927;
  assign n4312 = n4311 ^ n4304;
  assign n4313 = n4305 & n4312;
  assign n4314 = n4313 ^ x87;
  assign n4315 = n4314 ^ x88;
  assign n4316 = ~n4088 & ~n4138;
  assign n4317 = n4316 ^ n4090;
  assign n4318 = n4317 ^ n4314;
  assign n4319 = n4315 & ~n4318;
  assign n4320 = n4319 ^ x88;
  assign n4321 = n4320 ^ x89;
  assign n4322 = n4094 & ~n4138;
  assign n4323 = n4322 ^ n4096;
  assign n4324 = n4323 ^ n4320;
  assign n4325 = n4321 & ~n4324;
  assign n4326 = n4325 ^ x89;
  assign n4327 = n4326 ^ x90;
  assign n4328 = n4100 & ~n4138;
  assign n4329 = n4328 ^ n4102;
  assign n4330 = n4329 ^ n4326;
  assign n4331 = n4327 & ~n4330;
  assign n4332 = n4331 ^ x90;
  assign n4333 = n4332 ^ x91;
  assign n4334 = n4106 & ~n4138;
  assign n4335 = n4334 ^ n4108;
  assign n4336 = n4335 ^ n4332;
  assign n4337 = n4333 & ~n4336;
  assign n4338 = n4337 ^ x91;
  assign n4339 = n4338 ^ x92;
  assign n4340 = n4112 & ~n4138;
  assign n4341 = n4340 ^ n4114;
  assign n4342 = n4341 ^ n4338;
  assign n4343 = n4339 & ~n4342;
  assign n4344 = n4343 ^ x92;
  assign n4345 = n4344 ^ x93;
  assign n4346 = n4118 & ~n4138;
  assign n4347 = n4346 ^ n4120;
  assign n4348 = n4347 ^ n4344;
  assign n4349 = n4345 & n4348;
  assign n4350 = n4349 ^ x93;
  assign n4351 = n4350 ^ x94;
  assign n4352 = n4124 & ~n4138;
  assign n4353 = n4352 ^ n4126;
  assign n4354 = n4353 ^ n4350;
  assign n4355 = n4351 & ~n4354;
  assign n4356 = n4355 ^ x94;
  assign n4141 = n4130 & ~n4138;
  assign n4142 = n4141 ^ n4133;
  assign n4143 = ~x95 & n4142;
  assign n4139 = ~n3914 & n4138;
  assign n4140 = ~n240 & ~n4139;
  assign n4378 = ~x96 & ~n4140;
  assign n4379 = ~n4143 & ~n4378;
  assign n4380 = n4356 & n4379;
  assign n4381 = x95 & ~n4378;
  assign n4382 = ~n4142 & n4381;
  assign n241 = n155 & n157;
  assign n4358 = n156 & n241;
  assign n4383 = x96 & n4140;
  assign n4384 = n4358 & ~n4383;
  assign n4385 = ~n4382 & n4384;
  assign n4386 = ~n4380 & n4385;
  assign n4387 = n4386 ^ n4374;
  assign n4388 = n4374 & n4387;
  assign n4389 = n4388 ^ n4374;
  assign n4390 = n4377 & n4389;
  assign n4391 = n4390 ^ n4388;
  assign n4392 = n4391 ^ n4374;
  assign n4393 = n4392 ^ n4386;
  assign n4394 = ~n4376 & n4393;
  assign n4395 = n4394 ^ n4375;
  assign n4396 = n4395 ^ x32;
  assign n4397 = n4396 ^ x66;
  assign n4398 = x64 & n4386;
  assign n4399 = x30 & n4174;
  assign n4400 = n4399 ^ x31;
  assign n4401 = n4398 & n4400;
  assign n4402 = ~x30 & n4171;
  assign n4403 = ~x31 & x65;
  assign n4404 = ~n4402 & ~n4403;
  assign n4405 = ~n4386 & ~n4404;
  assign n4406 = ~x30 & x65;
  assign n4407 = n4406 ^ n4403;
  assign n4408 = x64 & n4407;
  assign n4409 = n4408 ^ n4403;
  assign n4410 = ~n4405 & ~n4409;
  assign n4411 = ~n4401 & n4410;
  assign n4412 = n4411 ^ n4396;
  assign n4413 = ~n4397 & ~n4412;
  assign n4414 = n4413 ^ x66;
  assign n4415 = n4414 ^ x67;
  assign n4416 = n4184 ^ x66;
  assign n4417 = n4386 & ~n4416;
  assign n4418 = n4417 ^ n4168;
  assign n4419 = n4418 ^ n4414;
  assign n4420 = n4415 & ~n4419;
  assign n4421 = n4420 ^ x67;
  assign n4422 = n4421 ^ x68;
  assign n4144 = x96 & ~n4143;
  assign n4357 = n4144 & n4356;
  assign n4359 = x95 & x96;
  assign n4360 = ~n4142 & n4359;
  assign n4361 = n4358 & ~n4360;
  assign n4362 = ~n4357 & n4361;
  assign n4363 = ~n4140 & ~n4362;
  assign n4364 = ~n240 & ~n4363;
  assign n4367 = ~x97 & ~n4364;
  assign n4423 = n4188 & n4386;
  assign n4424 = n4423 ^ n4191;
  assign n4425 = n4424 ^ n4421;
  assign n4426 = n4422 & n4425;
  assign n4427 = n4426 ^ x68;
  assign n4428 = n4427 ^ x69;
  assign n4429 = n4195 & n4386;
  assign n4430 = n4429 ^ n4197;
  assign n4431 = n4430 ^ n4427;
  assign n4432 = n4428 & n4431;
  assign n4433 = n4432 ^ x69;
  assign n4434 = n4433 ^ x70;
  assign n4435 = n4201 & n4386;
  assign n4436 = n4435 ^ n4203;
  assign n4437 = n4436 ^ n4433;
  assign n4438 = n4434 & n4437;
  assign n4439 = n4438 ^ x70;
  assign n4440 = n4439 ^ x71;
  assign n4441 = n4207 & n4386;
  assign n4442 = n4441 ^ n4209;
  assign n4443 = n4442 ^ n4439;
  assign n4444 = n4440 & ~n4443;
  assign n4445 = n4444 ^ x71;
  assign n4446 = n4445 ^ x72;
  assign n4447 = n4213 & n4386;
  assign n4448 = n4447 ^ n4215;
  assign n4449 = n4448 ^ n4445;
  assign n4450 = n4446 & n4449;
  assign n4451 = n4450 ^ x72;
  assign n4452 = n4451 ^ x73;
  assign n4453 = n4219 & n4386;
  assign n4454 = n4453 ^ n4221;
  assign n4455 = n4454 ^ n4451;
  assign n4456 = n4452 & ~n4455;
  assign n4457 = n4456 ^ x73;
  assign n4458 = n4457 ^ x74;
  assign n4459 = n4225 & n4386;
  assign n4460 = n4459 ^ n4227;
  assign n4461 = n4460 ^ n4457;
  assign n4462 = n4458 & ~n4461;
  assign n4463 = n4462 ^ x74;
  assign n4464 = n4463 ^ x75;
  assign n4465 = n4231 & n4386;
  assign n4466 = n4465 ^ n4233;
  assign n4467 = n4466 ^ n4463;
  assign n4468 = n4464 & ~n4467;
  assign n4469 = n4468 ^ x75;
  assign n4470 = n4469 ^ x76;
  assign n4471 = n4237 & n4386;
  assign n4472 = n4471 ^ n4239;
  assign n4473 = n4472 ^ n4469;
  assign n4474 = n4470 & ~n4473;
  assign n4475 = n4474 ^ x76;
  assign n4476 = n4475 ^ x77;
  assign n4477 = n4243 & n4386;
  assign n4478 = n4477 ^ n4245;
  assign n4479 = n4478 ^ n4475;
  assign n4480 = n4476 & ~n4479;
  assign n4481 = n4480 ^ x77;
  assign n4482 = n4481 ^ x78;
  assign n4483 = n4249 & n4386;
  assign n4484 = n4483 ^ n4251;
  assign n4485 = n4484 ^ n4481;
  assign n4486 = n4482 & ~n4485;
  assign n4487 = n4486 ^ x78;
  assign n4488 = n4487 ^ x79;
  assign n4489 = n4255 & n4386;
  assign n4490 = n4489 ^ n4257;
  assign n4491 = n4490 ^ n4487;
  assign n4492 = n4488 & ~n4491;
  assign n4493 = n4492 ^ x79;
  assign n4494 = n4493 ^ x80;
  assign n4495 = n4260 ^ x79;
  assign n4496 = n4386 & n4495;
  assign n4497 = n4496 ^ n4146;
  assign n4498 = n4497 ^ n4493;
  assign n4499 = n4494 & ~n4498;
  assign n4500 = n4499 ^ x80;
  assign n4501 = n4500 ^ x81;
  assign n4502 = n4260 ^ n4146;
  assign n4503 = n4495 & ~n4502;
  assign n4504 = n4503 ^ x79;
  assign n4505 = n4504 ^ x80;
  assign n4506 = n4386 & n4505;
  assign n4507 = n4506 ^ n4149;
  assign n4508 = n4507 ^ n4500;
  assign n4509 = n4501 & n4508;
  assign n4510 = n4509 ^ x81;
  assign n4511 = n4510 ^ x82;
  assign n4512 = ~n4268 & n4386;
  assign n4513 = n4512 ^ n4270;
  assign n4514 = n4513 ^ n4510;
  assign n4515 = n4511 & ~n4514;
  assign n4516 = n4515 ^ x82;
  assign n4517 = n4516 ^ x83;
  assign n4518 = n4274 & n4386;
  assign n4519 = n4518 ^ n4276;
  assign n4520 = n4519 ^ n4516;
  assign n4521 = n4517 & n4520;
  assign n4522 = n4521 ^ x83;
  assign n4523 = n4522 ^ x84;
  assign n4524 = n4280 & n4386;
  assign n4525 = n4524 ^ n4282;
  assign n4526 = n4525 ^ n4522;
  assign n4527 = n4523 & ~n4526;
  assign n4528 = n4527 ^ x84;
  assign n4529 = n4528 ^ x85;
  assign n4530 = n4286 & n4386;
  assign n4531 = n4530 ^ n4288;
  assign n4532 = n4531 ^ n4528;
  assign n4533 = n4529 & ~n4532;
  assign n4534 = n4533 ^ x85;
  assign n4535 = n4534 ^ x86;
  assign n4536 = n4292 & n4386;
  assign n4537 = n4536 ^ n4294;
  assign n4538 = n4537 ^ n4534;
  assign n4539 = n4535 & n4538;
  assign n4540 = n4539 ^ x86;
  assign n4541 = n4540 ^ x87;
  assign n4542 = n4298 & n4386;
  assign n4543 = n4542 ^ n4301;
  assign n4544 = n4543 ^ n4540;
  assign n4545 = n4541 & n4544;
  assign n4546 = n4545 ^ x87;
  assign n4547 = n4546 ^ x88;
  assign n4548 = n4305 & n4386;
  assign n4549 = n4548 ^ n4311;
  assign n4550 = n4549 ^ n4546;
  assign n4551 = n4547 & n4550;
  assign n4552 = n4551 ^ x88;
  assign n4553 = n4552 ^ x89;
  assign n4554 = n4315 & n4386;
  assign n4555 = n4554 ^ n4317;
  assign n4556 = n4555 ^ n4552;
  assign n4557 = n4553 & ~n4556;
  assign n4558 = n4557 ^ x89;
  assign n4559 = n4558 ^ x90;
  assign n4560 = n4321 & n4386;
  assign n4561 = n4560 ^ n4323;
  assign n4562 = n4561 ^ n4558;
  assign n4563 = n4559 & ~n4562;
  assign n4564 = n4563 ^ x90;
  assign n4565 = n4564 ^ x91;
  assign n4566 = n4327 & n4386;
  assign n4567 = n4566 ^ n4329;
  assign n4568 = n4567 ^ n4564;
  assign n4569 = n4565 & ~n4568;
  assign n4570 = n4569 ^ x91;
  assign n4571 = n4570 ^ x92;
  assign n4572 = n4333 & n4386;
  assign n4573 = n4572 ^ n4335;
  assign n4574 = n4573 ^ n4570;
  assign n4575 = n4571 & ~n4574;
  assign n4576 = n4575 ^ x92;
  assign n4577 = n4576 ^ x93;
  assign n4578 = n4339 & n4386;
  assign n4579 = n4578 ^ n4341;
  assign n4580 = n4579 ^ n4576;
  assign n4581 = n4577 & ~n4580;
  assign n4582 = n4581 ^ x93;
  assign n4583 = n4582 ^ x94;
  assign n4584 = n4345 & n4386;
  assign n4585 = n4584 ^ n4347;
  assign n4586 = n4585 ^ n4582;
  assign n4587 = n4583 & n4586;
  assign n4588 = n4587 ^ x94;
  assign n4589 = n4588 ^ x95;
  assign n4590 = n4351 & n4386;
  assign n4591 = n4590 ^ n4353;
  assign n4592 = n4591 ^ n4588;
  assign n4593 = n4589 & ~n4592;
  assign n4594 = n4593 ^ x95;
  assign n4595 = n4594 ^ x96;
  assign n4596 = n4356 ^ x95;
  assign n4597 = n4386 & n4596;
  assign n4598 = n4597 ^ n4142;
  assign n4599 = n4598 ^ n4594;
  assign n4600 = n4595 & ~n4599;
  assign n4601 = n4600 ^ n4594;
  assign n4602 = ~n4367 & n4601;
  assign n4606 = x97 & n4140;
  assign n4607 = ~x98 & n241;
  assign n4608 = ~n4606 & n4607;
  assign n4609 = ~n4602 & n4608;
  assign n4610 = n4422 & n4609;
  assign n4611 = n4610 ^ n4424;
  assign n4612 = n4611 ^ x69;
  assign n4613 = n4415 & n4609;
  assign n4614 = n4613 ^ n4418;
  assign n4615 = x68 & n4614;
  assign n4616 = n4615 ^ n4611;
  assign n4617 = n4616 ^ n4611;
  assign n4618 = ~x29 & ~x30;
  assign n4619 = ~n4609 & n4618;
  assign n4620 = ~x29 & x65;
  assign n4621 = ~n4619 & ~n4620;
  assign n4622 = x64 & ~n4621;
  assign n4623 = x64 & n4609;
  assign n4624 = x29 & ~x65;
  assign n4625 = x30 & ~n4624;
  assign n4626 = n4625 ^ n4406;
  assign n4627 = n4623 & n4626;
  assign n4628 = n4627 ^ n4406;
  assign n4629 = ~n4622 & ~n4628;
  assign n4630 = n4629 ^ x66;
  assign n4631 = n289 & ~n4386;
  assign n4632 = n4631 ^ x65;
  assign n4633 = ~x30 & n4632;
  assign n4634 = ~n202 & ~n4633;
  assign n4635 = x65 & n4386;
  assign n4636 = x30 & ~n4635;
  assign n4637 = x65 & n4636;
  assign n4638 = n4634 & ~n4637;
  assign n4639 = n4638 ^ n4398;
  assign n4640 = n4638 ^ n4636;
  assign n4641 = n4638 ^ n4609;
  assign n4642 = n4638 & n4641;
  assign n4643 = n4642 ^ n4638;
  assign n4644 = n4640 & n4643;
  assign n4645 = n4644 ^ n4642;
  assign n4646 = n4645 ^ n4638;
  assign n4647 = n4646 ^ n4609;
  assign n4648 = ~n4639 & n4647;
  assign n4649 = n4648 ^ n4398;
  assign n4650 = n4649 ^ x31;
  assign n4651 = n4650 ^ n4629;
  assign n4652 = ~n4630 & ~n4651;
  assign n4653 = n4652 ^ x66;
  assign n4654 = ~x67 & ~n4653;
  assign n4655 = x67 & ~n4629;
  assign n4656 = ~x66 & n4650;
  assign n4657 = n4655 & ~n4656;
  assign n4658 = n1864 & ~n4650;
  assign n4659 = n4411 ^ x66;
  assign n4660 = n4609 & ~n4659;
  assign n4661 = n4660 ^ n4396;
  assign n4662 = ~n4658 & n4661;
  assign n4663 = ~n4657 & n4662;
  assign n4664 = ~n4654 & ~n4663;
  assign n4665 = ~x68 & ~n4614;
  assign n4666 = n4664 & ~n4665;
  assign n4667 = n4666 ^ n4611;
  assign n4668 = n4667 ^ n4611;
  assign n4669 = ~n4617 & ~n4668;
  assign n4670 = n4669 ^ n4611;
  assign n4671 = ~n4612 & ~n4670;
  assign n4672 = n4671 ^ x69;
  assign n4673 = n4672 ^ x70;
  assign n4674 = n4428 & n4609;
  assign n4675 = n4674 ^ n4430;
  assign n4676 = n4675 ^ n4672;
  assign n4677 = n4673 & n4676;
  assign n4678 = n4677 ^ x70;
  assign n4679 = n4678 ^ x71;
  assign n4680 = n4434 & n4609;
  assign n4681 = n4680 ^ n4436;
  assign n4682 = n4681 ^ n4678;
  assign n4683 = n4679 & n4682;
  assign n4684 = n4683 ^ x71;
  assign n4685 = n4684 ^ x72;
  assign n4686 = n4440 & n4609;
  assign n4687 = n4686 ^ n4442;
  assign n4688 = n4687 ^ n4684;
  assign n4689 = n4685 & ~n4688;
  assign n4690 = n4689 ^ x72;
  assign n4691 = n4690 ^ x73;
  assign n4692 = n4446 & n4609;
  assign n4693 = n4692 ^ n4448;
  assign n4694 = n4693 ^ n4690;
  assign n4695 = n4691 & n4694;
  assign n4696 = n4695 ^ x73;
  assign n4697 = n4696 ^ x74;
  assign n4698 = n4452 & n4609;
  assign n4699 = n4698 ^ n4454;
  assign n4700 = n4699 ^ n4696;
  assign n4701 = n4697 & ~n4700;
  assign n4702 = n4701 ^ x74;
  assign n4703 = n4702 ^ x75;
  assign n4704 = n4458 & n4609;
  assign n4705 = n4704 ^ n4460;
  assign n4706 = n4705 ^ n4702;
  assign n4707 = n4703 & ~n4706;
  assign n4708 = n4707 ^ x75;
  assign n4709 = n4708 ^ x76;
  assign n4710 = n4464 & n4609;
  assign n4711 = n4710 ^ n4466;
  assign n4712 = n4711 ^ n4708;
  assign n4713 = n4709 & ~n4712;
  assign n4714 = n4713 ^ x76;
  assign n4715 = n4714 ^ x77;
  assign n4716 = n4470 & n4609;
  assign n4717 = n4716 ^ n4472;
  assign n4718 = n4717 ^ n4714;
  assign n4719 = n4715 & ~n4718;
  assign n4720 = n4719 ^ x77;
  assign n4721 = n4720 ^ x78;
  assign n4722 = n4476 & n4609;
  assign n4723 = n4722 ^ n4478;
  assign n4724 = n4723 ^ n4720;
  assign n4725 = n4721 & ~n4724;
  assign n4726 = n4725 ^ x78;
  assign n4727 = n4726 ^ x79;
  assign n4728 = n4482 & n4609;
  assign n4729 = n4728 ^ n4484;
  assign n4730 = n4729 ^ n4726;
  assign n4731 = n4727 & ~n4730;
  assign n4732 = n4731 ^ x79;
  assign n4733 = n4732 ^ x80;
  assign n4734 = n4488 & n4609;
  assign n4735 = n4734 ^ n4490;
  assign n4736 = n4735 ^ n4732;
  assign n4737 = n4733 & ~n4736;
  assign n4738 = n4737 ^ x80;
  assign n4739 = n4738 ^ x81;
  assign n4740 = n4494 & n4609;
  assign n4741 = n4740 ^ n4497;
  assign n4742 = n4741 ^ n4738;
  assign n4743 = n4739 & ~n4742;
  assign n4744 = n4743 ^ x81;
  assign n4745 = n4744 ^ x82;
  assign n4746 = n4501 & n4609;
  assign n4747 = n4746 ^ n4507;
  assign n4748 = n4747 ^ n4744;
  assign n4749 = n4745 & n4748;
  assign n4750 = n4749 ^ x82;
  assign n4751 = n4750 ^ x83;
  assign n4752 = n4511 & n4609;
  assign n4753 = n4752 ^ n4513;
  assign n4754 = n4753 ^ n4750;
  assign n4755 = n4751 & ~n4754;
  assign n4756 = n4755 ^ x83;
  assign n4757 = n4756 ^ x84;
  assign n4758 = n4517 & n4609;
  assign n4759 = n4758 ^ n4519;
  assign n4760 = n4759 ^ n4756;
  assign n4761 = n4757 & n4760;
  assign n4762 = n4761 ^ x84;
  assign n4763 = n4762 ^ x85;
  assign n4764 = n4523 & n4609;
  assign n4765 = n4764 ^ n4525;
  assign n4766 = n4765 ^ n4762;
  assign n4767 = n4763 & ~n4766;
  assign n4768 = n4767 ^ x85;
  assign n4769 = n4768 ^ x86;
  assign n4770 = n4529 & n4609;
  assign n4771 = n4770 ^ n4531;
  assign n4772 = n4771 ^ n4768;
  assign n4773 = n4769 & ~n4772;
  assign n4774 = n4773 ^ x86;
  assign n4775 = n4774 ^ x87;
  assign n4776 = n4535 & n4609;
  assign n4777 = n4776 ^ n4537;
  assign n4778 = n4777 ^ n4774;
  assign n4779 = n4775 & n4778;
  assign n4780 = n4779 ^ x87;
  assign n4781 = n4780 ^ x88;
  assign n4782 = n4541 & n4609;
  assign n4783 = n4782 ^ n4543;
  assign n4784 = n4783 ^ n4780;
  assign n4785 = n4781 & n4784;
  assign n4786 = n4785 ^ x88;
  assign n4787 = n4786 ^ x89;
  assign n4788 = n4547 & n4609;
  assign n4789 = n4788 ^ n4549;
  assign n4790 = n4789 ^ n4786;
  assign n4791 = n4787 & n4790;
  assign n4792 = n4791 ^ x89;
  assign n4793 = n4792 ^ x90;
  assign n4794 = n4553 & n4609;
  assign n4795 = n4794 ^ n4555;
  assign n4796 = n4795 ^ n4792;
  assign n4797 = n4793 & ~n4796;
  assign n4798 = n4797 ^ x90;
  assign n4799 = n4798 ^ x91;
  assign n4800 = n4559 & n4609;
  assign n4801 = n4800 ^ n4561;
  assign n4802 = n4801 ^ n4798;
  assign n4803 = n4799 & ~n4802;
  assign n4804 = n4803 ^ x91;
  assign n4805 = n4804 ^ x92;
  assign n4806 = n4565 & n4609;
  assign n4807 = n4806 ^ n4567;
  assign n4808 = n4807 ^ n4804;
  assign n4809 = n4805 & ~n4808;
  assign n4810 = n4809 ^ x92;
  assign n4811 = n4810 ^ x93;
  assign n4812 = n4571 & n4609;
  assign n4813 = n4812 ^ n4573;
  assign n4814 = n4813 ^ n4810;
  assign n4815 = n4811 & ~n4814;
  assign n4816 = n4815 ^ x93;
  assign n4817 = n4816 ^ x94;
  assign n4818 = n4577 & n4609;
  assign n4819 = n4818 ^ n4579;
  assign n4820 = n4819 ^ n4816;
  assign n4821 = n4817 & ~n4820;
  assign n4822 = n4821 ^ x94;
  assign n4823 = n4822 ^ x95;
  assign n4824 = n4583 & n4609;
  assign n4825 = n4824 ^ n4585;
  assign n4826 = n4825 ^ n4822;
  assign n4827 = n4823 & n4826;
  assign n4828 = n4827 ^ x95;
  assign n4829 = n4828 ^ x96;
  assign n4365 = x98 & n4364;
  assign n4366 = n241 & ~n4365;
  assign n4603 = ~n240 & ~n4602;
  assign n4604 = ~x98 & ~n4364;
  assign n4605 = ~n4603 & n4604;
  assign n4830 = n4589 & n4609;
  assign n4831 = n4830 ^ n4591;
  assign n4832 = n4831 ^ n4828;
  assign n4833 = n4829 & ~n4832;
  assign n4834 = n4833 ^ x96;
  assign n4835 = n4834 ^ x97;
  assign n4836 = n4595 & n4609;
  assign n4837 = n4836 ^ n4598;
  assign n4838 = n4837 ^ n4834;
  assign n4839 = n4835 & ~n4838;
  assign n4840 = n4839 ^ n4834;
  assign n4841 = ~n4605 & n4840;
  assign n4842 = n4366 & ~n4841;
  assign n4843 = n4829 & n4842;
  assign n4844 = n4843 ^ n4831;
  assign n4845 = ~x97 & ~n4844;
  assign n4846 = n4835 & n4842;
  assign n4847 = n4846 ^ n4837;
  assign n4848 = ~x98 & n4847;
  assign n4849 = ~n4845 & ~n4848;
  assign n4850 = n4805 & n4842;
  assign n4851 = n4850 ^ n4807;
  assign n4852 = ~x93 & ~n4851;
  assign n4853 = n4811 & n4842;
  assign n4854 = n4853 ^ n4813;
  assign n4855 = ~x94 & ~n4854;
  assign n4856 = ~n4852 & ~n4855;
  assign n4857 = n4664 ^ x68;
  assign n4858 = n4842 & n4857;
  assign n4859 = n4858 ^ n4614;
  assign n4860 = ~x69 & ~n4859;
  assign n4861 = ~n4615 & ~n4666;
  assign n4862 = n4861 ^ x69;
  assign n4863 = n4842 & ~n4862;
  assign n4864 = n4863 ^ n4611;
  assign n4865 = ~x70 & n4864;
  assign n4866 = ~n4860 & ~n4865;
  assign n4867 = ~x29 & n4842;
  assign n4868 = ~x28 & ~n4867;
  assign n4869 = ~x65 & ~n4868;
  assign n4870 = ~x28 & ~n4624;
  assign n4871 = ~n4842 & ~n4870;
  assign n4872 = x28 & ~x29;
  assign n4873 = x64 & ~n4872;
  assign n4874 = ~n4871 & n4873;
  assign n4875 = ~n4869 & n4874;
  assign n4876 = x64 & n4842;
  assign n4877 = n4620 & ~n4876;
  assign n4878 = ~n4875 & ~n4877;
  assign n4879 = n4878 ^ x66;
  assign n4880 = x65 & n4842;
  assign n4881 = ~n4623 & ~n4880;
  assign n4882 = x65 & n4609;
  assign n4883 = x29 & ~n4882;
  assign n4884 = n4876 & ~n4883;
  assign n4885 = ~n4881 & ~n4884;
  assign n4886 = n289 & ~n4609;
  assign n4887 = n4886 ^ x65;
  assign n4888 = n4867 & n4887;
  assign n4889 = ~n4885 & ~n4888;
  assign n4890 = n4889 ^ x30;
  assign n4891 = n4890 ^ n4878;
  assign n4892 = ~n4879 & n4891;
  assign n4893 = n4892 ^ x66;
  assign n4894 = n4893 ^ x67;
  assign n4895 = ~n4630 & n4842;
  assign n4896 = n4895 ^ n4650;
  assign n4897 = n4896 ^ n4893;
  assign n4898 = n4894 & n4897;
  assign n4899 = n4898 ^ x67;
  assign n4900 = n4899 ^ x68;
  assign n4901 = n4653 ^ x67;
  assign n4902 = n4842 & n4901;
  assign n4903 = n4902 ^ n4661;
  assign n4904 = n4903 ^ n4899;
  assign n4905 = n4900 & n4904;
  assign n4906 = n4905 ^ x68;
  assign n4907 = n4866 & n4906;
  assign n4908 = n4864 ^ x70;
  assign n4909 = x69 & n4859;
  assign n4910 = n4909 ^ n4864;
  assign n4911 = ~n4908 & n4910;
  assign n4912 = n4911 ^ x70;
  assign n4913 = ~n4907 & ~n4912;
  assign n4914 = n4913 ^ x71;
  assign n4915 = n4673 & n4842;
  assign n4916 = n4915 ^ n4675;
  assign n4917 = n4916 ^ n4913;
  assign n4918 = ~n4914 & ~n4917;
  assign n4919 = n4918 ^ x71;
  assign n4920 = n4919 ^ x72;
  assign n4921 = n4679 & n4842;
  assign n4922 = n4921 ^ n4681;
  assign n4923 = n4922 ^ n4919;
  assign n4924 = n4920 & n4923;
  assign n4925 = n4924 ^ x72;
  assign n4926 = n4925 ^ x73;
  assign n4927 = n4685 & n4842;
  assign n4928 = n4927 ^ n4687;
  assign n4929 = n4928 ^ n4925;
  assign n4930 = n4926 & ~n4929;
  assign n4931 = n4930 ^ x73;
  assign n4932 = n4931 ^ x74;
  assign n4933 = n4691 & n4842;
  assign n4934 = n4933 ^ n4693;
  assign n4935 = n4934 ^ n4931;
  assign n4936 = n4932 & n4935;
  assign n4937 = n4936 ^ x74;
  assign n4938 = n4937 ^ x75;
  assign n4939 = n4697 & n4842;
  assign n4940 = n4939 ^ n4699;
  assign n4941 = n4940 ^ n4937;
  assign n4942 = n4938 & ~n4941;
  assign n4943 = n4942 ^ x75;
  assign n4944 = n4943 ^ x76;
  assign n4945 = n4703 & n4842;
  assign n4946 = n4945 ^ n4705;
  assign n4947 = n4946 ^ n4943;
  assign n4948 = n4944 & ~n4947;
  assign n4949 = n4948 ^ x76;
  assign n4950 = n4949 ^ x77;
  assign n4951 = n4709 & n4842;
  assign n4952 = n4951 ^ n4711;
  assign n4953 = n4952 ^ n4949;
  assign n4954 = n4950 & ~n4953;
  assign n4955 = n4954 ^ x77;
  assign n4956 = n4955 ^ x78;
  assign n4957 = n4715 & n4842;
  assign n4958 = n4957 ^ n4717;
  assign n4959 = n4958 ^ n4955;
  assign n4960 = n4956 & ~n4959;
  assign n4961 = n4960 ^ x78;
  assign n4962 = n4961 ^ x79;
  assign n4963 = n4721 & n4842;
  assign n4964 = n4963 ^ n4723;
  assign n4965 = n4964 ^ n4961;
  assign n4966 = n4962 & ~n4965;
  assign n4967 = n4966 ^ x79;
  assign n4968 = n4967 ^ x80;
  assign n4969 = n4727 & n4842;
  assign n4970 = n4969 ^ n4729;
  assign n4971 = n4970 ^ n4967;
  assign n4972 = n4968 & ~n4971;
  assign n4973 = n4972 ^ x80;
  assign n4974 = n4973 ^ x81;
  assign n4975 = n4733 & n4842;
  assign n4976 = n4975 ^ n4735;
  assign n4977 = n4976 ^ n4973;
  assign n4978 = n4974 & ~n4977;
  assign n4979 = n4978 ^ x81;
  assign n4980 = n4979 ^ x82;
  assign n4981 = n4739 & n4842;
  assign n4982 = n4981 ^ n4741;
  assign n4983 = n4982 ^ n4979;
  assign n4984 = n4980 & ~n4983;
  assign n4985 = n4984 ^ x82;
  assign n4986 = n4985 ^ x83;
  assign n4987 = n4745 & n4842;
  assign n4988 = n4987 ^ n4747;
  assign n4989 = n4988 ^ n4985;
  assign n4990 = n4986 & n4989;
  assign n4991 = n4990 ^ x83;
  assign n4992 = n4991 ^ x84;
  assign n4993 = n4751 & n4842;
  assign n4994 = n4993 ^ n4753;
  assign n4995 = n4994 ^ n4991;
  assign n4996 = n4992 & ~n4995;
  assign n4997 = n4996 ^ x84;
  assign n4998 = n4997 ^ x85;
  assign n4999 = n4757 & n4842;
  assign n5000 = n4999 ^ n4759;
  assign n5001 = n5000 ^ n4997;
  assign n5002 = n4998 & n5001;
  assign n5003 = n5002 ^ x85;
  assign n5004 = n5003 ^ x86;
  assign n5005 = n4763 & n4842;
  assign n5006 = n5005 ^ n4765;
  assign n5007 = n5006 ^ n5003;
  assign n5008 = n5004 & ~n5007;
  assign n5009 = n5008 ^ x86;
  assign n5010 = n5009 ^ x87;
  assign n5011 = n4769 & n4842;
  assign n5012 = n5011 ^ n4771;
  assign n5013 = n5012 ^ n5009;
  assign n5014 = n5010 & ~n5013;
  assign n5015 = n5014 ^ x87;
  assign n5016 = n5015 ^ x88;
  assign n5017 = n4775 & n4842;
  assign n5018 = n5017 ^ n4777;
  assign n5019 = n5018 ^ n5015;
  assign n5020 = n5016 & n5019;
  assign n5021 = n5020 ^ x88;
  assign n5022 = n5021 ^ x89;
  assign n5023 = n4781 & n4842;
  assign n5024 = n5023 ^ n4783;
  assign n5025 = n5024 ^ n5021;
  assign n5026 = n5022 & n5025;
  assign n5027 = n5026 ^ x89;
  assign n5028 = n5027 ^ x90;
  assign n5029 = n4787 & n4842;
  assign n5030 = n5029 ^ n4789;
  assign n5031 = n5030 ^ n5027;
  assign n5032 = n5028 & n5031;
  assign n5033 = n5032 ^ x90;
  assign n5034 = n5033 ^ x91;
  assign n5035 = n4793 & n4842;
  assign n5036 = n5035 ^ n4795;
  assign n5037 = n5036 ^ n5033;
  assign n5038 = n5034 & ~n5037;
  assign n5039 = n5038 ^ x91;
  assign n5040 = n5039 ^ x92;
  assign n5041 = n4799 & n4842;
  assign n5042 = n5041 ^ n4801;
  assign n5043 = n5042 ^ n5039;
  assign n5044 = n5040 & ~n5043;
  assign n5045 = n5044 ^ x92;
  assign n5046 = n4856 & n5045;
  assign n5047 = n4854 ^ x94;
  assign n5048 = x93 & n4851;
  assign n5049 = n5048 ^ n4854;
  assign n5050 = n5047 & ~n5049;
  assign n5051 = n5050 ^ x94;
  assign n5052 = ~n5046 & ~n5051;
  assign n5053 = n5052 ^ x95;
  assign n5054 = n4817 & n4842;
  assign n5055 = n5054 ^ n4819;
  assign n5056 = n5055 ^ n5052;
  assign n5057 = ~n5053 & n5056;
  assign n5058 = n5057 ^ x95;
  assign n5059 = n5058 ^ x96;
  assign n5060 = n4823 & n4842;
  assign n5061 = n5060 ^ n4825;
  assign n5062 = n5061 ^ n5058;
  assign n5063 = n5059 & n5062;
  assign n5064 = n5063 ^ x96;
  assign n5065 = n4849 & n5064;
  assign n5066 = n4847 ^ x98;
  assign n5067 = x97 & n4844;
  assign n5068 = n5067 ^ n4847;
  assign n5069 = ~n5066 & n5068;
  assign n5070 = n5069 ^ x98;
  assign n5071 = ~n5065 & ~n5070;
  assign n5072 = x99 & ~n5071;
  assign n5073 = ~x100 & n155;
  assign n5074 = ~n5072 & n5073;
  assign n5075 = n4363 & ~n4609;
  assign n5076 = ~n4842 & n5075;
  assign n5077 = ~n240 & ~n5076;
  assign n5078 = ~n5074 & ~n5077;
  assign n5079 = ~n240 & ~n5078;
  assign n5080 = n5073 & ~n5079;
  assign n5081 = x100 & n5079;
  assign n5082 = n155 & ~n5081;
  assign n5083 = n5071 ^ x99;
  assign n5084 = n5077 ^ n5071;
  assign n5085 = ~n5083 & ~n5084;
  assign n5086 = n5085 ^ n5071;
  assign n5087 = n5073 & n5086;
  assign n5088 = n5034 & n5087;
  assign n5089 = n5088 ^ n5036;
  assign n5090 = ~x92 & ~n5089;
  assign n5091 = n5040 & n5087;
  assign n5092 = n5091 ^ n5042;
  assign n5093 = ~x93 & ~n5092;
  assign n5094 = ~n5090 & ~n5093;
  assign n5095 = n5004 & n5087;
  assign n5096 = n5095 ^ n5006;
  assign n5097 = ~x87 & ~n5096;
  assign n5098 = n5010 & n5087;
  assign n5099 = n5098 ^ n5012;
  assign n5100 = ~x88 & ~n5099;
  assign n5101 = ~n5097 & ~n5100;
  assign n5102 = n4974 & n5087;
  assign n5103 = n5102 ^ n4976;
  assign n5104 = ~x82 & ~n5103;
  assign n5105 = n4968 & n5087;
  assign n5106 = n5105 ^ n4970;
  assign n5107 = ~x81 & ~n5106;
  assign n5108 = ~n5104 & ~n5107;
  assign n5109 = n4950 & n5087;
  assign n5110 = n5109 ^ n4952;
  assign n5111 = n5110 ^ x78;
  assign n5112 = n4944 & n5087;
  assign n5113 = n5112 ^ n4946;
  assign n5114 = x77 & n5113;
  assign n5115 = n5114 ^ n5110;
  assign n5116 = n5115 ^ n5110;
  assign n5117 = ~x77 & ~n5113;
  assign n5118 = n289 & ~n4842;
  assign n5119 = n5118 ^ x65;
  assign n5120 = ~x28 & n5119;
  assign n5121 = ~n202 & ~n5120;
  assign n5122 = x28 & ~n4880;
  assign n5123 = x65 & n5122;
  assign n5124 = n5121 & ~n5123;
  assign n5125 = n5124 ^ n4876;
  assign n5126 = n5124 ^ n5122;
  assign n5127 = n5124 ^ n5087;
  assign n5128 = n5124 & n5127;
  assign n5129 = n5128 ^ n5124;
  assign n5130 = n5126 & n5129;
  assign n5131 = n5130 ^ n5128;
  assign n5132 = n5131 ^ n5124;
  assign n5133 = n5132 ^ n5087;
  assign n5134 = ~n5125 & n5133;
  assign n5135 = n5134 ^ n4876;
  assign n5136 = n5135 ^ x29;
  assign n5137 = n5136 ^ x66;
  assign n5138 = x64 & n5087;
  assign n5139 = x27 & ~x65;
  assign n5140 = x28 & ~n5139;
  assign n5141 = n5138 & n5140;
  assign n5143 = x65 ^ x28;
  assign n5150 = n5143 ^ x65;
  assign n5142 = x65 ^ x27;
  assign n5144 = n5143 ^ n5142;
  assign n5145 = n5144 ^ x65;
  assign n5146 = n5142 ^ x64;
  assign n5147 = n5146 ^ n5142;
  assign n5148 = n5147 ^ n5145;
  assign n5149 = ~n5145 & ~n5148;
  assign n5151 = n5150 ^ n5149;
  assign n5152 = n5151 ^ n5145;
  assign n5153 = n5087 ^ x65;
  assign n5154 = n5153 ^ x65;
  assign n5155 = n5149 ^ n5145;
  assign n5156 = ~n5154 & ~n5155;
  assign n5157 = n5156 ^ x65;
  assign n5158 = ~n5152 & n5157;
  assign n5159 = n5158 ^ x65;
  assign n5160 = n5159 ^ x65;
  assign n5161 = n5160 ^ x65;
  assign n5162 = ~n5141 & ~n5161;
  assign n5163 = n5162 ^ n5136;
  assign n5164 = ~n5137 & ~n5163;
  assign n5165 = n5164 ^ x66;
  assign n5166 = n5165 ^ x67;
  assign n5167 = ~n4879 & n5087;
  assign n5168 = n5167 ^ n4890;
  assign n5169 = n5168 ^ n5165;
  assign n5170 = n5166 & ~n5169;
  assign n5171 = n5170 ^ x67;
  assign n5172 = n5171 ^ x68;
  assign n5173 = n4894 & n5087;
  assign n5174 = n5173 ^ n4896;
  assign n5175 = n5174 ^ n5171;
  assign n5176 = n5172 & n5175;
  assign n5177 = n5176 ^ x68;
  assign n5178 = n5177 ^ x69;
  assign n5179 = n4900 & n5087;
  assign n5180 = n5179 ^ n4903;
  assign n5181 = n5180 ^ n5177;
  assign n5182 = n5178 & n5181;
  assign n5183 = n5182 ^ x69;
  assign n5184 = n5183 ^ x70;
  assign n5185 = n4906 ^ x69;
  assign n5186 = n5087 & n5185;
  assign n5187 = n5186 ^ n4859;
  assign n5188 = n5187 ^ n5183;
  assign n5189 = n5184 & ~n5188;
  assign n5190 = n5189 ^ x70;
  assign n5191 = n5190 ^ x71;
  assign n5192 = n4906 ^ n4859;
  assign n5193 = n5185 & ~n5192;
  assign n5194 = n5193 ^ x69;
  assign n5195 = n5194 ^ x70;
  assign n5196 = n5087 & n5195;
  assign n5197 = n5196 ^ n4864;
  assign n5198 = n5197 ^ n5190;
  assign n5199 = n5191 & n5198;
  assign n5200 = n5199 ^ x71;
  assign n5201 = n5200 ^ x72;
  assign n5202 = ~n4914 & n5087;
  assign n5203 = n5202 ^ n4916;
  assign n5204 = n5203 ^ n5200;
  assign n5205 = n5201 & n5204;
  assign n5206 = n5205 ^ x72;
  assign n5207 = n5206 ^ x73;
  assign n5208 = n4920 & n5087;
  assign n5209 = n5208 ^ n4922;
  assign n5210 = n5209 ^ n5206;
  assign n5211 = n5207 & n5210;
  assign n5212 = n5211 ^ x73;
  assign n5213 = n5212 ^ x74;
  assign n5214 = n4926 & n5087;
  assign n5215 = n5214 ^ n4928;
  assign n5216 = n5215 ^ n5212;
  assign n5217 = n5213 & ~n5216;
  assign n5218 = n5217 ^ x74;
  assign n5219 = n5218 ^ x75;
  assign n5220 = n4932 & n5087;
  assign n5221 = n5220 ^ n4934;
  assign n5222 = n5221 ^ n5218;
  assign n5223 = n5219 & n5222;
  assign n5224 = n5223 ^ x75;
  assign n5225 = n5224 ^ x76;
  assign n5226 = n4938 & n5087;
  assign n5227 = n5226 ^ n4940;
  assign n5228 = n5227 ^ n5224;
  assign n5229 = n5225 & ~n5228;
  assign n5230 = n5229 ^ x76;
  assign n5231 = ~n5117 & n5230;
  assign n5232 = n5231 ^ n5110;
  assign n5233 = n5232 ^ n5110;
  assign n5234 = ~n5116 & ~n5233;
  assign n5235 = n5234 ^ n5110;
  assign n5236 = n5111 & n5235;
  assign n5237 = n5236 ^ x78;
  assign n5238 = n5237 ^ x79;
  assign n5239 = n4958 ^ x78;
  assign n5240 = n5239 ^ n4955;
  assign n5241 = n5240 ^ n4958;
  assign n5242 = n5087 & n5241;
  assign n5243 = n5242 ^ n4958;
  assign n5244 = n5243 ^ n5237;
  assign n5245 = n5238 & ~n5244;
  assign n5246 = n5245 ^ x79;
  assign n5247 = n5246 ^ x80;
  assign n5248 = n4962 & n5087;
  assign n5249 = n5248 ^ n4964;
  assign n5250 = n5249 ^ n5246;
  assign n5251 = n5247 & ~n5250;
  assign n5252 = n5251 ^ x80;
  assign n5253 = n5108 & n5252;
  assign n5254 = n5103 ^ x82;
  assign n5255 = x81 & n5106;
  assign n5256 = n5255 ^ n5103;
  assign n5257 = n5254 & ~n5256;
  assign n5258 = n5257 ^ x82;
  assign n5259 = ~n5253 & ~n5258;
  assign n5260 = n4980 & n5087;
  assign n5261 = n5260 ^ n4982;
  assign n5262 = ~x83 & ~n5261;
  assign n5263 = n4986 & n5087;
  assign n5264 = n5263 ^ n4988;
  assign n5265 = ~x84 & n5264;
  assign n5266 = ~n5262 & ~n5265;
  assign n5267 = ~n5259 & n5266;
  assign n5268 = n5264 ^ x84;
  assign n5269 = x83 & n5261;
  assign n5270 = n5269 ^ n5264;
  assign n5271 = ~n5268 & n5270;
  assign n5272 = n5271 ^ x84;
  assign n5273 = ~n5267 & ~n5272;
  assign n5274 = n5273 ^ x85;
  assign n5275 = n4992 & n5087;
  assign n5276 = n5275 ^ n4994;
  assign n5277 = n5276 ^ n5273;
  assign n5278 = ~n5274 & n5277;
  assign n5279 = n5278 ^ x85;
  assign n5280 = n5279 ^ x86;
  assign n5281 = n4998 & n5087;
  assign n5282 = n5281 ^ n5000;
  assign n5283 = n5282 ^ n5279;
  assign n5284 = n5280 & n5283;
  assign n5285 = n5284 ^ x86;
  assign n5286 = n5101 & n5285;
  assign n5287 = n5099 ^ x88;
  assign n5288 = x87 & n5096;
  assign n5289 = n5288 ^ n5099;
  assign n5290 = n5287 & ~n5289;
  assign n5291 = n5290 ^ x88;
  assign n5292 = ~n5286 & ~n5291;
  assign n5293 = n5292 ^ x89;
  assign n5294 = n5016 & n5087;
  assign n5295 = n5294 ^ n5018;
  assign n5296 = n5295 ^ n5292;
  assign n5297 = ~n5293 & ~n5296;
  assign n5298 = n5297 ^ x89;
  assign n5299 = n5298 ^ x90;
  assign n5300 = n5022 & n5087;
  assign n5301 = n5300 ^ n5024;
  assign n5302 = n5301 ^ n5298;
  assign n5303 = n5299 & n5302;
  assign n5304 = n5303 ^ x90;
  assign n5305 = n5304 ^ x91;
  assign n5306 = n5028 & n5087;
  assign n5307 = n5306 ^ n5030;
  assign n5308 = n5307 ^ n5304;
  assign n5309 = n5305 & n5308;
  assign n5310 = n5309 ^ x91;
  assign n5311 = n5094 & n5310;
  assign n5312 = n5092 ^ x93;
  assign n5313 = x92 & n5089;
  assign n5314 = n5313 ^ n5092;
  assign n5315 = n5312 & ~n5314;
  assign n5316 = n5315 ^ x93;
  assign n5317 = ~n5311 & ~n5316;
  assign n5318 = n5317 ^ x94;
  assign n5319 = n5045 ^ x93;
  assign n5320 = n5087 & n5319;
  assign n5321 = n5320 ^ n4851;
  assign n5322 = n5321 ^ n5317;
  assign n5323 = ~n5318 & n5322;
  assign n5324 = n5323 ^ x94;
  assign n5325 = n5324 ^ x95;
  assign n5326 = n5045 ^ n4851;
  assign n5327 = n5319 & ~n5326;
  assign n5328 = n5327 ^ x93;
  assign n5329 = n5328 ^ x94;
  assign n5330 = n5087 & n5329;
  assign n5331 = n5330 ^ n4854;
  assign n5332 = n5331 ^ n5324;
  assign n5333 = n5325 & ~n5332;
  assign n5334 = n5333 ^ x95;
  assign n5335 = n5334 ^ x96;
  assign n5336 = ~n5053 & n5087;
  assign n5337 = n5336 ^ n5055;
  assign n5338 = n5337 ^ n5334;
  assign n5339 = n5335 & ~n5338;
  assign n5340 = n5339 ^ x96;
  assign n5341 = n5340 ^ x97;
  assign n5342 = n5059 & n5087;
  assign n5343 = n5342 ^ n5061;
  assign n5344 = n5343 ^ n5340;
  assign n5345 = n5341 & n5344;
  assign n5346 = n5345 ^ x97;
  assign n5347 = n5346 ^ x98;
  assign n5348 = n5064 ^ x97;
  assign n5349 = n5087 & n5348;
  assign n5350 = n5349 ^ n4844;
  assign n5351 = n5350 ^ n5346;
  assign n5352 = n5347 & ~n5351;
  assign n5353 = n5352 ^ x98;
  assign n5354 = n5353 ^ x99;
  assign n5355 = n5064 ^ n4844;
  assign n5356 = n5348 & ~n5355;
  assign n5357 = n5356 ^ x97;
  assign n5358 = n5357 ^ x98;
  assign n5359 = n5087 & n5358;
  assign n5360 = n5359 ^ n4847;
  assign n5361 = n5360 ^ n5353;
  assign n5362 = n5354 & ~n5361;
  assign n5363 = n5362 ^ n5353;
  assign n5364 = n5082 & ~n5363;
  assign n5365 = ~n5080 & ~n5364;
  assign n5366 = n5078 & n5365;
  assign n5367 = ~n240 & ~n5366;
  assign n5368 = ~x101 & ~n5367;
  assign n5369 = n5354 & ~n5365;
  assign n5370 = n5369 ^ n5360;
  assign n5371 = ~n5368 & ~n5370;
  assign n5372 = x100 & x101;
  assign n5373 = ~n5371 & ~n5372;
  assign n5374 = n5335 & ~n5365;
  assign n5375 = n5374 ^ n5337;
  assign n5376 = ~x97 & ~n5375;
  assign n5377 = n5325 & ~n5365;
  assign n5378 = n5377 ^ n5331;
  assign n5379 = ~x96 & ~n5378;
  assign n5380 = ~n5376 & ~n5379;
  assign n5381 = n5310 ^ x92;
  assign n5382 = n5310 ^ n5089;
  assign n5383 = n5381 & ~n5382;
  assign n5384 = n5383 ^ x92;
  assign n5385 = n5384 ^ x93;
  assign n5386 = ~n5365 & n5385;
  assign n5387 = n5386 ^ n5092;
  assign n5388 = n5387 ^ x94;
  assign n5389 = ~n5365 & n5381;
  assign n5390 = n5389 ^ n5089;
  assign n5391 = ~x93 & ~n5390;
  assign n5392 = n5391 ^ n5387;
  assign n5393 = n5392 ^ n5387;
  assign n5394 = x93 & n5390;
  assign n5395 = n5285 ^ x87;
  assign n5396 = n5285 ^ n5096;
  assign n5397 = n5395 & ~n5396;
  assign n5398 = n5397 ^ x87;
  assign n5399 = n5398 ^ x88;
  assign n5400 = ~n5365 & n5399;
  assign n5401 = n5400 ^ n5099;
  assign n5402 = ~x89 & ~n5401;
  assign n5403 = ~n5293 & ~n5365;
  assign n5404 = n5403 ^ n5295;
  assign n5405 = ~x90 & n5404;
  assign n5406 = ~n5402 & ~n5405;
  assign n5407 = n5225 & ~n5365;
  assign n5408 = n5407 ^ n5227;
  assign n5409 = ~x77 & ~n5408;
  assign n5410 = n5230 ^ x77;
  assign n5411 = ~n5365 & n5410;
  assign n5412 = n5411 ^ n5113;
  assign n5413 = ~x78 & ~n5412;
  assign n5414 = ~n5409 & ~n5413;
  assign n5415 = ~x27 & x64;
  assign n5416 = ~n5153 & n5415;
  assign n5417 = ~n202 & ~n5416;
  assign n5418 = x65 & n5087;
  assign n5419 = x27 & ~n5418;
  assign n5420 = x65 & n5419;
  assign n5421 = n5417 & ~n5420;
  assign n5422 = n5421 ^ n5138;
  assign n5423 = n5421 ^ n5419;
  assign n5424 = n5421 ^ n5365;
  assign n5425 = n5421 & ~n5424;
  assign n5426 = n5425 ^ n5421;
  assign n5427 = n5423 & n5426;
  assign n5428 = n5427 ^ n5425;
  assign n5429 = n5428 ^ n5421;
  assign n5430 = n5429 ^ n5365;
  assign n5431 = ~n5422 & ~n5430;
  assign n5432 = n5431 ^ n5138;
  assign n5433 = n5432 ^ x28;
  assign n5434 = n5433 ^ x66;
  assign n5435 = x64 & ~n5365;
  assign n5436 = x26 & n5139;
  assign n5437 = n5436 ^ x27;
  assign n5438 = n5435 & n5437;
  assign n5439 = ~x26 & n5415;
  assign n5440 = ~x27 & x65;
  assign n5441 = ~n5439 & ~n5440;
  assign n5442 = n5365 & ~n5441;
  assign n5443 = ~x26 & x65;
  assign n5444 = n5443 ^ n5440;
  assign n5445 = x64 & n5444;
  assign n5446 = n5445 ^ n5440;
  assign n5447 = ~n5442 & ~n5446;
  assign n5448 = ~n5438 & n5447;
  assign n5449 = n5448 ^ n5433;
  assign n5450 = ~n5434 & ~n5449;
  assign n5451 = n5450 ^ x66;
  assign n5452 = n5451 ^ x67;
  assign n5453 = n5162 ^ x66;
  assign n5454 = ~n5365 & ~n5453;
  assign n5455 = n5454 ^ n5136;
  assign n5456 = n5455 ^ n5451;
  assign n5457 = n5452 & n5456;
  assign n5458 = n5457 ^ x67;
  assign n5459 = n5458 ^ x68;
  assign n5460 = n5166 & ~n5365;
  assign n5461 = n5460 ^ n5168;
  assign n5462 = n5461 ^ n5458;
  assign n5463 = n5459 & ~n5462;
  assign n5464 = n5463 ^ x68;
  assign n5465 = n5464 ^ x69;
  assign n5466 = n5172 & ~n5365;
  assign n5467 = n5466 ^ n5174;
  assign n5468 = n5467 ^ n5464;
  assign n5469 = n5465 & n5468;
  assign n5470 = n5469 ^ x69;
  assign n5471 = n5470 ^ x70;
  assign n5472 = n5178 & ~n5365;
  assign n5473 = n5472 ^ n5180;
  assign n5474 = n5473 ^ n5470;
  assign n5475 = n5471 & n5474;
  assign n5476 = n5475 ^ x70;
  assign n5477 = n5476 ^ x71;
  assign n5478 = n5184 & ~n5365;
  assign n5479 = n5478 ^ n5187;
  assign n5480 = n5479 ^ n5476;
  assign n5481 = n5477 & ~n5480;
  assign n5482 = n5481 ^ x71;
  assign n5483 = n5482 ^ x72;
  assign n5484 = n5191 & ~n5365;
  assign n5485 = n5484 ^ n5197;
  assign n5486 = n5485 ^ n5482;
  assign n5487 = n5483 & n5486;
  assign n5488 = n5487 ^ x72;
  assign n5489 = n5488 ^ x73;
  assign n5490 = n5201 & ~n5365;
  assign n5491 = n5490 ^ n5203;
  assign n5492 = n5491 ^ n5488;
  assign n5493 = n5489 & n5492;
  assign n5494 = n5493 ^ x73;
  assign n5495 = n5494 ^ x74;
  assign n5496 = n5207 & ~n5365;
  assign n5497 = n5496 ^ n5209;
  assign n5498 = n5497 ^ n5494;
  assign n5499 = n5495 & n5498;
  assign n5500 = n5499 ^ x74;
  assign n5501 = n5500 ^ x75;
  assign n5502 = n5213 & ~n5365;
  assign n5503 = n5502 ^ n5215;
  assign n5504 = n5503 ^ n5500;
  assign n5505 = n5501 & ~n5504;
  assign n5506 = n5505 ^ x75;
  assign n5507 = n5506 ^ x76;
  assign n5508 = n5219 & ~n5365;
  assign n5509 = n5508 ^ n5221;
  assign n5510 = n5509 ^ n5506;
  assign n5511 = n5507 & n5510;
  assign n5512 = n5511 ^ x76;
  assign n5513 = n5414 & n5512;
  assign n5514 = n5412 ^ x78;
  assign n5515 = x77 & n5408;
  assign n5516 = n5515 ^ n5412;
  assign n5517 = n5514 & ~n5516;
  assign n5518 = n5517 ^ x78;
  assign n5519 = ~n5513 & ~n5518;
  assign n5520 = n5519 ^ x79;
  assign n5521 = ~n5114 & ~n5231;
  assign n5522 = n5521 ^ x78;
  assign n5523 = ~n5365 & ~n5522;
  assign n5524 = n5523 ^ n5110;
  assign n5525 = n5524 ^ n5519;
  assign n5526 = ~n5520 & n5525;
  assign n5527 = n5526 ^ x79;
  assign n5528 = n5527 ^ x80;
  assign n5529 = n5238 & ~n5365;
  assign n5530 = n5529 ^ n5243;
  assign n5531 = n5530 ^ n5527;
  assign n5532 = n5528 & ~n5531;
  assign n5533 = n5532 ^ x80;
  assign n5534 = n5533 ^ x81;
  assign n5535 = n5247 & ~n5365;
  assign n5536 = n5535 ^ n5249;
  assign n5537 = n5536 ^ n5533;
  assign n5538 = n5534 & ~n5537;
  assign n5539 = n5538 ^ x81;
  assign n5540 = n5539 ^ x82;
  assign n5541 = n5252 ^ x81;
  assign n5542 = ~n5365 & n5541;
  assign n5543 = n5542 ^ n5106;
  assign n5544 = n5543 ^ n5539;
  assign n5545 = n5540 & ~n5544;
  assign n5546 = n5545 ^ x82;
  assign n5547 = n5546 ^ x83;
  assign n5548 = n5252 ^ n5106;
  assign n5549 = n5541 & ~n5548;
  assign n5550 = n5549 ^ x81;
  assign n5551 = n5550 ^ x82;
  assign n5552 = ~n5365 & n5551;
  assign n5553 = n5552 ^ n5103;
  assign n5554 = n5553 ^ n5546;
  assign n5555 = n5547 & ~n5554;
  assign n5556 = n5555 ^ x83;
  assign n5557 = n5556 ^ x84;
  assign n5558 = n5259 ^ x83;
  assign n5559 = ~n5365 & ~n5558;
  assign n5560 = n5559 ^ n5261;
  assign n5561 = n5560 ^ n5556;
  assign n5562 = n5557 & ~n5561;
  assign n5563 = n5562 ^ x84;
  assign n5564 = n5563 ^ x85;
  assign n5565 = n5261 ^ n5259;
  assign n5566 = ~n5558 & n5565;
  assign n5567 = n5566 ^ x83;
  assign n5568 = n5567 ^ x84;
  assign n5569 = ~n5365 & n5568;
  assign n5570 = n5569 ^ n5264;
  assign n5571 = n5570 ^ n5563;
  assign n5572 = n5564 & n5571;
  assign n5573 = n5572 ^ x85;
  assign n5574 = n5573 ^ x86;
  assign n5575 = ~n5274 & ~n5365;
  assign n5576 = n5575 ^ n5276;
  assign n5577 = n5576 ^ n5573;
  assign n5578 = n5574 & ~n5577;
  assign n5579 = n5578 ^ x86;
  assign n5580 = n5579 ^ x87;
  assign n5581 = n5280 & ~n5365;
  assign n5582 = n5581 ^ n5282;
  assign n5583 = n5582 ^ n5579;
  assign n5584 = n5580 & n5583;
  assign n5585 = n5584 ^ x87;
  assign n5586 = n5585 ^ x88;
  assign n5587 = ~n5365 & n5395;
  assign n5588 = n5587 ^ n5096;
  assign n5589 = n5588 ^ n5585;
  assign n5590 = n5586 & ~n5589;
  assign n5591 = n5590 ^ x88;
  assign n5592 = n5406 & n5591;
  assign n5593 = n5404 ^ x90;
  assign n5594 = x89 & n5401;
  assign n5595 = n5594 ^ n5404;
  assign n5596 = ~n5593 & n5595;
  assign n5597 = n5596 ^ x90;
  assign n5598 = ~n5592 & ~n5597;
  assign n5599 = n5598 ^ x91;
  assign n5600 = n5299 & ~n5365;
  assign n5601 = n5600 ^ n5301;
  assign n5602 = n5601 ^ n5598;
  assign n5603 = ~n5599 & ~n5602;
  assign n5604 = n5603 ^ x91;
  assign n5605 = n5604 ^ x92;
  assign n5606 = n5305 & ~n5365;
  assign n5607 = n5606 ^ n5307;
  assign n5608 = n5607 ^ n5604;
  assign n5609 = n5605 & n5608;
  assign n5610 = n5609 ^ x92;
  assign n5611 = ~n5394 & ~n5610;
  assign n5612 = n5611 ^ n5387;
  assign n5613 = n5612 ^ n5387;
  assign n5614 = ~n5393 & ~n5613;
  assign n5615 = n5614 ^ n5387;
  assign n5616 = n5388 & ~n5615;
  assign n5617 = n5616 ^ x94;
  assign n5618 = n5617 ^ x95;
  assign n5619 = ~n5318 & ~n5365;
  assign n5620 = n5619 ^ n5321;
  assign n5621 = n5620 ^ n5617;
  assign n5622 = n5618 & ~n5621;
  assign n5623 = n5622 ^ x95;
  assign n5624 = n5380 & n5623;
  assign n5625 = n5375 ^ x97;
  assign n5626 = x96 & n5378;
  assign n5627 = n5626 ^ n5375;
  assign n5628 = n5625 & ~n5627;
  assign n5629 = n5628 ^ x97;
  assign n5630 = ~n5624 & ~n5629;
  assign n5631 = n5630 ^ x98;
  assign n5632 = n5341 & ~n5365;
  assign n5633 = n5632 ^ n5343;
  assign n5634 = n5633 ^ n5630;
  assign n5635 = ~n5631 & ~n5634;
  assign n5636 = n5635 ^ x98;
  assign n5637 = n5636 ^ x99;
  assign n5638 = n5347 & ~n5365;
  assign n5639 = n5638 ^ n5350;
  assign n5640 = n5639 ^ n5636;
  assign n5641 = n5637 & ~n5640;
  assign n5642 = n5641 ^ x99;
  assign n5643 = ~n5373 & n5642;
  assign n5644 = x100 & n5371;
  assign n5645 = x101 & n5367;
  assign n5646 = n154 & ~n5645;
  assign n5647 = ~n5644 & n5646;
  assign n5648 = ~n5643 & n5647;
  assign n5649 = x100 & n5367;
  assign n5650 = n5642 & n5649;
  assign n5651 = n5648 & ~n5650;
  assign n5652 = n5591 ^ x89;
  assign n5653 = n5651 & n5652;
  assign n5654 = n5653 ^ n5401;
  assign n5655 = ~x90 & ~n5654;
  assign n5656 = n5591 ^ n5401;
  assign n5657 = n5652 & ~n5656;
  assign n5658 = n5657 ^ x89;
  assign n5659 = n5658 ^ x90;
  assign n5660 = n5651 & n5659;
  assign n5661 = n5660 ^ n5404;
  assign n5662 = ~x91 & n5661;
  assign n5663 = ~n5655 & ~n5662;
  assign n5664 = n5651 ^ n288;
  assign n5665 = n5664 ^ n288;
  assign n5666 = n2322 & n5665;
  assign n5667 = n5666 ^ n288;
  assign n5668 = n5365 & n5667;
  assign n5669 = n5668 ^ n288;
  assign n5670 = x26 & n5669;
  assign n5671 = n5365 ^ x65;
  assign n5672 = n5671 ^ x65;
  assign n5673 = n289 & n5672;
  assign n5674 = n5673 ^ x65;
  assign n5675 = ~x26 & n5674;
  assign n5676 = ~n202 & ~n5675;
  assign n5677 = n5676 ^ n5435;
  assign n5678 = n5651 & ~n5677;
  assign n5679 = n5678 ^ n5435;
  assign n5680 = ~n5670 & ~n5679;
  assign n5681 = n5680 ^ x27;
  assign n5682 = n5681 ^ x66;
  assign n5683 = x64 & n5651;
  assign n5684 = x25 & ~x65;
  assign n5685 = x26 & ~n5684;
  assign n5686 = n5683 & n5685;
  assign n5687 = ~x25 & x64;
  assign n5688 = ~x26 & n5687;
  assign n5689 = ~n5443 & ~n5688;
  assign n5690 = ~n5651 & ~n5689;
  assign n5691 = ~x25 & x65;
  assign n5692 = x64 & n5691;
  assign n5693 = ~x26 & n202;
  assign n5694 = ~n5692 & ~n5693;
  assign n5695 = ~n5690 & n5694;
  assign n5696 = ~n5686 & n5695;
  assign n5697 = n5696 ^ n5681;
  assign n5698 = n5682 & n5697;
  assign n5699 = n5698 ^ x66;
  assign n5700 = n5699 ^ x67;
  assign n5701 = n5448 ^ x66;
  assign n5702 = n5651 & ~n5701;
  assign n5703 = n5702 ^ n5433;
  assign n5704 = n5703 ^ n5699;
  assign n5705 = n5700 & n5704;
  assign n5706 = n5705 ^ x67;
  assign n5707 = n5706 ^ x68;
  assign n5708 = n5452 & n5651;
  assign n5709 = n5708 ^ n5455;
  assign n5710 = n5709 ^ n5706;
  assign n5711 = n5707 & n5710;
  assign n5712 = n5711 ^ x68;
  assign n5713 = n5712 ^ x69;
  assign n5714 = n5459 & n5651;
  assign n5715 = n5714 ^ n5461;
  assign n5716 = n5715 ^ n5712;
  assign n5717 = n5713 & ~n5716;
  assign n5718 = n5717 ^ x69;
  assign n5719 = n5718 ^ x70;
  assign n5720 = n5465 & n5651;
  assign n5721 = n5720 ^ n5467;
  assign n5722 = n5721 ^ n5718;
  assign n5723 = n5719 & n5722;
  assign n5724 = n5723 ^ x70;
  assign n5725 = n5724 ^ x71;
  assign n5726 = n5471 & n5651;
  assign n5727 = n5726 ^ n5473;
  assign n5728 = n5727 ^ n5724;
  assign n5729 = n5725 & n5728;
  assign n5730 = n5729 ^ x71;
  assign n5731 = n5730 ^ x72;
  assign n5732 = n5477 & n5651;
  assign n5733 = n5732 ^ n5479;
  assign n5734 = n5733 ^ n5730;
  assign n5735 = n5731 & ~n5734;
  assign n5736 = n5735 ^ x72;
  assign n5737 = n5736 ^ x73;
  assign n5738 = n5483 & n5651;
  assign n5739 = n5738 ^ n5485;
  assign n5740 = n5739 ^ n5736;
  assign n5741 = n5737 & n5740;
  assign n5742 = n5741 ^ x73;
  assign n5743 = n5742 ^ x74;
  assign n5744 = n5489 & n5651;
  assign n5745 = n5744 ^ n5491;
  assign n5746 = n5745 ^ n5742;
  assign n5747 = n5743 & n5746;
  assign n5748 = n5747 ^ x74;
  assign n5749 = n5748 ^ x75;
  assign n5750 = n5495 & n5651;
  assign n5751 = n5750 ^ n5497;
  assign n5752 = n5751 ^ n5748;
  assign n5753 = n5749 & n5752;
  assign n5754 = n5753 ^ x75;
  assign n5755 = n5754 ^ x76;
  assign n5756 = n5501 & n5651;
  assign n5757 = n5756 ^ n5503;
  assign n5758 = n5757 ^ n5754;
  assign n5759 = n5755 & ~n5758;
  assign n5760 = n5759 ^ x76;
  assign n5761 = n5760 ^ x77;
  assign n5762 = n5507 & n5651;
  assign n5763 = n5762 ^ n5509;
  assign n5764 = n5763 ^ n5760;
  assign n5765 = n5761 & n5764;
  assign n5766 = n5765 ^ x77;
  assign n5767 = n5766 ^ x78;
  assign n5768 = n5512 ^ x77;
  assign n5769 = n5651 & n5768;
  assign n5770 = n5769 ^ n5408;
  assign n5771 = n5770 ^ n5766;
  assign n5772 = n5767 & ~n5771;
  assign n5773 = n5772 ^ x78;
  assign n5774 = n5773 ^ x79;
  assign n5775 = n5512 ^ n5408;
  assign n5776 = n5768 & ~n5775;
  assign n5777 = n5776 ^ x77;
  assign n5778 = n5777 ^ x78;
  assign n5779 = n5651 & n5778;
  assign n5780 = n5779 ^ n5412;
  assign n5781 = n5780 ^ n5773;
  assign n5782 = n5774 & ~n5781;
  assign n5783 = n5782 ^ x79;
  assign n5784 = n5783 ^ x80;
  assign n5785 = ~n5520 & n5651;
  assign n5786 = n5785 ^ n5524;
  assign n5787 = n5786 ^ n5783;
  assign n5788 = n5784 & ~n5787;
  assign n5789 = n5788 ^ x80;
  assign n5790 = n5789 ^ x81;
  assign n5791 = n5528 & n5651;
  assign n5792 = n5791 ^ n5530;
  assign n5793 = n5792 ^ n5789;
  assign n5794 = n5790 & ~n5793;
  assign n5795 = n5794 ^ x81;
  assign n5796 = n5795 ^ x82;
  assign n5797 = n5534 & n5651;
  assign n5798 = n5797 ^ n5536;
  assign n5799 = n5798 ^ n5795;
  assign n5800 = n5796 & ~n5799;
  assign n5801 = n5800 ^ x82;
  assign n5802 = n5801 ^ x83;
  assign n5803 = n5540 & n5651;
  assign n5804 = n5803 ^ n5543;
  assign n5805 = n5804 ^ n5801;
  assign n5806 = n5802 & ~n5805;
  assign n5807 = n5806 ^ x83;
  assign n5808 = n5807 ^ x84;
  assign n5809 = n5547 & n5651;
  assign n5810 = n5809 ^ n5553;
  assign n5811 = n5810 ^ n5807;
  assign n5812 = n5808 & ~n5811;
  assign n5813 = n5812 ^ x84;
  assign n5814 = n5813 ^ x85;
  assign n5815 = n5557 & n5651;
  assign n5816 = n5815 ^ n5560;
  assign n5817 = n5816 ^ n5813;
  assign n5818 = n5814 & ~n5817;
  assign n5819 = n5818 ^ x85;
  assign n5820 = n5819 ^ x86;
  assign n5821 = n5564 & n5651;
  assign n5822 = n5821 ^ n5570;
  assign n5823 = n5822 ^ n5819;
  assign n5824 = n5820 & n5823;
  assign n5825 = n5824 ^ x86;
  assign n5826 = n5825 ^ x87;
  assign n5827 = n5574 & n5651;
  assign n5828 = n5827 ^ n5576;
  assign n5829 = n5828 ^ n5825;
  assign n5830 = n5826 & ~n5829;
  assign n5831 = n5830 ^ x87;
  assign n5832 = n5831 ^ x88;
  assign n5833 = n5580 & n5651;
  assign n5834 = n5833 ^ n5582;
  assign n5835 = n5834 ^ n5831;
  assign n5836 = n5832 & n5835;
  assign n5837 = n5836 ^ x88;
  assign n5838 = n5837 ^ x89;
  assign n5839 = n5586 & n5651;
  assign n5840 = n5839 ^ n5588;
  assign n5841 = n5840 ^ n5837;
  assign n5842 = n5838 & ~n5841;
  assign n5843 = n5842 ^ x89;
  assign n5844 = n5663 & n5843;
  assign n5845 = n5661 ^ x91;
  assign n5846 = x90 & n5654;
  assign n5847 = n5846 ^ n5661;
  assign n5848 = ~n5845 & n5847;
  assign n5849 = n5848 ^ x91;
  assign n5850 = ~n5844 & ~n5849;
  assign n5851 = ~n5599 & n5651;
  assign n5852 = n5851 ^ n5601;
  assign n5853 = ~x92 & n5852;
  assign n5854 = n5605 & n5651;
  assign n5855 = n5854 ^ n5607;
  assign n5856 = ~x93 & n5855;
  assign n5857 = ~n5853 & ~n5856;
  assign n5858 = ~n5850 & n5857;
  assign n5859 = n5855 ^ x93;
  assign n5860 = x92 & ~n5852;
  assign n5861 = n5860 ^ n5855;
  assign n5862 = ~n5859 & n5861;
  assign n5863 = n5862 ^ x93;
  assign n5864 = ~n5858 & ~n5863;
  assign n5865 = n5864 ^ x94;
  assign n5866 = n5610 ^ x93;
  assign n5867 = n5651 & n5866;
  assign n5868 = n5867 ^ n5390;
  assign n5869 = n5868 ^ n5864;
  assign n5870 = ~n5865 & n5869;
  assign n5871 = n5870 ^ x94;
  assign n5872 = n5871 ^ x95;
  assign n5873 = ~n5391 & ~n5611;
  assign n5874 = n5873 ^ x94;
  assign n5875 = n5651 & n5874;
  assign n5876 = n5875 ^ n5387;
  assign n5877 = n5876 ^ n5871;
  assign n5878 = n5872 & ~n5877;
  assign n5879 = n5878 ^ x95;
  assign n5880 = n5879 ^ x96;
  assign n5881 = n5618 & n5651;
  assign n5882 = n5881 ^ n5620;
  assign n5883 = n5882 ^ n5879;
  assign n5884 = n5880 & ~n5883;
  assign n5885 = n5884 ^ x96;
  assign n5886 = n5885 ^ x97;
  assign n5887 = n5623 ^ x96;
  assign n5888 = n5651 & n5887;
  assign n5889 = n5888 ^ n5378;
  assign n5890 = n5889 ^ n5885;
  assign n5891 = n5886 & ~n5890;
  assign n5892 = n5891 ^ x97;
  assign n5893 = n5892 ^ x98;
  assign n5894 = n5623 ^ n5378;
  assign n5895 = n5887 & ~n5894;
  assign n5896 = n5895 ^ x96;
  assign n5897 = n5896 ^ x97;
  assign n5898 = n5651 & n5897;
  assign n5899 = n5898 ^ n5375;
  assign n5900 = n5899 ^ n5892;
  assign n5901 = n5893 & ~n5900;
  assign n5902 = n5901 ^ x98;
  assign n5903 = n5902 ^ x99;
  assign n5904 = ~n5631 & n5651;
  assign n5905 = n5904 ^ n5633;
  assign n5906 = n5905 ^ n5902;
  assign n5907 = n5903 & n5906;
  assign n5908 = n5907 ^ x99;
  assign n5909 = n5908 ^ x100;
  assign n5910 = n5637 & n5651;
  assign n5911 = n5910 ^ n5639;
  assign n5912 = n5911 ^ n5908;
  assign n5913 = n5909 & ~n5912;
  assign n5914 = n5913 ^ x100;
  assign n5915 = n5914 ^ x101;
  assign n5916 = n5642 ^ x100;
  assign n5917 = n5648 & n5916;
  assign n5918 = n5917 ^ n5370;
  assign n5919 = n5918 ^ n5914;
  assign n5920 = n5915 & n5919;
  assign n5921 = n5920 ^ x101;
  assign n5922 = n153 & ~n5921;
  assign n5923 = ~n154 & n5366;
  assign n5924 = ~n5922 & n5923;
  assign n5925 = ~n240 & n5648;
  assign n5926 = ~n5367 & ~n5925;
  assign n5927 = n5926 ^ x102;
  assign n5928 = n5921 ^ x102;
  assign n5929 = ~n5927 & n5928;
  assign n5930 = n5929 ^ x102;
  assign n5931 = n153 & ~n5930;
  assign n5932 = n5915 & n5931;
  assign n5933 = n5932 ^ n5918;
  assign n5934 = ~x102 & n5933;
  assign n5935 = ~n240 & ~n5924;
  assign n5936 = ~x103 & ~n5935;
  assign n5937 = ~n5934 & ~n5936;
  assign n5938 = n5886 & n5931;
  assign n5939 = n5938 ^ n5889;
  assign n5940 = n5939 ^ x98;
  assign n5941 = n5880 & n5931;
  assign n5942 = n5941 ^ n5882;
  assign n5943 = ~x97 & ~n5942;
  assign n5944 = n5719 & n5931;
  assign n5945 = n5944 ^ n5721;
  assign n5946 = ~x71 & n5945;
  assign n5947 = n5725 & n5931;
  assign n5948 = n5947 ^ n5727;
  assign n5949 = ~x72 & n5948;
  assign n5950 = ~n5946 & ~n5949;
  assign n5951 = x65 & ~n5651;
  assign n5952 = x25 & n5951;
  assign n5953 = n5931 & n5952;
  assign n5954 = n5683 & n5684;
  assign n5955 = ~n5953 & ~n5954;
  assign n5956 = n5651 ^ n1680;
  assign n5957 = n5687 ^ n5651;
  assign n5958 = n5651 ^ n202;
  assign n5959 = n5958 ^ n5651;
  assign n5960 = n5957 & ~n5959;
  assign n5961 = n5960 ^ n5651;
  assign n5962 = ~n5956 & n5961;
  assign n5963 = n5962 ^ n202;
  assign n5964 = n5963 ^ n5683;
  assign n5965 = n5931 & n5964;
  assign n5966 = n5965 ^ n5683;
  assign n5967 = n5955 & ~n5966;
  assign n5968 = n5967 ^ x26;
  assign n5969 = n5968 ^ x66;
  assign n5970 = x64 & n5931;
  assign n5971 = x24 & n5684;
  assign n5972 = n5971 ^ x25;
  assign n5973 = n5970 & n5972;
  assign n5974 = ~x24 & n5687;
  assign n5975 = ~n5691 & ~n5974;
  assign n5976 = ~n5931 & ~n5975;
  assign n5977 = ~x24 & x65;
  assign n5978 = n5977 ^ n5691;
  assign n5979 = x64 & n5978;
  assign n5980 = n5979 ^ n5691;
  assign n5981 = ~n5976 & ~n5980;
  assign n5982 = ~n5973 & n5981;
  assign n5983 = n5982 ^ n5968;
  assign n5984 = n5969 & n5983;
  assign n5985 = n5984 ^ x66;
  assign n5986 = n5985 ^ x67;
  assign n5987 = n5696 ^ x66;
  assign n5988 = n5931 & ~n5987;
  assign n5989 = n5988 ^ n5681;
  assign n5990 = n5989 ^ n5985;
  assign n5991 = n5986 & ~n5990;
  assign n5992 = n5991 ^ x67;
  assign n5993 = n5992 ^ x68;
  assign n5994 = n5700 & n5931;
  assign n5995 = n5994 ^ n5703;
  assign n5996 = n5995 ^ n5992;
  assign n5997 = n5993 & n5996;
  assign n5998 = n5997 ^ x68;
  assign n5999 = n5998 ^ x69;
  assign n6000 = n5707 & n5931;
  assign n6001 = n6000 ^ n5709;
  assign n6002 = n6001 ^ n5998;
  assign n6003 = n5999 & n6002;
  assign n6004 = n6003 ^ x69;
  assign n6005 = n6004 ^ x70;
  assign n6006 = n5713 & n5931;
  assign n6007 = n6006 ^ n5715;
  assign n6008 = n6007 ^ n6004;
  assign n6009 = n6005 & ~n6008;
  assign n6010 = n6009 ^ x70;
  assign n6011 = n5950 & n6010;
  assign n6012 = n5948 ^ x72;
  assign n6013 = x71 & ~n5945;
  assign n6014 = n6013 ^ n5948;
  assign n6015 = ~n6012 & n6014;
  assign n6016 = n6015 ^ x72;
  assign n6017 = ~n6011 & ~n6016;
  assign n6018 = n6017 ^ x73;
  assign n6019 = n5731 & n5931;
  assign n6020 = n6019 ^ n5733;
  assign n6021 = n6020 ^ n6017;
  assign n6022 = ~n6018 & n6021;
  assign n6023 = n6022 ^ x73;
  assign n6024 = n6023 ^ x74;
  assign n6025 = n5737 & n5931;
  assign n6026 = n6025 ^ n5739;
  assign n6027 = n6026 ^ n6023;
  assign n6028 = n6024 & n6027;
  assign n6029 = n6028 ^ x74;
  assign n6030 = n6029 ^ x75;
  assign n6031 = n5743 & n5931;
  assign n6032 = n6031 ^ n5745;
  assign n6033 = n6032 ^ n6029;
  assign n6034 = n6030 & n6033;
  assign n6035 = n6034 ^ x75;
  assign n6036 = n6035 ^ x76;
  assign n6037 = n5749 & n5931;
  assign n6038 = n6037 ^ n5751;
  assign n6039 = n6038 ^ n6035;
  assign n6040 = n6036 & n6039;
  assign n6041 = n6040 ^ x76;
  assign n6042 = n6041 ^ x77;
  assign n6043 = n5755 & n5931;
  assign n6044 = n6043 ^ n5757;
  assign n6045 = n6044 ^ n6041;
  assign n6046 = n6042 & ~n6045;
  assign n6047 = n6046 ^ x77;
  assign n6048 = n6047 ^ x78;
  assign n6049 = n5761 & n5931;
  assign n6050 = n6049 ^ n5763;
  assign n6051 = n6050 ^ n6047;
  assign n6052 = n6048 & n6051;
  assign n6053 = n6052 ^ x78;
  assign n6054 = n6053 ^ x79;
  assign n6055 = n5767 & n5931;
  assign n6056 = n6055 ^ n5770;
  assign n6057 = n6056 ^ n6053;
  assign n6058 = n6054 & ~n6057;
  assign n6059 = n6058 ^ x79;
  assign n6060 = n6059 ^ x80;
  assign n6061 = n5774 & n5931;
  assign n6062 = n6061 ^ n5780;
  assign n6063 = n6062 ^ n6059;
  assign n6064 = n6060 & ~n6063;
  assign n6065 = n6064 ^ x80;
  assign n6066 = n6065 ^ x81;
  assign n6067 = n5784 & n5931;
  assign n6068 = n6067 ^ n5786;
  assign n6069 = n6068 ^ n6065;
  assign n6070 = n6066 & ~n6069;
  assign n6071 = n6070 ^ x81;
  assign n6072 = n6071 ^ x82;
  assign n6073 = n5790 & n5931;
  assign n6074 = n6073 ^ n5792;
  assign n6075 = n6074 ^ n6071;
  assign n6076 = n6072 & ~n6075;
  assign n6077 = n6076 ^ x82;
  assign n6078 = n6077 ^ x83;
  assign n6079 = n5796 & n5931;
  assign n6080 = n6079 ^ n5798;
  assign n6081 = n6080 ^ n6077;
  assign n6082 = n6078 & ~n6081;
  assign n6083 = n6082 ^ x83;
  assign n6084 = n6083 ^ x84;
  assign n6085 = n5802 & n5931;
  assign n6086 = n6085 ^ n5804;
  assign n6087 = n6086 ^ n6083;
  assign n6088 = n6084 & ~n6087;
  assign n6089 = n6088 ^ x84;
  assign n6090 = n6089 ^ x85;
  assign n6091 = n5808 & n5931;
  assign n6092 = n6091 ^ n5810;
  assign n6093 = n6092 ^ n6089;
  assign n6094 = n6090 & ~n6093;
  assign n6095 = n6094 ^ x85;
  assign n6096 = n6095 ^ x86;
  assign n6097 = n5814 & n5931;
  assign n6098 = n6097 ^ n5816;
  assign n6099 = n6098 ^ n6095;
  assign n6100 = n6096 & ~n6099;
  assign n6101 = n6100 ^ x86;
  assign n6102 = n6101 ^ x87;
  assign n6103 = n5820 & n5931;
  assign n6104 = n6103 ^ n5822;
  assign n6105 = n6104 ^ n6101;
  assign n6106 = n6102 & n6105;
  assign n6107 = n6106 ^ x87;
  assign n6108 = n6107 ^ x88;
  assign n6109 = n5826 & n5931;
  assign n6110 = n6109 ^ n5828;
  assign n6111 = n6110 ^ n6107;
  assign n6112 = n6108 & ~n6111;
  assign n6113 = n6112 ^ x88;
  assign n6114 = n6113 ^ x89;
  assign n6115 = n5832 & n5931;
  assign n6116 = n6115 ^ n5834;
  assign n6117 = n6116 ^ n6113;
  assign n6118 = n6114 & n6117;
  assign n6119 = n6118 ^ x89;
  assign n6120 = n6119 ^ x90;
  assign n6121 = n5838 & n5931;
  assign n6122 = n6121 ^ n5840;
  assign n6123 = n6122 ^ n6119;
  assign n6124 = n6120 & ~n6123;
  assign n6125 = n6124 ^ x90;
  assign n6126 = n6125 ^ x91;
  assign n6127 = n5843 ^ x90;
  assign n6128 = n5931 & n6127;
  assign n6129 = n6128 ^ n5654;
  assign n6130 = n6129 ^ n6125;
  assign n6131 = n6126 & ~n6130;
  assign n6132 = n6131 ^ x91;
  assign n6133 = n6132 ^ x92;
  assign n6134 = n5843 ^ n5654;
  assign n6135 = n6127 & ~n6134;
  assign n6136 = n6135 ^ x90;
  assign n6137 = n6136 ^ x91;
  assign n6138 = n5931 & n6137;
  assign n6139 = n6138 ^ n5661;
  assign n6140 = n6139 ^ n6132;
  assign n6141 = n6133 & n6140;
  assign n6142 = n6141 ^ x92;
  assign n6143 = n6142 ^ x93;
  assign n6144 = n5850 ^ x92;
  assign n6145 = n5931 & ~n6144;
  assign n6146 = n6145 ^ n5852;
  assign n6147 = n6146 ^ n6142;
  assign n6148 = n6143 & n6147;
  assign n6149 = n6148 ^ x93;
  assign n6150 = n6149 ^ x94;
  assign n6151 = n5852 ^ n5850;
  assign n6152 = ~n6144 & ~n6151;
  assign n6153 = n6152 ^ x92;
  assign n6154 = n6153 ^ x93;
  assign n6155 = n5931 & n6154;
  assign n6156 = n6155 ^ n5855;
  assign n6157 = n6156 ^ n6149;
  assign n6158 = n6150 & n6157;
  assign n6159 = n6158 ^ x94;
  assign n6160 = n6159 ^ x95;
  assign n6161 = ~n5865 & n5931;
  assign n6162 = n6161 ^ n5868;
  assign n6163 = n6162 ^ n6159;
  assign n6164 = n6160 & ~n6163;
  assign n6165 = n6164 ^ x95;
  assign n6166 = n6165 ^ x96;
  assign n6167 = n5872 & n5931;
  assign n6168 = n6167 ^ n5876;
  assign n6169 = n6168 ^ n6165;
  assign n6170 = n6166 & ~n6169;
  assign n6171 = n6170 ^ x96;
  assign n6172 = ~n5943 & n6171;
  assign n6173 = n6172 ^ n5939;
  assign n6174 = n6173 ^ n5939;
  assign n6175 = x97 & n5942;
  assign n6176 = n6175 ^ n5939;
  assign n6177 = n6176 ^ n5939;
  assign n6178 = ~n6174 & ~n6177;
  assign n6179 = n6178 ^ n5939;
  assign n6180 = n5940 & n6179;
  assign n6181 = n6180 ^ x98;
  assign n6182 = n6181 ^ x99;
  assign n6183 = n5893 & n5931;
  assign n6184 = n6183 ^ n5899;
  assign n6185 = n6184 ^ n6181;
  assign n6186 = n6182 & ~n6185;
  assign n6187 = n6186 ^ x99;
  assign n6188 = n6187 ^ x100;
  assign n6189 = n5903 & n5931;
  assign n6190 = n6189 ^ n5905;
  assign n6191 = n6190 ^ n6187;
  assign n6192 = n6188 & n6191;
  assign n6193 = n6192 ^ x100;
  assign n6194 = n6193 ^ x101;
  assign n6195 = n5909 & n5931;
  assign n6196 = n6195 ^ n5911;
  assign n6197 = n6196 ^ n6193;
  assign n6198 = n6194 & ~n6197;
  assign n6199 = n6198 ^ x101;
  assign n6200 = n5937 & n6199;
  assign n6201 = x102 & ~n5936;
  assign n6202 = ~n5933 & n6201;
  assign n6203 = n152 & ~n5367;
  assign n6204 = ~n153 & ~n6203;
  assign n6205 = ~n6202 & ~n6204;
  assign n6206 = ~n6200 & n6205;
  assign n6207 = n5924 & ~n6206;
  assign n6208 = ~x108 & n147;
  assign n6209 = n150 & n6208;
  assign n6210 = ~x105 & n6209;
  assign n6211 = ~n240 & ~n6207;
  assign n6212 = n6211 ^ x104;
  assign n6213 = n6199 ^ x102;
  assign n6214 = n6206 & n6213;
  assign n6215 = n6214 ^ n5933;
  assign n6216 = x103 & ~n6215;
  assign n6217 = n6216 ^ n6211;
  assign n6218 = n6217 ^ n6211;
  assign n6219 = n6194 & n6206;
  assign n6220 = n6219 ^ n6196;
  assign n6221 = x102 & n6220;
  assign n6222 = n6166 & n6206;
  assign n6223 = n6222 ^ n6168;
  assign n6224 = n6223 ^ x97;
  assign n6225 = n6160 & n6206;
  assign n6226 = n6225 ^ n6162;
  assign n6227 = x96 & n6226;
  assign n6228 = n6227 ^ n6223;
  assign n6229 = n6228 ^ n6223;
  assign n6230 = ~x96 & ~n6226;
  assign n6231 = n6126 & n6206;
  assign n6232 = n6231 ^ n6129;
  assign n6233 = ~x92 & ~n6232;
  assign n6234 = n6133 & n6206;
  assign n6235 = n6234 ^ n6139;
  assign n6236 = ~x93 & n6235;
  assign n6237 = ~n6233 & ~n6236;
  assign n6238 = n6090 & n6206;
  assign n6239 = n6238 ^ n6092;
  assign n6240 = ~x86 & ~n6239;
  assign n6241 = n6096 & n6206;
  assign n6242 = n6241 ^ n6098;
  assign n6243 = ~x87 & ~n6242;
  assign n6244 = ~n6240 & ~n6243;
  assign n6245 = x65 & n5931;
  assign n6246 = n6245 ^ x24;
  assign n6247 = n6246 ^ n6245;
  assign n6248 = n289 & ~n5931;
  assign n6249 = n6248 ^ x65;
  assign n6250 = n6249 ^ n6245;
  assign n6251 = ~n6247 & ~n6250;
  assign n6252 = n6251 ^ n6245;
  assign n6253 = ~n202 & n6252;
  assign n6254 = n6253 ^ n5970;
  assign n6255 = ~x24 & n6249;
  assign n6256 = ~x65 & ~n6255;
  assign n6257 = n6256 ^ n6253;
  assign n6258 = n6253 ^ n6206;
  assign n6259 = ~n6253 & ~n6258;
  assign n6260 = n6259 ^ n6253;
  assign n6261 = ~n6257 & ~n6260;
  assign n6262 = n6261 ^ n6259;
  assign n6263 = n6262 ^ n6253;
  assign n6264 = n6263 ^ n6206;
  assign n6265 = ~n6254 & ~n6264;
  assign n6266 = n6265 ^ n5970;
  assign n6267 = n6266 ^ x25;
  assign n6268 = n6267 ^ x66;
  assign n6269 = x64 & n6206;
  assign n6270 = x24 & ~x65;
  assign n6271 = x23 & n6270;
  assign n6272 = n6271 ^ x24;
  assign n6273 = n6269 & n6272;
  assign n6275 = x65 ^ x24;
  assign n6282 = n6275 ^ x65;
  assign n6274 = x65 ^ x23;
  assign n6276 = n6275 ^ n6274;
  assign n6277 = n6276 ^ x65;
  assign n6278 = n6274 ^ x64;
  assign n6279 = n6278 ^ n6274;
  assign n6280 = n6279 ^ n6277;
  assign n6281 = ~n6277 & ~n6280;
  assign n6283 = n6282 ^ n6281;
  assign n6284 = n6283 ^ n6277;
  assign n6285 = n6206 ^ x65;
  assign n6286 = n6285 ^ x65;
  assign n6287 = n6281 ^ n6277;
  assign n6288 = ~n6286 & ~n6287;
  assign n6289 = n6288 ^ x65;
  assign n6290 = ~n6284 & n6289;
  assign n6291 = n6290 ^ x65;
  assign n6292 = n6291 ^ x65;
  assign n6293 = n6292 ^ x65;
  assign n6294 = ~n6273 & ~n6293;
  assign n6295 = n6294 ^ n6267;
  assign n6296 = ~n6268 & ~n6295;
  assign n6297 = n6296 ^ x66;
  assign n6298 = n6297 ^ x67;
  assign n6299 = n5982 ^ x66;
  assign n6300 = n6206 & ~n6299;
  assign n6301 = n6300 ^ n5968;
  assign n6302 = n6301 ^ n6297;
  assign n6303 = n6298 & ~n6302;
  assign n6304 = n6303 ^ x67;
  assign n6305 = n6304 ^ x68;
  assign n6306 = n5986 & n6206;
  assign n6307 = n6306 ^ n5989;
  assign n6308 = n6307 ^ n6304;
  assign n6309 = n6305 & ~n6308;
  assign n6310 = n6309 ^ x68;
  assign n6311 = n6310 ^ x69;
  assign n6312 = n5993 & n6206;
  assign n6313 = n6312 ^ n5995;
  assign n6314 = n6313 ^ n6310;
  assign n6315 = n6311 & n6314;
  assign n6316 = n6315 ^ x69;
  assign n6317 = n6316 ^ x70;
  assign n6318 = n5999 & n6206;
  assign n6319 = n6318 ^ n6001;
  assign n6320 = n6319 ^ n6316;
  assign n6321 = n6317 & n6320;
  assign n6322 = n6321 ^ x70;
  assign n6323 = n6322 ^ x71;
  assign n6324 = n6005 & n6206;
  assign n6325 = n6324 ^ n6007;
  assign n6326 = n6325 ^ n6322;
  assign n6327 = n6323 & ~n6326;
  assign n6328 = n6327 ^ x71;
  assign n6329 = n6328 ^ x72;
  assign n6330 = n6010 ^ x71;
  assign n6331 = n6206 & n6330;
  assign n6332 = n6331 ^ n5945;
  assign n6333 = n6332 ^ n6328;
  assign n6334 = n6329 & n6333;
  assign n6335 = n6334 ^ x72;
  assign n6336 = n6335 ^ x73;
  assign n6337 = n6010 ^ n5945;
  assign n6338 = n6330 & n6337;
  assign n6339 = n6338 ^ x71;
  assign n6340 = n6339 ^ x72;
  assign n6341 = n6206 & n6340;
  assign n6342 = n6341 ^ n5948;
  assign n6343 = n6342 ^ n6335;
  assign n6344 = n6336 & n6343;
  assign n6345 = n6344 ^ x73;
  assign n6346 = n6345 ^ x74;
  assign n6347 = ~n6018 & n6206;
  assign n6348 = n6347 ^ n6020;
  assign n6349 = n6348 ^ n6345;
  assign n6350 = n6346 & ~n6349;
  assign n6351 = n6350 ^ x74;
  assign n6352 = n6351 ^ x75;
  assign n6353 = n6024 & n6206;
  assign n6354 = n6353 ^ n6026;
  assign n6355 = n6354 ^ n6351;
  assign n6356 = n6352 & n6355;
  assign n6357 = n6356 ^ x75;
  assign n6358 = n6357 ^ x76;
  assign n6359 = n6030 & n6206;
  assign n6360 = n6359 ^ n6032;
  assign n6361 = n6360 ^ n6357;
  assign n6362 = n6358 & n6361;
  assign n6363 = n6362 ^ x76;
  assign n6364 = n6363 ^ x77;
  assign n6365 = n6036 & n6206;
  assign n6366 = n6365 ^ n6038;
  assign n6367 = n6366 ^ n6363;
  assign n6368 = n6364 & n6367;
  assign n6369 = n6368 ^ x77;
  assign n6370 = n6369 ^ x78;
  assign n6371 = n6042 & n6206;
  assign n6372 = n6371 ^ n6044;
  assign n6373 = n6372 ^ n6369;
  assign n6374 = n6370 & ~n6373;
  assign n6375 = n6374 ^ x78;
  assign n6376 = n6375 ^ x79;
  assign n6377 = n6048 & n6206;
  assign n6378 = n6377 ^ n6050;
  assign n6379 = n6378 ^ n6375;
  assign n6380 = n6376 & n6379;
  assign n6381 = n6380 ^ x79;
  assign n6382 = n6381 ^ x80;
  assign n6383 = n6054 & n6206;
  assign n6384 = n6383 ^ n6056;
  assign n6385 = n6384 ^ n6381;
  assign n6386 = n6382 & ~n6385;
  assign n6387 = n6386 ^ x80;
  assign n6388 = n6387 ^ x81;
  assign n6389 = n6060 & n6206;
  assign n6390 = n6389 ^ n6062;
  assign n6391 = n6390 ^ n6387;
  assign n6392 = n6388 & ~n6391;
  assign n6393 = n6392 ^ x81;
  assign n6394 = n6393 ^ x82;
  assign n6395 = n6066 & n6206;
  assign n6396 = n6395 ^ n6068;
  assign n6397 = n6396 ^ n6393;
  assign n6398 = n6394 & ~n6397;
  assign n6399 = n6398 ^ x82;
  assign n6400 = n6399 ^ x83;
  assign n6401 = n6072 & n6206;
  assign n6402 = n6401 ^ n6074;
  assign n6403 = n6402 ^ n6399;
  assign n6404 = n6400 & ~n6403;
  assign n6405 = n6404 ^ x83;
  assign n6406 = n6405 ^ x84;
  assign n6407 = n6078 & n6206;
  assign n6408 = n6407 ^ n6080;
  assign n6409 = n6408 ^ n6405;
  assign n6410 = n6406 & ~n6409;
  assign n6411 = n6410 ^ x84;
  assign n6412 = n6411 ^ x85;
  assign n6413 = n6084 & n6206;
  assign n6414 = n6413 ^ n6086;
  assign n6415 = n6414 ^ n6411;
  assign n6416 = n6412 & ~n6415;
  assign n6417 = n6416 ^ x85;
  assign n6418 = n6244 & n6417;
  assign n6419 = n6242 ^ x87;
  assign n6420 = x86 & n6239;
  assign n6421 = n6420 ^ n6242;
  assign n6422 = n6419 & ~n6421;
  assign n6423 = n6422 ^ x87;
  assign n6424 = ~n6418 & ~n6423;
  assign n6425 = n6102 & n6206;
  assign n6426 = n6425 ^ n6104;
  assign n6427 = ~x88 & n6426;
  assign n6428 = n6108 & n6206;
  assign n6429 = n6428 ^ n6110;
  assign n6430 = ~x89 & ~n6429;
  assign n6431 = ~n6427 & ~n6430;
  assign n6432 = ~n6424 & n6431;
  assign n6433 = n6429 ^ x89;
  assign n6434 = x88 & ~n6426;
  assign n6435 = n6434 ^ n6429;
  assign n6436 = n6433 & ~n6435;
  assign n6437 = n6436 ^ x89;
  assign n6438 = ~n6432 & ~n6437;
  assign n6439 = n6438 ^ x90;
  assign n6440 = n6114 & n6206;
  assign n6441 = n6440 ^ n6116;
  assign n6442 = n6441 ^ n6438;
  assign n6443 = ~n6439 & ~n6442;
  assign n6444 = n6443 ^ x90;
  assign n6445 = n6444 ^ x91;
  assign n6446 = n6120 & n6206;
  assign n6447 = n6446 ^ n6122;
  assign n6448 = n6447 ^ n6444;
  assign n6449 = n6445 & ~n6448;
  assign n6450 = n6449 ^ x91;
  assign n6451 = n6237 & n6450;
  assign n6452 = n6235 ^ x93;
  assign n6453 = x92 & n6232;
  assign n6454 = n6453 ^ n6235;
  assign n6455 = ~n6452 & n6454;
  assign n6456 = n6455 ^ x93;
  assign n6457 = ~n6451 & ~n6456;
  assign n6458 = n6457 ^ x94;
  assign n6459 = n6143 & n6206;
  assign n6460 = n6459 ^ n6146;
  assign n6461 = n6460 ^ n6457;
  assign n6462 = ~n6458 & ~n6461;
  assign n6463 = n6462 ^ x94;
  assign n6464 = n6463 ^ x95;
  assign n6465 = n6150 & n6206;
  assign n6466 = n6465 ^ n6156;
  assign n6467 = n6466 ^ n6463;
  assign n6468 = n6464 & n6467;
  assign n6469 = n6468 ^ x95;
  assign n6470 = ~n6230 & n6469;
  assign n6471 = n6470 ^ n6223;
  assign n6472 = n6471 ^ n6223;
  assign n6473 = ~n6229 & ~n6472;
  assign n6474 = n6473 ^ n6223;
  assign n6475 = n6224 & n6474;
  assign n6476 = n6475 ^ x97;
  assign n6477 = n6476 ^ x98;
  assign n6478 = n6171 ^ x97;
  assign n6479 = n6206 & n6478;
  assign n6480 = n6479 ^ n5942;
  assign n6481 = n6480 ^ n6476;
  assign n6482 = n6477 & ~n6481;
  assign n6483 = n6482 ^ x98;
  assign n6484 = n6483 ^ x99;
  assign n6485 = ~n6172 & ~n6175;
  assign n6486 = n6485 ^ x98;
  assign n6487 = n6206 & ~n6486;
  assign n6488 = n6487 ^ n5939;
  assign n6489 = n6488 ^ n6483;
  assign n6490 = n6484 & ~n6489;
  assign n6491 = n6490 ^ x99;
  assign n6492 = n6491 ^ x100;
  assign n6493 = n6182 & n6206;
  assign n6494 = n6493 ^ n6184;
  assign n6495 = n6494 ^ n6491;
  assign n6496 = n6492 & ~n6495;
  assign n6497 = n6496 ^ x100;
  assign n6498 = n6497 ^ x101;
  assign n6499 = n6188 & n6206;
  assign n6500 = n6499 ^ n6190;
  assign n6501 = n6500 ^ n6497;
  assign n6502 = n6498 & n6501;
  assign n6503 = n6502 ^ x101;
  assign n6504 = ~n6221 & ~n6503;
  assign n6505 = ~x102 & ~n6220;
  assign n6506 = ~x103 & n6215;
  assign n6507 = ~n6505 & ~n6506;
  assign n6508 = ~n6504 & n6507;
  assign n6509 = n6508 ^ n6211;
  assign n6510 = n6509 ^ n6211;
  assign n6511 = ~n6218 & ~n6510;
  assign n6512 = n6511 ^ n6211;
  assign n6513 = n6212 & n6512;
  assign n6514 = n6513 ^ x104;
  assign n6515 = n6210 & ~n6514;
  assign n6516 = n6207 & ~n6515;
  assign n6517 = ~n240 & ~n6516;
  assign n6518 = ~x107 & n6208;
  assign n6519 = n6317 & n6515;
  assign n6520 = n6519 ^ n6319;
  assign n6521 = ~x71 & n6520;
  assign n6522 = n6323 & n6515;
  assign n6523 = n6522 ^ n6325;
  assign n6524 = ~x72 & ~n6523;
  assign n6525 = ~n6521 & ~n6524;
  assign n6526 = n6206 ^ x64;
  assign n6527 = n6526 ^ x64;
  assign n6528 = n6515 ^ x64;
  assign n6529 = ~n6527 & n6528;
  assign n6530 = n6529 ^ x64;
  assign n6531 = n6285 & n6530;
  assign n6532 = x23 & n6531;
  assign n6533 = ~x65 & n6206;
  assign n6534 = ~x23 & x64;
  assign n6535 = x65 & ~n6206;
  assign n6536 = n6534 & ~n6535;
  assign n6537 = ~n202 & ~n6536;
  assign n6538 = ~n6533 & ~n6537;
  assign n6539 = n6538 ^ n6269;
  assign n6540 = n6515 & n6539;
  assign n6541 = n6540 ^ n6269;
  assign n6542 = ~n6532 & ~n6541;
  assign n6543 = n6542 ^ x24;
  assign n6544 = n6543 ^ x66;
  assign n6545 = x64 & n6515;
  assign n6546 = n6545 ^ x23;
  assign n6547 = n6546 ^ x65;
  assign n6548 = ~x22 & x64;
  assign n6549 = n6548 ^ n6546;
  assign n6550 = ~n6547 & n6549;
  assign n6551 = n6550 ^ x65;
  assign n6552 = n6551 ^ n6543;
  assign n6553 = n6544 & ~n6552;
  assign n6554 = n6553 ^ x66;
  assign n6555 = n6554 ^ x67;
  assign n6556 = n6294 ^ x66;
  assign n6557 = n6515 & ~n6556;
  assign n6558 = n6557 ^ n6267;
  assign n6559 = n6558 ^ n6554;
  assign n6560 = n6555 & n6559;
  assign n6561 = n6560 ^ x67;
  assign n6562 = n6561 ^ x68;
  assign n6563 = n6298 & n6515;
  assign n6564 = n6563 ^ n6301;
  assign n6565 = n6564 ^ n6561;
  assign n6566 = n6562 & ~n6565;
  assign n6567 = n6566 ^ x68;
  assign n6568 = n6567 ^ x69;
  assign n6569 = n6305 & n6515;
  assign n6570 = n6569 ^ n6307;
  assign n6571 = n6570 ^ n6567;
  assign n6572 = n6568 & ~n6571;
  assign n6573 = n6572 ^ x69;
  assign n6574 = n6573 ^ x70;
  assign n6575 = n6311 & n6515;
  assign n6576 = n6575 ^ n6313;
  assign n6577 = n6576 ^ n6573;
  assign n6578 = n6574 & n6577;
  assign n6579 = n6578 ^ x70;
  assign n6580 = n6525 & n6579;
  assign n6581 = n6523 ^ x72;
  assign n6582 = x71 & ~n6520;
  assign n6583 = n6582 ^ n6523;
  assign n6584 = n6581 & ~n6583;
  assign n6585 = n6584 ^ x72;
  assign n6586 = ~n6580 & ~n6585;
  assign n6587 = n6586 ^ x73;
  assign n6588 = n6329 & n6515;
  assign n6589 = n6588 ^ n6332;
  assign n6590 = n6589 ^ n6586;
  assign n6591 = ~n6587 & ~n6590;
  assign n6592 = n6591 ^ x73;
  assign n6593 = n6592 ^ x74;
  assign n6594 = n6336 & n6515;
  assign n6595 = n6594 ^ n6342;
  assign n6596 = n6595 ^ n6592;
  assign n6597 = n6593 & n6596;
  assign n6598 = n6597 ^ x74;
  assign n6599 = n6598 ^ x75;
  assign n6600 = n6346 & n6515;
  assign n6601 = n6600 ^ n6348;
  assign n6602 = n6601 ^ n6598;
  assign n6603 = n6599 & ~n6602;
  assign n6604 = n6603 ^ x75;
  assign n6605 = n6604 ^ x76;
  assign n6606 = n6352 & n6515;
  assign n6607 = n6606 ^ n6354;
  assign n6608 = n6607 ^ n6604;
  assign n6609 = n6605 & n6608;
  assign n6610 = n6609 ^ x76;
  assign n6611 = n6610 ^ x77;
  assign n6612 = n6358 & n6515;
  assign n6613 = n6612 ^ n6360;
  assign n6614 = n6613 ^ n6610;
  assign n6615 = n6611 & n6614;
  assign n6616 = n6615 ^ x77;
  assign n6617 = n6616 ^ x78;
  assign n6618 = n6364 & n6515;
  assign n6619 = n6618 ^ n6366;
  assign n6620 = n6619 ^ n6616;
  assign n6621 = n6617 & n6620;
  assign n6622 = n6621 ^ x78;
  assign n6623 = n6622 ^ x79;
  assign n6624 = n6370 & n6515;
  assign n6625 = n6624 ^ n6372;
  assign n6626 = n6625 ^ n6622;
  assign n6627 = n6623 & ~n6626;
  assign n6628 = n6627 ^ x79;
  assign n6629 = n6628 ^ x80;
  assign n6630 = n6376 & n6515;
  assign n6631 = n6630 ^ n6378;
  assign n6632 = n6631 ^ n6628;
  assign n6633 = n6629 & n6632;
  assign n6634 = n6633 ^ x80;
  assign n6635 = n6634 ^ x81;
  assign n6636 = n6382 & n6515;
  assign n6637 = n6636 ^ n6384;
  assign n6638 = n6637 ^ n6634;
  assign n6639 = n6635 & ~n6638;
  assign n6640 = n6639 ^ x81;
  assign n6641 = n6640 ^ x82;
  assign n6642 = n6388 & n6515;
  assign n6643 = n6642 ^ n6390;
  assign n6644 = n6643 ^ n6640;
  assign n6645 = n6641 & ~n6644;
  assign n6646 = n6645 ^ x82;
  assign n6647 = n6646 ^ x83;
  assign n6648 = n6394 & n6515;
  assign n6649 = n6648 ^ n6396;
  assign n6650 = n6649 ^ n6646;
  assign n6651 = n6647 & ~n6650;
  assign n6652 = n6651 ^ x83;
  assign n6653 = n6652 ^ x84;
  assign n6654 = n6400 & n6515;
  assign n6655 = n6654 ^ n6402;
  assign n6656 = n6655 ^ n6652;
  assign n6657 = n6653 & ~n6656;
  assign n6658 = n6657 ^ x84;
  assign n6659 = n6658 ^ x85;
  assign n6660 = n6406 & n6515;
  assign n6661 = n6660 ^ n6408;
  assign n6662 = n6661 ^ n6658;
  assign n6663 = n6659 & ~n6662;
  assign n6664 = n6663 ^ x85;
  assign n6665 = n6664 ^ x86;
  assign n6666 = n6412 & n6515;
  assign n6667 = n6666 ^ n6414;
  assign n6668 = n6667 ^ n6664;
  assign n6669 = n6665 & ~n6668;
  assign n6670 = n6669 ^ x86;
  assign n6671 = n6670 ^ x87;
  assign n6672 = n6417 ^ x86;
  assign n6673 = n6515 & n6672;
  assign n6674 = n6673 ^ n6239;
  assign n6675 = n6674 ^ n6670;
  assign n6676 = n6671 & ~n6675;
  assign n6677 = n6676 ^ x87;
  assign n6678 = n6677 ^ x88;
  assign n6679 = n6417 ^ n6239;
  assign n6680 = n6672 & ~n6679;
  assign n6681 = n6680 ^ x86;
  assign n6682 = n6681 ^ x87;
  assign n6683 = n6515 & n6682;
  assign n6684 = n6683 ^ n6242;
  assign n6685 = n6684 ^ n6677;
  assign n6686 = n6678 & ~n6685;
  assign n6687 = n6686 ^ x88;
  assign n6688 = n6687 ^ x89;
  assign n6689 = n6424 ^ x88;
  assign n6690 = n6515 & ~n6689;
  assign n6691 = n6690 ^ n6426;
  assign n6692 = n6691 ^ n6687;
  assign n6693 = n6688 & n6692;
  assign n6694 = n6693 ^ x89;
  assign n6695 = n6694 ^ x90;
  assign n6696 = n6426 ^ n6424;
  assign n6697 = ~n6689 & ~n6696;
  assign n6698 = n6697 ^ x88;
  assign n6699 = n6698 ^ x89;
  assign n6700 = n6515 & n6699;
  assign n6701 = n6700 ^ n6429;
  assign n6702 = n6701 ^ n6694;
  assign n6703 = n6695 & ~n6702;
  assign n6704 = n6703 ^ x90;
  assign n6705 = n6704 ^ x91;
  assign n6706 = ~n6439 & n6515;
  assign n6707 = n6706 ^ n6441;
  assign n6708 = n6707 ^ n6704;
  assign n6709 = n6705 & n6708;
  assign n6710 = n6709 ^ x91;
  assign n6711 = n6710 ^ x92;
  assign n6712 = n6445 & n6515;
  assign n6713 = n6712 ^ n6447;
  assign n6714 = n6713 ^ n6710;
  assign n6715 = n6711 & ~n6714;
  assign n6716 = n6715 ^ x92;
  assign n6717 = n6716 ^ x93;
  assign n6718 = n6450 ^ x92;
  assign n6719 = n6515 & n6718;
  assign n6720 = n6719 ^ n6232;
  assign n6721 = n6720 ^ n6716;
  assign n6722 = n6717 & ~n6721;
  assign n6723 = n6722 ^ x93;
  assign n6724 = n6723 ^ x94;
  assign n6725 = n6450 ^ n6232;
  assign n6726 = n6718 & ~n6725;
  assign n6727 = n6726 ^ x92;
  assign n6728 = n6727 ^ x93;
  assign n6729 = n6515 & n6728;
  assign n6730 = n6729 ^ n6235;
  assign n6731 = n6730 ^ n6723;
  assign n6732 = n6724 & n6731;
  assign n6733 = n6732 ^ x94;
  assign n6734 = n6733 ^ x95;
  assign n6735 = ~n6458 & n6515;
  assign n6736 = n6735 ^ n6460;
  assign n6737 = n6736 ^ n6733;
  assign n6738 = n6734 & n6737;
  assign n6739 = n6738 ^ x95;
  assign n6740 = n6739 ^ x96;
  assign n6741 = n6464 & n6515;
  assign n6742 = n6741 ^ n6466;
  assign n6743 = n6742 ^ n6739;
  assign n6744 = n6740 & n6743;
  assign n6745 = n6744 ^ x96;
  assign n6746 = n6745 ^ x97;
  assign n6747 = n6469 ^ x96;
  assign n6748 = n6515 & n6747;
  assign n6749 = n6748 ^ n6226;
  assign n6750 = n6749 ^ n6745;
  assign n6751 = n6746 & ~n6750;
  assign n6752 = n6751 ^ x97;
  assign n6753 = n6752 ^ x98;
  assign n6754 = x98 & n6752;
  assign n6755 = ~n6227 & ~n6470;
  assign n6756 = n6755 ^ x97;
  assign n6757 = n6515 & ~n6756;
  assign n6758 = n6757 ^ n6223;
  assign n6759 = x98 & n6758;
  assign n6760 = ~x99 & ~n6759;
  assign n6761 = ~n6754 & n6760;
  assign n6762 = n6477 & n6515;
  assign n6763 = n6762 ^ n6480;
  assign n6764 = ~n6761 & n6763;
  assign n6765 = x98 & x99;
  assign n6766 = n6765 ^ n6758;
  assign n6767 = ~x99 & ~n6763;
  assign n6768 = n6767 ^ n6765;
  assign n6769 = n6758 ^ n6752;
  assign n6770 = n6769 ^ n6767;
  assign n6771 = n6767 & ~n6770;
  assign n6772 = n6771 ^ n6767;
  assign n6773 = ~n6768 & n6772;
  assign n6774 = n6773 ^ n6771;
  assign n6775 = n6774 ^ n6767;
  assign n6776 = n6775 ^ n6769;
  assign n6777 = n6766 & ~n6776;
  assign n6778 = n6777 ^ n6765;
  assign n6779 = ~n6764 & ~n6778;
  assign n6780 = n6779 ^ x100;
  assign n6781 = n6484 & n6515;
  assign n6782 = n6781 ^ n6488;
  assign n6783 = n6782 ^ n6779;
  assign n6784 = ~n6780 & n6783;
  assign n6785 = n6784 ^ x100;
  assign n6786 = n6785 ^ x101;
  assign n6787 = n6492 & n6515;
  assign n6788 = n6787 ^ n6494;
  assign n6789 = n6788 ^ n6785;
  assign n6790 = n6786 & ~n6789;
  assign n6791 = n6790 ^ x101;
  assign n6792 = n6791 ^ x102;
  assign n6793 = n6498 & n6515;
  assign n6794 = n6793 ^ n6500;
  assign n6795 = n6794 ^ n6791;
  assign n6796 = n6792 & n6795;
  assign n6797 = n6796 ^ x102;
  assign n6798 = n6797 ^ x103;
  assign n6799 = n6503 ^ x102;
  assign n6800 = n6515 & n6799;
  assign n6801 = n6800 ^ n6220;
  assign n6802 = n6801 ^ n6797;
  assign n6803 = n6798 & ~n6802;
  assign n6804 = n6803 ^ x103;
  assign n6805 = n6804 ^ x104;
  assign n6806 = ~n6504 & ~n6505;
  assign n6807 = n6806 ^ x103;
  assign n6808 = n6515 & n6807;
  assign n6809 = n6808 ^ n6215;
  assign n6810 = n6809 ^ n6804;
  assign n6811 = n6805 & n6810;
  assign n6812 = n6811 ^ x104;
  assign n6813 = n6812 ^ x105;
  assign n6814 = n6517 ^ x105;
  assign n6815 = n6813 & n6814;
  assign n6816 = n6815 ^ x105;
  assign n6817 = n6209 & ~n6816;
  assign n6818 = n6753 & n6817;
  assign n6819 = n6818 ^ n6758;
  assign n6820 = x99 & n6819;
  assign n6821 = n6753 & ~n6769;
  assign n6822 = n6821 ^ x98;
  assign n6823 = n6822 ^ x99;
  assign n6824 = n6817 & n6823;
  assign n6825 = n6824 ^ n6763;
  assign n6826 = x100 & n6825;
  assign n6827 = ~n6820 & ~n6826;
  assign n6828 = n6705 & n6817;
  assign n6829 = n6828 ^ n6707;
  assign n6830 = ~x92 & n6829;
  assign n6831 = n6711 & n6817;
  assign n6832 = n6831 ^ n6713;
  assign n6833 = ~x93 & ~n6832;
  assign n6834 = ~n6830 & ~n6833;
  assign n6835 = x64 & n6817;
  assign n6836 = x21 & ~x65;
  assign n6837 = x22 & ~n6836;
  assign n6838 = ~n6547 & n6837;
  assign n6839 = n6835 & n6838;
  assign n6840 = ~x66 & ~n6839;
  assign n6841 = ~x21 & x65;
  assign n6842 = ~x21 & ~x22;
  assign n6843 = ~n6841 & ~n6842;
  assign n6844 = x64 & ~n6843;
  assign n6845 = ~x22 & n6841;
  assign n6846 = n6845 ^ n6817;
  assign n6847 = n6817 ^ n6546;
  assign n6848 = n6817 & ~n6847;
  assign n6849 = n6848 ^ n6817;
  assign n6850 = ~n6846 & n6849;
  assign n6851 = n6850 ^ n6848;
  assign n6852 = n6851 ^ n6817;
  assign n6853 = n6852 ^ n6546;
  assign n6854 = n6844 & ~n6853;
  assign n6855 = n6840 & ~n6854;
  assign n6856 = ~x22 & x65;
  assign n6857 = ~n6835 & n6856;
  assign n6858 = ~n6847 & n6857;
  assign n6859 = n6855 & ~n6858;
  assign n6860 = ~x21 & x64;
  assign n6861 = n6817 & n6860;
  assign n6862 = ~n6844 & ~n6856;
  assign n6863 = ~n6861 & n6862;
  assign n6864 = ~x65 & ~n6548;
  assign n6865 = n6817 & ~n6864;
  assign n6866 = n6546 & ~n6865;
  assign n6867 = n6863 & n6866;
  assign n6868 = n6548 & ~n6841;
  assign n6869 = ~n6547 & n6868;
  assign n6870 = x22 & n202;
  assign n6871 = ~n6546 & n6870;
  assign n6872 = ~n6869 & ~n6871;
  assign n6873 = n6817 & ~n6872;
  assign n6874 = ~n6867 & ~n6873;
  assign n6875 = ~n6859 & n6874;
  assign n6876 = n6875 ^ x67;
  assign n6877 = n6551 ^ x66;
  assign n6878 = n6817 & n6877;
  assign n6879 = n6878 ^ n6543;
  assign n6880 = n6879 ^ n6875;
  assign n6881 = n6876 & ~n6880;
  assign n6882 = n6881 ^ x67;
  assign n6883 = n6882 ^ x68;
  assign n6884 = n6555 & n6817;
  assign n6885 = n6884 ^ n6558;
  assign n6886 = n6885 ^ n6882;
  assign n6887 = n6883 & n6886;
  assign n6888 = n6887 ^ x68;
  assign n6889 = n6888 ^ x69;
  assign n6890 = n6562 & n6817;
  assign n6891 = n6890 ^ n6564;
  assign n6892 = n6891 ^ n6888;
  assign n6893 = n6889 & ~n6892;
  assign n6894 = n6893 ^ x69;
  assign n6895 = n6894 ^ x70;
  assign n6896 = n6568 & n6817;
  assign n6897 = n6896 ^ n6570;
  assign n6898 = n6897 ^ n6894;
  assign n6899 = n6895 & ~n6898;
  assign n6900 = n6899 ^ x70;
  assign n6901 = n6900 ^ x71;
  assign n6902 = n6574 & n6817;
  assign n6903 = n6902 ^ n6576;
  assign n6904 = n6903 ^ n6900;
  assign n6905 = n6901 & n6904;
  assign n6906 = n6905 ^ x71;
  assign n6907 = n6906 ^ x72;
  assign n6908 = n6579 ^ x71;
  assign n6909 = n6817 & n6908;
  assign n6910 = n6909 ^ n6520;
  assign n6911 = n6910 ^ n6906;
  assign n6912 = n6907 & n6911;
  assign n6913 = n6912 ^ x72;
  assign n6914 = n6913 ^ x73;
  assign n6915 = n6579 ^ n6520;
  assign n6916 = n6908 & n6915;
  assign n6917 = n6916 ^ x71;
  assign n6918 = n6917 ^ x72;
  assign n6919 = n6817 & n6918;
  assign n6920 = n6919 ^ n6523;
  assign n6921 = n6920 ^ n6913;
  assign n6922 = n6914 & ~n6921;
  assign n6923 = n6922 ^ x73;
  assign n6924 = n6923 ^ x74;
  assign n6925 = ~n6587 & n6817;
  assign n6926 = n6925 ^ n6589;
  assign n6927 = n6926 ^ n6923;
  assign n6928 = n6924 & n6927;
  assign n6929 = n6928 ^ x74;
  assign n6930 = n6929 ^ x75;
  assign n6931 = n6593 & n6817;
  assign n6932 = n6931 ^ n6595;
  assign n6933 = n6932 ^ n6929;
  assign n6934 = n6930 & n6933;
  assign n6935 = n6934 ^ x75;
  assign n6936 = n6935 ^ x76;
  assign n6937 = n6599 & n6817;
  assign n6938 = n6937 ^ n6601;
  assign n6939 = n6938 ^ n6935;
  assign n6940 = n6936 & ~n6939;
  assign n6941 = n6940 ^ x76;
  assign n6942 = n6941 ^ x77;
  assign n6943 = n6605 & n6817;
  assign n6944 = n6943 ^ n6607;
  assign n6945 = n6944 ^ n6941;
  assign n6946 = n6942 & n6945;
  assign n6947 = n6946 ^ x77;
  assign n6948 = n6947 ^ x78;
  assign n6949 = n6611 & n6817;
  assign n6950 = n6949 ^ n6613;
  assign n6951 = n6950 ^ n6947;
  assign n6952 = n6948 & n6951;
  assign n6953 = n6952 ^ x78;
  assign n6954 = n6953 ^ x79;
  assign n6955 = n6617 & n6817;
  assign n6956 = n6955 ^ n6619;
  assign n6957 = n6956 ^ n6953;
  assign n6958 = n6954 & n6957;
  assign n6959 = n6958 ^ x79;
  assign n6960 = n6959 ^ x80;
  assign n6961 = n6623 & n6817;
  assign n6962 = n6961 ^ n6625;
  assign n6963 = n6962 ^ n6959;
  assign n6964 = n6960 & ~n6963;
  assign n6965 = n6964 ^ x80;
  assign n6966 = n6965 ^ x81;
  assign n6967 = n6629 & n6817;
  assign n6968 = n6967 ^ n6631;
  assign n6969 = n6968 ^ n6965;
  assign n6970 = n6966 & n6969;
  assign n6971 = n6970 ^ x81;
  assign n6972 = n6971 ^ x82;
  assign n6973 = n6635 & n6817;
  assign n6974 = n6973 ^ n6637;
  assign n6975 = n6974 ^ n6971;
  assign n6976 = n6972 & ~n6975;
  assign n6977 = n6976 ^ x82;
  assign n6978 = n6977 ^ x83;
  assign n6979 = n6641 & n6817;
  assign n6980 = n6979 ^ n6643;
  assign n6981 = n6980 ^ n6977;
  assign n6982 = n6978 & ~n6981;
  assign n6983 = n6982 ^ x83;
  assign n6984 = n6983 ^ x84;
  assign n6985 = n6647 & n6817;
  assign n6986 = n6985 ^ n6649;
  assign n6987 = n6986 ^ n6983;
  assign n6988 = n6984 & ~n6987;
  assign n6989 = n6988 ^ x84;
  assign n6990 = n6989 ^ x85;
  assign n6991 = n6653 & n6817;
  assign n6992 = n6991 ^ n6655;
  assign n6993 = n6992 ^ n6989;
  assign n6994 = n6990 & ~n6993;
  assign n6995 = n6994 ^ x85;
  assign n6996 = n6995 ^ x86;
  assign n6997 = n6659 & n6817;
  assign n6998 = n6997 ^ n6661;
  assign n6999 = n6998 ^ n6995;
  assign n7000 = n6996 & ~n6999;
  assign n7001 = n7000 ^ x86;
  assign n7002 = n7001 ^ x87;
  assign n7003 = n6665 & n6817;
  assign n7004 = n7003 ^ n6667;
  assign n7005 = n7004 ^ n7001;
  assign n7006 = n7002 & ~n7005;
  assign n7007 = n7006 ^ x87;
  assign n7008 = n7007 ^ x88;
  assign n7009 = n6671 & n6817;
  assign n7010 = n7009 ^ n6674;
  assign n7011 = n7010 ^ n7007;
  assign n7012 = n7008 & ~n7011;
  assign n7013 = n7012 ^ x88;
  assign n7014 = n7013 ^ x89;
  assign n7015 = n6678 & n6817;
  assign n7016 = n7015 ^ n6684;
  assign n7017 = n7016 ^ n7013;
  assign n7018 = n7014 & ~n7017;
  assign n7019 = n7018 ^ x89;
  assign n7020 = n7019 ^ x90;
  assign n7021 = n6688 & n6817;
  assign n7022 = n7021 ^ n6691;
  assign n7023 = n7022 ^ n7019;
  assign n7024 = n7020 & n7023;
  assign n7025 = n7024 ^ x90;
  assign n7026 = n7025 ^ x91;
  assign n7027 = n6695 & n6817;
  assign n7028 = n7027 ^ n6701;
  assign n7029 = n7028 ^ n7025;
  assign n7030 = n7026 & ~n7029;
  assign n7031 = n7030 ^ x91;
  assign n7032 = n6834 & n7031;
  assign n7033 = n6832 ^ x93;
  assign n7034 = x92 & ~n6829;
  assign n7035 = n7034 ^ n6832;
  assign n7036 = n7033 & ~n7035;
  assign n7037 = n7036 ^ x93;
  assign n7038 = ~n7032 & ~n7037;
  assign n7039 = n6717 & n6817;
  assign n7040 = n7039 ^ n6720;
  assign n7041 = ~x94 & ~n7040;
  assign n7042 = n6724 & n6817;
  assign n7043 = n7042 ^ n6730;
  assign n7044 = ~x95 & n7043;
  assign n7045 = ~n7041 & ~n7044;
  assign n7046 = ~n7038 & n7045;
  assign n7047 = n7043 ^ x95;
  assign n7048 = x94 & n7040;
  assign n7049 = n7048 ^ n7043;
  assign n7050 = ~n7047 & n7049;
  assign n7051 = n7050 ^ x95;
  assign n7052 = ~n7046 & ~n7051;
  assign n7053 = n7052 ^ x96;
  assign n7054 = n6734 & n6817;
  assign n7055 = n7054 ^ n6736;
  assign n7056 = n7055 ^ n7052;
  assign n7057 = ~n7053 & ~n7056;
  assign n7058 = n7057 ^ x96;
  assign n7059 = n7058 ^ x97;
  assign n7060 = n6740 & n6817;
  assign n7061 = n7060 ^ n6742;
  assign n7062 = n7061 ^ n7058;
  assign n7063 = n7059 & n7062;
  assign n7064 = n7063 ^ x97;
  assign n7065 = n7064 ^ x98;
  assign n7066 = n6746 & n6817;
  assign n7067 = n7066 ^ n6749;
  assign n7068 = n7067 ^ n7064;
  assign n7069 = n7065 & ~n7068;
  assign n7070 = n7069 ^ x98;
  assign n7071 = n6827 & ~n7070;
  assign n7072 = n6825 ^ x100;
  assign n7073 = ~x99 & ~n6819;
  assign n7074 = n7073 ^ n6825;
  assign n7075 = n7072 & n7074;
  assign n7076 = n7075 ^ x100;
  assign n7077 = ~n7071 & n7076;
  assign n7078 = ~n6780 & n6817;
  assign n7079 = n7078 ^ n6782;
  assign n7080 = ~x101 & ~n7079;
  assign n7081 = n6786 & n6817;
  assign n7082 = n7081 ^ n6788;
  assign n7083 = ~x102 & ~n7082;
  assign n7084 = ~n7080 & ~n7083;
  assign n7085 = n7077 & n7084;
  assign n7086 = n7082 ^ x102;
  assign n7087 = x101 & n7079;
  assign n7088 = n7087 ^ n7082;
  assign n7089 = n7086 & ~n7088;
  assign n7090 = n7089 ^ x102;
  assign n7091 = ~n7085 & ~n7090;
  assign n7092 = n7091 ^ x103;
  assign n7093 = n6792 & n6817;
  assign n7094 = n7093 ^ n6794;
  assign n7095 = n7094 ^ n7091;
  assign n7096 = ~n7092 & ~n7095;
  assign n7097 = n7096 ^ x103;
  assign n7098 = n7097 ^ x104;
  assign n7099 = n6798 & n6817;
  assign n7100 = n7099 ^ n6801;
  assign n7101 = n7100 ^ n7097;
  assign n7102 = n7098 & ~n7101;
  assign n7103 = n7102 ^ x104;
  assign n7104 = n7103 ^ x105;
  assign n7105 = n6805 & n6817;
  assign n7106 = n7105 ^ n6809;
  assign n7107 = n7106 ^ n7103;
  assign n7108 = n7104 & n7107;
  assign n7109 = n7108 ^ x105;
  assign n7110 = n7109 ^ x106;
  assign n7111 = n7110 ^ x106;
  assign n7112 = ~x105 & ~n7103;
  assign n7113 = ~x105 & n7106;
  assign n7114 = ~n6812 & ~n7113;
  assign n7115 = ~n7112 & n7114;
  assign n7116 = ~x105 & n6812;
  assign n7117 = ~x106 & ~n7116;
  assign n7118 = ~n7115 & n7117;
  assign n7119 = n7118 ^ x106;
  assign n7120 = ~n7111 & n7119;
  assign n7121 = n7120 ^ x106;
  assign n7122 = n6518 & ~n7121;
  assign n7123 = ~n6517 & ~n7122;
  assign n7124 = ~x107 & n7123;
  assign n7125 = n7109 ^ n6517;
  assign n7126 = n7109 ^ n6813;
  assign n7127 = n6517 ^ x106;
  assign n7128 = n7127 ^ n6813;
  assign n7129 = n6813 & ~n7128;
  assign n7130 = n7129 ^ n6813;
  assign n7131 = n7126 & n7130;
  assign n7132 = n7131 ^ n7129;
  assign n7133 = n7132 ^ n6813;
  assign n7134 = n7133 ^ n7127;
  assign n7135 = n7125 & ~n7134;
  assign n7136 = n7135 ^ n7109;
  assign n7137 = n6518 & ~n7136;
  assign n7138 = ~n7092 & n7137;
  assign n7139 = n7138 ^ n7094;
  assign n7140 = ~x104 & n7139;
  assign n7141 = n7077 ^ x101;
  assign n7142 = n7079 ^ n7077;
  assign n7143 = n7141 & ~n7142;
  assign n7144 = n7143 ^ x101;
  assign n7145 = n7144 ^ x102;
  assign n7146 = n7137 & n7145;
  assign n7147 = n7146 ^ n7082;
  assign n7148 = n7147 ^ x103;
  assign n7149 = n7137 & n7141;
  assign n7150 = n7149 ^ n7079;
  assign n7151 = ~x102 & ~n7150;
  assign n7152 = n7151 ^ n7147;
  assign n7153 = n7152 ^ n7147;
  assign n7154 = x102 & n7150;
  assign n7155 = n7059 & n7137;
  assign n7156 = n7155 ^ n7061;
  assign n7157 = ~x98 & n7156;
  assign n7158 = n7065 & n7137;
  assign n7159 = n7158 ^ n7067;
  assign n7160 = ~x99 & ~n7159;
  assign n7161 = ~n7157 & ~n7160;
  assign n7162 = n6960 & n7137;
  assign n7163 = n7162 ^ n6962;
  assign n7164 = ~x81 & ~n7163;
  assign n7165 = n6966 & n7137;
  assign n7166 = n7165 ^ n6968;
  assign n7167 = ~x82 & n7166;
  assign n7168 = ~n7164 & ~n7167;
  assign n7169 = n6895 & n7137;
  assign n7170 = n7169 ^ n6897;
  assign n7171 = n7170 ^ x71;
  assign n7172 = n6889 & n7137;
  assign n7173 = n7172 ^ n6891;
  assign n7174 = x70 & n7173;
  assign n7175 = n7174 ^ n7170;
  assign n7176 = n7175 ^ n7170;
  assign n7177 = ~x70 & ~n7173;
  assign n7178 = x64 & n7137;
  assign n7179 = n7178 ^ x21;
  assign n7180 = n7179 ^ x65;
  assign n7181 = ~x20 & x64;
  assign n7182 = n7181 ^ n7179;
  assign n7183 = ~n7180 & n7182;
  assign n7184 = n7183 ^ x65;
  assign n7185 = n7184 ^ x66;
  assign n7186 = x65 & ~n6817;
  assign n7187 = x21 & n7186;
  assign n7188 = ~n202 & ~n7187;
  assign n7189 = n6817 ^ x65;
  assign n7190 = n6860 & ~n7189;
  assign n7191 = n7188 & ~n7190;
  assign n7192 = n7191 ^ n6835;
  assign n7193 = n7191 ^ n6836;
  assign n7194 = n7191 ^ n7137;
  assign n7195 = n7191 & n7194;
  assign n7196 = n7195 ^ n7191;
  assign n7197 = n7193 & n7196;
  assign n7198 = n7197 ^ n7195;
  assign n7199 = n7198 ^ n7191;
  assign n7200 = n7199 ^ n7137;
  assign n7201 = ~n7192 & n7200;
  assign n7202 = n7201 ^ n6835;
  assign n7203 = n7202 ^ x22;
  assign n7204 = n7203 ^ n7184;
  assign n7205 = n7185 & n7204;
  assign n7206 = n7205 ^ x66;
  assign n7207 = n7206 ^ x67;
  assign n7211 = n6837 ^ n6817;
  assign n7212 = n7211 ^ n6837;
  assign n7213 = n6842 ^ n6837;
  assign n7214 = ~n7212 & n7213;
  assign n7215 = n7214 ^ n6837;
  assign n7216 = ~n6841 & ~n7215;
  assign n7217 = x64 & ~n7216;
  assign n7218 = ~n6857 & ~n7217;
  assign n7219 = n7218 ^ x66;
  assign n7220 = n7137 & ~n7219;
  assign n7208 = x65 & n6548;
  assign n7209 = n6865 & ~n7208;
  assign n7210 = n7209 ^ n6546;
  assign n7221 = n7220 ^ n7210;
  assign n7222 = n7221 ^ n7206;
  assign n7223 = n7207 & n7222;
  assign n7224 = n7223 ^ x67;
  assign n7225 = n7224 ^ x68;
  assign n7226 = n6876 & n7137;
  assign n7227 = n7226 ^ n6879;
  assign n7228 = n7227 ^ n7224;
  assign n7229 = n7225 & ~n7228;
  assign n7230 = n7229 ^ x68;
  assign n7231 = n7230 ^ x69;
  assign n7232 = n6883 & n7137;
  assign n7233 = n7232 ^ n6885;
  assign n7234 = n7233 ^ n7230;
  assign n7235 = n7231 & n7234;
  assign n7236 = n7235 ^ x69;
  assign n7237 = ~n7177 & n7236;
  assign n7238 = n7237 ^ n7170;
  assign n7239 = n7238 ^ n7170;
  assign n7240 = ~n7176 & ~n7239;
  assign n7241 = n7240 ^ n7170;
  assign n7242 = n7171 & n7241;
  assign n7243 = n7242 ^ x71;
  assign n7244 = n7243 ^ x72;
  assign n7245 = n6901 & n7137;
  assign n7246 = n7245 ^ n6903;
  assign n7247 = n7246 ^ n7243;
  assign n7248 = n7244 & n7247;
  assign n7249 = n7248 ^ x72;
  assign n7250 = n7249 ^ x73;
  assign n7251 = n6907 & n7137;
  assign n7252 = n7251 ^ n6910;
  assign n7253 = n7252 ^ n7249;
  assign n7254 = n7250 & n7253;
  assign n7255 = n7254 ^ x73;
  assign n7256 = n7255 ^ x74;
  assign n7257 = n6914 & n7137;
  assign n7258 = n7257 ^ n6920;
  assign n7259 = n7258 ^ n7255;
  assign n7260 = n7256 & ~n7259;
  assign n7261 = n7260 ^ x74;
  assign n7262 = n7261 ^ x75;
  assign n7263 = n6924 & n7137;
  assign n7264 = n7263 ^ n6926;
  assign n7265 = n7264 ^ n7261;
  assign n7266 = n7262 & n7265;
  assign n7267 = n7266 ^ x75;
  assign n7268 = n7267 ^ x76;
  assign n7269 = n6930 & n7137;
  assign n7270 = n7269 ^ n6932;
  assign n7271 = n7270 ^ n7267;
  assign n7272 = n7268 & n7271;
  assign n7273 = n7272 ^ x76;
  assign n7274 = n7273 ^ x77;
  assign n7275 = n6936 & n7137;
  assign n7276 = n7275 ^ n6938;
  assign n7277 = n7276 ^ n7273;
  assign n7278 = n7274 & ~n7277;
  assign n7279 = n7278 ^ x77;
  assign n7280 = n7279 ^ x78;
  assign n7281 = n6942 & n7137;
  assign n7282 = n7281 ^ n6944;
  assign n7283 = n7282 ^ n7279;
  assign n7284 = n7280 & n7283;
  assign n7285 = n7284 ^ x78;
  assign n7286 = n7285 ^ x79;
  assign n7287 = n6948 & n7137;
  assign n7288 = n7287 ^ n6950;
  assign n7289 = n7288 ^ n7285;
  assign n7290 = n7286 & n7289;
  assign n7291 = n7290 ^ x79;
  assign n7292 = n7291 ^ x80;
  assign n7293 = n6954 & n7137;
  assign n7294 = n7293 ^ n6956;
  assign n7295 = n7294 ^ n7291;
  assign n7296 = n7292 & n7295;
  assign n7297 = n7296 ^ x80;
  assign n7298 = n7168 & n7297;
  assign n7299 = n7166 ^ x82;
  assign n7300 = x81 & n7163;
  assign n7301 = n7300 ^ n7166;
  assign n7302 = ~n7299 & n7301;
  assign n7303 = n7302 ^ x82;
  assign n7304 = ~n7298 & ~n7303;
  assign n7305 = n7304 ^ x83;
  assign n7306 = n6972 & n7137;
  assign n7307 = n7306 ^ n6974;
  assign n7308 = n7307 ^ n7304;
  assign n7309 = ~n7305 & n7308;
  assign n7310 = n7309 ^ x83;
  assign n7311 = n7310 ^ x84;
  assign n7312 = n6978 & n7137;
  assign n7313 = n7312 ^ n6980;
  assign n7314 = n7313 ^ n7310;
  assign n7315 = n7311 & ~n7314;
  assign n7316 = n7315 ^ x84;
  assign n7317 = n7316 ^ x85;
  assign n7318 = n6984 & n7137;
  assign n7319 = n7318 ^ n6986;
  assign n7320 = n7319 ^ n7316;
  assign n7321 = n7317 & ~n7320;
  assign n7322 = n7321 ^ x85;
  assign n7323 = n7322 ^ x86;
  assign n7324 = n6990 & n7137;
  assign n7325 = n7324 ^ n6992;
  assign n7326 = n7325 ^ n7322;
  assign n7327 = n7323 & ~n7326;
  assign n7328 = n7327 ^ x86;
  assign n7329 = n7328 ^ x87;
  assign n7330 = n6996 & n7137;
  assign n7331 = n7330 ^ n6998;
  assign n7332 = n7331 ^ n7328;
  assign n7333 = n7329 & ~n7332;
  assign n7334 = n7333 ^ x87;
  assign n7335 = n7334 ^ x88;
  assign n7336 = n7002 & n7137;
  assign n7337 = n7336 ^ n7004;
  assign n7338 = n7337 ^ n7334;
  assign n7339 = n7335 & ~n7338;
  assign n7340 = n7339 ^ x88;
  assign n7341 = n7340 ^ x89;
  assign n7342 = n7008 & n7137;
  assign n7343 = n7342 ^ n7010;
  assign n7344 = n7343 ^ n7340;
  assign n7345 = n7341 & ~n7344;
  assign n7346 = n7345 ^ x89;
  assign n7347 = n7346 ^ x90;
  assign n7348 = n7014 & n7137;
  assign n7349 = n7348 ^ n7016;
  assign n7350 = n7349 ^ n7346;
  assign n7351 = n7347 & ~n7350;
  assign n7352 = n7351 ^ x90;
  assign n7353 = n7352 ^ x91;
  assign n7354 = n7020 & n7137;
  assign n7355 = n7354 ^ n7022;
  assign n7356 = n7355 ^ n7352;
  assign n7357 = n7353 & n7356;
  assign n7358 = n7357 ^ x91;
  assign n7359 = n7358 ^ x92;
  assign n7360 = n7026 & n7137;
  assign n7361 = n7360 ^ n7028;
  assign n7362 = n7361 ^ n7358;
  assign n7363 = n7359 & ~n7362;
  assign n7364 = n7363 ^ x92;
  assign n7365 = n7364 ^ x93;
  assign n7366 = n7031 ^ x92;
  assign n7367 = n7137 & n7366;
  assign n7368 = n7367 ^ n6829;
  assign n7369 = n7368 ^ n7364;
  assign n7370 = n7365 & n7369;
  assign n7371 = n7370 ^ x93;
  assign n7372 = n7371 ^ x94;
  assign n7373 = n7031 ^ n6829;
  assign n7374 = n7366 & n7373;
  assign n7375 = n7374 ^ x92;
  assign n7376 = n7375 ^ x93;
  assign n7377 = n7137 & n7376;
  assign n7378 = n7377 ^ n6832;
  assign n7379 = n7378 ^ n7371;
  assign n7380 = n7372 & ~n7379;
  assign n7381 = n7380 ^ x94;
  assign n7382 = n7381 ^ x95;
  assign n7383 = n7038 ^ x94;
  assign n7384 = n7137 & ~n7383;
  assign n7385 = n7384 ^ n7040;
  assign n7386 = n7385 ^ n7381;
  assign n7387 = n7382 & ~n7386;
  assign n7388 = n7387 ^ x95;
  assign n7389 = n7388 ^ x96;
  assign n7390 = n7040 ^ n7038;
  assign n7391 = ~n7383 & n7390;
  assign n7392 = n7391 ^ x94;
  assign n7393 = n7392 ^ x95;
  assign n7394 = n7137 & n7393;
  assign n7395 = n7394 ^ n7043;
  assign n7396 = n7395 ^ n7388;
  assign n7397 = n7389 & n7396;
  assign n7398 = n7397 ^ x96;
  assign n7399 = n7398 ^ x97;
  assign n7400 = ~n7053 & n7137;
  assign n7401 = n7400 ^ n7055;
  assign n7402 = n7401 ^ n7398;
  assign n7403 = n7399 & n7402;
  assign n7404 = n7403 ^ x97;
  assign n7405 = n7161 & n7404;
  assign n7406 = n7159 ^ x99;
  assign n7407 = x98 & ~n7156;
  assign n7408 = n7407 ^ n7159;
  assign n7409 = n7406 & ~n7408;
  assign n7410 = n7409 ^ x99;
  assign n7411 = ~n7405 & ~n7410;
  assign n7412 = n7411 ^ x100;
  assign n7413 = n7070 ^ x99;
  assign n7414 = n7137 & n7413;
  assign n7415 = n7414 ^ n6819;
  assign n7416 = n7415 ^ n7411;
  assign n7417 = ~n7412 & n7416;
  assign n7418 = n7417 ^ x100;
  assign n7419 = n7418 ^ x101;
  assign n7420 = n7070 ^ n6819;
  assign n7421 = n7413 & ~n7420;
  assign n7422 = n7421 ^ x99;
  assign n7423 = n7422 ^ x100;
  assign n7424 = n7137 & n7423;
  assign n7425 = n7424 ^ n6825;
  assign n7426 = n7425 ^ n7418;
  assign n7427 = n7419 & ~n7426;
  assign n7428 = n7427 ^ x101;
  assign n7429 = ~n7154 & ~n7428;
  assign n7430 = n7429 ^ n7147;
  assign n7431 = n7430 ^ n7147;
  assign n7432 = ~n7153 & ~n7431;
  assign n7433 = n7432 ^ n7147;
  assign n7434 = n7148 & ~n7433;
  assign n7435 = n7434 ^ x103;
  assign n7436 = ~n7140 & n7435;
  assign n7437 = n7098 & n7137;
  assign n7438 = n7437 ^ n7100;
  assign n7439 = x104 & x105;
  assign n7440 = ~n7438 & ~n7439;
  assign n7441 = n7436 & ~n7440;
  assign n7442 = x105 & ~n7139;
  assign n7443 = n7435 & n7442;
  assign n7444 = n7438 ^ x105;
  assign n7445 = x104 & ~n7139;
  assign n7446 = n7445 ^ n7438;
  assign n7447 = n7444 & ~n7446;
  assign n7448 = n7447 ^ x105;
  assign n7449 = ~n7443 & ~n7448;
  assign n7450 = ~n7441 & n7449;
  assign n7451 = n7450 ^ x106;
  assign n7452 = n7104 & n7137;
  assign n7453 = n7452 ^ n7106;
  assign n7454 = n7453 ^ n7450;
  assign n7455 = ~n7451 & ~n7454;
  assign n7456 = n7455 ^ x106;
  assign n7457 = ~n7124 & n7456;
  assign n7458 = x107 & n6517;
  assign n7459 = n6208 & ~n7458;
  assign n7460 = ~n7457 & n7459;
  assign n7464 = x64 & n7460;
  assign n7465 = ~x20 & x65;
  assign n7466 = ~n7464 & n7465;
  assign n7467 = n7460 ^ n7179;
  assign n7468 = n7466 & ~n7467;
  assign n7469 = ~x66 & ~n7468;
  assign n7471 = ~x65 & n7460;
  assign n7472 = x20 & ~x65;
  assign n7473 = ~x19 & ~n7472;
  assign n7474 = ~n7471 & n7473;
  assign n7475 = ~n7179 & n7474;
  assign n7470 = x20 & n7460;
  assign n7476 = n7475 ^ n7470;
  assign n7477 = n7476 ^ n7475;
  assign n7478 = x19 & ~x65;
  assign n7479 = ~n7180 & ~n7478;
  assign n7480 = n7479 ^ n7475;
  assign n7481 = n7477 & n7480;
  assign n7482 = n7481 ^ n7475;
  assign n7483 = x64 & n7482;
  assign n7484 = n7469 & ~n7483;
  assign n7485 = n7179 & ~n7465;
  assign n7486 = ~x19 & x64;
  assign n7487 = n7486 ^ n7460;
  assign n7488 = ~x65 & ~n7181;
  assign n7489 = n7488 ^ n7486;
  assign n7490 = n7489 ^ n7488;
  assign n7491 = n7488 ^ n7472;
  assign n7492 = n7490 & ~n7491;
  assign n7493 = n7492 ^ n7488;
  assign n7494 = n7487 & n7493;
  assign n7495 = n7494 ^ n7460;
  assign n7496 = n7485 & ~n7495;
  assign n7497 = ~x21 & n202;
  assign n7498 = n7470 & n7497;
  assign n7499 = ~x19 & x65;
  assign n7500 = n7181 & ~n7499;
  assign n7501 = ~n7180 & n7500;
  assign n7502 = n7460 & n7501;
  assign n7503 = ~n7498 & ~n7502;
  assign n7504 = ~n7496 & n7503;
  assign n7505 = ~n7484 & n7504;
  assign n7506 = n7505 ^ x67;
  assign n7507 = n7185 & n7460;
  assign n7508 = n7507 ^ n7203;
  assign n7509 = n7508 ^ n7505;
  assign n7510 = n7506 & n7509;
  assign n7511 = n7510 ^ x67;
  assign n7512 = n7511 ^ x68;
  assign n7513 = n7207 & n7460;
  assign n7514 = n7513 ^ n7221;
  assign n7515 = n7514 ^ n7511;
  assign n7516 = n7512 & n7515;
  assign n7517 = n7516 ^ x68;
  assign n7518 = n7517 ^ x69;
  assign n7519 = n7225 & n7460;
  assign n7520 = n7519 ^ n7227;
  assign n7521 = n7520 ^ n7517;
  assign n7522 = n7518 & ~n7521;
  assign n7523 = n7522 ^ x69;
  assign n7524 = n7523 ^ x70;
  assign n7525 = n7231 & n7460;
  assign n7526 = n7525 ^ n7233;
  assign n7527 = n7526 ^ n7523;
  assign n7528 = n7524 & n7527;
  assign n7529 = n7528 ^ x70;
  assign n7530 = n7529 ^ x71;
  assign n7531 = n7236 ^ x70;
  assign n7532 = n7460 & n7531;
  assign n7533 = n7532 ^ n7173;
  assign n7534 = n7533 ^ n7529;
  assign n7535 = n7530 & ~n7534;
  assign n7536 = n7535 ^ x71;
  assign n7537 = n7536 ^ x72;
  assign n7538 = ~n7174 & ~n7237;
  assign n7539 = n7538 ^ x71;
  assign n7540 = n7460 & ~n7539;
  assign n7541 = n7540 ^ n7170;
  assign n7542 = n7541 ^ n7536;
  assign n7543 = n7537 & ~n7542;
  assign n7544 = n7543 ^ x72;
  assign n7545 = n7544 ^ x73;
  assign n7546 = n7244 & n7460;
  assign n7547 = n7546 ^ n7246;
  assign n7548 = n7547 ^ n7544;
  assign n7549 = n7545 & n7548;
  assign n7550 = n7549 ^ x73;
  assign n7551 = n7550 ^ x74;
  assign n7552 = n7250 & n7460;
  assign n7553 = n7552 ^ n7252;
  assign n7554 = n7553 ^ n7550;
  assign n7555 = n7551 & n7554;
  assign n7556 = n7555 ^ x74;
  assign n7557 = n7556 ^ x75;
  assign n7558 = n7256 & n7460;
  assign n7559 = n7558 ^ n7258;
  assign n7560 = n7559 ^ n7556;
  assign n7561 = n7557 & ~n7560;
  assign n7562 = n7561 ^ x75;
  assign n7563 = n7562 ^ x76;
  assign n7564 = n7262 & n7460;
  assign n7565 = n7564 ^ n7264;
  assign n7566 = n7565 ^ n7562;
  assign n7567 = n7563 & n7566;
  assign n7568 = n7567 ^ x76;
  assign n7569 = n7568 ^ x77;
  assign n7570 = n7268 & n7460;
  assign n7571 = n7570 ^ n7270;
  assign n7572 = n7571 ^ n7568;
  assign n7573 = n7569 & n7572;
  assign n7574 = n7573 ^ x77;
  assign n7575 = n7574 ^ x78;
  assign n7576 = n7274 & n7460;
  assign n7577 = n7576 ^ n7276;
  assign n7578 = n7577 ^ n7574;
  assign n7579 = n7575 & ~n7578;
  assign n7580 = n7579 ^ x78;
  assign n7581 = n7580 ^ x79;
  assign n7582 = n7280 & n7460;
  assign n7583 = n7582 ^ n7282;
  assign n7584 = n7583 ^ n7580;
  assign n7585 = n7581 & n7584;
  assign n7586 = n7585 ^ x79;
  assign n7587 = n7586 ^ x80;
  assign n7588 = n7286 & n7460;
  assign n7589 = n7588 ^ n7288;
  assign n7590 = n7589 ^ n7586;
  assign n7591 = n7587 & n7590;
  assign n7592 = n7591 ^ x80;
  assign n7593 = n7592 ^ x81;
  assign n7594 = n7292 & n7460;
  assign n7595 = n7594 ^ n7294;
  assign n7596 = n7595 ^ n7592;
  assign n7597 = n7593 & n7596;
  assign n7598 = n7597 ^ x81;
  assign n7599 = n7598 ^ x82;
  assign n7600 = n7297 ^ x81;
  assign n7601 = n7460 & n7600;
  assign n7602 = n7601 ^ n7163;
  assign n7603 = n7602 ^ n7598;
  assign n7604 = n7599 & ~n7603;
  assign n7605 = n7604 ^ x82;
  assign n7606 = n7605 ^ x83;
  assign n7607 = n7297 ^ n7163;
  assign n7608 = n7600 & ~n7607;
  assign n7609 = n7608 ^ x81;
  assign n7610 = n7609 ^ x82;
  assign n7611 = n7460 & n7610;
  assign n7612 = n7611 ^ n7166;
  assign n7613 = n7612 ^ n7605;
  assign n7614 = n7606 & n7613;
  assign n7615 = n7614 ^ x83;
  assign n7616 = n7615 ^ x84;
  assign n7617 = ~n7305 & n7460;
  assign n7618 = n7617 ^ n7307;
  assign n7619 = n7618 ^ n7615;
  assign n7620 = n7616 & ~n7619;
  assign n7621 = n7620 ^ x84;
  assign n7622 = n7621 ^ x85;
  assign n7623 = n7311 & n7460;
  assign n7624 = n7623 ^ n7313;
  assign n7625 = n7624 ^ n7621;
  assign n7626 = n7622 & ~n7625;
  assign n7627 = n7626 ^ x85;
  assign n7628 = n7627 ^ x86;
  assign n7629 = n7317 & n7460;
  assign n7630 = n7629 ^ n7319;
  assign n7631 = n7630 ^ n7627;
  assign n7632 = n7628 & ~n7631;
  assign n7633 = n7632 ^ x86;
  assign n7634 = n7633 ^ x87;
  assign n7635 = n7323 & n7460;
  assign n7636 = n7635 ^ n7325;
  assign n7637 = n7636 ^ n7633;
  assign n7638 = n7634 & ~n7637;
  assign n7639 = n7638 ^ x87;
  assign n7640 = n7639 ^ x88;
  assign n7641 = n7329 & n7460;
  assign n7642 = n7641 ^ n7331;
  assign n7643 = n7642 ^ n7639;
  assign n7644 = n7640 & ~n7643;
  assign n7645 = n7644 ^ x88;
  assign n7646 = n7645 ^ x89;
  assign n7647 = n7335 & n7460;
  assign n7648 = n7647 ^ n7337;
  assign n7649 = n7648 ^ n7645;
  assign n7650 = n7646 & ~n7649;
  assign n7651 = n7650 ^ x89;
  assign n7652 = n7651 ^ x90;
  assign n7653 = n7341 & n7460;
  assign n7654 = n7653 ^ n7343;
  assign n7655 = n7654 ^ n7651;
  assign n7656 = n7652 & ~n7655;
  assign n7657 = n7656 ^ x90;
  assign n7658 = n7657 ^ x91;
  assign n7659 = n7347 & n7460;
  assign n7660 = n7659 ^ n7349;
  assign n7661 = n7660 ^ n7657;
  assign n7662 = n7658 & ~n7661;
  assign n7663 = n7662 ^ x91;
  assign n7664 = n7663 ^ x92;
  assign n7665 = n7353 & n7460;
  assign n7666 = n7665 ^ n7355;
  assign n7667 = n7666 ^ n7663;
  assign n7668 = n7664 & n7667;
  assign n7669 = n7668 ^ x92;
  assign n7670 = n7669 ^ x93;
  assign n7671 = n7359 & n7460;
  assign n7672 = n7671 ^ n7361;
  assign n7673 = n7672 ^ n7669;
  assign n7674 = n7670 & ~n7673;
  assign n7675 = n7674 ^ x93;
  assign n7676 = n7675 ^ x94;
  assign n7677 = n7365 & n7460;
  assign n7678 = n7677 ^ n7368;
  assign n7679 = n7678 ^ n7675;
  assign n7680 = n7676 & n7679;
  assign n7681 = n7680 ^ x94;
  assign n7682 = n7681 ^ x95;
  assign n7683 = n7372 & n7460;
  assign n7684 = n7683 ^ n7378;
  assign n7685 = n7684 ^ n7681;
  assign n7686 = n7682 & ~n7685;
  assign n7687 = n7686 ^ x95;
  assign n7688 = n7687 ^ x96;
  assign n7689 = n7382 & n7460;
  assign n7690 = n7689 ^ n7385;
  assign n7691 = n7690 ^ n7687;
  assign n7692 = n7688 & ~n7691;
  assign n7693 = n7692 ^ x96;
  assign n7694 = n7693 ^ x97;
  assign n7695 = n7389 & n7460;
  assign n7696 = n7695 ^ n7395;
  assign n7697 = n7696 ^ n7693;
  assign n7698 = n7694 & n7697;
  assign n7699 = n7698 ^ x97;
  assign n7700 = n7699 ^ x98;
  assign n7701 = n7399 & n7460;
  assign n7702 = n7701 ^ n7401;
  assign n7703 = n7702 ^ n7699;
  assign n7704 = n7700 & n7703;
  assign n7705 = n7704 ^ x98;
  assign n7706 = n7705 ^ x99;
  assign n7707 = n7404 ^ x98;
  assign n7708 = n7460 & n7707;
  assign n7709 = n7708 ^ n7156;
  assign n7710 = n7709 ^ n7705;
  assign n7711 = n7706 & n7710;
  assign n7712 = n7711 ^ x99;
  assign n7713 = n7712 ^ x100;
  assign n7714 = n7404 ^ n7156;
  assign n7715 = n7707 & n7714;
  assign n7716 = n7715 ^ x98;
  assign n7717 = n7716 ^ x99;
  assign n7718 = n7460 & n7717;
  assign n7719 = n7718 ^ n7159;
  assign n7720 = n7719 ^ n7712;
  assign n7721 = n7713 & ~n7720;
  assign n7722 = n7721 ^ x100;
  assign n7723 = n7722 ^ x101;
  assign n7724 = ~n7412 & n7460;
  assign n7725 = n7724 ^ n7415;
  assign n7726 = n7725 ^ n7722;
  assign n7727 = n7723 & ~n7726;
  assign n7728 = n7727 ^ x101;
  assign n7729 = n7728 ^ x102;
  assign n7730 = n7419 & n7460;
  assign n7731 = n7730 ^ n7425;
  assign n7732 = n7731 ^ n7728;
  assign n7733 = n7729 & ~n7732;
  assign n7734 = n7733 ^ x102;
  assign n7735 = n7734 ^ x103;
  assign n7736 = n7428 ^ x102;
  assign n7737 = n7460 & n7736;
  assign n7738 = n7737 ^ n7150;
  assign n7739 = n7738 ^ n7734;
  assign n7740 = n7735 & ~n7739;
  assign n7741 = n7740 ^ x103;
  assign n7742 = n7741 ^ x104;
  assign n7743 = ~n7151 & ~n7429;
  assign n7744 = n7743 ^ x103;
  assign n7745 = n7460 & n7744;
  assign n7746 = n7745 ^ n7147;
  assign n7747 = n7746 ^ n7741;
  assign n7748 = n7742 & ~n7747;
  assign n7749 = n7748 ^ x104;
  assign n7750 = n7749 ^ x105;
  assign n7461 = ~n7451 & n7460;
  assign n7462 = n7461 ^ n7453;
  assign n7463 = x107 & ~n7462;
  assign n7751 = n7435 ^ x104;
  assign n7752 = n7460 & n7751;
  assign n7753 = n7752 ^ n7139;
  assign n7754 = n7753 ^ n7749;
  assign n7755 = n7750 & n7754;
  assign n7756 = n7755 ^ x105;
  assign n7757 = n7756 ^ x106;
  assign n7758 = ~n7436 & ~n7445;
  assign n7759 = n7758 ^ x105;
  assign n7760 = n7460 & ~n7759;
  assign n7761 = n7760 ^ n7438;
  assign n7762 = n7761 ^ n7756;
  assign n7763 = n7757 & ~n7762;
  assign n7764 = n7763 ^ x106;
  assign n7765 = ~n7463 & ~n7764;
  assign n7766 = ~x107 & n7462;
  assign n7768 = n7456 ^ x107;
  assign n7769 = ~x108 & ~n7768;
  assign n7775 = ~n7122 & n7769;
  assign n7776 = ~n7766 & ~n7775;
  assign n7777 = ~n7765 & n7776;
  assign n7778 = n147 & ~n6517;
  assign n7779 = ~n7777 & n7778;
  assign n7767 = ~n7765 & ~n7766;
  assign n7780 = n6208 & ~n7767;
  assign n7781 = ~n7779 & ~n7780;
  assign n7782 = n7750 & ~n7781;
  assign n7783 = n7782 ^ n7753;
  assign n7784 = ~x106 & n7783;
  assign n7785 = n7757 & ~n7781;
  assign n7786 = n7785 ^ n7761;
  assign n7787 = ~x107 & ~n7786;
  assign n7788 = ~n7784 & ~n7787;
  assign n7789 = n7688 & ~n7781;
  assign n7790 = n7789 ^ n7690;
  assign n7791 = x97 & n7790;
  assign n7792 = n7694 & ~n7781;
  assign n7793 = n7792 ^ n7696;
  assign n7794 = x98 & ~n7793;
  assign n7795 = ~n7791 & ~n7794;
  assign n7796 = n7581 & ~n7781;
  assign n7797 = n7796 ^ n7583;
  assign n7798 = x80 & ~n7797;
  assign n7799 = n7587 & ~n7781;
  assign n7800 = n7799 ^ n7589;
  assign n7801 = x81 & ~n7800;
  assign n7802 = ~n7798 & ~n7801;
  assign n7803 = n7781 ^ n7464;
  assign n7804 = n7803 ^ n7464;
  assign n7805 = n7464 ^ n7460;
  assign n7806 = n7805 ^ n7464;
  assign n7807 = ~n7804 & ~n7806;
  assign n7808 = n7807 ^ n7464;
  assign n7809 = x65 & n7808;
  assign n7810 = n7809 ^ n7464;
  assign n7811 = x19 & n7810;
  assign n7812 = x65 & ~n7460;
  assign n7813 = n7486 & ~n7812;
  assign n7814 = ~n202 & ~n7813;
  assign n7815 = ~n7471 & ~n7814;
  assign n7816 = n7815 ^ n7464;
  assign n7817 = ~n7781 & n7816;
  assign n7818 = n7817 ^ n7464;
  assign n7819 = ~n7811 & ~n7818;
  assign n7820 = n7819 ^ x20;
  assign n7821 = n7820 ^ x66;
  assign n7822 = x64 & ~n7781;
  assign n7823 = x18 & n7478;
  assign n7824 = n7823 ^ x19;
  assign n7825 = n7822 & n7824;
  assign n7826 = ~x18 & n7486;
  assign n7827 = ~n7499 & ~n7826;
  assign n7828 = n7781 & ~n7827;
  assign n7829 = ~x18 & x65;
  assign n7830 = n7829 ^ n7499;
  assign n7831 = x64 & n7830;
  assign n7832 = n7831 ^ n7499;
  assign n7833 = ~n7828 & ~n7832;
  assign n7834 = ~n7825 & n7833;
  assign n7835 = n7834 ^ n7820;
  assign n7836 = n7821 & n7835;
  assign n7837 = n7836 ^ x66;
  assign n7838 = n7837 ^ x67;
  assign n7842 = n7470 & ~n7478;
  assign n7843 = ~n7474 & ~n7842;
  assign n7844 = x64 & ~n7843;
  assign n7845 = ~n7466 & ~n7844;
  assign n7846 = n7845 ^ x66;
  assign n7847 = ~n7781 & ~n7846;
  assign n7839 = n7181 ^ x65;
  assign n7840 = n7460 & n7839;
  assign n7841 = n7840 ^ n7179;
  assign n7848 = n7847 ^ n7841;
  assign n7849 = n7848 ^ n7837;
  assign n7850 = n7838 & n7849;
  assign n7851 = n7850 ^ x67;
  assign n7852 = n7851 ^ x68;
  assign n7853 = n7506 & ~n7781;
  assign n7854 = n7853 ^ n7508;
  assign n7855 = n7854 ^ n7851;
  assign n7856 = n7852 & n7855;
  assign n7857 = n7856 ^ x68;
  assign n7858 = n7857 ^ x69;
  assign n7859 = n7512 & ~n7781;
  assign n7860 = n7859 ^ n7514;
  assign n7861 = n7860 ^ n7857;
  assign n7862 = n7858 & n7861;
  assign n7863 = n7862 ^ x69;
  assign n7864 = n7863 ^ x70;
  assign n7865 = n7518 & ~n7781;
  assign n7866 = n7865 ^ n7520;
  assign n7867 = n7866 ^ n7863;
  assign n7868 = n7864 & ~n7867;
  assign n7869 = n7868 ^ x70;
  assign n7870 = n7869 ^ x71;
  assign n7871 = n7524 & ~n7781;
  assign n7872 = n7871 ^ n7526;
  assign n7873 = n7872 ^ n7869;
  assign n7874 = n7870 & n7873;
  assign n7875 = n7874 ^ x71;
  assign n7876 = n7875 ^ x72;
  assign n7877 = n7530 & ~n7781;
  assign n7878 = n7877 ^ n7533;
  assign n7879 = n7878 ^ n7875;
  assign n7880 = n7876 & ~n7879;
  assign n7881 = n7880 ^ x72;
  assign n7882 = n7881 ^ x73;
  assign n7883 = n7537 & ~n7781;
  assign n7884 = n7883 ^ n7541;
  assign n7885 = n7884 ^ n7881;
  assign n7886 = n7882 & ~n7885;
  assign n7887 = n7886 ^ x73;
  assign n7888 = n7887 ^ x74;
  assign n7889 = n7545 & ~n7781;
  assign n7890 = n7889 ^ n7547;
  assign n7891 = n7890 ^ n7887;
  assign n7892 = n7888 & n7891;
  assign n7893 = n7892 ^ x74;
  assign n7894 = n7893 ^ x75;
  assign n7895 = n7551 & ~n7781;
  assign n7896 = n7895 ^ n7553;
  assign n7897 = n7896 ^ n7893;
  assign n7898 = n7894 & n7897;
  assign n7899 = n7898 ^ x75;
  assign n7900 = n7899 ^ x76;
  assign n7901 = n7557 & ~n7781;
  assign n7902 = n7901 ^ n7559;
  assign n7903 = n7902 ^ n7899;
  assign n7904 = n7900 & ~n7903;
  assign n7905 = n7904 ^ x76;
  assign n7906 = n7905 ^ x77;
  assign n7907 = n7563 & ~n7781;
  assign n7908 = n7907 ^ n7565;
  assign n7909 = n7908 ^ n7905;
  assign n7910 = n7906 & n7909;
  assign n7911 = n7910 ^ x77;
  assign n7912 = n7911 ^ x78;
  assign n7913 = n7569 & ~n7781;
  assign n7914 = n7913 ^ n7571;
  assign n7915 = n7914 ^ n7911;
  assign n7916 = n7912 & n7915;
  assign n7917 = n7916 ^ x78;
  assign n7918 = n7917 ^ x79;
  assign n7919 = n7575 & ~n7781;
  assign n7920 = n7919 ^ n7577;
  assign n7921 = n7920 ^ n7917;
  assign n7922 = n7918 & ~n7921;
  assign n7923 = n7922 ^ x79;
  assign n7924 = n7802 & ~n7923;
  assign n7925 = n7800 ^ x81;
  assign n7926 = ~x80 & n7797;
  assign n7927 = n7926 ^ n7800;
  assign n7928 = ~n7925 & ~n7927;
  assign n7929 = n7928 ^ x81;
  assign n7930 = ~n7924 & n7929;
  assign n7931 = n7930 ^ x82;
  assign n7932 = n7593 & ~n7781;
  assign n7933 = n7932 ^ n7595;
  assign n7934 = n7933 ^ n7930;
  assign n7935 = n7931 & n7934;
  assign n7936 = n7935 ^ x82;
  assign n7937 = n7936 ^ x83;
  assign n7938 = n7599 & ~n7781;
  assign n7939 = n7938 ^ n7602;
  assign n7940 = n7939 ^ n7936;
  assign n7941 = n7937 & ~n7940;
  assign n7942 = n7941 ^ x83;
  assign n7943 = n7942 ^ x84;
  assign n7944 = n7606 & ~n7781;
  assign n7945 = n7944 ^ n7612;
  assign n7946 = n7945 ^ n7942;
  assign n7947 = n7943 & n7946;
  assign n7948 = n7947 ^ x84;
  assign n7949 = n7948 ^ x85;
  assign n7950 = n7616 & ~n7781;
  assign n7951 = n7950 ^ n7618;
  assign n7952 = n7951 ^ n7948;
  assign n7953 = n7949 & ~n7952;
  assign n7954 = n7953 ^ x85;
  assign n7955 = n7954 ^ x86;
  assign n7956 = n7622 & ~n7781;
  assign n7957 = n7956 ^ n7624;
  assign n7958 = n7957 ^ n7954;
  assign n7959 = n7955 & ~n7958;
  assign n7960 = n7959 ^ x86;
  assign n7961 = n7960 ^ x87;
  assign n7962 = n7628 & ~n7781;
  assign n7963 = n7962 ^ n7630;
  assign n7964 = n7963 ^ n7960;
  assign n7965 = n7961 & ~n7964;
  assign n7966 = n7965 ^ x87;
  assign n7967 = n7966 ^ x88;
  assign n7968 = n7634 & ~n7781;
  assign n7969 = n7968 ^ n7636;
  assign n7970 = n7969 ^ n7966;
  assign n7971 = n7967 & ~n7970;
  assign n7972 = n7971 ^ x88;
  assign n7973 = n7972 ^ x89;
  assign n7974 = n7640 & ~n7781;
  assign n7975 = n7974 ^ n7642;
  assign n7976 = n7975 ^ n7972;
  assign n7977 = n7973 & ~n7976;
  assign n7978 = n7977 ^ x89;
  assign n7979 = n7978 ^ x90;
  assign n7980 = n7646 & ~n7781;
  assign n7981 = n7980 ^ n7648;
  assign n7982 = n7981 ^ n7978;
  assign n7983 = n7979 & ~n7982;
  assign n7984 = n7983 ^ x90;
  assign n7985 = n7984 ^ x91;
  assign n7986 = n7652 & ~n7781;
  assign n7987 = n7986 ^ n7654;
  assign n7988 = n7987 ^ n7984;
  assign n7989 = n7985 & ~n7988;
  assign n7990 = n7989 ^ x91;
  assign n7991 = n7990 ^ x92;
  assign n7992 = n7658 & ~n7781;
  assign n7993 = n7992 ^ n7660;
  assign n7994 = n7993 ^ n7990;
  assign n7995 = n7991 & ~n7994;
  assign n7996 = n7995 ^ x92;
  assign n7997 = n7996 ^ x93;
  assign n7998 = n7664 & ~n7781;
  assign n7999 = n7998 ^ n7666;
  assign n8000 = n7999 ^ n7996;
  assign n8001 = n7997 & n8000;
  assign n8002 = n8001 ^ x93;
  assign n8003 = n8002 ^ x94;
  assign n8004 = n7670 & ~n7781;
  assign n8005 = n8004 ^ n7672;
  assign n8006 = n8005 ^ n8002;
  assign n8007 = n8003 & ~n8006;
  assign n8008 = n8007 ^ x94;
  assign n8009 = n8008 ^ x95;
  assign n8010 = n7676 & ~n7781;
  assign n8011 = n8010 ^ n7678;
  assign n8012 = n8011 ^ n8008;
  assign n8013 = n8009 & n8012;
  assign n8014 = n8013 ^ x95;
  assign n8015 = n8014 ^ x96;
  assign n8016 = n7682 & ~n7781;
  assign n8017 = n8016 ^ n7684;
  assign n8018 = n8017 ^ n8014;
  assign n8019 = n8015 & ~n8018;
  assign n8020 = n8019 ^ x96;
  assign n8021 = n7795 & ~n8020;
  assign n8022 = n7793 ^ x98;
  assign n8023 = ~x97 & ~n7790;
  assign n8024 = n8023 ^ n7793;
  assign n8025 = ~n8022 & ~n8024;
  assign n8026 = n8025 ^ x98;
  assign n8027 = ~n8021 & n8026;
  assign n8028 = n7700 & ~n7781;
  assign n8029 = n8028 ^ n7702;
  assign n8030 = ~x99 & n8029;
  assign n8031 = n7706 & ~n7781;
  assign n8032 = n8031 ^ n7709;
  assign n8033 = ~x100 & n8032;
  assign n8034 = ~n8030 & ~n8033;
  assign n8035 = n8027 & n8034;
  assign n8036 = n8032 ^ x100;
  assign n8037 = x99 & ~n8029;
  assign n8038 = n8037 ^ n8032;
  assign n8039 = ~n8036 & n8038;
  assign n8040 = n8039 ^ x100;
  assign n8041 = ~n8035 & ~n8040;
  assign n8042 = n8041 ^ x101;
  assign n8043 = n7713 & ~n7781;
  assign n8044 = n8043 ^ n7719;
  assign n8045 = n8044 ^ n8041;
  assign n8046 = ~n8042 & n8045;
  assign n8047 = n8046 ^ x101;
  assign n8048 = n8047 ^ x102;
  assign n8049 = n7723 & ~n7781;
  assign n8050 = n8049 ^ n7725;
  assign n8051 = n8050 ^ n8047;
  assign n8052 = n8048 & ~n8051;
  assign n8053 = n8052 ^ x102;
  assign n8054 = n8053 ^ x103;
  assign n8055 = n7729 & ~n7781;
  assign n8056 = n8055 ^ n7731;
  assign n8057 = n8056 ^ n8053;
  assign n8058 = n8054 & ~n8057;
  assign n8059 = n8058 ^ x103;
  assign n8060 = n8059 ^ x104;
  assign n8061 = n7735 & ~n7781;
  assign n8062 = n8061 ^ n7738;
  assign n8063 = n8062 ^ n8059;
  assign n8064 = n8060 & ~n8063;
  assign n8065 = n8064 ^ x104;
  assign n8066 = n8065 ^ x105;
  assign n8067 = n7742 & ~n7781;
  assign n8068 = n8067 ^ n7746;
  assign n8069 = n8068 ^ n8065;
  assign n8070 = n8066 & ~n8069;
  assign n8071 = n8070 ^ x105;
  assign n8072 = n7788 & n8071;
  assign n8073 = n7786 ^ x107;
  assign n8074 = x106 & ~n7783;
  assign n8075 = n8074 ^ n7786;
  assign n8076 = n8073 & ~n8075;
  assign n8077 = n8076 ^ x107;
  assign n8078 = ~n8072 & ~n8077;
  assign n8079 = n8078 ^ x108;
  assign n8080 = n7764 ^ x107;
  assign n8081 = ~n7781 & n8080;
  assign n8082 = n8081 ^ n7462;
  assign n8083 = n8082 ^ n8078;
  assign n8084 = ~n8079 & ~n8083;
  assign n8085 = n8084 ^ x108;
  assign n7770 = n7769 ^ x108;
  assign n7771 = ~n7767 & n7770;
  assign n7772 = n7771 ^ x108;
  assign n7773 = n147 & ~n7772;
  assign n7774 = n7123 & ~n7773;
  assign n8089 = ~x109 & n7774;
  assign n8090 = n8085 & ~n8089;
  assign n8091 = x109 & n6517;
  assign n8092 = n146 & ~n8091;
  assign n8093 = ~n8090 & n8092;
  assign n8101 = n8093 ^ n7822;
  assign n8102 = n8101 ^ n7822;
  assign n8103 = n7822 ^ n7781;
  assign n8104 = n8103 ^ n7822;
  assign n8105 = n8102 & n8104;
  assign n8106 = n8105 ^ n7822;
  assign n8107 = x65 & n8106;
  assign n8108 = n8107 ^ n7822;
  assign n8109 = x18 & n8108;
  assign n8110 = ~n288 & n7781;
  assign n8111 = ~x18 & ~n8110;
  assign n8112 = ~n202 & ~n8111;
  assign n8113 = ~x65 & ~n7781;
  assign n8114 = ~n8112 & ~n8113;
  assign n8115 = n8114 ^ n7822;
  assign n8116 = n8093 & n8115;
  assign n8117 = n8116 ^ n7822;
  assign n8118 = ~n8109 & ~n8117;
  assign n8119 = n8118 ^ x19;
  assign n8120 = n8119 ^ x66;
  assign n8121 = x64 & n8093;
  assign n8122 = n8121 ^ x18;
  assign n8123 = n8122 ^ x65;
  assign n8124 = ~x17 & x64;
  assign n8125 = n8124 ^ n8122;
  assign n8126 = ~n8123 & n8125;
  assign n8127 = n8126 ^ x65;
  assign n8128 = n8127 ^ n8119;
  assign n8129 = n8120 & ~n8128;
  assign n8130 = n8129 ^ x66;
  assign n8131 = n8130 ^ x67;
  assign n8132 = n7834 ^ x66;
  assign n8133 = n8093 & ~n8132;
  assign n8134 = n8133 ^ n7820;
  assign n8135 = n8134 ^ n8130;
  assign n8136 = n8131 & ~n8135;
  assign n8137 = n8136 ^ x67;
  assign n8138 = n8137 ^ x68;
  assign n8139 = n7838 & n8093;
  assign n8140 = n8139 ^ n7848;
  assign n8141 = n8140 ^ n8137;
  assign n8142 = n8138 & n8141;
  assign n8143 = n8142 ^ x68;
  assign n8144 = n8143 ^ x69;
  assign n8094 = n7943 & n8093;
  assign n8095 = n8094 ^ n7945;
  assign n8096 = ~x85 & n8095;
  assign n8097 = n7949 & n8093;
  assign n8098 = n8097 ^ n7951;
  assign n8099 = ~x86 & ~n8098;
  assign n8100 = ~n8096 & ~n8099;
  assign n8145 = n7852 & n8093;
  assign n8146 = n8145 ^ n7854;
  assign n8147 = n8146 ^ n8143;
  assign n8148 = n8144 & n8147;
  assign n8149 = n8148 ^ x69;
  assign n8150 = n8149 ^ x70;
  assign n8151 = n7858 & n8093;
  assign n8152 = n8151 ^ n7860;
  assign n8153 = n8152 ^ n8149;
  assign n8154 = n8150 & n8153;
  assign n8155 = n8154 ^ x70;
  assign n8156 = n8155 ^ x71;
  assign n8157 = n7864 & n8093;
  assign n8158 = n8157 ^ n7866;
  assign n8159 = n8158 ^ n8155;
  assign n8160 = n8156 & ~n8159;
  assign n8161 = n8160 ^ x71;
  assign n8162 = n8161 ^ x72;
  assign n8163 = n7870 & n8093;
  assign n8164 = n8163 ^ n7872;
  assign n8165 = n8164 ^ n8161;
  assign n8166 = n8162 & n8165;
  assign n8167 = n8166 ^ x72;
  assign n8168 = n8167 ^ x73;
  assign n8169 = n7876 & n8093;
  assign n8170 = n8169 ^ n7878;
  assign n8171 = n8170 ^ n8167;
  assign n8172 = n8168 & ~n8171;
  assign n8173 = n8172 ^ x73;
  assign n8174 = n8173 ^ x74;
  assign n8175 = n7884 ^ x73;
  assign n8176 = n8175 ^ n7881;
  assign n8177 = n8176 ^ n7884;
  assign n8178 = n8093 & n8177;
  assign n8179 = n8178 ^ n7884;
  assign n8180 = n8179 ^ n8173;
  assign n8181 = n8174 & ~n8180;
  assign n8182 = n8181 ^ x74;
  assign n8183 = n8182 ^ x75;
  assign n8184 = n7888 & n8093;
  assign n8185 = n8184 ^ n7890;
  assign n8186 = n8185 ^ n8182;
  assign n8187 = n8183 & n8186;
  assign n8188 = n8187 ^ x75;
  assign n8189 = n8188 ^ x76;
  assign n8190 = n7894 & n8093;
  assign n8191 = n8190 ^ n7896;
  assign n8192 = n8191 ^ n8188;
  assign n8193 = n8189 & n8192;
  assign n8194 = n8193 ^ x76;
  assign n8195 = n8194 ^ x77;
  assign n8196 = n7900 & n8093;
  assign n8197 = n8196 ^ n7902;
  assign n8198 = n8197 ^ n8194;
  assign n8199 = n8195 & ~n8198;
  assign n8200 = n8199 ^ x77;
  assign n8201 = n8200 ^ x78;
  assign n8202 = n7906 & n8093;
  assign n8203 = n8202 ^ n7908;
  assign n8204 = n8203 ^ n8200;
  assign n8205 = n8201 & n8204;
  assign n8206 = n8205 ^ x78;
  assign n8207 = n8206 ^ x79;
  assign n8208 = n7912 & n8093;
  assign n8209 = n8208 ^ n7914;
  assign n8210 = n8209 ^ n8206;
  assign n8211 = n8207 & n8210;
  assign n8212 = n8211 ^ x79;
  assign n8213 = n8212 ^ x80;
  assign n8214 = n7918 & n8093;
  assign n8215 = n8214 ^ n7920;
  assign n8216 = n8215 ^ n8212;
  assign n8217 = n8213 & ~n8216;
  assign n8218 = n8217 ^ x80;
  assign n8219 = n8218 ^ x81;
  assign n8220 = n7923 ^ x80;
  assign n8221 = n8093 & n8220;
  assign n8222 = n8221 ^ n7797;
  assign n8223 = n8222 ^ n8218;
  assign n8224 = n8219 & n8223;
  assign n8225 = n8224 ^ x81;
  assign n8226 = n8225 ^ x82;
  assign n8227 = n7923 ^ n7797;
  assign n8228 = n8220 & n8227;
  assign n8229 = n8228 ^ x80;
  assign n8230 = n8229 ^ x81;
  assign n8231 = n8093 & n8230;
  assign n8232 = n8231 ^ n7800;
  assign n8233 = n8232 ^ n8225;
  assign n8234 = n8226 & n8233;
  assign n8235 = n8234 ^ x82;
  assign n8236 = n8235 ^ x83;
  assign n8237 = n7931 & n8093;
  assign n8238 = n8237 ^ n7933;
  assign n8239 = n8238 ^ n8235;
  assign n8240 = n8236 & n8239;
  assign n8241 = n8240 ^ x83;
  assign n8242 = n8241 ^ x84;
  assign n8243 = n7937 & n8093;
  assign n8244 = n8243 ^ n7939;
  assign n8245 = n8244 ^ n8241;
  assign n8246 = n8242 & ~n8245;
  assign n8247 = n8246 ^ x84;
  assign n8248 = n8100 & n8247;
  assign n8249 = n8098 ^ x86;
  assign n8250 = x85 & ~n8095;
  assign n8251 = n8250 ^ n8098;
  assign n8252 = n8249 & ~n8251;
  assign n8253 = n8252 ^ x86;
  assign n8254 = ~n8248 & ~n8253;
  assign n8255 = n8254 ^ x87;
  assign n8256 = n7955 & n8093;
  assign n8257 = n8256 ^ n7957;
  assign n8258 = n8257 ^ n8254;
  assign n8259 = ~n8255 & n8258;
  assign n8260 = n8259 ^ x87;
  assign n8261 = n8260 ^ x88;
  assign n8262 = n7961 & n8093;
  assign n8263 = n8262 ^ n7963;
  assign n8264 = n8263 ^ n8260;
  assign n8265 = n8261 & ~n8264;
  assign n8266 = n8265 ^ x88;
  assign n8267 = n8266 ^ x89;
  assign n8268 = n7967 & n8093;
  assign n8269 = n8268 ^ n7969;
  assign n8270 = n8269 ^ n8266;
  assign n8271 = n8267 & ~n8270;
  assign n8272 = n8271 ^ x89;
  assign n8273 = n8272 ^ x90;
  assign n8274 = n7973 & n8093;
  assign n8275 = n8274 ^ n7975;
  assign n8276 = n8275 ^ n8272;
  assign n8277 = n8273 & ~n8276;
  assign n8278 = n8277 ^ x90;
  assign n8279 = n8278 ^ x91;
  assign n8280 = n7979 & n8093;
  assign n8281 = n8280 ^ n7981;
  assign n8282 = n8281 ^ n8278;
  assign n8283 = n8279 & ~n8282;
  assign n8284 = n8283 ^ x91;
  assign n8285 = n8284 ^ x92;
  assign n8286 = n7985 & n8093;
  assign n8287 = n8286 ^ n7987;
  assign n8288 = n8287 ^ n8284;
  assign n8289 = n8285 & ~n8288;
  assign n8290 = n8289 ^ x92;
  assign n8291 = n8290 ^ x93;
  assign n8292 = n7991 & n8093;
  assign n8293 = n8292 ^ n7993;
  assign n8294 = n8293 ^ n8290;
  assign n8295 = n8291 & ~n8294;
  assign n8296 = n8295 ^ x93;
  assign n8297 = n8296 ^ x94;
  assign n8298 = n7997 & n8093;
  assign n8299 = n8298 ^ n7999;
  assign n8300 = n8299 ^ n8296;
  assign n8301 = n8297 & n8300;
  assign n8302 = n8301 ^ x94;
  assign n8303 = n8302 ^ x95;
  assign n8304 = n8003 & n8093;
  assign n8305 = n8304 ^ n8005;
  assign n8306 = n8305 ^ n8302;
  assign n8307 = n8303 & ~n8306;
  assign n8308 = n8307 ^ x95;
  assign n8309 = n8308 ^ x96;
  assign n8310 = n8009 & n8093;
  assign n8311 = n8310 ^ n8011;
  assign n8312 = n8311 ^ n8308;
  assign n8313 = n8309 & n8312;
  assign n8314 = n8313 ^ x96;
  assign n8315 = n8314 ^ x97;
  assign n8316 = n8015 & n8093;
  assign n8317 = n8316 ^ n8017;
  assign n8318 = n8317 ^ n8314;
  assign n8319 = n8315 & ~n8318;
  assign n8320 = n8319 ^ x97;
  assign n8321 = n8320 ^ x98;
  assign n8322 = n8020 ^ x97;
  assign n8323 = n8093 & n8322;
  assign n8324 = n8323 ^ n7790;
  assign n8325 = n8324 ^ n8320;
  assign n8326 = n8321 & ~n8325;
  assign n8327 = n8326 ^ x98;
  assign n8328 = n8327 ^ x99;
  assign n8329 = n8020 ^ n7790;
  assign n8330 = n8322 & ~n8329;
  assign n8331 = n8330 ^ x97;
  assign n8332 = n8331 ^ x98;
  assign n8333 = n8093 & n8332;
  assign n8334 = n8333 ^ n7793;
  assign n8335 = n8334 ^ n8327;
  assign n8336 = n8328 & n8335;
  assign n8337 = n8336 ^ x99;
  assign n8338 = n8337 ^ x100;
  assign n8339 = n8027 ^ x99;
  assign n8340 = n8093 & n8339;
  assign n8341 = n8340 ^ n8029;
  assign n8342 = n8341 ^ n8337;
  assign n8343 = n8338 & n8342;
  assign n8344 = n8343 ^ x100;
  assign n8345 = n8344 ^ x101;
  assign n8346 = n8029 ^ n8027;
  assign n8347 = n8339 & n8346;
  assign n8348 = n8347 ^ x99;
  assign n8349 = n8348 ^ x100;
  assign n8350 = n8093 & n8349;
  assign n8351 = n8350 ^ n8032;
  assign n8352 = n8351 ^ n8344;
  assign n8353 = n8345 & n8352;
  assign n8354 = n8353 ^ x101;
  assign n8355 = n8354 ^ x102;
  assign n8356 = ~n8042 & n8093;
  assign n8357 = n8356 ^ n8044;
  assign n8358 = n8357 ^ n8354;
  assign n8359 = n8355 & ~n8358;
  assign n8360 = n8359 ^ x102;
  assign n8361 = n8360 ^ x103;
  assign n8362 = n8048 & n8093;
  assign n8363 = n8362 ^ n8050;
  assign n8364 = n8363 ^ n8360;
  assign n8365 = n8361 & ~n8364;
  assign n8366 = n8365 ^ x103;
  assign n8367 = n8366 ^ x104;
  assign n8368 = n8054 & n8093;
  assign n8369 = n8368 ^ n8056;
  assign n8370 = n8369 ^ n8366;
  assign n8371 = n8367 & ~n8370;
  assign n8372 = n8371 ^ x104;
  assign n8373 = n8372 ^ x105;
  assign n8374 = n8060 & n8093;
  assign n8375 = n8374 ^ n8062;
  assign n8376 = n8375 ^ n8372;
  assign n8377 = n8373 & ~n8376;
  assign n8378 = n8377 ^ x105;
  assign n8379 = n8378 ^ x106;
  assign n8380 = n8066 & n8093;
  assign n8381 = n8380 ^ n8068;
  assign n8382 = n8381 ^ n8378;
  assign n8383 = n8379 & ~n8382;
  assign n8384 = n8383 ^ x106;
  assign n8385 = n8384 ^ x107;
  assign n8386 = n8071 ^ x106;
  assign n8387 = n8093 & n8386;
  assign n8388 = n8387 ^ n7783;
  assign n8389 = n8388 ^ n8384;
  assign n8390 = n8385 & n8389;
  assign n8391 = n8390 ^ x107;
  assign n8392 = n8391 ^ x108;
  assign n8393 = n8071 ^ n7783;
  assign n8394 = n8386 & n8393;
  assign n8395 = n8394 ^ x106;
  assign n8396 = n8395 ^ x107;
  assign n8397 = n8093 & n8396;
  assign n8398 = n8397 ^ n7786;
  assign n8399 = n8398 ^ n8391;
  assign n8400 = n8392 & ~n8399;
  assign n8401 = n8400 ^ x108;
  assign n8402 = n8401 ^ x109;
  assign n8403 = ~n8079 & n8093;
  assign n8404 = n8403 ^ n8082;
  assign n8405 = n8404 ^ n8401;
  assign n8406 = n8402 & n8405;
  assign n8407 = n8406 ^ x109;
  assign n8408 = n145 & ~n8407;
  assign n8409 = ~n146 & ~n8408;
  assign n8086 = n8085 ^ x109;
  assign n8087 = n146 & n8086;
  assign n8088 = n7774 & ~n8087;
  assign n8410 = ~x110 & ~n8407;
  assign n8414 = ~n8088 & ~n8410;
  assign n8415 = ~n8409 & ~n8414;
  assign n8440 = n8144 & n8415;
  assign n8441 = n8440 ^ n8146;
  assign n8442 = n8441 ^ x70;
  assign n8443 = n8138 & n8415;
  assign n8444 = n8443 ^ n8140;
  assign n8445 = x69 & ~n8444;
  assign n8446 = n8445 ^ n8441;
  assign n8447 = n8446 ^ n8441;
  assign n8448 = ~x69 & n8444;
  assign n8449 = ~n8122 & ~n8415;
  assign n8450 = ~x16 & x65;
  assign n8451 = n8449 & n8450;
  assign n8452 = x17 & n8415;
  assign n8453 = x16 & ~x65;
  assign n8454 = ~n8123 & ~n8453;
  assign n8455 = n8452 & n8454;
  assign n8456 = ~n8451 & ~n8455;
  assign n8457 = x64 & ~n8456;
  assign n8458 = x64 & n8415;
  assign n8459 = ~x17 & x65;
  assign n8460 = ~n8458 & n8459;
  assign n8461 = n8415 ^ n8122;
  assign n8462 = n8460 & ~n8461;
  assign n8463 = ~x65 & n8415;
  assign n8464 = ~x16 & x64;
  assign n8465 = ~x17 & n8464;
  assign n8466 = ~n8122 & n8465;
  assign n8467 = ~n8463 & n8466;
  assign n8468 = ~x66 & ~n8467;
  assign n8469 = ~n8462 & n8468;
  assign n8470 = ~n8457 & n8469;
  assign n8471 = x17 & ~x65;
  assign n8472 = ~n8415 & n8471;
  assign n8473 = n8464 & ~n8472;
  assign n8474 = ~x65 & ~n8124;
  assign n8475 = n8415 & ~n8474;
  assign n8476 = n8122 & ~n8459;
  assign n8477 = ~n8475 & n8476;
  assign n8478 = ~n8473 & n8477;
  assign n8479 = n8124 & ~n8450;
  assign n8480 = ~n8123 & n8479;
  assign n8481 = ~x18 & n202;
  assign n8482 = x17 & n8481;
  assign n8483 = ~n8480 & ~n8482;
  assign n8484 = n8415 & ~n8483;
  assign n8485 = ~n8478 & ~n8484;
  assign n8486 = ~n8470 & n8485;
  assign n8487 = n8486 ^ x67;
  assign n8488 = n8127 ^ x66;
  assign n8489 = n8415 & n8488;
  assign n8490 = n8489 ^ n8119;
  assign n8491 = n8490 ^ n8486;
  assign n8492 = n8487 & ~n8491;
  assign n8493 = n8492 ^ x67;
  assign n8494 = n8493 ^ x68;
  assign n8495 = n8131 & n8415;
  assign n8496 = n8495 ^ n8134;
  assign n8497 = n8496 ^ n8493;
  assign n8498 = n8494 & ~n8497;
  assign n8499 = n8498 ^ x68;
  assign n8500 = ~n8448 & n8499;
  assign n8501 = n8500 ^ n8441;
  assign n8502 = n8501 ^ n8441;
  assign n8503 = ~n8447 & ~n8502;
  assign n8504 = n8503 ^ n8441;
  assign n8505 = ~n8442 & ~n8504;
  assign n8506 = n8505 ^ x70;
  assign n8507 = n8506 ^ x71;
  assign n8508 = n8150 & n8415;
  assign n8509 = n8508 ^ n8152;
  assign n8510 = n8509 ^ n8506;
  assign n8511 = n8507 & n8510;
  assign n8512 = n8511 ^ x71;
  assign n8513 = n8512 ^ x72;
  assign n8514 = n8156 & n8415;
  assign n8515 = n8514 ^ n8158;
  assign n8516 = n8515 ^ n8512;
  assign n8517 = n8513 & ~n8516;
  assign n8518 = n8517 ^ x72;
  assign n8519 = n8518 ^ x73;
  assign n8520 = n8162 & n8415;
  assign n8521 = n8520 ^ n8164;
  assign n8522 = n8521 ^ n8518;
  assign n8523 = n8519 & n8522;
  assign n8524 = n8523 ^ x73;
  assign n8525 = n8524 ^ x74;
  assign n8526 = n8168 & n8415;
  assign n8527 = n8526 ^ n8170;
  assign n8528 = n8527 ^ n8524;
  assign n8529 = n8525 & ~n8528;
  assign n8530 = n8529 ^ x74;
  assign n8531 = n8530 ^ x75;
  assign n8532 = n8174 & n8415;
  assign n8533 = n8532 ^ n8179;
  assign n8534 = n8533 ^ n8530;
  assign n8535 = n8531 & ~n8534;
  assign n8536 = n8535 ^ x75;
  assign n8537 = n8536 ^ x76;
  assign n8538 = n8183 & n8415;
  assign n8539 = n8538 ^ n8185;
  assign n8540 = n8539 ^ n8536;
  assign n8541 = n8537 & n8540;
  assign n8542 = n8541 ^ x76;
  assign n8543 = n8542 ^ x77;
  assign n8544 = n8189 & n8415;
  assign n8545 = n8544 ^ n8191;
  assign n8546 = n8545 ^ n8542;
  assign n8547 = n8543 & n8546;
  assign n8548 = n8547 ^ x77;
  assign n8549 = n8548 ^ x78;
  assign n8550 = n8195 & n8415;
  assign n8551 = n8550 ^ n8197;
  assign n8552 = n8551 ^ n8548;
  assign n8553 = n8549 & ~n8552;
  assign n8554 = n8553 ^ x78;
  assign n8555 = n8554 ^ x79;
  assign n8556 = n8201 & n8415;
  assign n8557 = n8556 ^ n8203;
  assign n8558 = n8557 ^ n8554;
  assign n8559 = n8555 & n8558;
  assign n8560 = n8559 ^ x79;
  assign n8561 = n8560 ^ x80;
  assign n8416 = n8402 & n8415;
  assign n8417 = n8416 ^ n8404;
  assign n8418 = x110 & ~n8417;
  assign n8419 = n8379 & n8415;
  assign n8420 = n8419 ^ n8381;
  assign n8421 = n8420 ^ x107;
  assign n8422 = n8373 & n8415;
  assign n8423 = n8422 ^ n8375;
  assign n8424 = x106 & n8423;
  assign n8425 = n8338 & n8415;
  assign n8426 = n8425 ^ n8341;
  assign n8427 = n8426 ^ x101;
  assign n8428 = n8328 & n8415;
  assign n8429 = n8428 ^ n8334;
  assign n8430 = x100 & ~n8429;
  assign n8431 = n8430 ^ n8426;
  assign n8432 = n8431 ^ n8426;
  assign n8433 = ~x100 & n8429;
  assign n8434 = n8297 & n8415;
  assign n8435 = n8434 ^ n8299;
  assign n8436 = n8435 ^ x95;
  assign n8437 = n8291 & n8415;
  assign n8438 = n8437 ^ n8293;
  assign n8439 = x94 & n8438;
  assign n8562 = n8207 & n8415;
  assign n8563 = n8562 ^ n8209;
  assign n8564 = n8563 ^ n8560;
  assign n8565 = n8561 & n8564;
  assign n8566 = n8565 ^ x80;
  assign n8567 = n8566 ^ x81;
  assign n8568 = n8213 & n8415;
  assign n8569 = n8568 ^ n8215;
  assign n8570 = n8569 ^ n8566;
  assign n8571 = n8567 & ~n8570;
  assign n8572 = n8571 ^ x81;
  assign n8573 = n8572 ^ x82;
  assign n8574 = n8219 & n8415;
  assign n8575 = n8574 ^ n8222;
  assign n8576 = n8575 ^ n8572;
  assign n8577 = n8573 & n8576;
  assign n8578 = n8577 ^ x82;
  assign n8579 = n8578 ^ x83;
  assign n8580 = n8226 & n8415;
  assign n8581 = n8580 ^ n8232;
  assign n8582 = n8581 ^ n8578;
  assign n8583 = n8579 & n8582;
  assign n8584 = n8583 ^ x83;
  assign n8585 = n8584 ^ x84;
  assign n8586 = n8236 & n8415;
  assign n8587 = n8586 ^ n8238;
  assign n8588 = n8587 ^ n8584;
  assign n8589 = n8585 & n8588;
  assign n8590 = n8589 ^ x84;
  assign n8591 = n8590 ^ x85;
  assign n8592 = n8242 & n8415;
  assign n8593 = n8592 ^ n8244;
  assign n8594 = n8593 ^ n8590;
  assign n8595 = n8591 & ~n8594;
  assign n8596 = n8595 ^ x85;
  assign n8597 = n8596 ^ x86;
  assign n8598 = n8247 ^ x85;
  assign n8599 = n8415 & n8598;
  assign n8600 = n8599 ^ n8095;
  assign n8601 = n8600 ^ n8596;
  assign n8602 = n8597 & n8601;
  assign n8603 = n8602 ^ x86;
  assign n8604 = n8603 ^ x87;
  assign n8605 = n8247 ^ n8095;
  assign n8606 = n8598 & n8605;
  assign n8607 = n8606 ^ x85;
  assign n8608 = n8607 ^ x86;
  assign n8609 = n8415 & n8608;
  assign n8610 = n8609 ^ n8098;
  assign n8611 = n8610 ^ n8603;
  assign n8612 = n8604 & ~n8611;
  assign n8613 = n8612 ^ x87;
  assign n8614 = n8613 ^ x88;
  assign n8615 = ~n8255 & n8415;
  assign n8616 = n8615 ^ n8257;
  assign n8617 = n8616 ^ n8613;
  assign n8618 = n8614 & ~n8617;
  assign n8619 = n8618 ^ x88;
  assign n8620 = n8619 ^ x89;
  assign n8621 = n8261 & n8415;
  assign n8622 = n8621 ^ n8263;
  assign n8623 = n8622 ^ n8619;
  assign n8624 = n8620 & ~n8623;
  assign n8625 = n8624 ^ x89;
  assign n8626 = n8625 ^ x90;
  assign n8627 = n8267 & n8415;
  assign n8628 = n8627 ^ n8269;
  assign n8629 = n8628 ^ n8625;
  assign n8630 = n8626 & ~n8629;
  assign n8631 = n8630 ^ x90;
  assign n8632 = n8631 ^ x91;
  assign n8633 = n8273 & n8415;
  assign n8634 = n8633 ^ n8275;
  assign n8635 = n8634 ^ n8631;
  assign n8636 = n8632 & ~n8635;
  assign n8637 = n8636 ^ x91;
  assign n8638 = n8637 ^ x92;
  assign n8639 = n8279 & n8415;
  assign n8640 = n8639 ^ n8281;
  assign n8641 = n8640 ^ n8637;
  assign n8642 = n8638 & ~n8641;
  assign n8643 = n8642 ^ x92;
  assign n8644 = n8643 ^ x93;
  assign n8645 = n8285 & n8415;
  assign n8646 = n8645 ^ n8287;
  assign n8647 = n8646 ^ n8643;
  assign n8648 = n8644 & ~n8647;
  assign n8649 = n8648 ^ x93;
  assign n8650 = ~n8439 & ~n8649;
  assign n8651 = n8650 ^ n8435;
  assign n8652 = n8651 ^ n8435;
  assign n8653 = ~x94 & ~n8438;
  assign n8654 = n8653 ^ n8435;
  assign n8655 = n8654 ^ n8435;
  assign n8656 = ~n8652 & ~n8655;
  assign n8657 = n8656 ^ n8435;
  assign n8658 = ~n8436 & n8657;
  assign n8659 = n8658 ^ x95;
  assign n8660 = n8659 ^ x96;
  assign n8661 = n8303 & n8415;
  assign n8662 = n8661 ^ n8305;
  assign n8663 = n8662 ^ n8659;
  assign n8664 = n8660 & ~n8663;
  assign n8665 = n8664 ^ x96;
  assign n8666 = n8665 ^ x97;
  assign n8667 = n8309 & n8415;
  assign n8668 = n8667 ^ n8311;
  assign n8669 = n8668 ^ n8665;
  assign n8670 = n8666 & n8669;
  assign n8671 = n8670 ^ x97;
  assign n8672 = n8671 ^ x98;
  assign n8673 = n8315 & n8415;
  assign n8674 = n8673 ^ n8317;
  assign n8675 = n8674 ^ n8671;
  assign n8676 = n8672 & ~n8675;
  assign n8677 = n8676 ^ x98;
  assign n8678 = n8677 ^ x99;
  assign n8679 = n8321 & n8415;
  assign n8680 = n8679 ^ n8324;
  assign n8681 = n8680 ^ n8677;
  assign n8682 = n8678 & ~n8681;
  assign n8683 = n8682 ^ x99;
  assign n8684 = ~n8433 & n8683;
  assign n8685 = n8684 ^ n8426;
  assign n8686 = n8685 ^ n8426;
  assign n8687 = ~n8432 & ~n8686;
  assign n8688 = n8687 ^ n8426;
  assign n8689 = ~n8427 & ~n8688;
  assign n8690 = n8689 ^ x101;
  assign n8691 = n8690 ^ x102;
  assign n8692 = n8345 & n8415;
  assign n8693 = n8692 ^ n8351;
  assign n8694 = n8693 ^ n8690;
  assign n8695 = n8691 & n8694;
  assign n8696 = n8695 ^ x102;
  assign n8697 = n8696 ^ x103;
  assign n8698 = n8355 & n8415;
  assign n8699 = n8698 ^ n8357;
  assign n8700 = n8699 ^ n8696;
  assign n8701 = n8697 & ~n8700;
  assign n8702 = n8701 ^ x103;
  assign n8703 = n8702 ^ x104;
  assign n8704 = n8361 & n8415;
  assign n8705 = n8704 ^ n8363;
  assign n8706 = n8705 ^ n8702;
  assign n8707 = n8703 & ~n8706;
  assign n8708 = n8707 ^ x104;
  assign n8709 = n8708 ^ x105;
  assign n8710 = n8367 & n8415;
  assign n8711 = n8710 ^ n8369;
  assign n8712 = n8711 ^ n8708;
  assign n8713 = n8709 & ~n8712;
  assign n8714 = n8713 ^ x105;
  assign n8715 = ~n8424 & ~n8714;
  assign n8716 = n8715 ^ n8420;
  assign n8717 = n8716 ^ n8420;
  assign n8718 = ~x106 & ~n8423;
  assign n8719 = n8718 ^ n8420;
  assign n8720 = n8719 ^ n8420;
  assign n8721 = ~n8717 & ~n8720;
  assign n8722 = n8721 ^ n8420;
  assign n8723 = n8421 & ~n8722;
  assign n8724 = n8723 ^ x107;
  assign n8725 = n8724 ^ x108;
  assign n8726 = n8385 & n8415;
  assign n8727 = n8726 ^ n8388;
  assign n8728 = n8727 ^ n8724;
  assign n8729 = n8725 & n8728;
  assign n8730 = n8729 ^ x108;
  assign n8731 = n8730 ^ x109;
  assign n8732 = n8392 & n8415;
  assign n8733 = n8732 ^ n8398;
  assign n8734 = n8733 ^ n8730;
  assign n8735 = n8731 & ~n8734;
  assign n8736 = n8735 ^ x109;
  assign n8737 = ~n8418 & ~n8736;
  assign n8738 = ~x110 & n8417;
  assign n8739 = ~n8737 & ~n8738;
  assign n8740 = n8088 & ~n8739;
  assign n8411 = ~n8409 & ~n8410;
  assign n8412 = n8088 & ~n8411;
  assign n8741 = ~n8412 & ~n8738;
  assign n8742 = ~n8737 & n8741;
  assign n8743 = ~x111 & ~n8742;
  assign n8744 = ~n8740 & ~n8743;
  assign n8413 = n141 & n143;
  assign n8745 = ~x112 & n8413;
  assign n8746 = ~n8744 & n8745;
  assign n8766 = n8561 & n8746;
  assign n8767 = n8766 ^ n8563;
  assign n8768 = ~x81 & n8767;
  assign n8769 = n8567 & n8746;
  assign n8770 = n8769 ^ n8569;
  assign n8771 = ~x82 & ~n8770;
  assign n8772 = ~n8768 & ~n8771;
  assign n8773 = x65 & n8745;
  assign n8774 = x16 & n8773;
  assign n8775 = ~n8415 & n8774;
  assign n8776 = ~n8744 & n8775;
  assign n8777 = n8453 & n8458;
  assign n8778 = ~n8776 & ~n8777;
  assign n8779 = n8746 ^ n8458;
  assign n8780 = n8779 ^ n8458;
  assign n8781 = ~x16 & ~n8463;
  assign n8782 = ~n288 & ~n8415;
  assign n8783 = n8781 & ~n8782;
  assign n8784 = ~n202 & ~n8783;
  assign n8785 = n8784 ^ n8458;
  assign n8786 = n8780 & ~n8785;
  assign n8787 = n8786 ^ n8458;
  assign n8788 = n8778 & ~n8787;
  assign n8789 = n8788 ^ x17;
  assign n8790 = n8789 ^ x66;
  assign n8791 = x64 & n8746;
  assign n8792 = x15 & n8453;
  assign n8793 = n8792 ^ x16;
  assign n8794 = n8791 & n8793;
  assign n8795 = ~x15 & n8464;
  assign n8796 = ~n8450 & ~n8795;
  assign n8797 = ~n8746 & ~n8796;
  assign n8798 = ~x15 & x65;
  assign n8799 = n8798 ^ n8450;
  assign n8800 = x64 & n8799;
  assign n8801 = n8800 ^ n8450;
  assign n8802 = ~n8797 & ~n8801;
  assign n8803 = ~n8794 & n8802;
  assign n8804 = n8803 ^ n8789;
  assign n8805 = n8790 & n8804;
  assign n8806 = n8805 ^ x66;
  assign n8807 = n8806 ^ x67;
  assign n8811 = ~n8471 & n8781;
  assign n8812 = n8452 & ~n8453;
  assign n8813 = ~n8811 & ~n8812;
  assign n8814 = x64 & ~n8813;
  assign n8815 = ~n8460 & ~n8814;
  assign n8816 = n8815 ^ x66;
  assign n8817 = n8746 & ~n8816;
  assign n8808 = x65 & n8124;
  assign n8809 = n8475 & ~n8808;
  assign n8810 = n8809 ^ n8122;
  assign n8818 = n8817 ^ n8810;
  assign n8819 = n8818 ^ n8806;
  assign n8820 = n8807 & n8819;
  assign n8821 = n8820 ^ x67;
  assign n8822 = n8821 ^ x68;
  assign n8823 = n8487 & n8746;
  assign n8824 = n8823 ^ n8490;
  assign n8825 = n8824 ^ n8821;
  assign n8826 = n8822 & ~n8825;
  assign n8827 = n8826 ^ x68;
  assign n8828 = n8827 ^ x69;
  assign n8829 = n8494 & n8746;
  assign n8830 = n8829 ^ n8496;
  assign n8831 = n8830 ^ n8827;
  assign n8832 = n8828 & ~n8831;
  assign n8833 = n8832 ^ x69;
  assign n8834 = n8833 ^ x70;
  assign n8835 = n8499 ^ x69;
  assign n8836 = n8746 & n8835;
  assign n8837 = n8836 ^ n8444;
  assign n8838 = n8837 ^ n8833;
  assign n8839 = n8834 & n8838;
  assign n8840 = n8839 ^ x70;
  assign n8841 = n8840 ^ x71;
  assign n8842 = ~n8445 & ~n8500;
  assign n8843 = n8842 ^ x70;
  assign n8844 = n8746 & ~n8843;
  assign n8845 = n8844 ^ n8441;
  assign n8846 = n8845 ^ n8840;
  assign n8847 = n8841 & n8846;
  assign n8848 = n8847 ^ x71;
  assign n8849 = n8848 ^ x72;
  assign n8850 = n8507 & n8746;
  assign n8851 = n8850 ^ n8509;
  assign n8852 = n8851 ^ n8848;
  assign n8853 = n8849 & n8852;
  assign n8854 = n8853 ^ x72;
  assign n8855 = n8854 ^ x73;
  assign n8856 = n8513 & n8746;
  assign n8857 = n8856 ^ n8515;
  assign n8858 = n8857 ^ n8854;
  assign n8859 = n8855 & ~n8858;
  assign n8860 = n8859 ^ x73;
  assign n8861 = n8860 ^ x74;
  assign n8862 = n8519 & n8746;
  assign n8863 = n8862 ^ n8521;
  assign n8864 = n8863 ^ n8860;
  assign n8865 = n8861 & n8864;
  assign n8866 = n8865 ^ x74;
  assign n8867 = n8866 ^ x75;
  assign n8868 = n8525 & n8746;
  assign n8869 = n8868 ^ n8527;
  assign n8870 = n8869 ^ n8866;
  assign n8871 = n8867 & ~n8870;
  assign n8872 = n8871 ^ x75;
  assign n8873 = n8872 ^ x76;
  assign n8874 = n8531 & n8746;
  assign n8875 = n8874 ^ n8533;
  assign n8876 = n8875 ^ n8872;
  assign n8877 = n8873 & ~n8876;
  assign n8878 = n8877 ^ x76;
  assign n8879 = n8878 ^ x77;
  assign n8880 = n8537 & n8746;
  assign n8881 = n8880 ^ n8539;
  assign n8882 = n8881 ^ n8878;
  assign n8883 = n8879 & n8882;
  assign n8884 = n8883 ^ x77;
  assign n8885 = n8884 ^ x78;
  assign n8886 = n8543 & n8746;
  assign n8887 = n8886 ^ n8545;
  assign n8888 = n8887 ^ n8884;
  assign n8889 = n8885 & n8888;
  assign n8890 = n8889 ^ x78;
  assign n8891 = n8890 ^ x79;
  assign n8892 = n8549 & n8746;
  assign n8893 = n8892 ^ n8551;
  assign n8894 = n8893 ^ n8890;
  assign n8895 = n8891 & ~n8894;
  assign n8896 = n8895 ^ x79;
  assign n8897 = n8896 ^ x80;
  assign n8898 = n8555 & n8746;
  assign n8899 = n8898 ^ n8557;
  assign n8900 = n8899 ^ n8896;
  assign n8901 = n8897 & n8900;
  assign n8902 = n8901 ^ x80;
  assign n8903 = n8772 & n8902;
  assign n8904 = n8770 ^ x82;
  assign n8905 = x81 & ~n8767;
  assign n8906 = n8905 ^ n8770;
  assign n8907 = n8904 & ~n8906;
  assign n8908 = n8907 ^ x82;
  assign n8909 = ~n8903 & ~n8908;
  assign n8910 = n8909 ^ x83;
  assign n8911 = n8573 & n8746;
  assign n8912 = n8911 ^ n8575;
  assign n8913 = n8912 ^ n8909;
  assign n8914 = ~n8910 & ~n8913;
  assign n8915 = n8914 ^ x83;
  assign n8916 = n8915 ^ x84;
  assign n8917 = n8579 & n8746;
  assign n8918 = n8917 ^ n8581;
  assign n8919 = n8918 ^ n8915;
  assign n8920 = n8916 & n8919;
  assign n8921 = n8920 ^ x84;
  assign n8922 = n8921 ^ x85;
  assign n8923 = n8585 & n8746;
  assign n8924 = n8923 ^ n8587;
  assign n8925 = n8924 ^ n8921;
  assign n8926 = n8922 & n8925;
  assign n8927 = n8926 ^ x85;
  assign n8928 = n8927 ^ x86;
  assign n8929 = n8591 & n8746;
  assign n8930 = n8929 ^ n8593;
  assign n8931 = n8930 ^ n8927;
  assign n8932 = n8928 & ~n8931;
  assign n8933 = n8932 ^ x86;
  assign n8934 = n8933 ^ x87;
  assign n8747 = n8736 ^ x110;
  assign n8748 = n8746 & n8747;
  assign n8749 = n8748 ^ n8417;
  assign n8750 = n8731 & n8746;
  assign n8751 = n8750 ^ n8733;
  assign n8752 = n8751 ^ x110;
  assign n8753 = n8725 & n8746;
  assign n8754 = n8753 ^ n8727;
  assign n8755 = x109 & ~n8754;
  assign n8756 = n8755 ^ n8751;
  assign n8757 = n8756 ^ n8751;
  assign n8758 = ~x109 & n8754;
  assign n8759 = n8697 & n8746;
  assign n8760 = n8759 ^ n8699;
  assign n8761 = ~x104 & ~n8760;
  assign n8762 = n8703 & n8746;
  assign n8763 = n8762 ^ n8705;
  assign n8764 = ~x105 & ~n8763;
  assign n8765 = ~n8761 & ~n8764;
  assign n8935 = n8597 & n8746;
  assign n8936 = n8935 ^ n8600;
  assign n8937 = n8936 ^ n8933;
  assign n8938 = n8934 & n8937;
  assign n8939 = n8938 ^ x87;
  assign n8940 = n8939 ^ x88;
  assign n8941 = n8604 & n8746;
  assign n8942 = n8941 ^ n8610;
  assign n8943 = n8942 ^ n8939;
  assign n8944 = n8940 & ~n8943;
  assign n8945 = n8944 ^ x88;
  assign n8946 = n8945 ^ x89;
  assign n8947 = n8614 & n8746;
  assign n8948 = n8947 ^ n8616;
  assign n8949 = n8948 ^ n8945;
  assign n8950 = n8946 & ~n8949;
  assign n8951 = n8950 ^ x89;
  assign n8952 = n8951 ^ x90;
  assign n8953 = n8620 & n8746;
  assign n8954 = n8953 ^ n8622;
  assign n8955 = n8954 ^ n8951;
  assign n8956 = n8952 & ~n8955;
  assign n8957 = n8956 ^ x90;
  assign n8958 = n8957 ^ x91;
  assign n8959 = n8626 & n8746;
  assign n8960 = n8959 ^ n8628;
  assign n8961 = n8960 ^ n8957;
  assign n8962 = n8958 & ~n8961;
  assign n8963 = n8962 ^ x91;
  assign n8964 = n8963 ^ x92;
  assign n8965 = n8632 & n8746;
  assign n8966 = n8965 ^ n8634;
  assign n8967 = n8966 ^ n8963;
  assign n8968 = n8964 & ~n8967;
  assign n8969 = n8968 ^ x92;
  assign n8970 = n8969 ^ x93;
  assign n8971 = n8638 & n8746;
  assign n8972 = n8971 ^ n8640;
  assign n8973 = n8972 ^ n8969;
  assign n8974 = n8970 & ~n8973;
  assign n8975 = n8974 ^ x93;
  assign n8976 = n8975 ^ x94;
  assign n8977 = n8644 & n8746;
  assign n8978 = n8977 ^ n8646;
  assign n8979 = n8978 ^ n8975;
  assign n8980 = n8976 & ~n8979;
  assign n8981 = n8980 ^ x94;
  assign n8982 = n8981 ^ x95;
  assign n8983 = n8649 ^ x94;
  assign n8984 = n8746 & n8983;
  assign n8985 = n8984 ^ n8438;
  assign n8986 = n8985 ^ n8981;
  assign n8987 = n8982 & ~n8986;
  assign n8988 = n8987 ^ x95;
  assign n8989 = n8988 ^ x96;
  assign n8990 = ~n8650 & ~n8653;
  assign n8991 = n8990 ^ x95;
  assign n8992 = n8746 & n8991;
  assign n8993 = n8992 ^ n8435;
  assign n8994 = n8993 ^ n8988;
  assign n8995 = n8989 & n8994;
  assign n8996 = n8995 ^ x96;
  assign n8997 = n8996 ^ x97;
  assign n8998 = n8660 & n8746;
  assign n8999 = n8998 ^ n8662;
  assign n9000 = n8999 ^ n8996;
  assign n9001 = n8997 & ~n9000;
  assign n9002 = n9001 ^ x97;
  assign n9003 = n9002 ^ x98;
  assign n9004 = n8666 & n8746;
  assign n9005 = n9004 ^ n8668;
  assign n9006 = n9005 ^ n9002;
  assign n9007 = n9003 & n9006;
  assign n9008 = n9007 ^ x98;
  assign n9009 = n9008 ^ x99;
  assign n9010 = n8672 & n8746;
  assign n9011 = n9010 ^ n8674;
  assign n9012 = n9011 ^ n9008;
  assign n9013 = n9009 & ~n9012;
  assign n9014 = n9013 ^ x99;
  assign n9015 = n9014 ^ x100;
  assign n9016 = n8678 & n8746;
  assign n9017 = n9016 ^ n8680;
  assign n9018 = n9017 ^ n9014;
  assign n9019 = n9015 & ~n9018;
  assign n9020 = n9019 ^ x100;
  assign n9021 = n9020 ^ x101;
  assign n9022 = n8683 ^ x100;
  assign n9023 = n8746 & n9022;
  assign n9024 = n9023 ^ n8429;
  assign n9025 = n9024 ^ n9020;
  assign n9026 = n9021 & n9025;
  assign n9027 = n9026 ^ x101;
  assign n9028 = n9027 ^ x102;
  assign n9029 = ~n8430 & ~n8684;
  assign n9030 = n9029 ^ x101;
  assign n9031 = n8746 & ~n9030;
  assign n9032 = n9031 ^ n8426;
  assign n9033 = n9032 ^ n9027;
  assign n9034 = n9028 & n9033;
  assign n9035 = n9034 ^ x102;
  assign n9036 = n9035 ^ x103;
  assign n9037 = n8691 & n8746;
  assign n9038 = n9037 ^ n8693;
  assign n9039 = n9038 ^ n9035;
  assign n9040 = n9036 & n9039;
  assign n9041 = n9040 ^ x103;
  assign n9042 = n8765 & n9041;
  assign n9043 = n8763 ^ x105;
  assign n9044 = x104 & n8760;
  assign n9045 = n9044 ^ n8763;
  assign n9046 = n9043 & ~n9045;
  assign n9047 = n9046 ^ x105;
  assign n9048 = ~n9042 & ~n9047;
  assign n9049 = n9048 ^ x106;
  assign n9050 = n8709 & n8746;
  assign n9051 = n9050 ^ n8711;
  assign n9052 = n9051 ^ n9048;
  assign n9053 = ~n9049 & n9052;
  assign n9054 = n9053 ^ x106;
  assign n9055 = n9054 ^ x107;
  assign n9056 = n8714 ^ x106;
  assign n9057 = n8746 & n9056;
  assign n9058 = n9057 ^ n8423;
  assign n9059 = n9058 ^ n9054;
  assign n9060 = n9055 & ~n9059;
  assign n9061 = n9060 ^ x107;
  assign n9062 = n9061 ^ x108;
  assign n9063 = ~n8715 & ~n8718;
  assign n9064 = n9063 ^ x107;
  assign n9065 = n8746 & n9064;
  assign n9066 = n9065 ^ n8420;
  assign n9067 = n9066 ^ n9061;
  assign n9068 = n9062 & ~n9067;
  assign n9069 = n9068 ^ x108;
  assign n9070 = ~n8758 & n9069;
  assign n9071 = n9070 ^ n8751;
  assign n9072 = n9071 ^ n8751;
  assign n9073 = ~n8757 & ~n9072;
  assign n9074 = n9073 ^ n8751;
  assign n9075 = n8752 & n9074;
  assign n9076 = n9075 ^ x110;
  assign n9077 = ~n8749 & n9076;
  assign n9078 = ~x111 & ~n9077;
  assign n9080 = n8749 & ~n9076;
  assign n9081 = ~n9078 & ~n9080;
  assign n9088 = n7774 & n8413;
  assign n9089 = ~n9081 & n9088;
  assign n9090 = ~x111 & n8739;
  assign n9091 = n8746 & n9090;
  assign n9092 = n8412 & ~n9091;
  assign n9093 = n9077 & ~n9092;
  assign n9094 = n8745 & ~n9093;
  assign n9095 = ~n8739 & n8746;
  assign n9096 = n8412 & ~n9095;
  assign n9097 = x111 & ~n9096;
  assign n9098 = ~n9080 & n9097;
  assign n9099 = n9094 & ~n9098;
  assign n9100 = ~n9089 & ~n9099;
  assign n9101 = n8934 & ~n9100;
  assign n9102 = n9101 ^ n8936;
  assign n9103 = ~x88 & n9102;
  assign n9104 = n8940 & ~n9100;
  assign n9105 = n9104 ^ n8942;
  assign n9106 = ~x89 & ~n9105;
  assign n9107 = ~n9103 & ~n9106;
  assign n9108 = n8922 & ~n9100;
  assign n9109 = n9108 ^ n8924;
  assign n9110 = n9109 ^ x86;
  assign n9111 = n8916 & ~n9100;
  assign n9112 = n9111 ^ n8918;
  assign n9113 = x85 & ~n9112;
  assign n9114 = n8867 & ~n9100;
  assign n9115 = n9114 ^ n8869;
  assign n9116 = ~x76 & ~n9115;
  assign n9117 = n8873 & ~n9100;
  assign n9118 = n9117 ^ n8875;
  assign n9119 = ~x77 & ~n9118;
  assign n9120 = ~n9116 & ~n9119;
  assign n9121 = x64 & ~n9100;
  assign n9122 = n9121 ^ x15;
  assign n9123 = n9122 ^ x65;
  assign n9124 = ~x14 & x64;
  assign n9125 = n9124 ^ n9122;
  assign n9126 = ~n9123 & n9125;
  assign n9127 = n9126 ^ x65;
  assign n9128 = n9127 ^ x66;
  assign n9129 = ~n8744 & n8773;
  assign n9130 = n9129 ^ x15;
  assign n9131 = n9130 ^ n9129;
  assign n9132 = n288 & ~n8746;
  assign n9133 = ~n9129 & ~n9132;
  assign n9134 = n9133 ^ n9129;
  assign n9135 = ~n9131 & n9134;
  assign n9136 = n9135 ^ n9129;
  assign n9137 = ~n202 & n9136;
  assign n9138 = n9137 ^ n8791;
  assign n9139 = ~x15 & ~n9133;
  assign n9140 = ~x65 & ~n9139;
  assign n9141 = n9140 ^ n9137;
  assign n9142 = n9137 ^ n9100;
  assign n9143 = ~n9137 & n9142;
  assign n9144 = n9143 ^ n9137;
  assign n9145 = ~n9141 & ~n9144;
  assign n9146 = n9145 ^ n9143;
  assign n9147 = n9146 ^ n9137;
  assign n9148 = n9147 ^ n9100;
  assign n9149 = ~n9138 & n9148;
  assign n9150 = n9149 ^ n8791;
  assign n9151 = n9150 ^ x16;
  assign n9152 = n9151 ^ n9127;
  assign n9153 = n9128 & n9152;
  assign n9154 = n9153 ^ x66;
  assign n9155 = n9154 ^ x67;
  assign n9156 = n8803 ^ x66;
  assign n9157 = ~n9100 & ~n9156;
  assign n9158 = n9157 ^ n8789;
  assign n9159 = n9158 ^ n9154;
  assign n9160 = n9155 & ~n9159;
  assign n9161 = n9160 ^ x67;
  assign n9162 = n9161 ^ x68;
  assign n9163 = n8807 & ~n9100;
  assign n9164 = n9163 ^ n8818;
  assign n9165 = n9164 ^ n9161;
  assign n9166 = n9162 & n9165;
  assign n9167 = n9166 ^ x68;
  assign n9168 = n9167 ^ x69;
  assign n9169 = n8822 & ~n9100;
  assign n9170 = n9169 ^ n8824;
  assign n9171 = n9170 ^ n9167;
  assign n9172 = n9168 & ~n9171;
  assign n9173 = n9172 ^ x69;
  assign n9174 = n9173 ^ x70;
  assign n9175 = n8828 & ~n9100;
  assign n9176 = n9175 ^ n8830;
  assign n9177 = n9176 ^ n9173;
  assign n9178 = n9174 & ~n9177;
  assign n9179 = n9178 ^ x70;
  assign n9180 = n9179 ^ x71;
  assign n9181 = n8834 & ~n9100;
  assign n9182 = n9181 ^ n8837;
  assign n9183 = n9182 ^ n9179;
  assign n9184 = n9180 & n9183;
  assign n9185 = n9184 ^ x71;
  assign n9186 = n9185 ^ x72;
  assign n9187 = n8841 & ~n9100;
  assign n9188 = n9187 ^ n8845;
  assign n9189 = n9188 ^ n9185;
  assign n9190 = n9186 & n9189;
  assign n9191 = n9190 ^ x72;
  assign n9192 = n9191 ^ x73;
  assign n9193 = n8849 & ~n9100;
  assign n9194 = n9193 ^ n8851;
  assign n9195 = n9194 ^ n9191;
  assign n9196 = n9192 & n9195;
  assign n9197 = n9196 ^ x73;
  assign n9198 = n9197 ^ x74;
  assign n9199 = n8855 & ~n9100;
  assign n9200 = n9199 ^ n8857;
  assign n9201 = n9200 ^ n9197;
  assign n9202 = n9198 & ~n9201;
  assign n9203 = n9202 ^ x74;
  assign n9204 = n9203 ^ x75;
  assign n9205 = n8861 & ~n9100;
  assign n9206 = n9205 ^ n8863;
  assign n9207 = n9206 ^ n9203;
  assign n9208 = n9204 & n9207;
  assign n9209 = n9208 ^ x75;
  assign n9210 = n9120 & n9209;
  assign n9211 = n9118 ^ x77;
  assign n9212 = x76 & n9115;
  assign n9213 = n9212 ^ n9118;
  assign n9214 = n9211 & ~n9213;
  assign n9215 = n9214 ^ x77;
  assign n9216 = ~n9210 & ~n9215;
  assign n9217 = n9216 ^ x78;
  assign n9218 = n8879 & ~n9100;
  assign n9219 = n9218 ^ n8881;
  assign n9220 = n9219 ^ n9216;
  assign n9221 = ~n9217 & ~n9220;
  assign n9222 = n9221 ^ x78;
  assign n9223 = n9222 ^ x79;
  assign n9224 = n8885 & ~n9100;
  assign n9225 = n9224 ^ n8887;
  assign n9226 = n9225 ^ n9222;
  assign n9227 = n9223 & n9226;
  assign n9228 = n9227 ^ x79;
  assign n9229 = n9228 ^ x80;
  assign n9230 = n8891 & ~n9100;
  assign n9231 = n9230 ^ n8893;
  assign n9232 = n9231 ^ n9228;
  assign n9233 = n9229 & ~n9232;
  assign n9234 = n9233 ^ x80;
  assign n9235 = n9234 ^ x81;
  assign n9236 = n8897 & ~n9100;
  assign n9237 = n9236 ^ n8899;
  assign n9238 = n9237 ^ n9234;
  assign n9239 = n9235 & n9238;
  assign n9240 = n9239 ^ x81;
  assign n9241 = n9240 ^ x82;
  assign n9242 = n8902 ^ x81;
  assign n9243 = ~n9100 & n9242;
  assign n9244 = n9243 ^ n8767;
  assign n9245 = n9244 ^ n9240;
  assign n9246 = n9241 & n9245;
  assign n9247 = n9246 ^ x82;
  assign n9248 = n9247 ^ x83;
  assign n9249 = n8902 ^ n8767;
  assign n9250 = n9242 & n9249;
  assign n9251 = n9250 ^ x81;
  assign n9252 = n9251 ^ x82;
  assign n9253 = ~n9100 & n9252;
  assign n9254 = n9253 ^ n8770;
  assign n9255 = n9254 ^ n9247;
  assign n9256 = n9248 & ~n9255;
  assign n9257 = n9256 ^ x83;
  assign n9258 = n9257 ^ x84;
  assign n9259 = ~n8910 & ~n9100;
  assign n9260 = n9259 ^ n8912;
  assign n9261 = n9260 ^ n9257;
  assign n9262 = n9258 & n9261;
  assign n9263 = n9262 ^ x84;
  assign n9264 = ~n9113 & ~n9263;
  assign n9265 = n9264 ^ n9109;
  assign n9266 = n9265 ^ n9109;
  assign n9267 = ~x85 & n9112;
  assign n9268 = n9267 ^ n9109;
  assign n9269 = n9268 ^ n9109;
  assign n9270 = ~n9266 & ~n9269;
  assign n9271 = n9270 ^ n9109;
  assign n9272 = ~n9110 & n9271;
  assign n9273 = n9272 ^ x86;
  assign n9274 = n9273 ^ x87;
  assign n9275 = n8928 & ~n9100;
  assign n9276 = n9275 ^ n8930;
  assign n9277 = n9276 ^ n9273;
  assign n9278 = n9274 & ~n9277;
  assign n9279 = n9278 ^ x87;
  assign n9280 = n9107 & n9279;
  assign n9281 = n9105 ^ x89;
  assign n9282 = x88 & ~n9102;
  assign n9283 = n9282 ^ n9105;
  assign n9284 = n9281 & ~n9283;
  assign n9285 = n9284 ^ x89;
  assign n9286 = ~n9280 & ~n9285;
  assign n9287 = n8946 & ~n9100;
  assign n9288 = n9287 ^ n8948;
  assign n9289 = ~x90 & ~n9288;
  assign n9290 = n8952 & ~n9100;
  assign n9291 = n9290 ^ n8954;
  assign n9292 = ~x91 & ~n9291;
  assign n9293 = ~n9289 & ~n9292;
  assign n9294 = ~n9286 & n9293;
  assign n9295 = n9291 ^ x91;
  assign n9296 = x90 & n9288;
  assign n9297 = n9296 ^ n9291;
  assign n9298 = n9295 & ~n9297;
  assign n9299 = n9298 ^ x91;
  assign n9300 = ~n9294 & ~n9299;
  assign n9301 = n9300 ^ x92;
  assign n9302 = n8958 & ~n9100;
  assign n9303 = n9302 ^ n8960;
  assign n9304 = n9303 ^ n9300;
  assign n9305 = ~n9301 & n9304;
  assign n9306 = n9305 ^ x92;
  assign n9307 = n9306 ^ x93;
  assign n9308 = n8964 & ~n9100;
  assign n9309 = n9308 ^ n8966;
  assign n9310 = n9309 ^ n9306;
  assign n9311 = n9307 & ~n9310;
  assign n9312 = n9311 ^ x93;
  assign n9313 = n9312 ^ x94;
  assign n9314 = n8970 & ~n9100;
  assign n9315 = n9314 ^ n8972;
  assign n9316 = n9315 ^ n9312;
  assign n9317 = n9313 & ~n9316;
  assign n9318 = n9317 ^ x94;
  assign n9319 = n9318 ^ x95;
  assign n9320 = n8976 & ~n9100;
  assign n9321 = n9320 ^ n8978;
  assign n9322 = n9321 ^ n9318;
  assign n9323 = n9319 & ~n9322;
  assign n9324 = n9323 ^ x95;
  assign n9325 = n9324 ^ x96;
  assign n9326 = n8982 & ~n9100;
  assign n9327 = n9326 ^ n8985;
  assign n9328 = n9327 ^ n9324;
  assign n9329 = n9325 & ~n9328;
  assign n9330 = n9329 ^ x96;
  assign n9331 = n9330 ^ x97;
  assign n9332 = n8989 & ~n9100;
  assign n9333 = n9332 ^ n8993;
  assign n9334 = n9333 ^ n9330;
  assign n9335 = n9331 & n9334;
  assign n9336 = n9335 ^ x97;
  assign n9337 = n9336 ^ x98;
  assign n9338 = n8997 & ~n9100;
  assign n9339 = n9338 ^ n8999;
  assign n9340 = n9339 ^ n9336;
  assign n9341 = n9337 & ~n9340;
  assign n9342 = n9341 ^ x98;
  assign n9343 = n9342 ^ x99;
  assign n9344 = n9003 & ~n9100;
  assign n9345 = n9344 ^ n9005;
  assign n9346 = n9345 ^ n9342;
  assign n9347 = n9343 & n9346;
  assign n9348 = n9347 ^ x99;
  assign n9349 = n9348 ^ x100;
  assign n9350 = n9009 & ~n9100;
  assign n9351 = n9350 ^ n9011;
  assign n9352 = n9351 ^ n9348;
  assign n9353 = n9349 & ~n9352;
  assign n9354 = n9353 ^ x100;
  assign n9355 = n9354 ^ x101;
  assign n9356 = n9015 & ~n9100;
  assign n9357 = n9356 ^ n9017;
  assign n9358 = n9357 ^ n9354;
  assign n9359 = n9355 & ~n9358;
  assign n9360 = n9359 ^ x101;
  assign n9361 = n9360 ^ x102;
  assign n9362 = n9021 & ~n9100;
  assign n9363 = n9362 ^ n9024;
  assign n9364 = n9363 ^ n9360;
  assign n9365 = n9361 & n9364;
  assign n9366 = n9365 ^ x102;
  assign n9367 = n9366 ^ x103;
  assign n9368 = n9028 & ~n9100;
  assign n9369 = n9368 ^ n9032;
  assign n9370 = n9369 ^ n9366;
  assign n9371 = n9367 & n9370;
  assign n9372 = n9371 ^ x103;
  assign n9373 = n9372 ^ x104;
  assign n9374 = n9036 & ~n9100;
  assign n9375 = n9374 ^ n9038;
  assign n9376 = n9375 ^ n9372;
  assign n9377 = n9373 & n9376;
  assign n9378 = n9377 ^ x104;
  assign n9379 = n9378 ^ x105;
  assign n9380 = n9041 ^ x104;
  assign n9381 = ~n9100 & n9380;
  assign n9382 = n9381 ^ n8760;
  assign n9383 = n9382 ^ n9378;
  assign n9384 = n9379 & ~n9383;
  assign n9385 = n9384 ^ x105;
  assign n9386 = n9385 ^ x106;
  assign n9387 = n9041 ^ n8760;
  assign n9388 = n9380 & ~n9387;
  assign n9389 = n9388 ^ x104;
  assign n9390 = n9389 ^ x105;
  assign n9391 = ~n9100 & n9390;
  assign n9392 = n9391 ^ n8763;
  assign n9393 = n9392 ^ n9385;
  assign n9394 = n9386 & ~n9393;
  assign n9395 = n9394 ^ x106;
  assign n9396 = n9395 ^ x107;
  assign n9397 = ~n9049 & ~n9100;
  assign n9398 = n9397 ^ n9051;
  assign n9399 = n9398 ^ n9395;
  assign n9400 = n9396 & ~n9399;
  assign n9401 = n9400 ^ x107;
  assign n9402 = n9401 ^ x108;
  assign n9403 = n9055 & ~n9100;
  assign n9404 = n9403 ^ n9058;
  assign n9405 = n9404 ^ n9401;
  assign n9406 = n9402 & ~n9405;
  assign n9407 = n9406 ^ x108;
  assign n9408 = n9407 ^ x109;
  assign n9409 = n9062 & ~n9100;
  assign n9410 = n9409 ^ n9066;
  assign n9411 = n9410 ^ n9407;
  assign n9412 = n9408 & ~n9411;
  assign n9413 = n9412 ^ x109;
  assign n9414 = n9413 ^ x110;
  assign n9415 = n9069 ^ x109;
  assign n9416 = ~n9100 & n9415;
  assign n9417 = n9416 ^ n8754;
  assign n9418 = n9417 ^ n9413;
  assign n9419 = n9414 & n9418;
  assign n9420 = n9419 ^ x110;
  assign n9421 = n9420 ^ x111;
  assign n9422 = ~n8755 & ~n9070;
  assign n9423 = n9422 ^ x110;
  assign n9424 = ~n9100 & ~n9423;
  assign n9425 = n9424 ^ n8751;
  assign n9426 = n9425 ^ n9420;
  assign n9427 = n9421 & ~n9426;
  assign n9428 = n9427 ^ x111;
  assign n9429 = n9428 ^ x112;
  assign n9430 = n9076 ^ x111;
  assign n9431 = ~n9100 & n9430;
  assign n9432 = n9431 ^ n8749;
  assign n9433 = n9432 ^ n9428;
  assign n9434 = n9429 & n9433;
  assign n9435 = n9434 ^ x112;
  assign n9436 = n9435 ^ x113;
  assign n9439 = n9435 ^ n8088;
  assign n9440 = n9439 ^ n8088;
  assign n9079 = ~n8739 & n9078;
  assign n9082 = n9081 ^ n9079;
  assign n9083 = ~x112 & n9082;
  assign n9084 = n9083 ^ n9081;
  assign n9085 = n8413 & ~n9084;
  assign n9086 = n8412 & ~n9085;
  assign n9441 = n9086 ^ n8088;
  assign n9442 = n9440 & ~n9441;
  assign n9443 = n9442 ^ n8088;
  assign n9444 = n9436 & n9443;
  assign n9445 = n9444 ^ x113;
  assign n9446 = n9087 & ~n9445;
  assign n9470 = x64 & n9446;
  assign n9471 = ~x14 & x65;
  assign n9472 = ~n9470 & n9471;
  assign n9473 = n9446 ^ n9122;
  assign n9474 = n9472 & ~n9473;
  assign n9475 = ~n9122 & ~n9446;
  assign n9476 = x14 & ~x65;
  assign n9477 = ~x13 & x64;
  assign n9478 = ~n9476 & n9477;
  assign n9479 = n9475 & n9478;
  assign n9480 = ~x66 & ~n9479;
  assign n9481 = ~n9474 & n9480;
  assign n9482 = x13 & n9476;
  assign n9483 = n9482 ^ x14;
  assign n9484 = ~n9123 & n9483;
  assign n9485 = n9446 & n9484;
  assign n9486 = ~x13 & n9471;
  assign n9487 = ~n9122 & n9486;
  assign n9488 = ~n9485 & ~n9487;
  assign n9489 = x64 & ~n9488;
  assign n9490 = n9481 & ~n9489;
  assign n9497 = ~n9471 & ~n9478;
  assign n9498 = n9122 & n9497;
  assign n9491 = ~x13 & x65;
  assign n9492 = n9124 & ~n9491;
  assign n9493 = ~n9123 & n9492;
  assign n9494 = x14 & n202;
  assign n9495 = ~n9122 & n9494;
  assign n9496 = ~n9493 & ~n9495;
  assign n9499 = n9498 ^ n9496;
  assign n9500 = ~x65 & ~n9124;
  assign n9501 = ~n9477 & n9500;
  assign n9502 = n9501 ^ n9496;
  assign n9503 = n9496 ^ n9446;
  assign n9504 = n9496 & n9503;
  assign n9505 = n9504 ^ n9496;
  assign n9506 = n9502 & n9505;
  assign n9507 = n9506 ^ n9504;
  assign n9508 = n9507 ^ n9496;
  assign n9509 = n9508 ^ n9446;
  assign n9510 = ~n9499 & n9509;
  assign n9511 = n9510 ^ n9498;
  assign n9512 = ~n9490 & ~n9511;
  assign n9513 = n9512 ^ x67;
  assign n9514 = n9128 & n9446;
  assign n9515 = n9514 ^ n9151;
  assign n9516 = n9515 ^ n9512;
  assign n9517 = n9513 & n9516;
  assign n9518 = n9517 ^ x67;
  assign n9519 = n9518 ^ x68;
  assign n9520 = n9155 & n9446;
  assign n9521 = n9520 ^ n9158;
  assign n9522 = n9521 ^ n9518;
  assign n9523 = n9519 & ~n9522;
  assign n9524 = n9523 ^ x68;
  assign n9525 = n9524 ^ x69;
  assign n9526 = n9162 & n9446;
  assign n9527 = n9526 ^ n9164;
  assign n9528 = n9527 ^ n9524;
  assign n9529 = n9525 & n9528;
  assign n9530 = n9529 ^ x69;
  assign n9531 = n9530 ^ x70;
  assign n9532 = n9168 & n9446;
  assign n9533 = n9532 ^ n9170;
  assign n9534 = n9533 ^ n9530;
  assign n9535 = n9531 & ~n9534;
  assign n9536 = n9535 ^ x70;
  assign n9537 = n9536 ^ x71;
  assign n9538 = n9174 & n9446;
  assign n9539 = n9538 ^ n9176;
  assign n9540 = n9539 ^ n9536;
  assign n9541 = n9537 & ~n9540;
  assign n9542 = n9541 ^ x71;
  assign n9543 = n9542 ^ x72;
  assign n9544 = n9180 & n9446;
  assign n9545 = n9544 ^ n9182;
  assign n9546 = n9545 ^ n9542;
  assign n9547 = n9543 & n9546;
  assign n9548 = n9547 ^ x72;
  assign n9549 = n9548 ^ x73;
  assign n9550 = n9186 & n9446;
  assign n9551 = n9550 ^ n9188;
  assign n9552 = n9551 ^ n9548;
  assign n9553 = n9549 & n9552;
  assign n9554 = n9553 ^ x73;
  assign n9555 = n9554 ^ x74;
  assign n9447 = n9379 & n9446;
  assign n9448 = n9447 ^ n9382;
  assign n9449 = ~x106 & ~n9448;
  assign n9450 = n9386 & n9446;
  assign n9451 = n9450 ^ n9392;
  assign n9452 = ~x107 & ~n9451;
  assign n9453 = ~n9449 & ~n9452;
  assign n9454 = n9325 & n9446;
  assign n9455 = n9454 ^ n9327;
  assign n9456 = n9455 ^ x97;
  assign n9457 = n9319 & n9446;
  assign n9458 = n9457 ^ n9321;
  assign n9459 = x96 & n9458;
  assign n9460 = n9459 ^ n9455;
  assign n9461 = n9460 ^ n9455;
  assign n9462 = ~x96 & ~n9458;
  assign n9463 = n9248 & n9446;
  assign n9464 = n9463 ^ n9254;
  assign n9465 = ~x84 & ~n9464;
  assign n9466 = n9258 & n9446;
  assign n9467 = n9466 ^ n9260;
  assign n9468 = ~x85 & n9467;
  assign n9469 = ~n9465 & ~n9468;
  assign n9556 = n9192 & n9446;
  assign n9557 = n9556 ^ n9194;
  assign n9558 = n9557 ^ n9554;
  assign n9559 = n9555 & n9558;
  assign n9560 = n9559 ^ x74;
  assign n9561 = n9560 ^ x75;
  assign n9562 = n9198 & n9446;
  assign n9563 = n9562 ^ n9200;
  assign n9564 = n9563 ^ n9560;
  assign n9565 = n9561 & ~n9564;
  assign n9566 = n9565 ^ x75;
  assign n9567 = n9566 ^ x76;
  assign n9568 = n9204 & n9446;
  assign n9569 = n9568 ^ n9206;
  assign n9570 = n9569 ^ n9566;
  assign n9571 = n9567 & n9570;
  assign n9572 = n9571 ^ x76;
  assign n9573 = n9572 ^ x77;
  assign n9574 = n9209 ^ x76;
  assign n9575 = n9446 & n9574;
  assign n9576 = n9575 ^ n9115;
  assign n9577 = n9576 ^ n9572;
  assign n9578 = n9573 & ~n9577;
  assign n9579 = n9578 ^ x77;
  assign n9580 = n9579 ^ x78;
  assign n9581 = n9209 ^ n9115;
  assign n9582 = n9574 & ~n9581;
  assign n9583 = n9582 ^ x76;
  assign n9584 = n9583 ^ x77;
  assign n9585 = n9446 & n9584;
  assign n9586 = n9585 ^ n9118;
  assign n9587 = n9586 ^ n9579;
  assign n9588 = n9580 & ~n9587;
  assign n9589 = n9588 ^ x78;
  assign n9590 = n9589 ^ x79;
  assign n9591 = ~n9217 & n9446;
  assign n9592 = n9591 ^ n9219;
  assign n9593 = n9592 ^ n9589;
  assign n9594 = n9590 & n9593;
  assign n9595 = n9594 ^ x79;
  assign n9596 = n9595 ^ x80;
  assign n9597 = n9223 & n9446;
  assign n9598 = n9597 ^ n9225;
  assign n9599 = n9598 ^ n9595;
  assign n9600 = n9596 & n9599;
  assign n9601 = n9600 ^ x80;
  assign n9602 = n9601 ^ x81;
  assign n9603 = n9229 & n9446;
  assign n9604 = n9603 ^ n9231;
  assign n9605 = n9604 ^ n9601;
  assign n9606 = n9602 & ~n9605;
  assign n9607 = n9606 ^ x81;
  assign n9608 = n9607 ^ x82;
  assign n9609 = n9235 & n9446;
  assign n9610 = n9609 ^ n9237;
  assign n9611 = n9610 ^ n9607;
  assign n9612 = n9608 & n9611;
  assign n9613 = n9612 ^ x82;
  assign n9614 = n9613 ^ x83;
  assign n9615 = n9241 & n9446;
  assign n9616 = n9615 ^ n9244;
  assign n9617 = n9616 ^ n9613;
  assign n9618 = n9614 & n9617;
  assign n9619 = n9618 ^ x83;
  assign n9620 = n9469 & n9619;
  assign n9621 = n9467 ^ x85;
  assign n9622 = x84 & n9464;
  assign n9623 = n9622 ^ n9467;
  assign n9624 = ~n9621 & n9623;
  assign n9625 = n9624 ^ x85;
  assign n9626 = ~n9620 & ~n9625;
  assign n9627 = n9626 ^ x86;
  assign n9628 = n9263 ^ x85;
  assign n9629 = n9446 & n9628;
  assign n9630 = n9629 ^ n9112;
  assign n9631 = n9630 ^ n9626;
  assign n9632 = ~n9627 & ~n9631;
  assign n9633 = n9632 ^ x86;
  assign n9634 = n9633 ^ x87;
  assign n9635 = ~n9264 & ~n9267;
  assign n9636 = n9635 ^ x86;
  assign n9637 = n9446 & n9636;
  assign n9638 = n9637 ^ n9109;
  assign n9639 = n9638 ^ n9633;
  assign n9640 = n9634 & n9639;
  assign n9641 = n9640 ^ x87;
  assign n9642 = n9641 ^ x88;
  assign n9643 = n9274 & n9446;
  assign n9644 = n9643 ^ n9276;
  assign n9645 = n9644 ^ n9641;
  assign n9646 = n9642 & ~n9645;
  assign n9647 = n9646 ^ x88;
  assign n9648 = n9647 ^ x89;
  assign n9649 = n9279 ^ x88;
  assign n9650 = n9446 & n9649;
  assign n9651 = n9650 ^ n9102;
  assign n9652 = n9651 ^ n9647;
  assign n9653 = n9648 & n9652;
  assign n9654 = n9653 ^ x89;
  assign n9655 = n9654 ^ x90;
  assign n9656 = n9279 ^ n9102;
  assign n9657 = n9649 & n9656;
  assign n9658 = n9657 ^ x88;
  assign n9659 = n9658 ^ x89;
  assign n9660 = n9446 & n9659;
  assign n9661 = n9660 ^ n9105;
  assign n9662 = n9661 ^ n9654;
  assign n9663 = n9655 & ~n9662;
  assign n9664 = n9663 ^ x90;
  assign n9665 = n9664 ^ x91;
  assign n9666 = n9286 ^ x90;
  assign n9667 = n9446 & ~n9666;
  assign n9668 = n9667 ^ n9288;
  assign n9669 = n9668 ^ n9664;
  assign n9670 = n9665 & ~n9669;
  assign n9671 = n9670 ^ x91;
  assign n9672 = n9671 ^ x92;
  assign n9673 = n9288 ^ n9286;
  assign n9674 = ~n9666 & n9673;
  assign n9675 = n9674 ^ x90;
  assign n9676 = n9675 ^ x91;
  assign n9677 = n9446 & n9676;
  assign n9678 = n9677 ^ n9291;
  assign n9679 = n9678 ^ n9671;
  assign n9680 = n9672 & ~n9679;
  assign n9681 = n9680 ^ x92;
  assign n9682 = n9681 ^ x93;
  assign n9683 = ~n9301 & n9446;
  assign n9684 = n9683 ^ n9303;
  assign n9685 = n9684 ^ n9681;
  assign n9686 = n9682 & ~n9685;
  assign n9687 = n9686 ^ x93;
  assign n9688 = n9687 ^ x94;
  assign n9689 = n9307 & n9446;
  assign n9690 = n9689 ^ n9309;
  assign n9691 = n9690 ^ n9687;
  assign n9692 = n9688 & ~n9691;
  assign n9693 = n9692 ^ x94;
  assign n9694 = n9693 ^ x95;
  assign n9695 = n9313 & n9446;
  assign n9696 = n9695 ^ n9315;
  assign n9697 = n9696 ^ n9693;
  assign n9698 = n9694 & ~n9697;
  assign n9699 = n9698 ^ x95;
  assign n9700 = ~n9462 & n9699;
  assign n9701 = n9700 ^ n9455;
  assign n9702 = n9701 ^ n9455;
  assign n9703 = ~n9461 & ~n9702;
  assign n9704 = n9703 ^ n9455;
  assign n9705 = n9456 & n9704;
  assign n9706 = n9705 ^ x97;
  assign n9707 = n9706 ^ x98;
  assign n9708 = n9331 & n9446;
  assign n9709 = n9708 ^ n9333;
  assign n9710 = n9709 ^ n9706;
  assign n9711 = n9707 & n9710;
  assign n9712 = n9711 ^ x98;
  assign n9713 = n9712 ^ x99;
  assign n9714 = n9337 & n9446;
  assign n9715 = n9714 ^ n9339;
  assign n9716 = n9715 ^ n9712;
  assign n9717 = n9713 & ~n9716;
  assign n9718 = n9717 ^ x99;
  assign n9719 = n9718 ^ x100;
  assign n9720 = n9343 & n9446;
  assign n9721 = n9720 ^ n9345;
  assign n9722 = n9721 ^ n9718;
  assign n9723 = n9719 & n9722;
  assign n9724 = n9723 ^ x100;
  assign n9725 = n9724 ^ x101;
  assign n9726 = n9349 & n9446;
  assign n9727 = n9726 ^ n9351;
  assign n9728 = n9727 ^ n9724;
  assign n9729 = n9725 & ~n9728;
  assign n9730 = n9729 ^ x101;
  assign n9731 = n9730 ^ x102;
  assign n9732 = n9355 & n9446;
  assign n9733 = n9732 ^ n9357;
  assign n9734 = n9733 ^ n9730;
  assign n9735 = n9731 & ~n9734;
  assign n9736 = n9735 ^ x102;
  assign n9737 = n9736 ^ x103;
  assign n9738 = n9361 & n9446;
  assign n9739 = n9738 ^ n9363;
  assign n9740 = n9739 ^ n9736;
  assign n9741 = n9737 & n9740;
  assign n9742 = n9741 ^ x103;
  assign n9743 = n9742 ^ x104;
  assign n9744 = n9367 & n9446;
  assign n9745 = n9744 ^ n9369;
  assign n9746 = n9745 ^ n9742;
  assign n9747 = n9743 & n9746;
  assign n9748 = n9747 ^ x104;
  assign n9749 = n9748 ^ x105;
  assign n9750 = n9373 & n9446;
  assign n9751 = n9750 ^ n9375;
  assign n9752 = n9751 ^ n9748;
  assign n9753 = n9749 & n9752;
  assign n9754 = n9753 ^ x105;
  assign n9755 = n9453 & n9754;
  assign n9756 = n9451 ^ x107;
  assign n9757 = x106 & n9448;
  assign n9758 = n9757 ^ n9451;
  assign n9759 = n9756 & ~n9758;
  assign n9760 = n9759 ^ x107;
  assign n9761 = ~n9755 & ~n9760;
  assign n9762 = n9761 ^ x108;
  assign n9763 = n9396 & n9446;
  assign n9764 = n9763 ^ n9398;
  assign n9765 = n9764 ^ n9761;
  assign n9766 = ~n9762 & n9765;
  assign n9767 = n9766 ^ x108;
  assign n9768 = n9767 ^ x109;
  assign n9769 = n9402 & n9446;
  assign n9770 = n9769 ^ n9404;
  assign n9771 = n9770 ^ n9767;
  assign n9772 = n9768 & ~n9771;
  assign n9773 = n9772 ^ x109;
  assign n9774 = n9773 ^ x110;
  assign n9775 = n9408 & n9446;
  assign n9776 = n9775 ^ n9410;
  assign n9777 = n9776 ^ n9773;
  assign n9778 = n9774 & ~n9777;
  assign n9779 = n9778 ^ x110;
  assign n9780 = n9779 ^ x111;
  assign n9781 = n9414 & n9446;
  assign n9782 = n9781 ^ n9417;
  assign n9783 = n9782 ^ n9779;
  assign n9784 = n9780 & n9783;
  assign n9785 = n9784 ^ x111;
  assign n9786 = n9785 ^ x112;
  assign n9787 = n9421 & n9446;
  assign n9788 = n9787 ^ n9425;
  assign n9789 = n9788 ^ n9785;
  assign n9790 = n9786 & ~n9789;
  assign n9791 = n9790 ^ x112;
  assign n9792 = n9791 ^ x113;
  assign n9793 = n9429 & n9446;
  assign n9794 = n9793 ^ n9432;
  assign n9795 = n9794 ^ n9791;
  assign n9796 = n9792 & n9795;
  assign n9797 = n9796 ^ x113;
  assign n9798 = n9797 ^ x114;
  assign n9437 = n9087 & n9436;
  assign n9438 = n9086 & ~n9437;
  assign n9805 = n9797 ^ n9438;
  assign n9806 = n9798 & n9805;
  assign n9807 = n9806 ^ x114;
  assign n9808 = n141 & ~n9807;
  assign n9821 = n9555 & n9808;
  assign n9822 = n9821 ^ n9557;
  assign n9823 = ~x75 & n9822;
  assign n9824 = n9561 & n9808;
  assign n9825 = n9824 ^ n9563;
  assign n9826 = ~x76 & ~n9825;
  assign n9827 = ~n9823 & ~n9826;
  assign n9828 = x65 & n141;
  assign n9829 = ~n9446 & n9828;
  assign n9830 = ~n9807 & n9829;
  assign n9831 = ~x65 & n9446;
  assign n9832 = x64 & n9831;
  assign n9833 = ~n9830 & ~n9832;
  assign n9834 = x13 & ~n9833;
  assign n9835 = ~n288 & ~n9446;
  assign n9836 = ~x13 & ~n9835;
  assign n9837 = ~n202 & ~n9836;
  assign n9838 = ~n9831 & ~n9837;
  assign n9839 = n9838 ^ n9470;
  assign n9840 = n9808 & n9839;
  assign n9841 = n9840 ^ n9470;
  assign n9842 = ~n9834 & ~n9841;
  assign n9843 = n9842 ^ x14;
  assign n9844 = n9843 ^ x66;
  assign n9845 = x64 & n9808;
  assign n9846 = x13 & ~x65;
  assign n9847 = x12 & n9846;
  assign n9848 = n9847 ^ x13;
  assign n9849 = n9845 & n9848;
  assign n9850 = ~x12 & n9477;
  assign n9851 = ~n9491 & ~n9850;
  assign n9852 = ~n9808 & ~n9851;
  assign n9853 = x13 ^ x12;
  assign n9854 = x64 ^ x13;
  assign n9855 = n9854 ^ x13;
  assign n9856 = n9853 & n9855;
  assign n9857 = n9856 ^ x13;
  assign n9858 = x65 & ~n9857;
  assign n9859 = ~n9852 & ~n9858;
  assign n9860 = ~n9849 & n9859;
  assign n9861 = n9860 ^ n9843;
  assign n9862 = n9844 & n9861;
  assign n9863 = n9862 ^ x66;
  assign n9864 = n9863 ^ x67;
  assign n9868 = n9478 & ~n9831;
  assign n9869 = n9483 ^ n9471;
  assign n9870 = n9470 & n9869;
  assign n9871 = n9870 ^ n9471;
  assign n9872 = ~n9868 & ~n9871;
  assign n9873 = n9872 ^ x66;
  assign n9874 = n9808 & ~n9873;
  assign n9865 = n9124 ^ x65;
  assign n9866 = n9446 & n9865;
  assign n9867 = n9866 ^ n9122;
  assign n9875 = n9874 ^ n9867;
  assign n9876 = n9875 ^ n9863;
  assign n9877 = n9864 & n9876;
  assign n9878 = n9877 ^ x67;
  assign n9879 = n9878 ^ x68;
  assign n9880 = n9513 & n9808;
  assign n9881 = n9880 ^ n9515;
  assign n9882 = n9881 ^ n9878;
  assign n9883 = n9879 & n9882;
  assign n9884 = n9883 ^ x68;
  assign n9885 = n9884 ^ x69;
  assign n9886 = n9519 & n9808;
  assign n9887 = n9886 ^ n9521;
  assign n9888 = n9887 ^ n9884;
  assign n9889 = n9885 & ~n9888;
  assign n9890 = n9889 ^ x69;
  assign n9891 = n9890 ^ x70;
  assign n9892 = n9525 & n9808;
  assign n9893 = n9892 ^ n9527;
  assign n9894 = n9893 ^ n9890;
  assign n9895 = n9891 & n9894;
  assign n9896 = n9895 ^ x70;
  assign n9897 = n9896 ^ x71;
  assign n9898 = n9531 & n9808;
  assign n9899 = n9898 ^ n9533;
  assign n9900 = n9899 ^ n9896;
  assign n9901 = n9897 & ~n9900;
  assign n9902 = n9901 ^ x71;
  assign n9903 = n9902 ^ x72;
  assign n9904 = n9537 & n9808;
  assign n9905 = n9904 ^ n9539;
  assign n9906 = n9905 ^ n9902;
  assign n9907 = n9903 & ~n9906;
  assign n9908 = n9907 ^ x72;
  assign n9909 = n9908 ^ x73;
  assign n9910 = n9543 & n9808;
  assign n9911 = n9910 ^ n9545;
  assign n9912 = n9911 ^ n9908;
  assign n9913 = n9909 & n9912;
  assign n9914 = n9913 ^ x73;
  assign n9915 = n9914 ^ x74;
  assign n9916 = n9549 & n9808;
  assign n9917 = n9916 ^ n9551;
  assign n9918 = n9917 ^ n9914;
  assign n9919 = n9915 & n9918;
  assign n9920 = n9919 ^ x74;
  assign n9921 = n9827 & n9920;
  assign n9922 = n9825 ^ x76;
  assign n9923 = x75 & ~n9822;
  assign n9924 = n9923 ^ n9825;
  assign n9925 = n9922 & ~n9924;
  assign n9926 = n9925 ^ x76;
  assign n9927 = ~n9921 & ~n9926;
  assign n9928 = n9927 ^ x77;
  assign n9929 = n9567 & n9808;
  assign n9930 = n9929 ^ n9569;
  assign n9931 = n9930 ^ n9927;
  assign n9932 = ~n9928 & ~n9931;
  assign n9933 = n9932 ^ x77;
  assign n9934 = n9933 ^ x78;
  assign n9935 = n9573 & n9808;
  assign n9936 = n9935 ^ n9576;
  assign n9937 = n9936 ^ n9933;
  assign n9938 = n9934 & ~n9937;
  assign n9939 = n9938 ^ x78;
  assign n9940 = n9939 ^ x79;
  assign n9941 = n9580 & n9808;
  assign n9942 = n9941 ^ n9586;
  assign n9943 = n9942 ^ n9939;
  assign n9944 = n9940 & ~n9943;
  assign n9945 = n9944 ^ x79;
  assign n9946 = n9945 ^ x80;
  assign n9947 = n9590 & n9808;
  assign n9948 = n9947 ^ n9592;
  assign n9949 = n9948 ^ n9945;
  assign n9950 = n9946 & n9949;
  assign n9951 = n9950 ^ x80;
  assign n9952 = n9951 ^ x81;
  assign n9953 = n9596 & n9808;
  assign n9954 = n9953 ^ n9598;
  assign n9955 = n9954 ^ n9951;
  assign n9956 = n9952 & n9955;
  assign n9957 = n9956 ^ x81;
  assign n9958 = n9957 ^ x82;
  assign n9959 = n9602 & n9808;
  assign n9960 = n9959 ^ n9604;
  assign n9961 = n9960 ^ n9957;
  assign n9962 = n9958 & ~n9961;
  assign n9963 = n9962 ^ x82;
  assign n9964 = n9963 ^ x83;
  assign n9965 = n9608 & n9808;
  assign n9966 = n9965 ^ n9610;
  assign n9967 = n9966 ^ n9963;
  assign n9968 = n9964 & n9967;
  assign n9969 = n9968 ^ x83;
  assign n9970 = n9969 ^ x84;
  assign n9971 = n9614 & n9808;
  assign n9972 = n9971 ^ n9616;
  assign n9973 = n9972 ^ n9969;
  assign n9974 = n9970 & n9973;
  assign n9975 = n9974 ^ x84;
  assign n9976 = n9975 ^ x85;
  assign n9977 = n9619 ^ x84;
  assign n9978 = n9808 & n9977;
  assign n9979 = n9978 ^ n9464;
  assign n9980 = n9979 ^ n9975;
  assign n9981 = n9976 & ~n9980;
  assign n9982 = n9981 ^ x85;
  assign n9983 = n9982 ^ x86;
  assign n9984 = n9619 ^ n9464;
  assign n9985 = n9977 & ~n9984;
  assign n9986 = n9985 ^ x84;
  assign n9987 = n9986 ^ x85;
  assign n9988 = n9808 & n9987;
  assign n9989 = n9988 ^ n9467;
  assign n9990 = n9989 ^ n9982;
  assign n9991 = n9983 & n9990;
  assign n9992 = n9991 ^ x86;
  assign n9993 = n9992 ^ x87;
  assign n9994 = ~n9627 & n9808;
  assign n9995 = n9994 ^ n9630;
  assign n9996 = n9995 ^ n9992;
  assign n9997 = n9993 & n9996;
  assign n9998 = n9997 ^ x87;
  assign n9999 = n9998 ^ x88;
  assign n10000 = n9634 & n9808;
  assign n10001 = n10000 ^ n9638;
  assign n10002 = n10001 ^ n9998;
  assign n10003 = n9999 & n10002;
  assign n10004 = n10003 ^ x88;
  assign n10005 = n10004 ^ x89;
  assign n10006 = n9642 & n9808;
  assign n10007 = n10006 ^ n9644;
  assign n10008 = n10007 ^ n10004;
  assign n10009 = n10005 & ~n10008;
  assign n10010 = n10009 ^ x89;
  assign n10011 = n10010 ^ x90;
  assign n10012 = n9648 & n9808;
  assign n10013 = n10012 ^ n9651;
  assign n10014 = n10013 ^ n10010;
  assign n10015 = n10011 & n10014;
  assign n10016 = n10015 ^ x90;
  assign n10017 = n10016 ^ x91;
  assign n10018 = n9655 & n9808;
  assign n10019 = n10018 ^ n9661;
  assign n10020 = n10019 ^ n10016;
  assign n10021 = n10017 & ~n10020;
  assign n10022 = n10021 ^ x91;
  assign n10023 = n10022 ^ x92;
  assign n10024 = n9665 & n9808;
  assign n10025 = n10024 ^ n9668;
  assign n10026 = n10025 ^ n10022;
  assign n10027 = n10023 & ~n10026;
  assign n10028 = n10027 ^ x92;
  assign n10029 = n10028 ^ x93;
  assign n10030 = n9672 & n9808;
  assign n10031 = n10030 ^ n9678;
  assign n10032 = n10031 ^ n10028;
  assign n10033 = n10029 & ~n10032;
  assign n10034 = n10033 ^ x93;
  assign n10035 = n10034 ^ x94;
  assign n10036 = n9682 & n9808;
  assign n10037 = n10036 ^ n9684;
  assign n10038 = n10037 ^ n10034;
  assign n10039 = n10035 & ~n10038;
  assign n10040 = n10039 ^ x94;
  assign n10041 = n10040 ^ x95;
  assign n10042 = n9688 & n9808;
  assign n10043 = n10042 ^ n9690;
  assign n10044 = n10043 ^ n10040;
  assign n10045 = n10041 & ~n10044;
  assign n10046 = n10045 ^ x95;
  assign n10047 = n10046 ^ x96;
  assign n10048 = n9694 & n9808;
  assign n10049 = n10048 ^ n9696;
  assign n10050 = n10049 ^ n10046;
  assign n10051 = n10047 & ~n10050;
  assign n10052 = n10051 ^ x96;
  assign n10053 = n10052 ^ x97;
  assign n10054 = n9699 ^ x96;
  assign n10055 = n9808 & n10054;
  assign n10056 = n10055 ^ n9458;
  assign n10057 = n10056 ^ n10052;
  assign n10058 = n10053 & ~n10057;
  assign n10059 = n10058 ^ x97;
  assign n10060 = n10059 ^ x98;
  assign n10061 = ~n9459 & ~n9700;
  assign n10062 = n10061 ^ x97;
  assign n10063 = n9808 & ~n10062;
  assign n10064 = n10063 ^ n9455;
  assign n10065 = n10064 ^ n10059;
  assign n10066 = n10060 & ~n10065;
  assign n10067 = n10066 ^ x98;
  assign n10068 = n10067 ^ x99;
  assign n9809 = n9792 & n9808;
  assign n9810 = n9809 ^ n9794;
  assign n9811 = ~x114 & n9810;
  assign n9799 = n141 & n9798;
  assign n9800 = n9438 & ~n9799;
  assign n9812 = ~x115 & n9800;
  assign n9813 = ~n9811 & ~n9812;
  assign n9814 = n9713 & n9808;
  assign n9815 = n9814 ^ n9715;
  assign n9816 = ~x100 & ~n9815;
  assign n9817 = n9719 & n9808;
  assign n9818 = n9817 ^ n9721;
  assign n9819 = ~x101 & n9818;
  assign n9820 = ~n9816 & ~n9819;
  assign n10069 = n9707 & n9808;
  assign n10070 = n10069 ^ n9709;
  assign n10071 = n10070 ^ n10067;
  assign n10072 = n10068 & n10071;
  assign n10073 = n10072 ^ x99;
  assign n10074 = n9820 & n10073;
  assign n10075 = n9818 ^ x101;
  assign n10076 = x100 & n9815;
  assign n10077 = n10076 ^ n9818;
  assign n10078 = ~n10075 & n10077;
  assign n10079 = n10078 ^ x101;
  assign n10080 = ~n10074 & ~n10079;
  assign n10081 = n10080 ^ x102;
  assign n10082 = n9725 & n9808;
  assign n10083 = n10082 ^ n9727;
  assign n10084 = n10083 ^ n10080;
  assign n10085 = ~n10081 & n10084;
  assign n10086 = n10085 ^ x102;
  assign n10087 = n10086 ^ x103;
  assign n10088 = n9731 & n9808;
  assign n10089 = n10088 ^ n9733;
  assign n10090 = n10089 ^ n10086;
  assign n10091 = n10087 & ~n10090;
  assign n10092 = n10091 ^ x103;
  assign n10093 = n10092 ^ x104;
  assign n10094 = n9737 & n9808;
  assign n10095 = n10094 ^ n9739;
  assign n10096 = n10095 ^ n10092;
  assign n10097 = n10093 & n10096;
  assign n10098 = n10097 ^ x104;
  assign n10099 = n10098 ^ x105;
  assign n10100 = n9743 & n9808;
  assign n10101 = n10100 ^ n9745;
  assign n10102 = n10101 ^ n10098;
  assign n10103 = n10099 & n10102;
  assign n10104 = n10103 ^ x105;
  assign n10105 = n10104 ^ x106;
  assign n10106 = n9749 & n9808;
  assign n10107 = n10106 ^ n9751;
  assign n10108 = n10107 ^ n10104;
  assign n10109 = n10105 & n10108;
  assign n10110 = n10109 ^ x106;
  assign n10111 = n10110 ^ x107;
  assign n10112 = n9754 ^ x106;
  assign n10113 = n9808 & n10112;
  assign n10114 = n10113 ^ n9448;
  assign n10115 = n10114 ^ n10110;
  assign n10116 = n10111 & ~n10115;
  assign n10117 = n10116 ^ x107;
  assign n10118 = n10117 ^ x108;
  assign n10119 = n9754 ^ n9448;
  assign n10120 = n10112 & ~n10119;
  assign n10121 = n10120 ^ x106;
  assign n10122 = n10121 ^ x107;
  assign n10123 = n9808 & n10122;
  assign n10124 = n10123 ^ n9451;
  assign n10125 = n10124 ^ n10117;
  assign n10126 = n10118 & ~n10125;
  assign n10127 = n10126 ^ x108;
  assign n10128 = n10127 ^ x109;
  assign n10129 = ~n9762 & n9808;
  assign n10130 = n10129 ^ n9764;
  assign n10131 = n10130 ^ n10127;
  assign n10132 = n10128 & ~n10131;
  assign n10133 = n10132 ^ x109;
  assign n10134 = n10133 ^ x110;
  assign n10135 = n9768 & n9808;
  assign n10136 = n10135 ^ n9770;
  assign n10137 = n10136 ^ n10133;
  assign n10138 = n10134 & ~n10137;
  assign n10139 = n10138 ^ x110;
  assign n10140 = n10139 ^ x111;
  assign n10141 = n9774 & n9808;
  assign n10142 = n10141 ^ n9776;
  assign n10143 = n10142 ^ n10139;
  assign n10144 = n10140 & ~n10143;
  assign n10145 = n10144 ^ x111;
  assign n10146 = n10145 ^ x112;
  assign n10147 = n9780 & n9808;
  assign n10148 = n10147 ^ n9782;
  assign n10149 = n10148 ^ n10145;
  assign n10150 = n10146 & n10149;
  assign n10151 = n10150 ^ x112;
  assign n10152 = n10151 ^ x113;
  assign n10153 = n9786 & n9808;
  assign n10154 = n10153 ^ n9788;
  assign n10155 = n10154 ^ n10151;
  assign n10156 = n10152 & ~n10155;
  assign n10157 = n10156 ^ x113;
  assign n10158 = n9813 & n10157;
  assign n10159 = n9800 ^ x115;
  assign n10160 = x114 & ~n9810;
  assign n10161 = n10160 ^ x115;
  assign n10162 = ~n10159 & n10161;
  assign n10163 = n10162 ^ x115;
  assign n10164 = n140 & ~n10163;
  assign n10165 = ~n10158 & n10164;
  assign n10170 = n10068 & n10165;
  assign n10171 = n10170 ^ n10070;
  assign n10172 = ~x100 & n10171;
  assign n10173 = n10073 ^ x100;
  assign n10174 = n10165 & n10173;
  assign n10175 = n10174 ^ n9815;
  assign n10176 = ~x101 & ~n10175;
  assign n10177 = ~n10172 & ~n10176;
  assign n10178 = n9920 ^ x75;
  assign n10179 = n10165 & n10178;
  assign n10180 = n10179 ^ n9822;
  assign n10181 = n9903 & n10165;
  assign n10182 = n10181 ^ n9905;
  assign n10183 = n10182 ^ x73;
  assign n10184 = n9897 & n10165;
  assign n10185 = n10184 ^ n9899;
  assign n10186 = x72 & n10185;
  assign n10187 = n10186 ^ n10182;
  assign n10188 = n10187 ^ n10182;
  assign n10189 = ~x72 & ~n10185;
  assign n10190 = x65 & n9808;
  assign n10191 = n10190 ^ x12;
  assign n10192 = n10191 ^ n10190;
  assign n10193 = n289 & ~n9808;
  assign n10194 = n10193 ^ x65;
  assign n10195 = n10194 ^ n10190;
  assign n10196 = ~n10192 & ~n10195;
  assign n10197 = n10196 ^ n10190;
  assign n10198 = ~n202 & n10197;
  assign n10199 = n10198 ^ n9845;
  assign n10200 = ~x12 & n10194;
  assign n10201 = ~x65 & ~n10200;
  assign n10202 = n10201 ^ n10198;
  assign n10203 = n10198 ^ n10165;
  assign n10204 = ~n10198 & ~n10203;
  assign n10205 = n10204 ^ n10198;
  assign n10206 = ~n10202 & ~n10205;
  assign n10207 = n10206 ^ n10204;
  assign n10208 = n10207 ^ n10198;
  assign n10209 = n10208 ^ n10165;
  assign n10210 = ~n10199 & ~n10209;
  assign n10211 = n10210 ^ n9845;
  assign n10212 = n10211 ^ x13;
  assign n10213 = n10212 ^ x66;
  assign n10214 = x12 & x64;
  assign n10215 = x11 & ~x65;
  assign n10216 = n10214 & ~n10215;
  assign n10217 = n10165 & n10216;
  assign n10219 = x65 ^ x12;
  assign n10226 = n10219 ^ x65;
  assign n10218 = x65 ^ x11;
  assign n10220 = n10219 ^ n10218;
  assign n10221 = n10220 ^ x65;
  assign n10222 = n10218 ^ x64;
  assign n10223 = n10222 ^ n10218;
  assign n10224 = n10223 ^ n10221;
  assign n10225 = ~n10221 & ~n10224;
  assign n10227 = n10226 ^ n10225;
  assign n10228 = n10227 ^ n10221;
  assign n10229 = n10165 ^ x65;
  assign n10230 = n10229 ^ x65;
  assign n10231 = n10225 ^ n10221;
  assign n10232 = ~n10230 & ~n10231;
  assign n10233 = n10232 ^ x65;
  assign n10234 = ~n10228 & n10233;
  assign n10235 = n10234 ^ x65;
  assign n10236 = n10235 ^ x65;
  assign n10237 = n10236 ^ x65;
  assign n10238 = ~n10217 & ~n10237;
  assign n10239 = n10238 ^ n10212;
  assign n10240 = ~n10213 & ~n10239;
  assign n10241 = n10240 ^ x66;
  assign n10242 = n10241 ^ x67;
  assign n10243 = n9860 ^ x66;
  assign n10244 = n10165 & ~n10243;
  assign n10245 = n10244 ^ n9843;
  assign n10246 = n10245 ^ n10241;
  assign n10247 = n10242 & ~n10246;
  assign n10248 = n10247 ^ x67;
  assign n10249 = n10248 ^ x68;
  assign n10250 = n9864 & n10165;
  assign n10251 = n10250 ^ n9875;
  assign n10252 = n10251 ^ n10248;
  assign n10253 = n10249 & n10252;
  assign n10254 = n10253 ^ x68;
  assign n10255 = n10254 ^ x69;
  assign n10256 = n9879 & n10165;
  assign n10257 = n10256 ^ n9881;
  assign n10258 = n10257 ^ n10254;
  assign n10259 = n10255 & n10258;
  assign n10260 = n10259 ^ x69;
  assign n10261 = n10260 ^ x70;
  assign n10262 = n9885 & n10165;
  assign n10263 = n10262 ^ n9887;
  assign n10264 = n10263 ^ n10260;
  assign n10265 = n10261 & ~n10264;
  assign n10266 = n10265 ^ x70;
  assign n10267 = n10266 ^ x71;
  assign n10268 = n9891 & n10165;
  assign n10269 = n10268 ^ n9893;
  assign n10270 = n10269 ^ n10266;
  assign n10271 = n10267 & n10270;
  assign n10272 = n10271 ^ x71;
  assign n10273 = ~n10189 & n10272;
  assign n10274 = n10273 ^ n10182;
  assign n10275 = n10274 ^ n10182;
  assign n10276 = ~n10188 & ~n10275;
  assign n10277 = n10276 ^ n10182;
  assign n10278 = n10183 & n10277;
  assign n10279 = n10278 ^ x73;
  assign n10280 = n10279 ^ x74;
  assign n10281 = n9909 & n10165;
  assign n10282 = n10281 ^ n9911;
  assign n10283 = n10282 ^ n10279;
  assign n10284 = n10280 & n10283;
  assign n10285 = n10284 ^ x74;
  assign n10286 = n10285 ^ x75;
  assign n10287 = n9915 & n10165;
  assign n10288 = n10287 ^ n9917;
  assign n10289 = n10288 ^ n10285;
  assign n10290 = n10286 & n10289;
  assign n10291 = n10290 ^ x75;
  assign n10292 = ~n10180 & n10291;
  assign n10293 = x76 & n10291;
  assign n10294 = ~n10292 & ~n10293;
  assign n10295 = n9920 ^ n9822;
  assign n10296 = n10178 & n10295;
  assign n10297 = n10296 ^ x75;
  assign n10298 = n10297 ^ x76;
  assign n10299 = n10165 & n10298;
  assign n10300 = n10299 ^ n9825;
  assign n10301 = x76 & x77;
  assign n10302 = ~n10300 & ~n10301;
  assign n10303 = ~n10294 & ~n10302;
  assign n10304 = x77 & n10292;
  assign n10305 = n10300 ^ x77;
  assign n10306 = n10300 ^ x76;
  assign n10307 = n10306 ^ n10300;
  assign n10308 = n10300 ^ n10180;
  assign n10309 = n10308 ^ n10300;
  assign n10310 = n10307 & ~n10309;
  assign n10311 = n10310 ^ n10300;
  assign n10312 = n10305 & ~n10311;
  assign n10313 = n10312 ^ x77;
  assign n10314 = ~n10304 & ~n10313;
  assign n10315 = ~n10303 & n10314;
  assign n10316 = ~n9928 & n10165;
  assign n10317 = n10316 ^ n9930;
  assign n10318 = ~x78 & n10317;
  assign n10319 = n9934 & n10165;
  assign n10320 = n10319 ^ n9936;
  assign n10321 = ~x79 & ~n10320;
  assign n10322 = ~n10318 & ~n10321;
  assign n10323 = ~n10315 & n10322;
  assign n10324 = n10320 ^ x79;
  assign n10325 = x78 & ~n10317;
  assign n10326 = n10325 ^ n10320;
  assign n10327 = n10324 & ~n10326;
  assign n10328 = n10327 ^ x79;
  assign n10329 = ~n10323 & ~n10328;
  assign n10330 = n10329 ^ x80;
  assign n10331 = n9940 & n10165;
  assign n10332 = n10331 ^ n9942;
  assign n10333 = n10332 ^ n10329;
  assign n10334 = ~n10330 & n10333;
  assign n10335 = n10334 ^ x80;
  assign n10336 = n10335 ^ x81;
  assign n10337 = n9946 & n10165;
  assign n10338 = n10337 ^ n9948;
  assign n10339 = n10338 ^ n10335;
  assign n10340 = n10336 & n10339;
  assign n10341 = n10340 ^ x81;
  assign n10342 = n10341 ^ x82;
  assign n10343 = n9952 & n10165;
  assign n10344 = n10343 ^ n9954;
  assign n10345 = n10344 ^ n10341;
  assign n10346 = n10342 & n10345;
  assign n10347 = n10346 ^ x82;
  assign n10348 = n10347 ^ x83;
  assign n10349 = n9958 & n10165;
  assign n10350 = n10349 ^ n9960;
  assign n10351 = n10350 ^ n10347;
  assign n10352 = n10348 & ~n10351;
  assign n10353 = n10352 ^ x83;
  assign n10354 = n10353 ^ x84;
  assign n10355 = n9964 & n10165;
  assign n10356 = n10355 ^ n9966;
  assign n10357 = n10356 ^ n10353;
  assign n10358 = n10354 & n10357;
  assign n10359 = n10358 ^ x84;
  assign n10360 = n10359 ^ x85;
  assign n10361 = n9970 & n10165;
  assign n10362 = n10361 ^ n9972;
  assign n10363 = n10362 ^ n10359;
  assign n10364 = n10360 & n10363;
  assign n10365 = n10364 ^ x85;
  assign n10366 = n10365 ^ x86;
  assign n10367 = n9976 & n10165;
  assign n10368 = n10367 ^ n9979;
  assign n10369 = n10368 ^ n10365;
  assign n10370 = n10366 & ~n10369;
  assign n10371 = n10370 ^ x86;
  assign n10372 = n10371 ^ x87;
  assign n10373 = n9983 & n10165;
  assign n10374 = n10373 ^ n9989;
  assign n10375 = n10374 ^ n10371;
  assign n10376 = n10372 & n10375;
  assign n10377 = n10376 ^ x87;
  assign n10378 = n10377 ^ x88;
  assign n10379 = n9993 & n10165;
  assign n10380 = n10379 ^ n9995;
  assign n10381 = n10380 ^ n10377;
  assign n10382 = n10378 & n10381;
  assign n10383 = n10382 ^ x88;
  assign n10384 = n10383 ^ x89;
  assign n10385 = n9999 & n10165;
  assign n10386 = n10385 ^ n10001;
  assign n10387 = n10386 ^ n10383;
  assign n10388 = n10384 & n10387;
  assign n10389 = n10388 ^ x89;
  assign n10390 = n10389 ^ x90;
  assign n10391 = n10005 & n10165;
  assign n10392 = n10391 ^ n10007;
  assign n10393 = n10392 ^ n10389;
  assign n10394 = n10390 & ~n10393;
  assign n10395 = n10394 ^ x90;
  assign n10396 = n10395 ^ x91;
  assign n10397 = n10011 & n10165;
  assign n10398 = n10397 ^ n10013;
  assign n10399 = n10398 ^ n10395;
  assign n10400 = n10396 & n10399;
  assign n10401 = n10400 ^ x91;
  assign n10402 = n10401 ^ x92;
  assign n10403 = n10017 & n10165;
  assign n10404 = n10403 ^ n10019;
  assign n10405 = n10404 ^ n10401;
  assign n10406 = n10402 & ~n10405;
  assign n10407 = n10406 ^ x92;
  assign n10408 = n10407 ^ x93;
  assign n10409 = n10023 & n10165;
  assign n10410 = n10409 ^ n10025;
  assign n10411 = n10410 ^ n10407;
  assign n10412 = n10408 & ~n10411;
  assign n10413 = n10412 ^ x93;
  assign n10414 = n10413 ^ x94;
  assign n10415 = n10029 & n10165;
  assign n10416 = n10415 ^ n10031;
  assign n10417 = n10416 ^ n10413;
  assign n10418 = n10414 & ~n10417;
  assign n10419 = n10418 ^ x94;
  assign n10420 = n10419 ^ x95;
  assign n10421 = n10035 & n10165;
  assign n10422 = n10421 ^ n10037;
  assign n10423 = n10422 ^ n10419;
  assign n10424 = n10420 & ~n10423;
  assign n10425 = n10424 ^ x95;
  assign n10426 = n10425 ^ x96;
  assign n10427 = n10041 & n10165;
  assign n10428 = n10427 ^ n10043;
  assign n10429 = n10428 ^ n10425;
  assign n10430 = n10426 & ~n10429;
  assign n10431 = n10430 ^ x96;
  assign n10432 = n10431 ^ x97;
  assign n10433 = n10047 & n10165;
  assign n10434 = n10433 ^ n10049;
  assign n10435 = n10434 ^ n10431;
  assign n10436 = n10432 & ~n10435;
  assign n10437 = n10436 ^ x97;
  assign n10438 = n10437 ^ x98;
  assign n10439 = n10053 & n10165;
  assign n10440 = n10439 ^ n10056;
  assign n10441 = n10440 ^ n10437;
  assign n10442 = n10438 & ~n10441;
  assign n10443 = n10442 ^ x98;
  assign n10444 = n10443 ^ x99;
  assign n10445 = n10060 & n10165;
  assign n10446 = n10445 ^ n10064;
  assign n10447 = n10446 ^ n10443;
  assign n10448 = n10444 & ~n10447;
  assign n10449 = n10448 ^ x99;
  assign n10450 = n10177 & n10449;
  assign n10451 = n10175 ^ x101;
  assign n10452 = x100 & ~n10171;
  assign n10453 = n10452 ^ n10175;
  assign n10454 = n10451 & ~n10453;
  assign n10455 = n10454 ^ x101;
  assign n10456 = ~n10450 & ~n10455;
  assign n10457 = n10456 ^ x102;
  assign n10458 = n10073 ^ n9815;
  assign n10459 = n10173 & ~n10458;
  assign n10460 = n10459 ^ x100;
  assign n10461 = n10460 ^ x101;
  assign n10462 = n10165 & n10461;
  assign n10463 = n10462 ^ n9818;
  assign n10464 = n10463 ^ n10456;
  assign n10465 = ~n10457 & ~n10464;
  assign n10466 = n10465 ^ x102;
  assign n10467 = n10466 ^ x103;
  assign n10468 = ~n10081 & n10165;
  assign n10469 = n10468 ^ n10083;
  assign n10470 = n10469 ^ n10466;
  assign n10471 = n10467 & ~n10470;
  assign n10472 = n10471 ^ x103;
  assign n10473 = n10472 ^ x104;
  assign n10474 = n10087 & n10165;
  assign n10475 = n10474 ^ n10089;
  assign n10476 = n10475 ^ n10472;
  assign n10477 = n10473 & ~n10476;
  assign n10478 = n10477 ^ x104;
  assign n10479 = n10478 ^ x105;
  assign n10480 = n10093 & n10165;
  assign n10481 = n10480 ^ n10095;
  assign n10482 = n10481 ^ n10478;
  assign n10483 = n10479 & n10482;
  assign n10484 = n10483 ^ x105;
  assign n10485 = n10484 ^ x106;
  assign n10486 = n10099 & n10165;
  assign n10487 = n10486 ^ n10101;
  assign n10488 = n10487 ^ n10484;
  assign n10489 = n10485 & n10488;
  assign n10490 = n10489 ^ x106;
  assign n10491 = n10490 ^ x107;
  assign n10492 = n10105 & n10165;
  assign n10493 = n10492 ^ n10107;
  assign n10494 = n10493 ^ n10490;
  assign n10495 = n10491 & n10494;
  assign n10496 = n10495 ^ x107;
  assign n10497 = n10496 ^ x108;
  assign n10498 = n10111 & n10165;
  assign n10499 = n10498 ^ n10114;
  assign n10500 = n10499 ^ n10496;
  assign n10501 = n10497 & ~n10500;
  assign n10502 = n10501 ^ x108;
  assign n10503 = n10502 ^ x109;
  assign n10504 = n10118 & n10165;
  assign n10505 = n10504 ^ n10124;
  assign n10506 = n10505 ^ n10502;
  assign n10507 = n10503 & ~n10506;
  assign n10508 = n10507 ^ x109;
  assign n10509 = n10508 ^ x110;
  assign n10510 = n10128 & n10165;
  assign n10511 = n10510 ^ n10130;
  assign n10512 = n10511 ^ n10508;
  assign n10513 = n10509 & ~n10512;
  assign n10514 = n10513 ^ x110;
  assign n10515 = n10514 ^ x111;
  assign n9804 = ~x117 & n9803;
  assign n10166 = n10157 ^ x114;
  assign n10167 = n10165 & n10166;
  assign n10168 = n10167 ^ n9810;
  assign n10169 = x115 & ~n10168;
  assign n10516 = n10134 & n10165;
  assign n10517 = n10516 ^ n10136;
  assign n10518 = n10517 ^ n10514;
  assign n10519 = n10515 & ~n10518;
  assign n10520 = n10519 ^ x111;
  assign n10521 = n10520 ^ x112;
  assign n10522 = n10140 & n10165;
  assign n10523 = n10522 ^ n10142;
  assign n10524 = n10523 ^ n10520;
  assign n10525 = n10521 & ~n10524;
  assign n10526 = n10525 ^ x112;
  assign n10527 = n10526 ^ x113;
  assign n10528 = n10146 & n10165;
  assign n10529 = n10528 ^ n10148;
  assign n10530 = n10529 ^ n10526;
  assign n10531 = n10527 & n10530;
  assign n10532 = n10531 ^ x113;
  assign n10533 = n10532 ^ x114;
  assign n10534 = n10152 & n10165;
  assign n10535 = n10534 ^ n10154;
  assign n10536 = n10535 ^ n10532;
  assign n10537 = n10533 & ~n10536;
  assign n10538 = n10537 ^ x114;
  assign n10539 = ~n10169 & ~n10538;
  assign n10540 = ~x115 & n10168;
  assign n10543 = n10157 ^ n9810;
  assign n10544 = n10166 & n10543;
  assign n10545 = n10544 ^ x114;
  assign n10546 = n10545 ^ x115;
  assign n10552 = n9800 & ~n10546;
  assign n10553 = ~n10540 & ~n10552;
  assign n10554 = ~n10539 & n10553;
  assign n10555 = ~x116 & ~n10554;
  assign n10541 = ~n10539 & ~n10540;
  assign n10556 = n9800 & ~n10541;
  assign n10557 = ~n10555 & ~n10556;
  assign n10558 = n9804 & ~n10557;
  assign n10559 = n10515 & n10558;
  assign n10560 = n10559 ^ n10517;
  assign n10561 = ~x112 & ~n10560;
  assign n10562 = n10521 & n10558;
  assign n10563 = n10562 ^ n10523;
  assign n10564 = ~x113 & ~n10563;
  assign n10565 = ~n10561 & ~n10564;
  assign n10566 = n10286 & n10558;
  assign n10567 = n10566 ^ n10288;
  assign n10568 = ~x76 & n10567;
  assign n10569 = n10291 ^ x76;
  assign n10570 = n10558 & n10569;
  assign n10571 = n10570 ^ n10180;
  assign n10572 = ~x77 & n10571;
  assign n10573 = ~n10568 & ~n10572;
  assign n10574 = n10255 & n10558;
  assign n10575 = n10574 ^ n10257;
  assign n10576 = n10575 ^ x70;
  assign n10577 = n10249 & n10558;
  assign n10578 = n10577 ^ n10251;
  assign n10579 = x69 & ~n10578;
  assign n10580 = n10579 ^ n10575;
  assign n10581 = n10580 ^ n10575;
  assign n10582 = ~x69 & n10578;
  assign n10583 = n10165 ^ x64;
  assign n10584 = n10583 ^ x64;
  assign n10585 = n10558 ^ x64;
  assign n10586 = ~n10584 & n10585;
  assign n10587 = n10586 ^ x64;
  assign n10588 = n10229 & n10587;
  assign n10589 = x11 & n10588;
  assign n10591 = ~x65 & n10165;
  assign n10592 = ~x11 & x64;
  assign n10593 = x65 & ~n10165;
  assign n10594 = n10592 & ~n10593;
  assign n10595 = ~n202 & ~n10594;
  assign n10596 = ~n10591 & ~n10595;
  assign n10590 = x64 & n10165;
  assign n10597 = n10596 ^ n10590;
  assign n10598 = ~n10558 & n10597;
  assign n10599 = n10598 ^ n10596;
  assign n10600 = ~n10589 & ~n10599;
  assign n10601 = n10600 ^ x12;
  assign n10602 = n10601 ^ x66;
  assign n10603 = x64 & n10558;
  assign n10604 = x11 & n10603;
  assign n10605 = x10 & ~x65;
  assign n10606 = n10604 & ~n10605;
  assign n10607 = ~x10 & x64;
  assign n10608 = ~x65 & ~n10607;
  assign n10609 = ~x11 & ~n10608;
  assign n10610 = ~n10558 & n10609;
  assign n10611 = ~x11 & n202;
  assign n10612 = ~x10 & x65;
  assign n10613 = x64 & n10612;
  assign n10614 = ~n10611 & ~n10613;
  assign n10615 = ~n10610 & n10614;
  assign n10616 = ~n10606 & n10615;
  assign n10617 = n10616 ^ n10601;
  assign n10618 = n10602 & n10617;
  assign n10619 = n10618 ^ x66;
  assign n10620 = n10619 ^ x67;
  assign n10621 = n10238 ^ x66;
  assign n10622 = n10558 & ~n10621;
  assign n10623 = n10622 ^ n10212;
  assign n10624 = n10623 ^ n10619;
  assign n10625 = n10620 & n10624;
  assign n10626 = n10625 ^ x67;
  assign n10627 = n10626 ^ x68;
  assign n10628 = n10242 & n10558;
  assign n10629 = n10628 ^ n10245;
  assign n10630 = n10629 ^ n10626;
  assign n10631 = n10627 & ~n10630;
  assign n10632 = n10631 ^ x68;
  assign n10633 = ~n10582 & n10632;
  assign n10634 = n10633 ^ n10575;
  assign n10635 = n10634 ^ n10575;
  assign n10636 = ~n10581 & ~n10635;
  assign n10637 = n10636 ^ n10575;
  assign n10638 = ~n10576 & ~n10637;
  assign n10639 = n10638 ^ x70;
  assign n10640 = n10639 ^ x71;
  assign n10641 = n10261 & n10558;
  assign n10642 = n10641 ^ n10263;
  assign n10643 = n10642 ^ n10639;
  assign n10644 = n10640 & ~n10643;
  assign n10645 = n10644 ^ x71;
  assign n10646 = n10645 ^ x72;
  assign n10647 = n10267 & n10558;
  assign n10648 = n10647 ^ n10269;
  assign n10649 = n10648 ^ n10645;
  assign n10650 = n10646 & n10649;
  assign n10651 = n10650 ^ x72;
  assign n10652 = n10651 ^ x73;
  assign n10653 = n10272 ^ x72;
  assign n10654 = n10558 & n10653;
  assign n10655 = n10654 ^ n10185;
  assign n10656 = n10655 ^ n10651;
  assign n10657 = n10652 & ~n10656;
  assign n10658 = n10657 ^ x73;
  assign n10659 = n10658 ^ x74;
  assign n10660 = ~n10186 & ~n10273;
  assign n10661 = n10660 ^ x73;
  assign n10662 = n10558 & ~n10661;
  assign n10663 = n10662 ^ n10182;
  assign n10664 = n10663 ^ n10658;
  assign n10665 = n10659 & ~n10664;
  assign n10666 = n10665 ^ x74;
  assign n10667 = n10666 ^ x75;
  assign n10668 = n10280 & n10558;
  assign n10669 = n10668 ^ n10282;
  assign n10670 = n10669 ^ n10666;
  assign n10671 = n10667 & n10670;
  assign n10672 = n10671 ^ x75;
  assign n10673 = n10573 & n10672;
  assign n10674 = n10571 ^ x77;
  assign n10675 = x76 & ~n10567;
  assign n10676 = n10675 ^ n10571;
  assign n10677 = ~n10674 & n10676;
  assign n10678 = n10677 ^ x77;
  assign n10679 = ~n10673 & ~n10678;
  assign n10680 = n10679 ^ x78;
  assign n10681 = n10291 ^ n10180;
  assign n10682 = n10569 & n10681;
  assign n10683 = n10682 ^ x76;
  assign n10684 = n10683 ^ x77;
  assign n10685 = n10558 & n10684;
  assign n10686 = n10685 ^ n10300;
  assign n10687 = n10686 ^ n10679;
  assign n10688 = ~n10680 & n10687;
  assign n10689 = n10688 ^ x78;
  assign n10690 = n10689 ^ x79;
  assign n10691 = n10315 ^ x78;
  assign n10692 = n10558 & ~n10691;
  assign n10693 = n10692 ^ n10317;
  assign n10694 = n10693 ^ n10689;
  assign n10695 = n10690 & n10694;
  assign n10696 = n10695 ^ x79;
  assign n10697 = n10696 ^ x80;
  assign n10698 = n10317 ^ n10315;
  assign n10699 = ~n10691 & ~n10698;
  assign n10700 = n10699 ^ x78;
  assign n10701 = n10700 ^ x79;
  assign n10702 = n10558 & n10701;
  assign n10703 = n10702 ^ n10320;
  assign n10704 = n10703 ^ n10696;
  assign n10705 = n10697 & ~n10704;
  assign n10706 = n10705 ^ x80;
  assign n10707 = n10706 ^ x81;
  assign n10708 = ~n10330 & n10558;
  assign n10709 = n10708 ^ n10332;
  assign n10710 = n10709 ^ n10706;
  assign n10711 = n10707 & ~n10710;
  assign n10712 = n10711 ^ x81;
  assign n10713 = n10712 ^ x82;
  assign n10714 = n10336 & n10558;
  assign n10715 = n10714 ^ n10338;
  assign n10716 = n10715 ^ n10712;
  assign n10717 = n10713 & n10716;
  assign n10718 = n10717 ^ x82;
  assign n10719 = n10718 ^ x83;
  assign n10720 = n10342 & n10558;
  assign n10721 = n10720 ^ n10344;
  assign n10722 = n10721 ^ n10718;
  assign n10723 = n10719 & n10722;
  assign n10724 = n10723 ^ x83;
  assign n10725 = n10724 ^ x84;
  assign n10726 = n10348 & n10558;
  assign n10727 = n10726 ^ n10350;
  assign n10728 = n10727 ^ n10724;
  assign n10729 = n10725 & ~n10728;
  assign n10730 = n10729 ^ x84;
  assign n10731 = n10730 ^ x85;
  assign n10732 = n10354 & n10558;
  assign n10733 = n10732 ^ n10356;
  assign n10734 = n10733 ^ n10730;
  assign n10735 = n10731 & n10734;
  assign n10736 = n10735 ^ x85;
  assign n10737 = n10736 ^ x86;
  assign n10738 = n10360 & n10558;
  assign n10739 = n10738 ^ n10362;
  assign n10740 = n10739 ^ n10736;
  assign n10741 = n10737 & n10740;
  assign n10742 = n10741 ^ x86;
  assign n10743 = n10742 ^ x87;
  assign n10744 = n10366 & n10558;
  assign n10745 = n10744 ^ n10368;
  assign n10746 = n10745 ^ n10742;
  assign n10747 = n10743 & ~n10746;
  assign n10748 = n10747 ^ x87;
  assign n10749 = n10748 ^ x88;
  assign n10750 = n10372 & n10558;
  assign n10751 = n10750 ^ n10374;
  assign n10752 = n10751 ^ n10748;
  assign n10753 = n10749 & n10752;
  assign n10754 = n10753 ^ x88;
  assign n10755 = n10754 ^ x89;
  assign n10756 = n10378 & n10558;
  assign n10757 = n10756 ^ n10380;
  assign n10758 = n10757 ^ n10754;
  assign n10759 = n10755 & n10758;
  assign n10760 = n10759 ^ x89;
  assign n10761 = n10760 ^ x90;
  assign n10762 = n10384 & n10558;
  assign n10763 = n10762 ^ n10386;
  assign n10764 = n10763 ^ n10760;
  assign n10765 = n10761 & n10764;
  assign n10766 = n10765 ^ x90;
  assign n10767 = n10766 ^ x91;
  assign n10768 = n10390 & n10558;
  assign n10769 = n10768 ^ n10392;
  assign n10770 = n10769 ^ n10766;
  assign n10771 = n10767 & ~n10770;
  assign n10772 = n10771 ^ x91;
  assign n10773 = n10772 ^ x92;
  assign n10774 = n10396 & n10558;
  assign n10775 = n10774 ^ n10398;
  assign n10776 = n10775 ^ n10772;
  assign n10777 = n10773 & n10776;
  assign n10778 = n10777 ^ x92;
  assign n10779 = n10778 ^ x93;
  assign n10780 = n10402 & n10558;
  assign n10781 = n10780 ^ n10404;
  assign n10782 = n10781 ^ n10778;
  assign n10783 = n10779 & ~n10782;
  assign n10784 = n10783 ^ x93;
  assign n10785 = n10784 ^ x94;
  assign n10786 = n10408 & n10558;
  assign n10787 = n10786 ^ n10410;
  assign n10788 = n10787 ^ n10784;
  assign n10789 = n10785 & ~n10788;
  assign n10790 = n10789 ^ x94;
  assign n10791 = n10790 ^ x95;
  assign n10792 = n10414 & n10558;
  assign n10793 = n10792 ^ n10416;
  assign n10794 = n10793 ^ n10790;
  assign n10795 = n10791 & ~n10794;
  assign n10796 = n10795 ^ x95;
  assign n10797 = n10796 ^ x96;
  assign n10798 = n10420 & n10558;
  assign n10799 = n10798 ^ n10422;
  assign n10800 = n10799 ^ n10796;
  assign n10801 = n10797 & ~n10800;
  assign n10802 = n10801 ^ x96;
  assign n10803 = n10802 ^ x97;
  assign n10804 = n10426 & n10558;
  assign n10805 = n10804 ^ n10428;
  assign n10806 = n10805 ^ n10802;
  assign n10807 = n10803 & ~n10806;
  assign n10808 = n10807 ^ x97;
  assign n10809 = n10808 ^ x98;
  assign n10810 = n10432 & n10558;
  assign n10811 = n10810 ^ n10434;
  assign n10812 = n10811 ^ n10808;
  assign n10813 = n10809 & ~n10812;
  assign n10814 = n10813 ^ x98;
  assign n10815 = n10814 ^ x99;
  assign n10816 = n10438 & n10558;
  assign n10817 = n10816 ^ n10440;
  assign n10818 = n10817 ^ n10814;
  assign n10819 = n10815 & ~n10818;
  assign n10820 = n10819 ^ x99;
  assign n10821 = n10820 ^ x100;
  assign n10822 = n10444 & n10558;
  assign n10823 = n10822 ^ n10446;
  assign n10824 = n10823 ^ n10820;
  assign n10825 = n10821 & ~n10824;
  assign n10826 = n10825 ^ x100;
  assign n10827 = n10826 ^ x101;
  assign n10828 = n10449 ^ x100;
  assign n10829 = n10558 & n10828;
  assign n10830 = n10829 ^ n10171;
  assign n10831 = n10830 ^ n10826;
  assign n10832 = n10827 & n10831;
  assign n10833 = n10832 ^ x101;
  assign n10834 = n10833 ^ x102;
  assign n10835 = n10449 ^ n10171;
  assign n10836 = n10828 & n10835;
  assign n10837 = n10836 ^ x100;
  assign n10838 = n10837 ^ x101;
  assign n10839 = n10558 & n10838;
  assign n10840 = n10839 ^ n10175;
  assign n10841 = n10840 ^ n10833;
  assign n10842 = n10834 & ~n10841;
  assign n10843 = n10842 ^ x102;
  assign n10844 = n10843 ^ x103;
  assign n10845 = ~n10457 & n10558;
  assign n10846 = n10845 ^ n10463;
  assign n10847 = n10846 ^ n10843;
  assign n10848 = n10844 & n10847;
  assign n10849 = n10848 ^ x103;
  assign n10850 = n10849 ^ x104;
  assign n10851 = n10467 & n10558;
  assign n10852 = n10851 ^ n10469;
  assign n10853 = n10852 ^ n10849;
  assign n10854 = n10850 & ~n10853;
  assign n10855 = n10854 ^ x104;
  assign n10856 = n10855 ^ x105;
  assign n10857 = n10473 & n10558;
  assign n10858 = n10857 ^ n10475;
  assign n10859 = n10858 ^ n10855;
  assign n10860 = n10856 & ~n10859;
  assign n10861 = n10860 ^ x105;
  assign n10862 = n10861 ^ x106;
  assign n10863 = n10479 & n10558;
  assign n10864 = n10863 ^ n10481;
  assign n10865 = n10864 ^ n10861;
  assign n10866 = n10862 & n10865;
  assign n10867 = n10866 ^ x106;
  assign n10868 = n10867 ^ x107;
  assign n10869 = n10485 & n10558;
  assign n10870 = n10869 ^ n10487;
  assign n10871 = n10870 ^ n10867;
  assign n10872 = n10868 & n10871;
  assign n10873 = n10872 ^ x107;
  assign n10874 = n10873 ^ x108;
  assign n10875 = n10491 & n10558;
  assign n10876 = n10875 ^ n10493;
  assign n10877 = n10876 ^ n10873;
  assign n10878 = n10874 & n10877;
  assign n10879 = n10878 ^ x108;
  assign n10880 = n10879 ^ x109;
  assign n10881 = n10497 & n10558;
  assign n10882 = n10881 ^ n10499;
  assign n10883 = n10882 ^ n10879;
  assign n10884 = n10880 & ~n10883;
  assign n10885 = n10884 ^ x109;
  assign n10886 = n10885 ^ x110;
  assign n10887 = n10503 & n10558;
  assign n10888 = n10887 ^ n10505;
  assign n10889 = n10888 ^ n10885;
  assign n10890 = n10886 & ~n10889;
  assign n10891 = n10890 ^ x110;
  assign n10892 = n10891 ^ x111;
  assign n10893 = n10509 & n10558;
  assign n10894 = n10893 ^ n10511;
  assign n10895 = n10894 ^ n10891;
  assign n10896 = n10892 & ~n10895;
  assign n10897 = n10896 ^ x111;
  assign n10898 = n10565 & n10897;
  assign n10899 = n10563 ^ x113;
  assign n10900 = x112 & n10560;
  assign n10901 = n10900 ^ n10563;
  assign n10902 = n10899 & ~n10901;
  assign n10903 = n10902 ^ x113;
  assign n10904 = ~n10898 & ~n10903;
  assign n10905 = n10904 ^ x114;
  assign n10906 = n10527 & n10558;
  assign n10907 = n10906 ^ n10529;
  assign n10908 = n10907 ^ n10904;
  assign n10909 = ~n10905 & ~n10908;
  assign n10910 = n10909 ^ x114;
  assign n10911 = n10910 ^ x115;
  assign n10912 = n10533 & n10558;
  assign n10913 = n10912 ^ n10535;
  assign n10914 = n10913 ^ n10910;
  assign n10915 = n10911 & ~n10914;
  assign n10916 = n10915 ^ x115;
  assign n10917 = n10916 ^ x116;
  assign n10918 = n10538 ^ x115;
  assign n10919 = n10558 & n10918;
  assign n10920 = n10919 ^ n10168;
  assign n10921 = n10920 ^ n10916;
  assign n10922 = n10917 & n10921;
  assign n10923 = n10922 ^ x116;
  assign n10924 = n10923 ^ x117;
  assign n10542 = n10541 ^ x116;
  assign n10547 = ~n10541 & n10546;
  assign n10548 = ~n10542 & n10547;
  assign n10549 = n10548 ^ n10542;
  assign n10550 = n9804 & n10549;
  assign n10551 = n9800 & ~n10550;
  assign n10925 = n10551 ^ x117;
  assign n10926 = n10924 & ~n10925;
  assign n10927 = n10926 ^ x117;
  assign n10928 = n9803 & ~n10927;
  assign n10950 = n10603 ^ x11;
  assign n10951 = ~n10928 & ~n10950;
  assign n10952 = ~x9 & ~n10605;
  assign n10953 = n10951 & n10952;
  assign n10954 = n10950 ^ x65;
  assign n10955 = x9 & n10605;
  assign n10956 = n10955 ^ x10;
  assign n10957 = ~n10954 & n10956;
  assign n10958 = n10928 & n10957;
  assign n10959 = ~x9 & n10612;
  assign n10960 = ~n10950 & n10959;
  assign n10961 = ~n10958 & ~n10960;
  assign n10962 = ~n10953 & n10961;
  assign n10963 = x64 & ~n10962;
  assign n10964 = x64 & n10928;
  assign n10965 = n10612 & ~n10964;
  assign n10966 = n10950 ^ n10928;
  assign n10967 = n10965 & ~n10966;
  assign n10968 = ~x66 & ~n10967;
  assign n10969 = ~n10963 & n10968;
  assign n10975 = ~x9 & x64;
  assign n10976 = ~n10605 & n10975;
  assign n10977 = ~n10612 & ~n10976;
  assign n10978 = n10950 & n10977;
  assign n10970 = ~x9 & x65;
  assign n10971 = n10607 & ~n10970;
  assign n10972 = ~n10954 & n10971;
  assign n10973 = x10 & n10611;
  assign n10974 = ~n10972 & ~n10973;
  assign n10979 = n10978 ^ n10974;
  assign n10980 = n10608 & ~n10975;
  assign n10981 = n10980 ^ n10974;
  assign n10982 = n10974 ^ n10928;
  assign n10983 = n10974 & n10982;
  assign n10984 = n10983 ^ n10974;
  assign n10985 = n10981 & n10984;
  assign n10986 = n10985 ^ n10983;
  assign n10987 = n10986 ^ n10974;
  assign n10988 = n10987 ^ n10928;
  assign n10989 = ~n10979 & n10988;
  assign n10990 = n10989 ^ n10978;
  assign n10991 = ~n10969 & ~n10990;
  assign n10992 = n10991 ^ x67;
  assign n10993 = n10616 ^ x66;
  assign n10994 = n10928 & ~n10993;
  assign n10995 = n10994 ^ n10601;
  assign n10996 = n10995 ^ n10991;
  assign n10997 = n10992 & ~n10996;
  assign n10998 = n10997 ^ x67;
  assign n10999 = n10998 ^ x68;
  assign n11000 = n10620 & n10928;
  assign n11001 = n11000 ^ n10623;
  assign n11002 = n11001 ^ n10998;
  assign n11003 = n10999 & n11002;
  assign n11004 = n11003 ^ x68;
  assign n11005 = n11004 ^ x69;
  assign n11006 = n10627 & n10928;
  assign n11007 = n11006 ^ n10629;
  assign n11008 = n11007 ^ n11004;
  assign n11009 = n11005 & ~n11008;
  assign n11010 = n11009 ^ x69;
  assign n11011 = ~x70 & ~n11010;
  assign n11012 = ~n10579 & ~n10633;
  assign n11013 = n11012 ^ x70;
  assign n11014 = n10928 & ~n11013;
  assign n11015 = n11014 ^ n10575;
  assign n11016 = n10632 ^ x69;
  assign n11017 = n10928 & n11016;
  assign n11018 = n11017 ^ n10578;
  assign n11019 = ~n11015 & ~n11018;
  assign n11020 = ~n11011 & n11019;
  assign n11021 = n11015 ^ x71;
  assign n11023 = n11015 ^ n11010;
  assign n11022 = n11015 ^ x70;
  assign n11024 = n11023 ^ n11022;
  assign n11025 = n11024 ^ n11021;
  assign n11026 = n11018 ^ n11015;
  assign n11027 = n11015 & n11026;
  assign n11028 = n11027 ^ n11022;
  assign n11029 = n11028 ^ n11015;
  assign n11030 = ~n11025 & n11029;
  assign n11031 = n11030 ^ n11027;
  assign n11032 = n11031 ^ n11015;
  assign n11033 = ~n11021 & n11032;
  assign n11034 = n11033 ^ x71;
  assign n11035 = ~n11020 & ~n11034;
  assign n11036 = n11035 ^ x72;
  assign n11037 = n10640 & n10928;
  assign n11038 = n11037 ^ n10642;
  assign n11039 = n11038 ^ n11035;
  assign n11040 = ~n11036 & n11039;
  assign n11041 = n11040 ^ x72;
  assign n11042 = n11041 ^ x73;
  assign n11043 = n10646 & n10928;
  assign n11044 = n11043 ^ n10648;
  assign n11045 = n11044 ^ n11041;
  assign n11046 = n11042 & n11045;
  assign n11047 = n11046 ^ x73;
  assign n11048 = n11047 ^ x74;
  assign n11049 = n10652 & n10928;
  assign n11050 = n11049 ^ n10655;
  assign n11051 = n11050 ^ n11047;
  assign n11052 = n11048 & ~n11051;
  assign n11053 = n11052 ^ x74;
  assign n11054 = n11053 ^ x75;
  assign n11055 = n10659 & n10928;
  assign n11056 = n11055 ^ n10663;
  assign n11057 = n11056 ^ n11053;
  assign n11058 = n11054 & ~n11057;
  assign n11059 = n11058 ^ x75;
  assign n11060 = n11059 ^ x76;
  assign n11061 = n10667 & n10928;
  assign n11062 = n11061 ^ n10669;
  assign n11063 = n11062 ^ n11059;
  assign n11064 = n11060 & n11063;
  assign n11065 = n11064 ^ x76;
  assign n11066 = n11065 ^ x77;
  assign n11067 = n10672 ^ x76;
  assign n11068 = n10928 & n11067;
  assign n11069 = n11068 ^ n10567;
  assign n11070 = n11069 ^ n11065;
  assign n11071 = n11066 & n11070;
  assign n11072 = n11071 ^ x77;
  assign n11073 = n11072 ^ x78;
  assign n11074 = n10672 ^ n10567;
  assign n11075 = n11067 & n11074;
  assign n11076 = n11075 ^ x76;
  assign n11077 = n11076 ^ x77;
  assign n11078 = n10928 & n11077;
  assign n11079 = n11078 ^ n10571;
  assign n11080 = n11079 ^ n11072;
  assign n11081 = n11073 & n11080;
  assign n11082 = n11081 ^ x78;
  assign n11083 = n11082 ^ x79;
  assign n11084 = ~n10680 & n10928;
  assign n11085 = n11084 ^ n10686;
  assign n11086 = n11085 ^ n11082;
  assign n11087 = n11083 & ~n11086;
  assign n11088 = n11087 ^ x79;
  assign n11089 = n11088 ^ x80;
  assign n11090 = n10690 & n10928;
  assign n11091 = n11090 ^ n10693;
  assign n11092 = n11091 ^ n11088;
  assign n11093 = n11089 & n11092;
  assign n11094 = n11093 ^ x80;
  assign n11095 = n11094 ^ x81;
  assign n11096 = n10697 & n10928;
  assign n11097 = n11096 ^ n10703;
  assign n11098 = n11097 ^ n11094;
  assign n11099 = n11095 & ~n11098;
  assign n11100 = n11099 ^ x81;
  assign n11101 = n11100 ^ x82;
  assign n11102 = n10707 & n10928;
  assign n11103 = n11102 ^ n10709;
  assign n11104 = n11103 ^ n11100;
  assign n11105 = n11101 & ~n11104;
  assign n11106 = n11105 ^ x82;
  assign n11107 = n11106 ^ x83;
  assign n11108 = n10713 & n10928;
  assign n11109 = n11108 ^ n10715;
  assign n11110 = n11109 ^ n11106;
  assign n11111 = n11107 & n11110;
  assign n11112 = n11111 ^ x83;
  assign n11113 = n11112 ^ x84;
  assign n11114 = n10719 & n10928;
  assign n11115 = n11114 ^ n10721;
  assign n11116 = n11115 ^ n11112;
  assign n11117 = n11113 & n11116;
  assign n11118 = n11117 ^ x84;
  assign n11119 = n11118 ^ x85;
  assign n11120 = n10725 & n10928;
  assign n11121 = n11120 ^ n10727;
  assign n11122 = n11121 ^ n11118;
  assign n11123 = n11119 & ~n11122;
  assign n11124 = n11123 ^ x85;
  assign n11125 = n11124 ^ x86;
  assign n11126 = n10731 & n10928;
  assign n11127 = n11126 ^ n10733;
  assign n11128 = n11127 ^ n11124;
  assign n11129 = n11125 & n11128;
  assign n11130 = n11129 ^ x86;
  assign n11131 = n11130 ^ x87;
  assign n11132 = n10737 & n10928;
  assign n11133 = n11132 ^ n10739;
  assign n11134 = n11133 ^ n11130;
  assign n11135 = n11131 & n11134;
  assign n11136 = n11135 ^ x87;
  assign n11137 = n11136 ^ x88;
  assign n11138 = n10743 & n10928;
  assign n11139 = n11138 ^ n10745;
  assign n11140 = n11139 ^ n11136;
  assign n11141 = n11137 & ~n11140;
  assign n11142 = n11141 ^ x88;
  assign n11143 = n11142 ^ x89;
  assign n11144 = n10749 & n10928;
  assign n11145 = n11144 ^ n10751;
  assign n11146 = n11145 ^ n11142;
  assign n11147 = n11143 & n11146;
  assign n11148 = n11147 ^ x89;
  assign n11149 = n11148 ^ x90;
  assign n11150 = n10755 & n10928;
  assign n11151 = n11150 ^ n10757;
  assign n11152 = n11151 ^ n11148;
  assign n11153 = n11149 & n11152;
  assign n11154 = n11153 ^ x90;
  assign n11155 = n11154 ^ x91;
  assign n11156 = n10761 & n10928;
  assign n11157 = n11156 ^ n10763;
  assign n11158 = n11157 ^ n11154;
  assign n11159 = n11155 & n11158;
  assign n11160 = n11159 ^ x91;
  assign n11161 = n11160 ^ x92;
  assign n11162 = n10767 & n10928;
  assign n11163 = n11162 ^ n10769;
  assign n11164 = n11163 ^ n11160;
  assign n11165 = n11161 & ~n11164;
  assign n11166 = n11165 ^ x92;
  assign n11167 = n11166 ^ x93;
  assign n10929 = n10924 & n10928;
  assign n10930 = n10551 & ~n10929;
  assign n10931 = n10897 ^ x112;
  assign n10932 = n10897 ^ n10560;
  assign n10933 = n10931 & ~n10932;
  assign n10934 = n10933 ^ x112;
  assign n10935 = n10934 ^ x113;
  assign n10936 = n10928 & n10935;
  assign n10937 = n10936 ^ n10563;
  assign n10938 = ~x114 & ~n10937;
  assign n10939 = n10928 & n10931;
  assign n10940 = n10939 ^ n10560;
  assign n10941 = ~x113 & ~n10940;
  assign n10942 = ~n10938 & ~n10941;
  assign n10943 = n10862 & n10928;
  assign n10944 = n10943 ^ n10864;
  assign n10945 = ~x107 & n10944;
  assign n10946 = n10868 & n10928;
  assign n10947 = n10946 ^ n10870;
  assign n10948 = ~x108 & n10947;
  assign n10949 = ~n10945 & ~n10948;
  assign n11168 = n10773 & n10928;
  assign n11169 = n11168 ^ n10775;
  assign n11170 = n11169 ^ n11166;
  assign n11171 = n11167 & n11170;
  assign n11172 = n11171 ^ x93;
  assign n11173 = n11172 ^ x94;
  assign n11174 = n10779 & n10928;
  assign n11175 = n11174 ^ n10781;
  assign n11176 = n11175 ^ n11172;
  assign n11177 = n11173 & ~n11176;
  assign n11178 = n11177 ^ x94;
  assign n11179 = n11178 ^ x95;
  assign n11180 = n10785 & n10928;
  assign n11181 = n11180 ^ n10787;
  assign n11182 = n11181 ^ n11178;
  assign n11183 = n11179 & ~n11182;
  assign n11184 = n11183 ^ x95;
  assign n11185 = n11184 ^ x96;
  assign n11186 = n10791 & n10928;
  assign n11187 = n11186 ^ n10793;
  assign n11188 = n11187 ^ n11184;
  assign n11189 = n11185 & ~n11188;
  assign n11190 = n11189 ^ x96;
  assign n11191 = n11190 ^ x97;
  assign n11192 = n10797 & n10928;
  assign n11193 = n11192 ^ n10799;
  assign n11194 = n11193 ^ n11190;
  assign n11195 = n11191 & ~n11194;
  assign n11196 = n11195 ^ x97;
  assign n11197 = n11196 ^ x98;
  assign n11198 = n10803 & n10928;
  assign n11199 = n11198 ^ n10805;
  assign n11200 = n11199 ^ n11196;
  assign n11201 = n11197 & ~n11200;
  assign n11202 = n11201 ^ x98;
  assign n11203 = n11202 ^ x99;
  assign n11204 = n10809 & n10928;
  assign n11205 = n11204 ^ n10811;
  assign n11206 = n11205 ^ n11202;
  assign n11207 = n11203 & ~n11206;
  assign n11208 = n11207 ^ x99;
  assign n11209 = n11208 ^ x100;
  assign n11210 = n10815 & n10928;
  assign n11211 = n11210 ^ n10817;
  assign n11212 = n11211 ^ n11208;
  assign n11213 = n11209 & ~n11212;
  assign n11214 = n11213 ^ x100;
  assign n11215 = n11214 ^ x101;
  assign n11216 = n10821 & n10928;
  assign n11217 = n11216 ^ n10823;
  assign n11218 = n11217 ^ n11214;
  assign n11219 = n11215 & ~n11218;
  assign n11220 = n11219 ^ x101;
  assign n11221 = n11220 ^ x102;
  assign n11222 = n10827 & n10928;
  assign n11223 = n11222 ^ n10830;
  assign n11224 = n11223 ^ n11220;
  assign n11225 = n11221 & n11224;
  assign n11226 = n11225 ^ x102;
  assign n11227 = n11226 ^ x103;
  assign n11228 = n10834 & n10928;
  assign n11229 = n11228 ^ n10840;
  assign n11230 = n11229 ^ n11226;
  assign n11231 = n11227 & ~n11230;
  assign n11232 = n11231 ^ x103;
  assign n11233 = n11232 ^ x104;
  assign n11234 = n10844 & n10928;
  assign n11235 = n11234 ^ n10846;
  assign n11236 = n11235 ^ n11232;
  assign n11237 = n11233 & n11236;
  assign n11238 = n11237 ^ x104;
  assign n11239 = n11238 ^ x105;
  assign n11240 = n10850 & n10928;
  assign n11241 = n11240 ^ n10852;
  assign n11242 = n11241 ^ n11238;
  assign n11243 = n11239 & ~n11242;
  assign n11244 = n11243 ^ x105;
  assign n11245 = n11244 ^ x106;
  assign n11246 = n10856 & n10928;
  assign n11247 = n11246 ^ n10858;
  assign n11248 = n11247 ^ n11244;
  assign n11249 = n11245 & ~n11248;
  assign n11250 = n11249 ^ x106;
  assign n11251 = n10949 & n11250;
  assign n11252 = n10947 ^ x108;
  assign n11253 = x107 & ~n10944;
  assign n11254 = n11253 ^ n10947;
  assign n11255 = ~n11252 & n11254;
  assign n11256 = n11255 ^ x108;
  assign n11257 = ~n11251 & ~n11256;
  assign n11258 = n11257 ^ x109;
  assign n11259 = n10874 & n10928;
  assign n11260 = n11259 ^ n10876;
  assign n11261 = n11260 ^ n11257;
  assign n11262 = ~n11258 & ~n11261;
  assign n11263 = n11262 ^ x109;
  assign n11264 = n11263 ^ x110;
  assign n11265 = n10880 & n10928;
  assign n11266 = n11265 ^ n10882;
  assign n11267 = n11266 ^ n11263;
  assign n11268 = n11264 & ~n11267;
  assign n11269 = n11268 ^ x110;
  assign n11270 = n11269 ^ x111;
  assign n11271 = n10886 & n10928;
  assign n11272 = n11271 ^ n10888;
  assign n11273 = n11272 ^ n11269;
  assign n11274 = n11270 & ~n11273;
  assign n11275 = n11274 ^ x111;
  assign n11276 = n11275 ^ x112;
  assign n11277 = n10892 & n10928;
  assign n11278 = n11277 ^ n10894;
  assign n11279 = n11278 ^ n11275;
  assign n11280 = n11276 & ~n11279;
  assign n11281 = n11280 ^ x112;
  assign n11282 = n10942 & n11281;
  assign n11283 = n10937 ^ x114;
  assign n11284 = x113 & n10940;
  assign n11285 = n11284 ^ n10937;
  assign n11286 = n11283 & ~n11285;
  assign n11287 = n11286 ^ x114;
  assign n11288 = ~n11282 & ~n11287;
  assign n11289 = ~n10905 & n10928;
  assign n11290 = n11289 ^ n10907;
  assign n11291 = ~x115 & n11290;
  assign n11292 = n10911 & n10928;
  assign n11293 = n11292 ^ n10913;
  assign n11294 = ~x116 & ~n11293;
  assign n11295 = ~n11291 & ~n11294;
  assign n11296 = ~n11288 & n11295;
  assign n11297 = n11293 ^ x116;
  assign n11298 = x115 & ~n11290;
  assign n11299 = n11298 ^ n11293;
  assign n11300 = n11297 & ~n11299;
  assign n11301 = n11300 ^ x116;
  assign n11302 = ~n11296 & ~n11301;
  assign n11312 = x117 & ~n11302;
  assign n11313 = ~n10930 & n11312;
  assign n11304 = n10917 & n10928;
  assign n11305 = n11304 ^ n10920;
  assign n11314 = ~x118 & n10930;
  assign n11315 = ~n11305 & ~n11314;
  assign n11316 = x117 & x118;
  assign n11317 = ~n11315 & ~n11316;
  assign n11318 = ~n11302 & ~n11317;
  assign n11319 = x117 & n11315;
  assign n11320 = x118 & ~n10930;
  assign n11321 = n9802 & ~n11320;
  assign n11322 = ~n11319 & n11321;
  assign n11323 = ~n11318 & n11322;
  assign n11324 = ~n11313 & n11323;
  assign n11337 = n11167 & n11324;
  assign n11338 = n11337 ^ n11169;
  assign n11339 = ~x94 & n11338;
  assign n11340 = n11161 & n11324;
  assign n11341 = n11340 ^ n11163;
  assign n11342 = ~x93 & ~n11341;
  assign n11343 = ~n11339 & ~n11342;
  assign n11344 = n10928 ^ x65;
  assign n11345 = n10975 & ~n11344;
  assign n11346 = ~n202 & ~n11345;
  assign n11347 = x65 & n10928;
  assign n11348 = x9 & ~n11347;
  assign n11349 = x65 & n11348;
  assign n11350 = n11346 & ~n11349;
  assign n11351 = n11350 ^ n10964;
  assign n11352 = n11350 ^ n11348;
  assign n11353 = n11350 ^ n11324;
  assign n11354 = n11350 & n11353;
  assign n11355 = n11354 ^ n11350;
  assign n11356 = n11352 & n11355;
  assign n11357 = n11356 ^ n11354;
  assign n11358 = n11357 ^ n11350;
  assign n11359 = n11358 ^ n11324;
  assign n11360 = ~n11351 & n11359;
  assign n11361 = n11360 ^ n10964;
  assign n11362 = n11361 ^ x10;
  assign n11363 = n11362 ^ x66;
  assign n11364 = x64 & n11324;
  assign n11365 = x9 & ~x65;
  assign n11366 = x8 & n11365;
  assign n11367 = n11366 ^ x9;
  assign n11368 = n11364 & n11367;
  assign n11369 = ~x8 & n10975;
  assign n11370 = ~n10970 & ~n11369;
  assign n11371 = ~n11324 & ~n11370;
  assign n11372 = x9 ^ x8;
  assign n11373 = x64 ^ x9;
  assign n11374 = n11373 ^ x9;
  assign n11375 = n11372 & n11374;
  assign n11376 = n11375 ^ x9;
  assign n11377 = x65 & ~n11376;
  assign n11378 = ~n11371 & ~n11377;
  assign n11379 = ~n11368 & n11378;
  assign n11380 = n11379 ^ n11362;
  assign n11381 = ~n11363 & ~n11380;
  assign n11382 = n11381 ^ x66;
  assign n11383 = n11382 ^ x67;
  assign n11387 = ~x65 & n10928;
  assign n11388 = n10976 & ~n11387;
  assign n11389 = n10964 ^ n10956;
  assign n11390 = n11389 ^ n10956;
  assign n11391 = n10956 ^ n10612;
  assign n11392 = ~n11390 & n11391;
  assign n11393 = n11392 ^ n10956;
  assign n11394 = ~n11388 & ~n11393;
  assign n11395 = n11394 ^ x66;
  assign n11396 = n11324 & ~n11395;
  assign n11384 = n10607 ^ x65;
  assign n11385 = n10928 & n11384;
  assign n11386 = n11385 ^ n10950;
  assign n11397 = n11396 ^ n11386;
  assign n11398 = n11397 ^ n11382;
  assign n11399 = n11383 & n11398;
  assign n11400 = n11399 ^ x67;
  assign n11401 = n11400 ^ x68;
  assign n11402 = n10992 & n11324;
  assign n11403 = n11402 ^ n10995;
  assign n11404 = n11403 ^ n11400;
  assign n11405 = n11401 & ~n11404;
  assign n11406 = n11405 ^ x68;
  assign n11407 = n11406 ^ x69;
  assign n11408 = n10999 & n11324;
  assign n11409 = n11408 ^ n11001;
  assign n11410 = n11409 ^ n11406;
  assign n11411 = n11407 & n11410;
  assign n11412 = n11411 ^ x69;
  assign n11413 = n11412 ^ x70;
  assign n11414 = n11005 & n11324;
  assign n11415 = n11414 ^ n11007;
  assign n11416 = n11415 ^ n11412;
  assign n11417 = n11413 & ~n11416;
  assign n11418 = n11417 ^ x70;
  assign n11419 = n11418 ^ x71;
  assign n11420 = n11010 ^ x70;
  assign n11421 = n11324 & n11420;
  assign n11422 = n11421 ^ n11018;
  assign n11423 = n11422 ^ n11418;
  assign n11424 = n11419 & n11423;
  assign n11425 = n11424 ^ x71;
  assign n11426 = n11425 ^ x72;
  assign n11427 = x70 & ~n11018;
  assign n11428 = ~x70 & n11018;
  assign n11429 = n11010 & ~n11428;
  assign n11430 = ~n11427 & ~n11429;
  assign n11431 = n11430 ^ x71;
  assign n11432 = n11324 & ~n11431;
  assign n11433 = n11432 ^ n11015;
  assign n11434 = n11433 ^ n11425;
  assign n11435 = n11426 & n11434;
  assign n11436 = n11435 ^ x72;
  assign n11437 = n11436 ^ x73;
  assign n11438 = ~n11036 & n11324;
  assign n11439 = n11438 ^ n11038;
  assign n11440 = n11439 ^ n11436;
  assign n11441 = n11437 & ~n11440;
  assign n11442 = n11441 ^ x73;
  assign n11443 = n11442 ^ x74;
  assign n11444 = n11042 & n11324;
  assign n11445 = n11444 ^ n11044;
  assign n11446 = n11445 ^ n11442;
  assign n11447 = n11443 & n11446;
  assign n11448 = n11447 ^ x74;
  assign n11449 = n11448 ^ x75;
  assign n11450 = n11048 & n11324;
  assign n11451 = n11450 ^ n11050;
  assign n11452 = n11451 ^ n11448;
  assign n11453 = n11449 & ~n11452;
  assign n11454 = n11453 ^ x75;
  assign n11455 = n11454 ^ x76;
  assign n11456 = n11054 & n11324;
  assign n11457 = n11456 ^ n11056;
  assign n11458 = n11457 ^ n11454;
  assign n11459 = n11455 & ~n11458;
  assign n11460 = n11459 ^ x76;
  assign n11461 = n11460 ^ x77;
  assign n11462 = n11060 & n11324;
  assign n11463 = n11462 ^ n11062;
  assign n11464 = n11463 ^ n11460;
  assign n11465 = n11461 & n11464;
  assign n11466 = n11465 ^ x77;
  assign n11467 = n11466 ^ x78;
  assign n11468 = n11066 & n11324;
  assign n11469 = n11468 ^ n11069;
  assign n11470 = n11469 ^ n11466;
  assign n11471 = n11467 & n11470;
  assign n11472 = n11471 ^ x78;
  assign n11473 = n11472 ^ x79;
  assign n11474 = n11073 & n11324;
  assign n11475 = n11474 ^ n11079;
  assign n11476 = n11475 ^ n11472;
  assign n11477 = n11473 & n11476;
  assign n11478 = n11477 ^ x79;
  assign n11479 = n11478 ^ x80;
  assign n11480 = n11083 & n11324;
  assign n11481 = n11480 ^ n11085;
  assign n11482 = n11481 ^ n11478;
  assign n11483 = n11479 & ~n11482;
  assign n11484 = n11483 ^ x80;
  assign n11485 = n11484 ^ x81;
  assign n11486 = n11089 & n11324;
  assign n11487 = n11486 ^ n11091;
  assign n11488 = n11487 ^ n11484;
  assign n11489 = n11485 & n11488;
  assign n11490 = n11489 ^ x81;
  assign n11491 = n11490 ^ x82;
  assign n11492 = n11095 & n11324;
  assign n11493 = n11492 ^ n11097;
  assign n11494 = n11493 ^ n11490;
  assign n11495 = n11491 & ~n11494;
  assign n11496 = n11495 ^ x82;
  assign n11497 = n11496 ^ x83;
  assign n11498 = n11101 & n11324;
  assign n11499 = n11498 ^ n11103;
  assign n11500 = n11499 ^ n11496;
  assign n11501 = n11497 & ~n11500;
  assign n11502 = n11501 ^ x83;
  assign n11503 = n11502 ^ x84;
  assign n11504 = n11107 & n11324;
  assign n11505 = n11504 ^ n11109;
  assign n11506 = n11505 ^ n11502;
  assign n11507 = n11503 & n11506;
  assign n11508 = n11507 ^ x84;
  assign n11509 = n11508 ^ x85;
  assign n11510 = n11113 & n11324;
  assign n11511 = n11510 ^ n11115;
  assign n11512 = n11511 ^ n11508;
  assign n11513 = n11509 & n11512;
  assign n11514 = n11513 ^ x85;
  assign n11515 = n11514 ^ x86;
  assign n11516 = n11119 & n11324;
  assign n11517 = n11516 ^ n11121;
  assign n11518 = n11517 ^ n11514;
  assign n11519 = n11515 & ~n11518;
  assign n11520 = n11519 ^ x86;
  assign n11521 = n11520 ^ x87;
  assign n11522 = n11125 & n11324;
  assign n11523 = n11522 ^ n11127;
  assign n11524 = n11523 ^ n11520;
  assign n11525 = n11521 & n11524;
  assign n11526 = n11525 ^ x87;
  assign n11527 = n11526 ^ x88;
  assign n11528 = n11131 & n11324;
  assign n11529 = n11528 ^ n11133;
  assign n11530 = n11529 ^ n11526;
  assign n11531 = n11527 & n11530;
  assign n11532 = n11531 ^ x88;
  assign n11533 = n11532 ^ x89;
  assign n11534 = n11137 & n11324;
  assign n11535 = n11534 ^ n11139;
  assign n11536 = n11535 ^ n11532;
  assign n11537 = n11533 & ~n11536;
  assign n11538 = n11537 ^ x89;
  assign n11539 = n11538 ^ x90;
  assign n11540 = n11143 & n11324;
  assign n11541 = n11540 ^ n11145;
  assign n11542 = n11541 ^ n11538;
  assign n11543 = n11539 & n11542;
  assign n11544 = n11543 ^ x90;
  assign n11545 = n11544 ^ x91;
  assign n11546 = n11149 & n11324;
  assign n11547 = n11546 ^ n11151;
  assign n11548 = n11547 ^ n11544;
  assign n11549 = n11545 & n11548;
  assign n11550 = n11549 ^ x91;
  assign n11551 = n11550 ^ x92;
  assign n11552 = n11155 & n11324;
  assign n11553 = n11552 ^ n11157;
  assign n11554 = n11553 ^ n11550;
  assign n11555 = n11551 & n11554;
  assign n11556 = n11555 ^ x92;
  assign n11557 = n11343 & n11556;
  assign n11558 = n11338 ^ x94;
  assign n11559 = x93 & n11341;
  assign n11560 = n11559 ^ n11338;
  assign n11561 = ~n11558 & n11560;
  assign n11562 = n11561 ^ x94;
  assign n11563 = ~n11557 & ~n11562;
  assign n11564 = n11563 ^ x95;
  assign n11565 = n11173 & n11324;
  assign n11566 = n11565 ^ n11175;
  assign n11567 = n11566 ^ n11563;
  assign n11568 = ~n11564 & n11567;
  assign n11569 = n11568 ^ x95;
  assign n11570 = n11569 ^ x96;
  assign n11571 = n11179 & n11324;
  assign n11572 = n11571 ^ n11181;
  assign n11573 = n11572 ^ n11569;
  assign n11574 = n11570 & ~n11573;
  assign n11575 = n11574 ^ x96;
  assign n11576 = n11575 ^ x97;
  assign n11577 = n11185 & n11324;
  assign n11578 = n11577 ^ n11187;
  assign n11579 = n11578 ^ n11575;
  assign n11580 = n11576 & ~n11579;
  assign n11581 = n11580 ^ x97;
  assign n11582 = n11581 ^ x98;
  assign n11583 = n11191 & n11324;
  assign n11584 = n11583 ^ n11193;
  assign n11585 = n11584 ^ n11581;
  assign n11586 = n11582 & ~n11585;
  assign n11587 = n11586 ^ x98;
  assign n11588 = n11587 ^ x99;
  assign n11589 = n11197 & n11324;
  assign n11590 = n11589 ^ n11199;
  assign n11591 = n11590 ^ n11587;
  assign n11592 = n11588 & ~n11591;
  assign n11593 = n11592 ^ x99;
  assign n11594 = n11593 ^ x100;
  assign n11595 = n11203 & n11324;
  assign n11596 = n11595 ^ n11205;
  assign n11597 = n11596 ^ n11593;
  assign n11598 = n11594 & ~n11597;
  assign n11599 = n11598 ^ x100;
  assign n11600 = n11599 ^ x101;
  assign n11601 = n11209 & n11324;
  assign n11602 = n11601 ^ n11211;
  assign n11603 = n11602 ^ n11599;
  assign n11604 = n11600 & ~n11603;
  assign n11605 = n11604 ^ x101;
  assign n11606 = n11605 ^ x102;
  assign n11607 = n11215 & n11324;
  assign n11608 = n11607 ^ n11217;
  assign n11609 = n11608 ^ n11605;
  assign n11610 = n11606 & ~n11609;
  assign n11611 = n11610 ^ x102;
  assign n11612 = n11611 ^ x103;
  assign n11613 = n11221 & n11324;
  assign n11614 = n11613 ^ n11223;
  assign n11615 = n11614 ^ n11611;
  assign n11616 = n11612 & n11615;
  assign n11617 = n11616 ^ x103;
  assign n11618 = n11617 ^ x104;
  assign n11619 = n11227 & n11324;
  assign n11620 = n11619 ^ n11229;
  assign n11621 = n11620 ^ n11617;
  assign n11622 = n11618 & ~n11621;
  assign n11623 = n11622 ^ x104;
  assign n11624 = n11623 ^ x105;
  assign n11625 = n11233 & n11324;
  assign n11626 = n11625 ^ n11235;
  assign n11627 = n11626 ^ n11623;
  assign n11628 = n11624 & n11627;
  assign n11629 = n11628 ^ x105;
  assign n11630 = n11629 ^ x106;
  assign n11631 = n11239 & n11324;
  assign n11632 = n11631 ^ n11241;
  assign n11633 = n11632 ^ n11629;
  assign n11634 = n11630 & ~n11633;
  assign n11635 = n11634 ^ x106;
  assign n11636 = n11635 ^ x107;
  assign n11325 = n11288 ^ x115;
  assign n11326 = n11290 ^ n11288;
  assign n11327 = ~n11325 & ~n11326;
  assign n11328 = n11327 ^ x115;
  assign n11329 = n11328 ^ x116;
  assign n11330 = n11324 & n11329;
  assign n11331 = n11330 ^ n11293;
  assign n11332 = ~x117 & ~n11331;
  assign n11303 = n11302 ^ x117;
  assign n11333 = ~n11303 & n11323;
  assign n11334 = n11333 ^ n11305;
  assign n11335 = ~x118 & n11334;
  assign n11336 = ~n11332 & ~n11335;
  assign n11637 = n11245 & n11324;
  assign n11638 = n11637 ^ n11247;
  assign n11639 = n11638 ^ n11635;
  assign n11640 = n11636 & ~n11639;
  assign n11641 = n11640 ^ x107;
  assign n11642 = n11641 ^ x108;
  assign n11643 = n11250 ^ x107;
  assign n11644 = n11324 & n11643;
  assign n11645 = n11644 ^ n10944;
  assign n11646 = n11645 ^ n11641;
  assign n11647 = n11642 & n11646;
  assign n11648 = n11647 ^ x108;
  assign n11649 = n11648 ^ x109;
  assign n11650 = n11250 ^ n10944;
  assign n11651 = n11643 & n11650;
  assign n11652 = n11651 ^ x107;
  assign n11653 = n11652 ^ x108;
  assign n11654 = n11324 & n11653;
  assign n11655 = n11654 ^ n10947;
  assign n11656 = n11655 ^ n11648;
  assign n11657 = n11649 & n11656;
  assign n11658 = n11657 ^ x109;
  assign n11659 = n11658 ^ x110;
  assign n11660 = ~n11258 & n11324;
  assign n11661 = n11660 ^ n11260;
  assign n11662 = n11661 ^ n11658;
  assign n11663 = n11659 & n11662;
  assign n11664 = n11663 ^ x110;
  assign n11665 = n11664 ^ x111;
  assign n11666 = n11264 & n11324;
  assign n11667 = n11666 ^ n11266;
  assign n11668 = n11667 ^ n11664;
  assign n11669 = n11665 & ~n11668;
  assign n11670 = n11669 ^ x111;
  assign n11671 = n11670 ^ x112;
  assign n11672 = n11270 & n11324;
  assign n11673 = n11672 ^ n11272;
  assign n11674 = n11673 ^ n11670;
  assign n11675 = n11671 & ~n11674;
  assign n11676 = n11675 ^ x112;
  assign n11677 = n11676 ^ x113;
  assign n11678 = n11276 & n11324;
  assign n11679 = n11678 ^ n11278;
  assign n11680 = n11679 ^ n11676;
  assign n11681 = n11677 & ~n11680;
  assign n11682 = n11681 ^ x113;
  assign n11683 = n11682 ^ x114;
  assign n11684 = n11281 ^ x113;
  assign n11685 = n11324 & n11684;
  assign n11686 = n11685 ^ n10940;
  assign n11687 = n11686 ^ n11682;
  assign n11688 = n11683 & ~n11687;
  assign n11689 = n11688 ^ x114;
  assign n11690 = n11689 ^ x115;
  assign n11691 = n11281 ^ n10940;
  assign n11692 = n11684 & ~n11691;
  assign n11693 = n11692 ^ x113;
  assign n11694 = n11693 ^ x114;
  assign n11695 = n11324 & n11694;
  assign n11696 = n11695 ^ n10937;
  assign n11697 = n11696 ^ n11689;
  assign n11698 = n11690 & ~n11697;
  assign n11699 = n11698 ^ x115;
  assign n11700 = n11699 ^ x116;
  assign n11701 = n11324 & ~n11325;
  assign n11702 = n11701 ^ n11290;
  assign n11703 = n11702 ^ n11699;
  assign n11704 = n11700 & n11703;
  assign n11705 = n11704 ^ x116;
  assign n11706 = n11336 & n11705;
  assign n11707 = n11334 ^ x118;
  assign n11708 = x117 & n11331;
  assign n11709 = n11708 ^ n11334;
  assign n11710 = ~n11707 & n11709;
  assign n11711 = n11710 ^ x118;
  assign n11712 = ~n11706 & ~n11711;
  assign n11716 = x119 & ~n10551;
  assign n11717 = n9801 & ~n11716;
  assign n11718 = n11712 & n11717;
  assign n11306 = n11305 ^ n11302;
  assign n11307 = ~n11303 & ~n11306;
  assign n11308 = n11307 ^ x117;
  assign n11309 = n11308 ^ x118;
  assign n11310 = n9802 & n11309;
  assign n11311 = n10930 & ~n11310;
  assign n11719 = n9802 & n11311;
  assign n11720 = ~n11718 & ~n11719;
  assign n11733 = n11636 & ~n11720;
  assign n11734 = n11733 ^ n11638;
  assign n11735 = ~x108 & ~n11734;
  assign n11736 = n11630 & ~n11720;
  assign n11737 = n11736 ^ n11632;
  assign n11738 = ~x107 & ~n11737;
  assign n11739 = ~n11735 & ~n11738;
  assign n11740 = n11576 & ~n11720;
  assign n11741 = n11740 ^ n11578;
  assign n11742 = n11741 ^ x98;
  assign n11743 = n11570 & ~n11720;
  assign n11744 = n11743 ^ n11572;
  assign n11745 = x97 & n11744;
  assign n11746 = n11745 ^ n11741;
  assign n11747 = n11746 ^ n11741;
  assign n11748 = ~x97 & ~n11744;
  assign n11749 = n11467 & ~n11720;
  assign n11750 = n11749 ^ n11469;
  assign n11751 = ~x79 & n11750;
  assign n11752 = n11473 & ~n11720;
  assign n11753 = n11752 ^ n11475;
  assign n11754 = ~x80 & n11753;
  assign n11755 = ~n11751 & ~n11754;
  assign n11756 = n11426 & ~n11720;
  assign n11757 = n11756 ^ n11433;
  assign n11758 = n11757 ^ x73;
  assign n11759 = n11419 & ~n11720;
  assign n11760 = n11759 ^ n11422;
  assign n11761 = x72 & ~n11760;
  assign n11762 = n11761 ^ n11757;
  assign n11763 = n11762 ^ n11757;
  assign n11764 = ~x72 & n11760;
  assign n11765 = ~x65 & n11720;
  assign n11766 = ~x7 & x64;
  assign n11767 = n11765 & ~n11766;
  assign n11768 = x8 & x64;
  assign n11769 = x7 & ~x65;
  assign n11770 = n11768 & ~n11769;
  assign n11771 = n11770 ^ x8;
  assign n11772 = ~n11720 & ~n11771;
  assign n11773 = n11772 ^ x8;
  assign n11774 = ~n11767 & ~n11773;
  assign n11775 = x8 ^ x7;
  assign n11776 = ~x64 & n11775;
  assign n11777 = n11776 ^ x7;
  assign n11778 = x65 & ~n11777;
  assign n11779 = ~n11774 & ~n11778;
  assign n11780 = n11779 ^ x66;
  assign n11781 = n289 & ~n11324;
  assign n11782 = n11781 ^ x65;
  assign n11783 = ~x8 & n11782;
  assign n11784 = ~n202 & ~n11783;
  assign n11785 = x65 & n11324;
  assign n11786 = x8 & ~n11785;
  assign n11787 = x65 & n11786;
  assign n11788 = n11784 & ~n11787;
  assign n11789 = n11788 ^ n11364;
  assign n11790 = n11788 ^ n11786;
  assign n11791 = n11788 ^ n11720;
  assign n11792 = n11788 & ~n11791;
  assign n11793 = n11792 ^ n11788;
  assign n11794 = n11790 & n11793;
  assign n11795 = n11794 ^ n11792;
  assign n11796 = n11795 ^ n11788;
  assign n11797 = n11796 ^ n11720;
  assign n11798 = ~n11789 & ~n11797;
  assign n11799 = n11798 ^ n11364;
  assign n11800 = n11799 ^ x9;
  assign n11801 = n11800 ^ n11779;
  assign n11802 = ~n11780 & ~n11801;
  assign n11803 = n11802 ^ x66;
  assign n11804 = n11803 ^ x67;
  assign n11805 = n11379 ^ x66;
  assign n11806 = ~n11720 & ~n11805;
  assign n11807 = n11806 ^ n11362;
  assign n11808 = n11807 ^ n11803;
  assign n11809 = n11804 & n11808;
  assign n11810 = n11809 ^ x67;
  assign n11811 = n11810 ^ x68;
  assign n11812 = n11383 & ~n11720;
  assign n11813 = n11812 ^ n11397;
  assign n11814 = n11813 ^ n11810;
  assign n11815 = n11811 & n11814;
  assign n11816 = n11815 ^ x68;
  assign n11817 = n11816 ^ x69;
  assign n11818 = n11401 & ~n11720;
  assign n11819 = n11818 ^ n11403;
  assign n11820 = n11819 ^ n11816;
  assign n11821 = n11817 & ~n11820;
  assign n11822 = n11821 ^ x69;
  assign n11823 = n11822 ^ x70;
  assign n11824 = n11407 & ~n11720;
  assign n11825 = n11824 ^ n11409;
  assign n11826 = n11825 ^ n11822;
  assign n11827 = n11823 & n11826;
  assign n11828 = n11827 ^ x70;
  assign n11829 = n11828 ^ x71;
  assign n11830 = n11413 & ~n11720;
  assign n11831 = n11830 ^ n11415;
  assign n11832 = n11831 ^ n11828;
  assign n11833 = n11829 & ~n11832;
  assign n11834 = n11833 ^ x71;
  assign n11835 = ~n11764 & n11834;
  assign n11836 = n11835 ^ n11757;
  assign n11837 = n11836 ^ n11757;
  assign n11838 = ~n11763 & ~n11837;
  assign n11839 = n11838 ^ n11757;
  assign n11840 = ~n11758 & ~n11839;
  assign n11841 = n11840 ^ x73;
  assign n11842 = n11841 ^ x74;
  assign n11843 = n11437 & ~n11720;
  assign n11844 = n11843 ^ n11439;
  assign n11845 = n11844 ^ n11841;
  assign n11846 = n11842 & ~n11845;
  assign n11847 = n11846 ^ x74;
  assign n11848 = n11847 ^ x75;
  assign n11849 = n11443 & ~n11720;
  assign n11850 = n11849 ^ n11445;
  assign n11851 = n11850 ^ n11847;
  assign n11852 = n11848 & n11851;
  assign n11853 = n11852 ^ x75;
  assign n11854 = n11853 ^ x76;
  assign n11855 = n11449 & ~n11720;
  assign n11856 = n11855 ^ n11451;
  assign n11857 = n11856 ^ n11853;
  assign n11858 = n11854 & ~n11857;
  assign n11859 = n11858 ^ x76;
  assign n11860 = n11859 ^ x77;
  assign n11861 = n11455 & ~n11720;
  assign n11862 = n11861 ^ n11457;
  assign n11863 = n11862 ^ n11859;
  assign n11864 = n11860 & ~n11863;
  assign n11865 = n11864 ^ x77;
  assign n11866 = n11865 ^ x78;
  assign n11867 = n11461 & ~n11720;
  assign n11868 = n11867 ^ n11463;
  assign n11869 = n11868 ^ n11865;
  assign n11870 = n11866 & n11869;
  assign n11871 = n11870 ^ x78;
  assign n11872 = n11755 & n11871;
  assign n11873 = n11753 ^ x80;
  assign n11874 = x79 & ~n11750;
  assign n11875 = n11874 ^ n11753;
  assign n11876 = ~n11873 & n11875;
  assign n11877 = n11876 ^ x80;
  assign n11878 = ~n11872 & ~n11877;
  assign n11879 = n11878 ^ x81;
  assign n11880 = n11479 & ~n11720;
  assign n11881 = n11880 ^ n11481;
  assign n11882 = n11881 ^ n11878;
  assign n11883 = ~n11879 & n11882;
  assign n11884 = n11883 ^ x81;
  assign n11885 = n11884 ^ x82;
  assign n11886 = n11485 & ~n11720;
  assign n11887 = n11886 ^ n11487;
  assign n11888 = n11887 ^ n11884;
  assign n11889 = n11885 & n11888;
  assign n11890 = n11889 ^ x82;
  assign n11891 = n11890 ^ x83;
  assign n11892 = n11491 & ~n11720;
  assign n11893 = n11892 ^ n11493;
  assign n11894 = n11893 ^ n11890;
  assign n11895 = n11891 & ~n11894;
  assign n11896 = n11895 ^ x83;
  assign n11897 = n11896 ^ x84;
  assign n11898 = n11497 & ~n11720;
  assign n11899 = n11898 ^ n11499;
  assign n11900 = n11899 ^ n11896;
  assign n11901 = n11897 & ~n11900;
  assign n11902 = n11901 ^ x84;
  assign n11903 = n11902 ^ x85;
  assign n11904 = n11503 & ~n11720;
  assign n11905 = n11904 ^ n11505;
  assign n11906 = n11905 ^ n11902;
  assign n11907 = n11903 & n11906;
  assign n11908 = n11907 ^ x85;
  assign n11909 = n11908 ^ x86;
  assign n11910 = n11509 & ~n11720;
  assign n11911 = n11910 ^ n11511;
  assign n11912 = n11911 ^ n11908;
  assign n11913 = n11909 & n11912;
  assign n11914 = n11913 ^ x86;
  assign n11915 = n11914 ^ x87;
  assign n11916 = n11515 & ~n11720;
  assign n11917 = n11916 ^ n11517;
  assign n11918 = n11917 ^ n11914;
  assign n11919 = n11915 & ~n11918;
  assign n11920 = n11919 ^ x87;
  assign n11921 = n11920 ^ x88;
  assign n11922 = n11521 & ~n11720;
  assign n11923 = n11922 ^ n11523;
  assign n11924 = n11923 ^ n11920;
  assign n11925 = n11921 & n11924;
  assign n11926 = n11925 ^ x88;
  assign n11927 = n11926 ^ x89;
  assign n11928 = n11527 & ~n11720;
  assign n11929 = n11928 ^ n11529;
  assign n11930 = n11929 ^ n11926;
  assign n11931 = n11927 & n11930;
  assign n11932 = n11931 ^ x89;
  assign n11933 = n11932 ^ x90;
  assign n11934 = n11533 & ~n11720;
  assign n11935 = n11934 ^ n11535;
  assign n11936 = n11935 ^ n11932;
  assign n11937 = n11933 & ~n11936;
  assign n11938 = n11937 ^ x90;
  assign n11939 = n11938 ^ x91;
  assign n11940 = n11539 & ~n11720;
  assign n11941 = n11940 ^ n11541;
  assign n11942 = n11941 ^ n11938;
  assign n11943 = n11939 & n11942;
  assign n11944 = n11943 ^ x91;
  assign n11945 = n11944 ^ x92;
  assign n11946 = n11545 & ~n11720;
  assign n11947 = n11946 ^ n11547;
  assign n11948 = n11947 ^ n11944;
  assign n11949 = n11945 & n11948;
  assign n11950 = n11949 ^ x92;
  assign n11951 = n11950 ^ x93;
  assign n11952 = n11551 & ~n11720;
  assign n11953 = n11952 ^ n11553;
  assign n11954 = n11953 ^ n11950;
  assign n11955 = n11951 & n11954;
  assign n11956 = n11955 ^ x93;
  assign n11957 = n11956 ^ x94;
  assign n11958 = n11556 ^ x93;
  assign n11959 = ~n11720 & n11958;
  assign n11960 = n11959 ^ n11341;
  assign n11961 = n11960 ^ n11956;
  assign n11962 = n11957 & ~n11961;
  assign n11963 = n11962 ^ x94;
  assign n11964 = n11963 ^ x95;
  assign n11965 = n11556 ^ n11341;
  assign n11966 = n11958 & ~n11965;
  assign n11967 = n11966 ^ x93;
  assign n11968 = n11967 ^ x94;
  assign n11969 = ~n11720 & n11968;
  assign n11970 = n11969 ^ n11338;
  assign n11971 = n11970 ^ n11963;
  assign n11972 = n11964 & n11971;
  assign n11973 = n11972 ^ x95;
  assign n11974 = n11973 ^ x96;
  assign n11975 = ~n11564 & ~n11720;
  assign n11976 = n11975 ^ n11566;
  assign n11977 = n11976 ^ n11973;
  assign n11978 = n11974 & ~n11977;
  assign n11979 = n11978 ^ x96;
  assign n11980 = ~n11748 & n11979;
  assign n11981 = n11980 ^ n11741;
  assign n11982 = n11981 ^ n11741;
  assign n11983 = ~n11747 & ~n11982;
  assign n11984 = n11983 ^ n11741;
  assign n11985 = n11742 & n11984;
  assign n11986 = n11985 ^ x98;
  assign n11987 = n11986 ^ x99;
  assign n11988 = n11582 & ~n11720;
  assign n11989 = n11988 ^ n11584;
  assign n11990 = n11989 ^ n11986;
  assign n11991 = n11987 & ~n11990;
  assign n11992 = n11991 ^ x99;
  assign n11993 = n11992 ^ x100;
  assign n11994 = n11588 & ~n11720;
  assign n11995 = n11994 ^ n11590;
  assign n11996 = n11995 ^ n11992;
  assign n11997 = n11993 & ~n11996;
  assign n11998 = n11997 ^ x100;
  assign n11999 = n11998 ^ x101;
  assign n12000 = n11594 & ~n11720;
  assign n12001 = n12000 ^ n11596;
  assign n12002 = n12001 ^ n11998;
  assign n12003 = n11999 & ~n12002;
  assign n12004 = n12003 ^ x101;
  assign n12005 = n12004 ^ x102;
  assign n12006 = n11600 & ~n11720;
  assign n12007 = n12006 ^ n11602;
  assign n12008 = n12007 ^ n12004;
  assign n12009 = n12005 & ~n12008;
  assign n12010 = n12009 ^ x102;
  assign n12011 = n12010 ^ x103;
  assign n12012 = n11606 & ~n11720;
  assign n12013 = n12012 ^ n11608;
  assign n12014 = n12013 ^ n12010;
  assign n12015 = n12011 & ~n12014;
  assign n12016 = n12015 ^ x103;
  assign n12017 = n12016 ^ x104;
  assign n12018 = n11612 & ~n11720;
  assign n12019 = n12018 ^ n11614;
  assign n12020 = n12019 ^ n12016;
  assign n12021 = n12017 & n12020;
  assign n12022 = n12021 ^ x104;
  assign n12023 = n12022 ^ x105;
  assign n12024 = n11618 & ~n11720;
  assign n12025 = n12024 ^ n11620;
  assign n12026 = n12025 ^ n12022;
  assign n12027 = n12023 & ~n12026;
  assign n12028 = n12027 ^ x105;
  assign n12029 = n12028 ^ x106;
  assign n12030 = n11624 & ~n11720;
  assign n12031 = n12030 ^ n11626;
  assign n12032 = n12031 ^ n12028;
  assign n12033 = n12029 & n12032;
  assign n12034 = n12033 ^ x106;
  assign n12035 = n11739 & n12034;
  assign n12036 = n11734 ^ x108;
  assign n12037 = x107 & n11737;
  assign n12038 = n12037 ^ n11734;
  assign n12039 = n12036 & ~n12038;
  assign n12040 = n12039 ^ x108;
  assign n12041 = ~n12035 & ~n12040;
  assign n12042 = n12041 ^ x109;
  assign n12043 = n11645 ^ x108;
  assign n12044 = n12043 ^ n11641;
  assign n12045 = n12044 ^ n11645;
  assign n12046 = ~n11720 & n12045;
  assign n12047 = n12046 ^ n11645;
  assign n12048 = n12047 ^ n12041;
  assign n12049 = ~n12042 & ~n12048;
  assign n12050 = n12049 ^ x109;
  assign n12051 = n12050 ^ x110;
  assign n12052 = n11649 & ~n11720;
  assign n12053 = n12052 ^ n11655;
  assign n12054 = n12053 ^ n12050;
  assign n12055 = n12051 & n12054;
  assign n12056 = n12055 ^ x110;
  assign n12057 = n12056 ^ x111;
  assign n12058 = n11659 & ~n11720;
  assign n12059 = n12058 ^ n11661;
  assign n12060 = n12059 ^ n12056;
  assign n12061 = n12057 & n12060;
  assign n12062 = n12061 ^ x111;
  assign n12063 = n12062 ^ x112;
  assign n11721 = n11705 ^ x117;
  assign n11722 = ~n11720 & n11721;
  assign n11723 = n11722 ^ n11331;
  assign n11724 = ~x118 & ~n11723;
  assign n11725 = n11705 ^ n11331;
  assign n11726 = n11721 & ~n11725;
  assign n11727 = n11726 ^ x117;
  assign n11728 = n11727 ^ x118;
  assign n11729 = ~n11720 & n11728;
  assign n11730 = n11729 ^ n11334;
  assign n11731 = ~x119 & n11730;
  assign n11732 = ~n11724 & ~n11731;
  assign n12064 = n11665 & ~n11720;
  assign n12065 = n12064 ^ n11667;
  assign n12066 = n12065 ^ n12062;
  assign n12067 = n12063 & ~n12066;
  assign n12068 = n12067 ^ x112;
  assign n12069 = n12068 ^ x113;
  assign n12070 = n11671 & ~n11720;
  assign n12071 = n12070 ^ n11673;
  assign n12072 = n12071 ^ n12068;
  assign n12073 = n12069 & ~n12072;
  assign n12074 = n12073 ^ x113;
  assign n12075 = n12074 ^ x114;
  assign n12076 = n11677 & ~n11720;
  assign n12077 = n12076 ^ n11679;
  assign n12078 = n12077 ^ n12074;
  assign n12079 = n12075 & ~n12078;
  assign n12080 = n12079 ^ x114;
  assign n12081 = n12080 ^ x115;
  assign n12082 = n11683 & ~n11720;
  assign n12083 = n12082 ^ n11686;
  assign n12084 = n12083 ^ n12080;
  assign n12085 = n12081 & ~n12084;
  assign n12086 = n12085 ^ x115;
  assign n12087 = n12086 ^ x116;
  assign n12088 = n11690 & ~n11720;
  assign n12089 = n12088 ^ n11696;
  assign n12090 = n12089 ^ n12086;
  assign n12091 = n12087 & ~n12090;
  assign n12092 = n12091 ^ x116;
  assign n12093 = n12092 ^ x117;
  assign n12094 = n11700 & ~n11720;
  assign n12095 = n12094 ^ n11702;
  assign n12096 = n12095 ^ n12092;
  assign n12097 = n12093 & n12096;
  assign n12098 = n12097 ^ x117;
  assign n12099 = n11732 & n12098;
  assign n12100 = n11730 ^ x119;
  assign n12101 = x118 & n11723;
  assign n12102 = n12101 ^ n11730;
  assign n12103 = ~n12100 & n12102;
  assign n12104 = n12103 ^ x119;
  assign n12105 = ~n12099 & ~n12104;
  assign n11713 = n11712 ^ x119;
  assign n11714 = n9801 & ~n11713;
  assign n11715 = n11311 & ~n11714;
  assign n12110 = ~x120 & n11715;
  assign n12111 = ~n12105 & ~n12110;
  assign n12112 = x120 & ~n10930;
  assign n12113 = n135 & ~n12112;
  assign n12114 = ~n12111 & n12113;
  assign n12115 = n12063 & n12114;
  assign n12116 = n12115 ^ n12065;
  assign n12117 = ~x113 & ~n12116;
  assign n12118 = n12057 & n12114;
  assign n12119 = n12118 ^ n12059;
  assign n12120 = ~x112 & n12119;
  assign n12121 = ~n12117 & ~n12120;
  assign n12122 = n12034 ^ x107;
  assign n12123 = n12114 & n12122;
  assign n12124 = n12123 ^ n11737;
  assign n12125 = ~x108 & ~n12124;
  assign n12126 = n12034 ^ n11737;
  assign n12127 = n12122 & ~n12126;
  assign n12128 = n12127 ^ x107;
  assign n12129 = n12128 ^ x108;
  assign n12130 = n12114 & n12129;
  assign n12131 = n12130 ^ n11734;
  assign n12132 = ~x109 & ~n12131;
  assign n12133 = ~n12125 & ~n12132;
  assign n12134 = n11987 & n12114;
  assign n12135 = n12134 ^ n11989;
  assign n12136 = n12135 ^ x100;
  assign n12137 = ~n11745 & ~n11980;
  assign n12138 = n12137 ^ x98;
  assign n12139 = n12114 & ~n12138;
  assign n12140 = n12139 ^ n11741;
  assign n12141 = x99 & n12140;
  assign n12142 = n12141 ^ n12135;
  assign n12143 = n12142 ^ n12135;
  assign n12144 = ~x99 & ~n12140;
  assign n12145 = n11964 & n12114;
  assign n12146 = n12145 ^ n11970;
  assign n12147 = n12146 ^ x96;
  assign n12148 = n11957 & n12114;
  assign n12149 = n12148 ^ n11960;
  assign n12150 = x95 & n12149;
  assign n12151 = n12150 ^ n12146;
  assign n12152 = n12151 ^ n12146;
  assign n12153 = ~x95 & ~n12149;
  assign n12154 = n11927 & n12114;
  assign n12155 = n12154 ^ n11929;
  assign n12156 = n12155 ^ x90;
  assign n12157 = n11921 & n12114;
  assign n12158 = n12157 ^ n11923;
  assign n12159 = x89 & ~n12158;
  assign n12160 = n12159 ^ n12155;
  assign n12161 = n12160 ^ n12155;
  assign n12162 = ~x89 & n12158;
  assign n12163 = n11848 & n12114;
  assign n12164 = n12163 ^ n11850;
  assign n12165 = ~x76 & n12164;
  assign n12166 = n11854 & n12114;
  assign n12167 = n12166 ^ n11856;
  assign n12168 = ~x77 & ~n12167;
  assign n12169 = ~n12165 & ~n12168;
  assign n12176 = x64 & ~n11720;
  assign n12170 = x7 & n11720;
  assign n12171 = ~n11765 & n12170;
  assign n12172 = ~n202 & ~n12171;
  assign n12173 = n11720 ^ x65;
  assign n12174 = n11766 & n12173;
  assign n12175 = n12172 & ~n12174;
  assign n12177 = n12176 ^ n12175;
  assign n12178 = n12175 ^ n11769;
  assign n12179 = n12175 ^ n12114;
  assign n12180 = n12175 & n12179;
  assign n12181 = n12180 ^ n12175;
  assign n12182 = n12178 & n12181;
  assign n12183 = n12182 ^ n12180;
  assign n12184 = n12183 ^ n12175;
  assign n12185 = n12184 ^ n12114;
  assign n12186 = ~n12177 & n12185;
  assign n12187 = n12186 ^ n12176;
  assign n12188 = n12187 ^ x8;
  assign n12189 = n12188 ^ x66;
  assign n12190 = x64 & n12114;
  assign n12191 = x6 & n11769;
  assign n12192 = n12191 ^ x7;
  assign n12193 = n12190 & n12192;
  assign n12194 = ~x6 & n288;
  assign n12195 = n12194 ^ x65;
  assign n12196 = ~x7 & n12195;
  assign n12197 = ~n12114 & n12196;
  assign n12198 = x64 ^ x7;
  assign n12199 = n12198 ^ x7;
  assign n12200 = x7 ^ x6;
  assign n12201 = n12199 & n12200;
  assign n12202 = n12201 ^ x7;
  assign n12203 = x65 & ~n12202;
  assign n12204 = ~n12197 & ~n12203;
  assign n12205 = ~n12193 & n12204;
  assign n12206 = n12205 ^ n12188;
  assign n12207 = ~n12189 & ~n12206;
  assign n12208 = n12207 ^ x66;
  assign n12209 = n12208 ^ x67;
  assign n12210 = ~n11780 & n12114;
  assign n12211 = n12210 ^ n11800;
  assign n12212 = n12211 ^ n12208;
  assign n12213 = n12209 & n12212;
  assign n12214 = n12213 ^ x67;
  assign n12215 = n12214 ^ x68;
  assign n12216 = n11804 & n12114;
  assign n12217 = n12216 ^ n11807;
  assign n12218 = n12217 ^ n12214;
  assign n12219 = n12215 & n12218;
  assign n12220 = n12219 ^ x68;
  assign n12221 = n12220 ^ x69;
  assign n12222 = n11811 & n12114;
  assign n12223 = n12222 ^ n11813;
  assign n12224 = n12223 ^ n12220;
  assign n12225 = n12221 & n12224;
  assign n12226 = n12225 ^ x69;
  assign n12227 = n12226 ^ x70;
  assign n12228 = n11817 & n12114;
  assign n12229 = n12228 ^ n11819;
  assign n12230 = n12229 ^ n12226;
  assign n12231 = n12227 & ~n12230;
  assign n12232 = n12231 ^ x70;
  assign n12233 = n12232 ^ x71;
  assign n12234 = n11823 & n12114;
  assign n12235 = n12234 ^ n11825;
  assign n12236 = n12235 ^ n12232;
  assign n12237 = n12233 & n12236;
  assign n12238 = n12237 ^ x71;
  assign n12239 = n12238 ^ x72;
  assign n12240 = n11829 & n12114;
  assign n12241 = n12240 ^ n11831;
  assign n12242 = n12241 ^ n12238;
  assign n12243 = n12239 & ~n12242;
  assign n12244 = n12243 ^ x72;
  assign n12245 = n12244 ^ x73;
  assign n12246 = n11834 ^ x72;
  assign n12247 = n12114 & n12246;
  assign n12248 = n12247 ^ n11760;
  assign n12249 = n12248 ^ n12244;
  assign n12250 = n12245 & n12249;
  assign n12251 = n12250 ^ x73;
  assign n12252 = n12251 ^ x74;
  assign n12253 = ~n11761 & ~n11835;
  assign n12254 = n12253 ^ x73;
  assign n12255 = n12114 & ~n12254;
  assign n12256 = n12255 ^ n11757;
  assign n12257 = n12256 ^ n12251;
  assign n12258 = n12252 & n12257;
  assign n12259 = n12258 ^ x74;
  assign n12260 = n12259 ^ x75;
  assign n12261 = n11842 & n12114;
  assign n12262 = n12261 ^ n11844;
  assign n12263 = n12262 ^ n12259;
  assign n12264 = n12260 & ~n12263;
  assign n12265 = n12264 ^ x75;
  assign n12266 = n12169 & n12265;
  assign n12267 = n12167 ^ x77;
  assign n12268 = x76 & ~n12164;
  assign n12269 = n12268 ^ n12167;
  assign n12270 = n12267 & ~n12269;
  assign n12271 = n12270 ^ x77;
  assign n12272 = ~n12266 & ~n12271;
  assign n12273 = n12272 ^ x78;
  assign n12274 = n11860 & n12114;
  assign n12275 = n12274 ^ n11862;
  assign n12276 = n12275 ^ n12272;
  assign n12277 = ~n12273 & n12276;
  assign n12278 = n12277 ^ x78;
  assign n12279 = n12278 ^ x79;
  assign n12280 = n11866 & n12114;
  assign n12281 = n12280 ^ n11868;
  assign n12282 = n12281 ^ n12278;
  assign n12283 = n12279 & n12282;
  assign n12284 = n12283 ^ x79;
  assign n12285 = n12284 ^ x80;
  assign n12286 = n11871 ^ x79;
  assign n12287 = n12114 & n12286;
  assign n12288 = n12287 ^ n11750;
  assign n12289 = n12288 ^ n12284;
  assign n12290 = n12285 & n12289;
  assign n12291 = n12290 ^ x80;
  assign n12292 = n12291 ^ x81;
  assign n12293 = n11871 ^ n11750;
  assign n12294 = n12286 & n12293;
  assign n12295 = n12294 ^ x79;
  assign n12296 = n12295 ^ x80;
  assign n12297 = n12114 & n12296;
  assign n12298 = n12297 ^ n11753;
  assign n12299 = n12298 ^ n12291;
  assign n12300 = n12292 & n12299;
  assign n12301 = n12300 ^ x81;
  assign n12302 = n12301 ^ x82;
  assign n12303 = ~n11879 & n12114;
  assign n12304 = n12303 ^ n11881;
  assign n12305 = n12304 ^ n12301;
  assign n12306 = n12302 & ~n12305;
  assign n12307 = n12306 ^ x82;
  assign n12308 = n12307 ^ x83;
  assign n12309 = n11885 & n12114;
  assign n12310 = n12309 ^ n11887;
  assign n12311 = n12310 ^ n12307;
  assign n12312 = n12308 & n12311;
  assign n12313 = n12312 ^ x83;
  assign n12314 = n12313 ^ x84;
  assign n12315 = n11891 & n12114;
  assign n12316 = n12315 ^ n11893;
  assign n12317 = n12316 ^ n12313;
  assign n12318 = n12314 & ~n12317;
  assign n12319 = n12318 ^ x84;
  assign n12320 = n12319 ^ x85;
  assign n12321 = n11897 & n12114;
  assign n12322 = n12321 ^ n11899;
  assign n12323 = n12322 ^ n12319;
  assign n12324 = n12320 & ~n12323;
  assign n12325 = n12324 ^ x85;
  assign n12326 = n12325 ^ x86;
  assign n12327 = n11903 & n12114;
  assign n12328 = n12327 ^ n11905;
  assign n12329 = n12328 ^ n12325;
  assign n12330 = n12326 & n12329;
  assign n12331 = n12330 ^ x86;
  assign n12332 = n12331 ^ x87;
  assign n12333 = n11909 & n12114;
  assign n12334 = n12333 ^ n11911;
  assign n12335 = n12334 ^ n12331;
  assign n12336 = n12332 & n12335;
  assign n12337 = n12336 ^ x87;
  assign n12338 = n12337 ^ x88;
  assign n12339 = n11915 & n12114;
  assign n12340 = n12339 ^ n11917;
  assign n12341 = n12340 ^ n12337;
  assign n12342 = n12338 & ~n12341;
  assign n12343 = n12342 ^ x88;
  assign n12344 = ~n12162 & n12343;
  assign n12345 = n12344 ^ n12155;
  assign n12346 = n12345 ^ n12155;
  assign n12347 = ~n12161 & ~n12346;
  assign n12348 = n12347 ^ n12155;
  assign n12349 = ~n12156 & ~n12348;
  assign n12350 = n12349 ^ x90;
  assign n12351 = n12350 ^ x91;
  assign n12352 = n11933 & n12114;
  assign n12353 = n12352 ^ n11935;
  assign n12354 = n12353 ^ n12350;
  assign n12355 = n12351 & ~n12354;
  assign n12356 = n12355 ^ x91;
  assign n12357 = n12356 ^ x92;
  assign n12358 = n11939 & n12114;
  assign n12359 = n12358 ^ n11941;
  assign n12360 = n12359 ^ n12356;
  assign n12361 = n12357 & n12360;
  assign n12362 = n12361 ^ x92;
  assign n12363 = n12362 ^ x93;
  assign n12364 = n11945 & n12114;
  assign n12365 = n12364 ^ n11947;
  assign n12366 = n12365 ^ n12362;
  assign n12367 = n12363 & n12366;
  assign n12368 = n12367 ^ x93;
  assign n12369 = n12368 ^ x94;
  assign n12370 = n11951 & n12114;
  assign n12371 = n12370 ^ n11953;
  assign n12372 = n12371 ^ n12368;
  assign n12373 = n12369 & n12372;
  assign n12374 = n12373 ^ x94;
  assign n12375 = ~n12153 & n12374;
  assign n12376 = n12375 ^ n12146;
  assign n12377 = n12376 ^ n12146;
  assign n12378 = ~n12152 & ~n12377;
  assign n12379 = n12378 ^ n12146;
  assign n12380 = ~n12147 & ~n12379;
  assign n12381 = n12380 ^ x96;
  assign n12382 = n12381 ^ x97;
  assign n12383 = n11974 & n12114;
  assign n12384 = n12383 ^ n11976;
  assign n12385 = n12384 ^ n12381;
  assign n12386 = n12382 & ~n12385;
  assign n12387 = n12386 ^ x97;
  assign n12388 = n12387 ^ x98;
  assign n12389 = n11979 ^ x97;
  assign n12390 = n12114 & n12389;
  assign n12391 = n12390 ^ n11744;
  assign n12392 = n12391 ^ n12387;
  assign n12393 = n12388 & ~n12392;
  assign n12394 = n12393 ^ x98;
  assign n12395 = ~n12144 & n12394;
  assign n12396 = n12395 ^ n12135;
  assign n12397 = n12396 ^ n12135;
  assign n12398 = ~n12143 & ~n12397;
  assign n12399 = n12398 ^ n12135;
  assign n12400 = n12136 & n12399;
  assign n12401 = n12400 ^ x100;
  assign n12402 = n12401 ^ x101;
  assign n12403 = n11993 & n12114;
  assign n12404 = n12403 ^ n11995;
  assign n12405 = n12404 ^ n12401;
  assign n12406 = n12402 & ~n12405;
  assign n12407 = n12406 ^ x101;
  assign n12408 = n12407 ^ x102;
  assign n12409 = n11999 & n12114;
  assign n12410 = n12409 ^ n12001;
  assign n12411 = n12410 ^ n12407;
  assign n12412 = n12408 & ~n12411;
  assign n12413 = n12412 ^ x102;
  assign n12414 = n12413 ^ x103;
  assign n12415 = n12005 & n12114;
  assign n12416 = n12415 ^ n12007;
  assign n12417 = n12416 ^ n12413;
  assign n12418 = n12414 & ~n12417;
  assign n12419 = n12418 ^ x103;
  assign n12420 = n12419 ^ x104;
  assign n12421 = n12011 & n12114;
  assign n12422 = n12421 ^ n12013;
  assign n12423 = n12422 ^ n12419;
  assign n12424 = n12420 & ~n12423;
  assign n12425 = n12424 ^ x104;
  assign n12426 = n12425 ^ x105;
  assign n12427 = n12017 & n12114;
  assign n12428 = n12427 ^ n12019;
  assign n12429 = n12428 ^ n12425;
  assign n12430 = n12426 & n12429;
  assign n12431 = n12430 ^ x105;
  assign n12432 = n12431 ^ x106;
  assign n12433 = n12023 & n12114;
  assign n12434 = n12433 ^ n12025;
  assign n12435 = n12434 ^ n12431;
  assign n12436 = n12432 & ~n12435;
  assign n12437 = n12436 ^ x106;
  assign n12438 = n12437 ^ x107;
  assign n12439 = n12029 & n12114;
  assign n12440 = n12439 ^ n12031;
  assign n12441 = n12440 ^ n12437;
  assign n12442 = n12438 & n12441;
  assign n12443 = n12442 ^ x107;
  assign n12444 = n12133 & n12443;
  assign n12445 = n12131 ^ x109;
  assign n12446 = x108 & n12124;
  assign n12447 = n12446 ^ n12131;
  assign n12448 = n12445 & ~n12447;
  assign n12449 = n12448 ^ x109;
  assign n12450 = ~n12444 & ~n12449;
  assign n12451 = n12450 ^ x110;
  assign n12452 = ~n12042 & n12114;
  assign n12453 = n12452 ^ n12047;
  assign n12454 = n12453 ^ n12450;
  assign n12455 = ~n12451 & ~n12454;
  assign n12456 = n12455 ^ x110;
  assign n12457 = n12456 ^ x111;
  assign n12458 = n12051 & n12114;
  assign n12459 = n12458 ^ n12053;
  assign n12460 = n12459 ^ n12456;
  assign n12461 = n12457 & n12460;
  assign n12462 = n12461 ^ x111;
  assign n12463 = n12121 & n12462;
  assign n12464 = n12116 ^ x113;
  assign n12465 = x112 & ~n12119;
  assign n12466 = n12465 ^ n12116;
  assign n12467 = n12464 & ~n12466;
  assign n12468 = n12467 ^ x113;
  assign n12469 = ~n12463 & ~n12468;
  assign n12470 = n12469 ^ x114;
  assign n12471 = n12069 & n12114;
  assign n12472 = n12471 ^ n12071;
  assign n12473 = n12472 ^ n12469;
  assign n12474 = ~n12470 & n12473;
  assign n12475 = n12474 ^ x114;
  assign n12476 = n12475 ^ x115;
  assign n12477 = n12075 & n12114;
  assign n12478 = n12477 ^ n12077;
  assign n12479 = n12478 ^ n12475;
  assign n12480 = n12476 & ~n12479;
  assign n12481 = n12480 ^ x115;
  assign n12482 = n12481 ^ x116;
  assign n12483 = n12081 & n12114;
  assign n12484 = n12483 ^ n12083;
  assign n12485 = n12484 ^ n12481;
  assign n12486 = n12482 & ~n12485;
  assign n12487 = n12486 ^ x116;
  assign n12488 = n12487 ^ x117;
  assign n12489 = n12087 & n12114;
  assign n12490 = n12489 ^ n12089;
  assign n12491 = n12490 ^ n12487;
  assign n12492 = n12488 & ~n12491;
  assign n12493 = n12492 ^ x117;
  assign n12494 = n12493 ^ x118;
  assign n12495 = n12093 & n12114;
  assign n12496 = n12495 ^ n12095;
  assign n12497 = n12496 ^ n12493;
  assign n12498 = n12494 & n12497;
  assign n12499 = n12498 ^ x118;
  assign n12500 = n12499 ^ x119;
  assign n12106 = n12105 ^ x120;
  assign n12107 = n135 & ~n12106;
  assign n12108 = n11715 & ~n12107;
  assign n12109 = ~x121 & n12108;
  assign n12501 = n12098 ^ x118;
  assign n12502 = n12114 & n12501;
  assign n12503 = n12502 ^ n11723;
  assign n12504 = n12503 ^ n12499;
  assign n12505 = n12500 & ~n12504;
  assign n12506 = n12505 ^ x119;
  assign n12507 = n12506 ^ x120;
  assign n12508 = n12098 ^ n11723;
  assign n12509 = n12501 & ~n12508;
  assign n12510 = n12509 ^ x118;
  assign n12511 = n12510 ^ x119;
  assign n12512 = n12114 & n12511;
  assign n12513 = n12512 ^ n11730;
  assign n12514 = n12513 ^ n12506;
  assign n12515 = n12507 & n12514;
  assign n12516 = n12515 ^ x120;
  assign n12517 = ~n12109 & n12516;
  assign n12518 = x121 & ~n11311;
  assign n12519 = n134 & ~n12518;
  assign n12520 = ~n12517 & n12519;
  assign n12521 = n12500 & n12520;
  assign n12522 = n12521 ^ n12503;
  assign n12523 = n12522 ^ x120;
  assign n12524 = n12488 & n12520;
  assign n12525 = n12524 ^ n12490;
  assign n12526 = ~x118 & ~n12525;
  assign n12527 = ~n12470 & n12520;
  assign n12528 = n12527 ^ n12472;
  assign n12529 = n12528 ^ x115;
  assign n12530 = n12462 ^ x112;
  assign n12531 = n12462 ^ n12119;
  assign n12532 = n12530 & n12531;
  assign n12533 = n12532 ^ x112;
  assign n12534 = n12533 ^ x113;
  assign n12535 = n12520 & n12534;
  assign n12536 = n12535 ^ n12116;
  assign n12537 = x114 & n12536;
  assign n12538 = n12537 ^ n12528;
  assign n12539 = n12538 ^ n12528;
  assign n12540 = ~x114 & ~n12536;
  assign n12541 = n12432 & n12520;
  assign n12542 = n12541 ^ n12434;
  assign n12543 = ~x107 & ~n12542;
  assign n12544 = n12438 & n12520;
  assign n12545 = n12544 ^ n12440;
  assign n12546 = ~x108 & n12545;
  assign n12547 = ~n12543 & ~n12546;
  assign n12548 = n12363 & n12520;
  assign n12549 = n12548 ^ n12365;
  assign n12550 = n12549 ^ x94;
  assign n12551 = n12357 & n12520;
  assign n12552 = n12551 ^ n12359;
  assign n12553 = x93 & ~n12552;
  assign n12554 = n12553 ^ n12549;
  assign n12555 = n12554 ^ n12549;
  assign n12556 = ~x93 & n12552;
  assign n12557 = n12332 & n12520;
  assign n12558 = n12557 ^ n12334;
  assign n12559 = n12558 ^ x88;
  assign n12560 = n12326 & n12520;
  assign n12561 = n12560 ^ n12328;
  assign n12562 = x87 & ~n12561;
  assign n12563 = n12562 ^ n12558;
  assign n12564 = n12563 ^ n12558;
  assign n12565 = ~x87 & n12561;
  assign n12566 = n12265 ^ x76;
  assign n12567 = n12520 & n12566;
  assign n12568 = n12567 ^ n12164;
  assign n12569 = n12568 ^ x77;
  assign n12570 = n12260 & n12520;
  assign n12571 = n12570 ^ n12262;
  assign n12572 = x76 & n12571;
  assign n12573 = n12572 ^ n12568;
  assign n12574 = n12573 ^ n12568;
  assign n12575 = ~x76 & ~n12571;
  assign n12576 = n12520 ^ n288;
  assign n12577 = n12576 ^ n288;
  assign n12578 = n2322 & n12577;
  assign n12579 = n12578 ^ n288;
  assign n12580 = ~n12114 & n12579;
  assign n12581 = n12580 ^ n288;
  assign n12582 = x6 & n12581;
  assign n12583 = n289 & ~n12114;
  assign n12584 = n12583 ^ x65;
  assign n12585 = ~x6 & n12584;
  assign n12586 = ~n202 & ~n12585;
  assign n12587 = n12586 ^ n12190;
  assign n12588 = n12520 & ~n12587;
  assign n12589 = n12588 ^ n12190;
  assign n12590 = ~n12582 & ~n12589;
  assign n12591 = n12590 ^ x7;
  assign n12592 = n12591 ^ x66;
  assign n12593 = x6 & x64;
  assign n12594 = x5 & ~x65;
  assign n12595 = n12593 & ~n12594;
  assign n12596 = n12520 & n12595;
  assign n12598 = x65 ^ x6;
  assign n12605 = n12598 ^ x65;
  assign n12597 = x65 ^ x5;
  assign n12599 = n12598 ^ n12597;
  assign n12600 = n12599 ^ x65;
  assign n12601 = n12597 ^ x64;
  assign n12602 = n12601 ^ n12597;
  assign n12603 = n12602 ^ n12600;
  assign n12604 = ~n12600 & ~n12603;
  assign n12606 = n12605 ^ n12604;
  assign n12607 = n12606 ^ n12600;
  assign n12608 = n12520 ^ x65;
  assign n12609 = n12608 ^ x65;
  assign n12610 = n12604 ^ n12600;
  assign n12611 = ~n12609 & ~n12610;
  assign n12612 = n12611 ^ x65;
  assign n12613 = ~n12607 & n12612;
  assign n12614 = n12613 ^ x65;
  assign n12615 = n12614 ^ x65;
  assign n12616 = n12615 ^ x65;
  assign n12617 = ~n12596 & ~n12616;
  assign n12618 = n12617 ^ n12591;
  assign n12619 = n12592 & n12618;
  assign n12620 = n12619 ^ x66;
  assign n12621 = n12620 ^ x67;
  assign n12622 = n12205 ^ x66;
  assign n12623 = n12520 & ~n12622;
  assign n12624 = n12623 ^ n12188;
  assign n12625 = n12624 ^ n12620;
  assign n12626 = n12621 & n12625;
  assign n12627 = n12626 ^ x67;
  assign n12628 = n12627 ^ x68;
  assign n12629 = n12209 & n12520;
  assign n12630 = n12629 ^ n12211;
  assign n12631 = n12630 ^ n12627;
  assign n12632 = n12628 & n12631;
  assign n12633 = n12632 ^ x68;
  assign n12634 = n12633 ^ x69;
  assign n12635 = n12215 & n12520;
  assign n12636 = n12635 ^ n12217;
  assign n12637 = n12636 ^ n12633;
  assign n12638 = n12634 & n12637;
  assign n12639 = n12638 ^ x69;
  assign n12640 = n12639 ^ x70;
  assign n12641 = n12221 & n12520;
  assign n12642 = n12641 ^ n12223;
  assign n12643 = n12642 ^ n12639;
  assign n12644 = n12640 & n12643;
  assign n12645 = n12644 ^ x70;
  assign n12646 = n12645 ^ x71;
  assign n12647 = n12227 & n12520;
  assign n12648 = n12647 ^ n12229;
  assign n12649 = n12648 ^ n12645;
  assign n12650 = n12646 & ~n12649;
  assign n12651 = n12650 ^ x71;
  assign n12652 = n12651 ^ x72;
  assign n12653 = n12233 & n12520;
  assign n12654 = n12653 ^ n12235;
  assign n12655 = n12654 ^ n12651;
  assign n12656 = n12652 & n12655;
  assign n12657 = n12656 ^ x72;
  assign n12658 = n12657 ^ x73;
  assign n12659 = n12239 & n12520;
  assign n12660 = n12659 ^ n12241;
  assign n12661 = n12660 ^ n12657;
  assign n12662 = n12658 & ~n12661;
  assign n12663 = n12662 ^ x73;
  assign n12664 = n12663 ^ x74;
  assign n12665 = n12245 & n12520;
  assign n12666 = n12665 ^ n12248;
  assign n12667 = n12666 ^ n12663;
  assign n12668 = n12664 & n12667;
  assign n12669 = n12668 ^ x74;
  assign n12670 = n12669 ^ x75;
  assign n12671 = n12252 & n12520;
  assign n12672 = n12671 ^ n12256;
  assign n12673 = n12672 ^ n12669;
  assign n12674 = n12670 & n12673;
  assign n12675 = n12674 ^ x75;
  assign n12676 = ~n12575 & n12675;
  assign n12677 = n12676 ^ n12568;
  assign n12678 = n12677 ^ n12568;
  assign n12679 = ~n12574 & ~n12678;
  assign n12680 = n12679 ^ n12568;
  assign n12681 = ~n12569 & ~n12680;
  assign n12682 = n12681 ^ x77;
  assign n12683 = n12682 ^ x78;
  assign n12684 = n12265 ^ n12164;
  assign n12685 = n12566 & n12684;
  assign n12686 = n12685 ^ x76;
  assign n12687 = n12686 ^ x77;
  assign n12688 = n12520 & n12687;
  assign n12689 = n12688 ^ n12167;
  assign n12690 = n12689 ^ n12682;
  assign n12691 = n12683 & ~n12690;
  assign n12692 = n12691 ^ x78;
  assign n12693 = n12692 ^ x79;
  assign n12694 = ~n12273 & n12520;
  assign n12695 = n12694 ^ n12275;
  assign n12696 = n12695 ^ n12692;
  assign n12697 = n12693 & ~n12696;
  assign n12698 = n12697 ^ x79;
  assign n12699 = n12698 ^ x80;
  assign n12700 = n12279 & n12520;
  assign n12701 = n12700 ^ n12281;
  assign n12702 = n12701 ^ n12698;
  assign n12703 = n12699 & n12702;
  assign n12704 = n12703 ^ x80;
  assign n12705 = n12704 ^ x81;
  assign n12706 = n12285 & n12520;
  assign n12707 = n12706 ^ n12288;
  assign n12708 = n12707 ^ n12704;
  assign n12709 = n12705 & n12708;
  assign n12710 = n12709 ^ x81;
  assign n12711 = n12710 ^ x82;
  assign n12712 = n12292 & n12520;
  assign n12713 = n12712 ^ n12298;
  assign n12714 = n12713 ^ n12710;
  assign n12715 = n12711 & n12714;
  assign n12716 = n12715 ^ x82;
  assign n12717 = n12716 ^ x83;
  assign n12718 = n12302 & n12520;
  assign n12719 = n12718 ^ n12304;
  assign n12720 = n12719 ^ n12716;
  assign n12721 = n12717 & ~n12720;
  assign n12722 = n12721 ^ x83;
  assign n12723 = n12722 ^ x84;
  assign n12724 = n12308 & n12520;
  assign n12725 = n12724 ^ n12310;
  assign n12726 = n12725 ^ n12722;
  assign n12727 = n12723 & n12726;
  assign n12728 = n12727 ^ x84;
  assign n12729 = n12728 ^ x85;
  assign n12730 = n12314 & n12520;
  assign n12731 = n12730 ^ n12316;
  assign n12732 = n12731 ^ n12728;
  assign n12733 = n12729 & ~n12732;
  assign n12734 = n12733 ^ x85;
  assign n12735 = n12734 ^ x86;
  assign n12736 = n12320 & n12520;
  assign n12737 = n12736 ^ n12322;
  assign n12738 = n12737 ^ n12734;
  assign n12739 = n12735 & ~n12738;
  assign n12740 = n12739 ^ x86;
  assign n12741 = ~n12565 & n12740;
  assign n12742 = n12741 ^ n12558;
  assign n12743 = n12742 ^ n12558;
  assign n12744 = ~n12564 & ~n12743;
  assign n12745 = n12744 ^ n12558;
  assign n12746 = ~n12559 & ~n12745;
  assign n12747 = n12746 ^ x88;
  assign n12748 = n12747 ^ x89;
  assign n12749 = n12338 & n12520;
  assign n12750 = n12749 ^ n12340;
  assign n12751 = n12750 ^ n12747;
  assign n12752 = n12748 & ~n12751;
  assign n12753 = n12752 ^ x89;
  assign n12754 = n12753 ^ x90;
  assign n12755 = n12343 ^ x89;
  assign n12756 = n12520 & n12755;
  assign n12757 = n12756 ^ n12158;
  assign n12758 = n12757 ^ n12753;
  assign n12759 = n12754 & n12758;
  assign n12760 = n12759 ^ x90;
  assign n12761 = n12760 ^ x91;
  assign n12762 = ~n12159 & ~n12344;
  assign n12763 = n12762 ^ x90;
  assign n12764 = n12520 & ~n12763;
  assign n12765 = n12764 ^ n12155;
  assign n12766 = n12765 ^ n12760;
  assign n12767 = n12761 & n12766;
  assign n12768 = n12767 ^ x91;
  assign n12769 = n12768 ^ x92;
  assign n12770 = n12351 & n12520;
  assign n12771 = n12770 ^ n12353;
  assign n12772 = n12771 ^ n12768;
  assign n12773 = n12769 & ~n12772;
  assign n12774 = n12773 ^ x92;
  assign n12775 = ~n12556 & n12774;
  assign n12776 = n12775 ^ n12549;
  assign n12777 = n12776 ^ n12549;
  assign n12778 = ~n12555 & ~n12777;
  assign n12779 = n12778 ^ n12549;
  assign n12780 = ~n12550 & ~n12779;
  assign n12781 = n12780 ^ x94;
  assign n12782 = n12781 ^ x95;
  assign n12783 = n12369 & n12520;
  assign n12784 = n12783 ^ n12371;
  assign n12785 = n12784 ^ n12781;
  assign n12786 = n12782 & n12785;
  assign n12787 = n12786 ^ x95;
  assign n12788 = n12787 ^ x96;
  assign n12789 = n12374 ^ x95;
  assign n12790 = n12520 & n12789;
  assign n12791 = n12790 ^ n12149;
  assign n12792 = n12791 ^ n12787;
  assign n12793 = n12788 & ~n12792;
  assign n12794 = n12793 ^ x96;
  assign n12795 = n12794 ^ x97;
  assign n12796 = ~n12150 & ~n12375;
  assign n12797 = n12796 ^ x96;
  assign n12798 = n12520 & ~n12797;
  assign n12799 = n12798 ^ n12146;
  assign n12800 = n12799 ^ n12794;
  assign n12801 = n12795 & n12800;
  assign n12802 = n12801 ^ x97;
  assign n12803 = n12802 ^ x98;
  assign n12804 = n12382 & n12520;
  assign n12805 = n12804 ^ n12384;
  assign n12806 = n12805 ^ n12802;
  assign n12807 = n12803 & ~n12806;
  assign n12808 = n12807 ^ x98;
  assign n12809 = n12808 ^ x99;
  assign n12810 = n12388 & n12520;
  assign n12811 = n12810 ^ n12391;
  assign n12812 = n12811 ^ n12808;
  assign n12813 = n12809 & ~n12812;
  assign n12814 = n12813 ^ x99;
  assign n12815 = n12814 ^ x100;
  assign n12816 = n12394 ^ x99;
  assign n12817 = n12520 & n12816;
  assign n12818 = n12817 ^ n12140;
  assign n12819 = n12818 ^ n12814;
  assign n12820 = n12815 & ~n12819;
  assign n12821 = n12820 ^ x100;
  assign n12822 = n12821 ^ x101;
  assign n12823 = ~n12141 & ~n12395;
  assign n12824 = n12823 ^ x100;
  assign n12825 = n12520 & ~n12824;
  assign n12826 = n12825 ^ n12135;
  assign n12827 = n12826 ^ n12821;
  assign n12828 = n12822 & ~n12827;
  assign n12829 = n12828 ^ x101;
  assign n12830 = n12829 ^ x102;
  assign n12831 = n12402 & n12520;
  assign n12832 = n12831 ^ n12404;
  assign n12833 = n12832 ^ n12829;
  assign n12834 = n12830 & ~n12833;
  assign n12835 = n12834 ^ x102;
  assign n12836 = n12835 ^ x103;
  assign n12837 = n12408 & n12520;
  assign n12838 = n12837 ^ n12410;
  assign n12839 = n12838 ^ n12835;
  assign n12840 = n12836 & ~n12839;
  assign n12841 = n12840 ^ x103;
  assign n12842 = n12841 ^ x104;
  assign n12843 = n12414 & n12520;
  assign n12844 = n12843 ^ n12416;
  assign n12845 = n12844 ^ n12841;
  assign n12846 = n12842 & ~n12845;
  assign n12847 = n12846 ^ x104;
  assign n12848 = n12847 ^ x105;
  assign n12849 = n12420 & n12520;
  assign n12850 = n12849 ^ n12422;
  assign n12851 = n12850 ^ n12847;
  assign n12852 = n12848 & ~n12851;
  assign n12853 = n12852 ^ x105;
  assign n12854 = n12853 ^ x106;
  assign n12855 = n12426 & n12520;
  assign n12856 = n12855 ^ n12428;
  assign n12857 = n12856 ^ n12853;
  assign n12858 = n12854 & n12857;
  assign n12859 = n12858 ^ x106;
  assign n12860 = n12547 & n12859;
  assign n12861 = n12545 ^ x108;
  assign n12862 = x107 & n12542;
  assign n12863 = n12862 ^ n12545;
  assign n12864 = ~n12861 & n12863;
  assign n12865 = n12864 ^ x108;
  assign n12866 = ~n12860 & ~n12865;
  assign n12867 = n12866 ^ x109;
  assign n12868 = n12443 ^ x108;
  assign n12869 = n12520 & n12868;
  assign n12870 = n12869 ^ n12124;
  assign n12871 = n12870 ^ n12866;
  assign n12872 = ~n12867 & n12871;
  assign n12873 = n12872 ^ x109;
  assign n12874 = n12873 ^ x110;
  assign n12875 = n12443 ^ n12124;
  assign n12876 = n12868 & ~n12875;
  assign n12877 = n12876 ^ x108;
  assign n12878 = n12877 ^ x109;
  assign n12879 = n12520 & n12878;
  assign n12880 = n12879 ^ n12131;
  assign n12881 = n12880 ^ n12873;
  assign n12882 = n12874 & ~n12881;
  assign n12883 = n12882 ^ x110;
  assign n12884 = n12883 ^ x111;
  assign n12885 = ~n12451 & n12520;
  assign n12886 = n12885 ^ n12453;
  assign n12887 = n12886 ^ n12883;
  assign n12888 = n12884 & n12887;
  assign n12889 = n12888 ^ x111;
  assign n12890 = n12889 ^ x112;
  assign n12891 = n12457 & n12520;
  assign n12892 = n12891 ^ n12459;
  assign n12893 = n12892 ^ n12889;
  assign n12894 = n12890 & n12893;
  assign n12895 = n12894 ^ x112;
  assign n12896 = n12895 ^ x113;
  assign n12897 = n12520 & n12530;
  assign n12898 = n12897 ^ n12119;
  assign n12899 = n12898 ^ n12895;
  assign n12900 = n12896 & n12899;
  assign n12901 = n12900 ^ x113;
  assign n12902 = ~n12540 & n12901;
  assign n12903 = n12902 ^ n12528;
  assign n12904 = n12903 ^ n12528;
  assign n12905 = ~n12539 & ~n12904;
  assign n12906 = n12905 ^ n12528;
  assign n12907 = n12529 & n12906;
  assign n12908 = n12907 ^ x115;
  assign n12909 = n12908 ^ x116;
  assign n12910 = n12476 & n12520;
  assign n12911 = n12910 ^ n12478;
  assign n12912 = n12911 ^ n12908;
  assign n12913 = n12909 & ~n12912;
  assign n12914 = n12913 ^ x116;
  assign n12915 = n12914 ^ x117;
  assign n12916 = n12482 & n12520;
  assign n12917 = n12916 ^ n12484;
  assign n12918 = n12917 ^ n12914;
  assign n12919 = n12915 & ~n12918;
  assign n12920 = n12919 ^ x117;
  assign n12921 = ~n12526 & n12920;
  assign n12922 = n12494 & n12520;
  assign n12923 = n12922 ^ n12496;
  assign n12924 = x119 & ~n12923;
  assign n12925 = x118 & n12525;
  assign n12926 = ~n12924 & ~n12925;
  assign n12927 = ~n12921 & n12926;
  assign n12928 = n12927 ^ n12522;
  assign n12929 = n12928 ^ n12522;
  assign n12930 = ~x119 & n12923;
  assign n12931 = n12930 ^ n12522;
  assign n12932 = n12931 ^ n12522;
  assign n12933 = ~n12929 & ~n12932;
  assign n12934 = n12933 ^ n12522;
  assign n12935 = n12523 & ~n12934;
  assign n12936 = n12935 ^ x120;
  assign n12937 = n12936 ^ x121;
  assign n12938 = n12507 & n12520;
  assign n12939 = n12938 ^ n12513;
  assign n12940 = n12939 ^ n12936;
  assign n12941 = n12937 & n12940;
  assign n12942 = n12941 ^ x121;
  assign n12943 = n133 & ~n12942;
  assign n12944 = n12109 & ~n12516;
  assign n12945 = ~n134 & n12108;
  assign n12946 = ~n12944 & ~n12945;
  assign n12947 = ~n12943 & ~n12946;
  assign n12948 = x127 & ~n12947;
  assign n13427 = ~x3 & x65;
  assign n12949 = x122 & ~n11715;
  assign n12950 = n132 & ~n12949;
  assign n12951 = ~n12942 & n12950;
  assign n12952 = n12516 ^ x121;
  assign n12953 = n12108 & ~n12952;
  assign n12954 = n134 & n12953;
  assign n12955 = ~n12951 & ~n12954;
  assign n12956 = n12937 & ~n12955;
  assign n12957 = n12956 ^ n12939;
  assign n12958 = x122 & ~n12957;
  assign n12959 = n12901 ^ x114;
  assign n12960 = ~n12955 & n12959;
  assign n12961 = n12960 ^ n12536;
  assign n12962 = n12961 ^ x115;
  assign n12963 = n12896 & ~n12955;
  assign n12964 = n12963 ^ n12898;
  assign n12965 = x114 & ~n12964;
  assign n12966 = n12859 ^ x107;
  assign n12967 = n12859 ^ n12542;
  assign n12968 = n12966 & ~n12967;
  assign n12969 = n12968 ^ x107;
  assign n12970 = n12969 ^ x108;
  assign n12971 = ~n12955 & n12970;
  assign n12972 = n12971 ^ n12545;
  assign n12973 = ~x109 & n12972;
  assign n12974 = ~n12955 & n12966;
  assign n12975 = n12974 ^ n12542;
  assign n12976 = ~x108 & ~n12975;
  assign n12977 = ~n12973 & ~n12976;
  assign n12978 = n12815 & ~n12955;
  assign n12979 = n12978 ^ n12818;
  assign n12980 = n12979 ^ x101;
  assign n12981 = n12809 & ~n12955;
  assign n12982 = n12981 ^ n12811;
  assign n12983 = x100 & n12982;
  assign n12984 = n12983 ^ n12979;
  assign n12985 = n12984 ^ n12979;
  assign n12986 = ~x100 & ~n12982;
  assign n12987 = n12761 & ~n12955;
  assign n12988 = n12987 ^ n12765;
  assign n12989 = ~x92 & n12988;
  assign n12990 = n12754 & ~n12955;
  assign n12991 = n12990 ^ n12757;
  assign n12992 = ~x91 & n12991;
  assign n12993 = ~n12989 & ~n12992;
  assign n12994 = n12705 & ~n12955;
  assign n12995 = n12994 ^ n12707;
  assign n12996 = ~x82 & n12995;
  assign n12997 = n12711 & ~n12955;
  assign n12998 = n12997 ^ n12713;
  assign n12999 = ~x83 & n12998;
  assign n13000 = ~n12996 & ~n12999;
  assign n13001 = n12699 & ~n12955;
  assign n13002 = n13001 ^ n12701;
  assign n13003 = n13002 ^ x81;
  assign n13004 = n12693 & ~n12955;
  assign n13005 = n13004 ^ n12695;
  assign n13006 = ~x80 & ~n13005;
  assign n13007 = n13006 ^ n13002;
  assign n13008 = n13007 ^ n13002;
  assign n13009 = x80 & n13005;
  assign n13010 = n12658 & ~n12955;
  assign n13011 = n13010 ^ n12660;
  assign n13012 = n13011 ^ x74;
  assign n13013 = n12652 & ~n12955;
  assign n13014 = n13013 ^ n12654;
  assign n13015 = ~x73 & n13014;
  assign n13016 = n12955 ^ n288;
  assign n13017 = n13016 ^ n288;
  assign n13018 = n2322 & ~n13017;
  assign n13019 = n13018 ^ n288;
  assign n13020 = ~n12520 & n13019;
  assign n13021 = n13020 ^ n288;
  assign n13022 = x5 & n13021;
  assign n13027 = x64 & n12520;
  assign n13023 = n289 & ~n12520;
  assign n13024 = n13023 ^ x65;
  assign n13025 = ~x5 & n13024;
  assign n13026 = ~n202 & ~n13025;
  assign n13028 = n13027 ^ n13026;
  assign n13029 = ~n12955 & ~n13028;
  assign n13030 = n13029 ^ n13027;
  assign n13031 = ~n13022 & ~n13030;
  assign n13032 = n13031 ^ x6;
  assign n13033 = n13032 ^ x66;
  assign n13038 = x4 & ~x65;
  assign n13039 = x5 & x64;
  assign n13040 = ~n13038 & n13039;
  assign n13034 = ~x5 & x64;
  assign n13035 = ~x4 & n13034;
  assign n13036 = ~x5 & x65;
  assign n13037 = ~n13035 & ~n13036;
  assign n13041 = n13040 ^ n13037;
  assign n13042 = n12955 & ~n13041;
  assign n13043 = n13042 ^ n13040;
  assign n13044 = ~x4 & x65;
  assign n13045 = n13044 ^ n13036;
  assign n13046 = x64 & n13045;
  assign n13047 = n13046 ^ n13036;
  assign n13048 = ~n13043 & ~n13047;
  assign n13049 = n13048 ^ n13032;
  assign n13050 = n13033 & n13049;
  assign n13051 = n13050 ^ x66;
  assign n13052 = n13051 ^ x67;
  assign n13053 = n12617 ^ x66;
  assign n13054 = ~n12955 & ~n13053;
  assign n13055 = n13054 ^ n12591;
  assign n13056 = n13055 ^ n13051;
  assign n13057 = n13052 & ~n13056;
  assign n13058 = n13057 ^ x67;
  assign n13059 = n13058 ^ x68;
  assign n13060 = n12621 & ~n12955;
  assign n13061 = n13060 ^ n12624;
  assign n13062 = n13061 ^ n13058;
  assign n13063 = n13059 & n13062;
  assign n13064 = n13063 ^ x68;
  assign n13065 = n13064 ^ x69;
  assign n13066 = n12628 & ~n12955;
  assign n13067 = n13066 ^ n12630;
  assign n13068 = n13067 ^ n13064;
  assign n13069 = n13065 & n13068;
  assign n13070 = n13069 ^ x69;
  assign n13071 = n13070 ^ x70;
  assign n13072 = n12634 & ~n12955;
  assign n13073 = n13072 ^ n12636;
  assign n13074 = n13073 ^ n13070;
  assign n13075 = n13071 & n13074;
  assign n13076 = n13075 ^ x70;
  assign n13077 = n13076 ^ x71;
  assign n13078 = n12640 & ~n12955;
  assign n13079 = n13078 ^ n12642;
  assign n13080 = n13079 ^ n13076;
  assign n13081 = n13077 & n13080;
  assign n13082 = n13081 ^ x71;
  assign n13083 = n13082 ^ x72;
  assign n13084 = n12646 & ~n12955;
  assign n13085 = n13084 ^ n12648;
  assign n13086 = n13085 ^ n13082;
  assign n13087 = n13083 & ~n13086;
  assign n13088 = n13087 ^ x72;
  assign n13089 = ~n13015 & n13088;
  assign n13090 = n13089 ^ n13011;
  assign n13091 = n13090 ^ n13011;
  assign n13092 = x73 & ~n13014;
  assign n13093 = n13092 ^ n13011;
  assign n13094 = n13093 ^ n13011;
  assign n13095 = ~n13091 & ~n13094;
  assign n13096 = n13095 ^ n13011;
  assign n13097 = n13012 & n13096;
  assign n13098 = n13097 ^ x74;
  assign n13099 = n13098 ^ x75;
  assign n13100 = n12664 & ~n12955;
  assign n13101 = n13100 ^ n12666;
  assign n13102 = n13101 ^ n13098;
  assign n13103 = n13099 & n13102;
  assign n13104 = n13103 ^ x75;
  assign n13105 = n13104 ^ x76;
  assign n13106 = n12670 & ~n12955;
  assign n13107 = n13106 ^ n12672;
  assign n13108 = n13107 ^ n13104;
  assign n13109 = n13105 & n13108;
  assign n13110 = n13109 ^ x76;
  assign n13111 = n13110 ^ x77;
  assign n13112 = n12675 ^ x76;
  assign n13113 = ~n12955 & n13112;
  assign n13114 = n13113 ^ n12571;
  assign n13115 = n13114 ^ n13110;
  assign n13116 = n13111 & ~n13115;
  assign n13117 = n13116 ^ x77;
  assign n13118 = n13117 ^ x78;
  assign n13119 = ~n12572 & ~n12676;
  assign n13120 = n13119 ^ x77;
  assign n13121 = ~n12955 & ~n13120;
  assign n13122 = n13121 ^ n12568;
  assign n13123 = n13122 ^ n13117;
  assign n13124 = n13118 & n13123;
  assign n13125 = n13124 ^ x78;
  assign n13126 = n13125 ^ x79;
  assign n13127 = n12683 & ~n12955;
  assign n13128 = n13127 ^ n12689;
  assign n13129 = n13128 ^ n13125;
  assign n13130 = n13126 & ~n13129;
  assign n13131 = n13130 ^ x79;
  assign n13132 = ~n13009 & ~n13131;
  assign n13133 = n13132 ^ n13002;
  assign n13134 = n13133 ^ n13002;
  assign n13135 = ~n13008 & ~n13134;
  assign n13136 = n13135 ^ n13002;
  assign n13137 = ~n13003 & n13136;
  assign n13138 = n13137 ^ x81;
  assign n13139 = n13000 & n13138;
  assign n13140 = n12998 ^ x83;
  assign n13141 = x82 & ~n12995;
  assign n13142 = n13141 ^ n12998;
  assign n13143 = ~n13140 & n13142;
  assign n13144 = n13143 ^ x83;
  assign n13145 = ~n13139 & ~n13144;
  assign n13146 = n12717 & ~n12955;
  assign n13147 = n13146 ^ n12719;
  assign n13148 = ~x84 & ~n13147;
  assign n13149 = n12723 & ~n12955;
  assign n13150 = n13149 ^ n12725;
  assign n13151 = ~x85 & n13150;
  assign n13152 = ~n13148 & ~n13151;
  assign n13153 = ~n13145 & n13152;
  assign n13154 = n13150 ^ x85;
  assign n13155 = x84 & n13147;
  assign n13156 = n13155 ^ n13150;
  assign n13157 = ~n13154 & n13156;
  assign n13158 = n13157 ^ x85;
  assign n13159 = ~n13153 & ~n13158;
  assign n13160 = n13159 ^ x86;
  assign n13161 = n12729 & ~n12955;
  assign n13162 = n13161 ^ n12731;
  assign n13163 = n13162 ^ n13159;
  assign n13164 = ~n13160 & n13163;
  assign n13165 = n13164 ^ x86;
  assign n13166 = n13165 ^ x87;
  assign n13167 = n12735 & ~n12955;
  assign n13168 = n13167 ^ n12737;
  assign n13169 = n13168 ^ n13165;
  assign n13170 = n13166 & ~n13169;
  assign n13171 = n13170 ^ x87;
  assign n13172 = n13171 ^ x88;
  assign n13173 = n12740 ^ x87;
  assign n13174 = ~n12955 & n13173;
  assign n13175 = n13174 ^ n12561;
  assign n13176 = n13175 ^ n13171;
  assign n13177 = n13172 & n13176;
  assign n13178 = n13177 ^ x88;
  assign n13179 = n13178 ^ x89;
  assign n13180 = ~n12562 & ~n12741;
  assign n13181 = n13180 ^ x88;
  assign n13182 = ~n12955 & ~n13181;
  assign n13183 = n13182 ^ n12558;
  assign n13184 = n13183 ^ n13178;
  assign n13185 = n13179 & n13184;
  assign n13186 = n13185 ^ x89;
  assign n13187 = n13186 ^ x90;
  assign n13188 = n12748 & ~n12955;
  assign n13189 = n13188 ^ n12750;
  assign n13190 = n13189 ^ n13186;
  assign n13191 = n13187 & ~n13190;
  assign n13192 = n13191 ^ x90;
  assign n13193 = n12993 & n13192;
  assign n13194 = n12988 ^ x92;
  assign n13195 = x91 & ~n12991;
  assign n13196 = n13195 ^ n12988;
  assign n13197 = ~n13194 & n13196;
  assign n13198 = n13197 ^ x92;
  assign n13199 = ~n13193 & ~n13198;
  assign n13200 = n13199 ^ x93;
  assign n13201 = n12769 & ~n12955;
  assign n13202 = n13201 ^ n12771;
  assign n13203 = n13202 ^ n13199;
  assign n13204 = ~n13200 & n13203;
  assign n13205 = n13204 ^ x93;
  assign n13206 = n13205 ^ x94;
  assign n13207 = n12774 ^ x93;
  assign n13208 = ~n12955 & n13207;
  assign n13209 = n13208 ^ n12552;
  assign n13210 = n13209 ^ n13205;
  assign n13211 = n13206 & n13210;
  assign n13212 = n13211 ^ x94;
  assign n13213 = n13212 ^ x95;
  assign n13214 = ~n12553 & ~n12775;
  assign n13215 = n13214 ^ x94;
  assign n13216 = ~n12955 & ~n13215;
  assign n13217 = n13216 ^ n12549;
  assign n13218 = n13217 ^ n13212;
  assign n13219 = n13213 & n13218;
  assign n13220 = n13219 ^ x95;
  assign n13221 = n13220 ^ x96;
  assign n13222 = n12782 & ~n12955;
  assign n13223 = n13222 ^ n12784;
  assign n13224 = n13223 ^ n13220;
  assign n13225 = n13221 & n13224;
  assign n13226 = n13225 ^ x96;
  assign n13227 = n13226 ^ x97;
  assign n13228 = n12788 & ~n12955;
  assign n13229 = n13228 ^ n12791;
  assign n13230 = n13229 ^ n13226;
  assign n13231 = n13227 & ~n13230;
  assign n13232 = n13231 ^ x97;
  assign n13233 = n13232 ^ x98;
  assign n13234 = n12795 & ~n12955;
  assign n13235 = n13234 ^ n12799;
  assign n13236 = n13235 ^ n13232;
  assign n13237 = n13233 & n13236;
  assign n13238 = n13237 ^ x98;
  assign n13239 = n13238 ^ x99;
  assign n13240 = n12803 & ~n12955;
  assign n13241 = n13240 ^ n12805;
  assign n13242 = n13241 ^ n13238;
  assign n13243 = n13239 & ~n13242;
  assign n13244 = n13243 ^ x99;
  assign n13245 = ~n12986 & n13244;
  assign n13246 = n13245 ^ n12979;
  assign n13247 = n13246 ^ n12979;
  assign n13248 = ~n12985 & ~n13247;
  assign n13249 = n13248 ^ n12979;
  assign n13250 = n12980 & n13249;
  assign n13251 = n13250 ^ x101;
  assign n13252 = n13251 ^ x102;
  assign n13253 = n12822 & ~n12955;
  assign n13254 = n13253 ^ n12826;
  assign n13255 = n13254 ^ n13251;
  assign n13256 = n13252 & ~n13255;
  assign n13257 = n13256 ^ x102;
  assign n13258 = n13257 ^ x103;
  assign n13259 = n12830 & ~n12955;
  assign n13260 = n13259 ^ n12832;
  assign n13261 = n13260 ^ n13257;
  assign n13262 = n13258 & ~n13261;
  assign n13263 = n13262 ^ x103;
  assign n13264 = n13263 ^ x104;
  assign n13265 = n12836 & ~n12955;
  assign n13266 = n13265 ^ n12838;
  assign n13267 = n13266 ^ n13263;
  assign n13268 = n13264 & ~n13267;
  assign n13269 = n13268 ^ x104;
  assign n13270 = n13269 ^ x105;
  assign n13271 = n12842 & ~n12955;
  assign n13272 = n13271 ^ n12844;
  assign n13273 = n13272 ^ n13269;
  assign n13274 = n13270 & ~n13273;
  assign n13275 = n13274 ^ x105;
  assign n13276 = n13275 ^ x106;
  assign n13277 = n12848 & ~n12955;
  assign n13278 = n13277 ^ n12850;
  assign n13279 = n13278 ^ n13275;
  assign n13280 = n13276 & ~n13279;
  assign n13281 = n13280 ^ x106;
  assign n13282 = n13281 ^ x107;
  assign n13283 = n12854 & ~n12955;
  assign n13284 = n13283 ^ n12856;
  assign n13285 = n13284 ^ n13281;
  assign n13286 = n13282 & n13285;
  assign n13287 = n13286 ^ x107;
  assign n13288 = n12977 & n13287;
  assign n13289 = n12972 ^ x109;
  assign n13290 = x108 & n12975;
  assign n13291 = n13290 ^ n12972;
  assign n13292 = ~n13289 & n13291;
  assign n13293 = n13292 ^ x109;
  assign n13294 = ~n13288 & ~n13293;
  assign n13295 = n13294 ^ x110;
  assign n13296 = ~n12867 & ~n12955;
  assign n13297 = n13296 ^ n12870;
  assign n13298 = n13297 ^ n13294;
  assign n13299 = ~n13295 & n13298;
  assign n13300 = n13299 ^ x110;
  assign n13301 = n13300 ^ x111;
  assign n13302 = n12874 & ~n12955;
  assign n13303 = n13302 ^ n12880;
  assign n13304 = n13303 ^ n13300;
  assign n13305 = n13301 & ~n13304;
  assign n13306 = n13305 ^ x111;
  assign n13307 = n13306 ^ x112;
  assign n13308 = n12884 & ~n12955;
  assign n13309 = n13308 ^ n12886;
  assign n13310 = n13309 ^ n13306;
  assign n13311 = n13307 & n13310;
  assign n13312 = n13311 ^ x112;
  assign n13313 = n13312 ^ x113;
  assign n13314 = n12890 & ~n12955;
  assign n13315 = n13314 ^ n12892;
  assign n13316 = n13315 ^ n13312;
  assign n13317 = n13313 & n13316;
  assign n13318 = n13317 ^ x113;
  assign n13319 = ~n12965 & ~n13318;
  assign n13320 = n13319 ^ n12961;
  assign n13321 = n13320 ^ n12961;
  assign n13322 = ~x114 & n12964;
  assign n13323 = n13322 ^ n12961;
  assign n13324 = n13323 ^ n12961;
  assign n13325 = ~n13321 & ~n13324;
  assign n13326 = n13325 ^ n12961;
  assign n13327 = n12962 & ~n13326;
  assign n13328 = n13327 ^ x115;
  assign n13329 = n13328 ^ x116;
  assign n13330 = ~n12537 & ~n12902;
  assign n13331 = n13330 ^ x115;
  assign n13332 = ~n12955 & ~n13331;
  assign n13333 = n13332 ^ n12528;
  assign n13334 = n13333 ^ n13328;
  assign n13335 = n13329 & ~n13334;
  assign n13336 = n13335 ^ x116;
  assign n13337 = n13336 ^ x117;
  assign n13338 = n12909 & ~n12955;
  assign n13339 = n13338 ^ n12911;
  assign n13340 = n13339 ^ n13336;
  assign n13341 = n13337 & ~n13340;
  assign n13342 = n13341 ^ x117;
  assign n13343 = n13342 ^ x118;
  assign n13344 = n12915 & ~n12955;
  assign n13345 = n13344 ^ n12917;
  assign n13346 = n13345 ^ n13342;
  assign n13347 = n13343 & ~n13346;
  assign n13348 = n13347 ^ x118;
  assign n13349 = n13348 ^ x119;
  assign n13350 = n12920 ^ x118;
  assign n13351 = ~n12955 & n13350;
  assign n13352 = n13351 ^ n12525;
  assign n13353 = n13352 ^ n13348;
  assign n13354 = n13349 & ~n13353;
  assign n13355 = n13354 ^ x119;
  assign n13356 = n13355 ^ x120;
  assign n13357 = ~n12921 & ~n12925;
  assign n13358 = n13357 ^ x119;
  assign n13359 = ~n12955 & ~n13358;
  assign n13360 = n13359 ^ n12923;
  assign n13361 = n13360 ^ n13355;
  assign n13362 = n13356 & n13361;
  assign n13363 = n13362 ^ x120;
  assign n13364 = n13363 ^ x121;
  assign n13365 = ~n12927 & ~n12930;
  assign n13366 = n13365 ^ x120;
  assign n13367 = ~n12955 & n13366;
  assign n13368 = n13367 ^ n12522;
  assign n13369 = n13368 ^ n13363;
  assign n13370 = n13364 & ~n13369;
  assign n13371 = n13370 ^ x121;
  assign n13372 = ~n12958 & ~n13371;
  assign n13373 = ~x122 & n12957;
  assign n13374 = ~n13372 & ~n13373;
  assign n13375 = n13374 ^ x123;
  assign n13376 = n12947 & n13375;
  assign n13377 = n131 & n13376;
  assign n13378 = n13377 ^ n12947;
  assign n13379 = ~x124 & n13378;
  assign n13380 = n11715 & ~n13374;
  assign n13381 = ~n12947 & ~n13373;
  assign n13382 = ~n13372 & n13381;
  assign n13383 = ~x123 & ~n13382;
  assign n13384 = ~n13380 & ~n13383;
  assign n13385 = n131 & ~n13384;
  assign n13386 = n13307 & n13385;
  assign n13387 = n13386 ^ n13309;
  assign n13388 = n13387 ^ x113;
  assign n13389 = n13301 & n13385;
  assign n13390 = n13389 ^ n13303;
  assign n13391 = x112 & n13390;
  assign n13392 = n13391 ^ n13387;
  assign n13393 = n13392 ^ n13387;
  assign n13394 = ~x112 & ~n13390;
  assign n13395 = n13206 & n13385;
  assign n13396 = n13395 ^ n13209;
  assign n13397 = ~x95 & n13396;
  assign n13398 = n13213 & n13385;
  assign n13399 = n13398 ^ n13217;
  assign n13400 = ~x96 & n13399;
  assign n13401 = ~n13397 & ~n13400;
  assign n13402 = n13166 & n13385;
  assign n13403 = n13402 ^ n13168;
  assign n13404 = ~x88 & ~n13403;
  assign n13405 = n13172 & n13385;
  assign n13406 = n13405 ^ n13175;
  assign n13407 = ~x89 & n13406;
  assign n13408 = ~n13404 & ~n13407;
  assign n13409 = n13088 ^ x73;
  assign n13410 = n13385 & n13409;
  assign n13411 = n13410 ^ n13014;
  assign n13412 = ~x74 & n13411;
  assign n13413 = ~n13089 & ~n13092;
  assign n13414 = n13413 ^ x74;
  assign n13415 = n13385 & ~n13414;
  assign n13416 = n13415 ^ n13011;
  assign n13417 = ~x75 & ~n13416;
  assign n13418 = ~n13412 & ~n13417;
  assign n13419 = x64 & n13385;
  assign n13420 = x4 & n13419;
  assign n13421 = x3 & ~x65;
  assign n13422 = n13420 & ~n13421;
  assign n13423 = ~x3 & x64;
  assign n13424 = ~x65 & ~n13423;
  assign n13425 = ~x4 & ~n13424;
  assign n13426 = ~n13385 & n13425;
  assign n13428 = x64 & n13427;
  assign n13429 = ~x64 & n13044;
  assign n13430 = ~n13428 & ~n13429;
  assign n13431 = ~n13426 & n13430;
  assign n13432 = ~n13422 & n13431;
  assign n13433 = n13432 ^ x66;
  assign n13434 = x65 & n131;
  assign n13435 = n13434 ^ n288;
  assign n13436 = n13435 ^ n288;
  assign n13437 = n13384 ^ n288;
  assign n13438 = n13437 ^ n288;
  assign n13439 = n13436 & ~n13438;
  assign n13440 = n13439 ^ n288;
  assign n13441 = n12955 & n13440;
  assign n13442 = n13441 ^ n288;
  assign n13443 = x4 & n13442;
  assign n13444 = ~x4 & n288;
  assign n13445 = n12955 & n13444;
  assign n13446 = ~n202 & ~n13445;
  assign n13447 = n13385 & ~n13446;
  assign n13448 = ~n13044 & ~n13384;
  assign n13449 = x64 & ~n12955;
  assign n13450 = ~n13448 & n13449;
  assign n13451 = ~n13447 & ~n13450;
  assign n13452 = ~n13443 & n13451;
  assign n13453 = n13452 ^ x5;
  assign n13454 = n13453 ^ n13432;
  assign n13455 = ~n13433 & n13454;
  assign n13456 = n13455 ^ x66;
  assign n13457 = ~x67 & ~n13456;
  assign n13458 = ~x66 & ~n13453;
  assign n13459 = x67 & ~n13432;
  assign n13460 = ~n13458 & n13459;
  assign n13461 = n1864 & n13453;
  assign n13462 = n13048 ^ x66;
  assign n13463 = n13385 & ~n13462;
  assign n13464 = n13463 ^ n13032;
  assign n13465 = ~n13461 & ~n13464;
  assign n13466 = ~n13460 & n13465;
  assign n13467 = ~n13457 & ~n13466;
  assign n13468 = n13467 ^ x68;
  assign n13469 = n13052 & n13385;
  assign n13470 = n13469 ^ n13055;
  assign n13471 = n13470 ^ n13467;
  assign n13472 = n13468 & ~n13471;
  assign n13473 = n13472 ^ x68;
  assign n13474 = n13473 ^ x69;
  assign n13475 = n13059 & n13385;
  assign n13476 = n13475 ^ n13061;
  assign n13477 = n13476 ^ n13473;
  assign n13478 = n13474 & n13477;
  assign n13479 = n13478 ^ x69;
  assign n13480 = n13479 ^ x70;
  assign n13481 = n13065 & n13385;
  assign n13482 = n13481 ^ n13067;
  assign n13483 = n13482 ^ n13479;
  assign n13484 = n13480 & n13483;
  assign n13485 = n13484 ^ x70;
  assign n13486 = n13485 ^ x71;
  assign n13487 = n13071 & n13385;
  assign n13488 = n13487 ^ n13073;
  assign n13489 = n13488 ^ n13485;
  assign n13490 = n13486 & n13489;
  assign n13491 = n13490 ^ x71;
  assign n13492 = n13491 ^ x72;
  assign n13493 = n13077 & n13385;
  assign n13494 = n13493 ^ n13079;
  assign n13495 = n13494 ^ n13491;
  assign n13496 = n13492 & n13495;
  assign n13497 = n13496 ^ x72;
  assign n13498 = n13497 ^ x73;
  assign n13499 = n13083 & n13385;
  assign n13500 = n13499 ^ n13085;
  assign n13501 = n13500 ^ n13497;
  assign n13502 = n13498 & ~n13501;
  assign n13503 = n13502 ^ x73;
  assign n13504 = n13418 & n13503;
  assign n13505 = n13416 ^ x75;
  assign n13506 = x74 & ~n13411;
  assign n13507 = n13506 ^ n13416;
  assign n13508 = n13505 & ~n13507;
  assign n13509 = n13508 ^ x75;
  assign n13510 = ~n13504 & ~n13509;
  assign n13511 = n13510 ^ x76;
  assign n13512 = n13099 & n13385;
  assign n13513 = n13512 ^ n13101;
  assign n13514 = n13513 ^ n13510;
  assign n13515 = ~n13511 & ~n13514;
  assign n13516 = n13515 ^ x76;
  assign n13517 = n13516 ^ x77;
  assign n13518 = n13105 & n13385;
  assign n13519 = n13518 ^ n13107;
  assign n13520 = n13519 ^ n13516;
  assign n13521 = n13517 & n13520;
  assign n13522 = n13521 ^ x77;
  assign n13523 = n13522 ^ x78;
  assign n13524 = n13111 & n13385;
  assign n13525 = n13524 ^ n13114;
  assign n13526 = n13525 ^ n13522;
  assign n13527 = n13523 & ~n13526;
  assign n13528 = n13527 ^ x78;
  assign n13529 = n13528 ^ x79;
  assign n13530 = n13118 & n13385;
  assign n13531 = n13530 ^ n13122;
  assign n13532 = n13531 ^ n13528;
  assign n13533 = n13529 & n13532;
  assign n13534 = n13533 ^ x79;
  assign n13535 = n13534 ^ x80;
  assign n13536 = n13126 & n13385;
  assign n13537 = n13536 ^ n13128;
  assign n13538 = n13537 ^ n13534;
  assign n13539 = n13535 & ~n13538;
  assign n13540 = n13539 ^ x80;
  assign n13541 = n13540 ^ x81;
  assign n13542 = n13131 ^ x80;
  assign n13543 = n13385 & n13542;
  assign n13544 = n13543 ^ n13005;
  assign n13545 = n13544 ^ n13540;
  assign n13546 = n13541 & ~n13545;
  assign n13547 = n13546 ^ x81;
  assign n13548 = n13547 ^ x82;
  assign n13549 = ~n13006 & ~n13132;
  assign n13550 = n13549 ^ x81;
  assign n13551 = n13385 & n13550;
  assign n13552 = n13551 ^ n13002;
  assign n13553 = n13552 ^ n13547;
  assign n13554 = n13548 & n13553;
  assign n13555 = n13554 ^ x82;
  assign n13556 = n13555 ^ x83;
  assign n13557 = n13138 ^ x82;
  assign n13558 = n13385 & n13557;
  assign n13559 = n13558 ^ n12995;
  assign n13560 = n13559 ^ n13555;
  assign n13561 = n13556 & n13560;
  assign n13562 = n13561 ^ x83;
  assign n13563 = n13562 ^ x84;
  assign n13564 = n13138 ^ n12995;
  assign n13565 = n13557 & n13564;
  assign n13566 = n13565 ^ x82;
  assign n13567 = n13566 ^ x83;
  assign n13568 = n13385 & n13567;
  assign n13569 = n13568 ^ n12998;
  assign n13570 = n13569 ^ n13562;
  assign n13571 = n13563 & n13570;
  assign n13572 = n13571 ^ x84;
  assign n13573 = n13572 ^ x85;
  assign n13574 = n13145 ^ x84;
  assign n13575 = n13385 & ~n13574;
  assign n13576 = n13575 ^ n13147;
  assign n13577 = n13576 ^ n13572;
  assign n13578 = n13573 & ~n13577;
  assign n13579 = n13578 ^ x85;
  assign n13580 = n13579 ^ x86;
  assign n13581 = n13147 ^ n13145;
  assign n13582 = ~n13574 & n13581;
  assign n13583 = n13582 ^ x84;
  assign n13584 = n13583 ^ x85;
  assign n13585 = n13385 & n13584;
  assign n13586 = n13585 ^ n13150;
  assign n13587 = n13586 ^ n13579;
  assign n13588 = n13580 & n13587;
  assign n13589 = n13588 ^ x86;
  assign n13590 = n13589 ^ x87;
  assign n13591 = ~n13160 & n13385;
  assign n13592 = n13591 ^ n13162;
  assign n13593 = n13592 ^ n13589;
  assign n13594 = n13590 & ~n13593;
  assign n13595 = n13594 ^ x87;
  assign n13596 = n13408 & n13595;
  assign n13597 = n13406 ^ x89;
  assign n13598 = x88 & n13403;
  assign n13599 = n13598 ^ n13406;
  assign n13600 = ~n13597 & n13599;
  assign n13601 = n13600 ^ x89;
  assign n13602 = ~n13596 & ~n13601;
  assign n13603 = n13602 ^ x90;
  assign n13604 = n13179 & n13385;
  assign n13605 = n13604 ^ n13183;
  assign n13606 = n13605 ^ n13602;
  assign n13607 = ~n13603 & ~n13606;
  assign n13608 = n13607 ^ x90;
  assign n13609 = n13608 ^ x91;
  assign n13610 = n13187 & n13385;
  assign n13611 = n13610 ^ n13189;
  assign n13612 = n13611 ^ n13608;
  assign n13613 = n13609 & ~n13612;
  assign n13614 = n13613 ^ x91;
  assign n13615 = n13614 ^ x92;
  assign n13616 = n13192 ^ x91;
  assign n13617 = n13385 & n13616;
  assign n13618 = n13617 ^ n12991;
  assign n13619 = n13618 ^ n13614;
  assign n13620 = n13615 & n13619;
  assign n13621 = n13620 ^ x92;
  assign n13622 = n13621 ^ x93;
  assign n13623 = n13192 ^ n12991;
  assign n13624 = n13616 & n13623;
  assign n13625 = n13624 ^ x91;
  assign n13626 = n13625 ^ x92;
  assign n13627 = n13385 & n13626;
  assign n13628 = n13627 ^ n12988;
  assign n13629 = n13628 ^ n13621;
  assign n13630 = n13622 & n13629;
  assign n13631 = n13630 ^ x93;
  assign n13632 = n13631 ^ x94;
  assign n13633 = ~n13200 & n13385;
  assign n13634 = n13633 ^ n13202;
  assign n13635 = n13634 ^ n13631;
  assign n13636 = n13632 & ~n13635;
  assign n13637 = n13636 ^ x94;
  assign n13638 = n13401 & n13637;
  assign n13639 = n13399 ^ x96;
  assign n13640 = x95 & ~n13396;
  assign n13641 = n13640 ^ n13399;
  assign n13642 = ~n13639 & n13641;
  assign n13643 = n13642 ^ x96;
  assign n13644 = ~n13638 & ~n13643;
  assign n13645 = n13644 ^ x97;
  assign n13646 = n13221 & n13385;
  assign n13647 = n13646 ^ n13223;
  assign n13648 = n13647 ^ n13644;
  assign n13649 = ~n13645 & ~n13648;
  assign n13650 = n13649 ^ x97;
  assign n13651 = n13650 ^ x98;
  assign n13652 = n13227 & n13385;
  assign n13653 = n13652 ^ n13229;
  assign n13654 = n13653 ^ n13650;
  assign n13655 = n13651 & ~n13654;
  assign n13656 = n13655 ^ x98;
  assign n13657 = n13656 ^ x99;
  assign n13658 = n13233 & n13385;
  assign n13659 = n13658 ^ n13235;
  assign n13660 = n13659 ^ n13656;
  assign n13661 = n13657 & n13660;
  assign n13662 = n13661 ^ x99;
  assign n13663 = n13662 ^ x100;
  assign n13664 = n13239 & n13385;
  assign n13665 = n13664 ^ n13241;
  assign n13666 = n13665 ^ n13662;
  assign n13667 = n13663 & ~n13666;
  assign n13668 = n13667 ^ x100;
  assign n13669 = n13668 ^ x101;
  assign n13670 = n13244 ^ x100;
  assign n13671 = n13385 & n13670;
  assign n13672 = n13671 ^ n12982;
  assign n13673 = n13672 ^ n13668;
  assign n13674 = n13669 & ~n13673;
  assign n13675 = n13674 ^ x101;
  assign n13676 = n13675 ^ x102;
  assign n13677 = ~n12983 & ~n13245;
  assign n13678 = n13677 ^ x101;
  assign n13679 = n13385 & ~n13678;
  assign n13680 = n13679 ^ n12979;
  assign n13681 = n13680 ^ n13675;
  assign n13682 = n13676 & ~n13681;
  assign n13683 = n13682 ^ x102;
  assign n13684 = n13683 ^ x103;
  assign n13685 = n13252 & n13385;
  assign n13686 = n13685 ^ n13254;
  assign n13687 = n13686 ^ n13683;
  assign n13688 = n13684 & ~n13687;
  assign n13689 = n13688 ^ x103;
  assign n13690 = n13689 ^ x104;
  assign n13691 = n13258 & n13385;
  assign n13692 = n13691 ^ n13260;
  assign n13693 = n13692 ^ n13689;
  assign n13694 = n13690 & ~n13693;
  assign n13695 = n13694 ^ x104;
  assign n13696 = n13695 ^ x105;
  assign n13697 = n13264 & n13385;
  assign n13698 = n13697 ^ n13266;
  assign n13699 = n13698 ^ n13695;
  assign n13700 = n13696 & ~n13699;
  assign n13701 = n13700 ^ x105;
  assign n13702 = n13701 ^ x106;
  assign n13703 = n13270 & n13385;
  assign n13704 = n13703 ^ n13272;
  assign n13705 = n13704 ^ n13701;
  assign n13706 = n13702 & ~n13705;
  assign n13707 = n13706 ^ x106;
  assign n13708 = n13707 ^ x107;
  assign n13709 = n13276 & n13385;
  assign n13710 = n13709 ^ n13278;
  assign n13711 = n13710 ^ n13707;
  assign n13712 = n13708 & ~n13711;
  assign n13713 = n13712 ^ x107;
  assign n13714 = n13713 ^ x108;
  assign n13715 = n13282 & n13385;
  assign n13716 = n13715 ^ n13284;
  assign n13717 = n13716 ^ n13713;
  assign n13718 = n13714 & n13717;
  assign n13719 = n13718 ^ x108;
  assign n13720 = n13719 ^ x109;
  assign n13721 = n13287 ^ x108;
  assign n13722 = n13385 & n13721;
  assign n13723 = n13722 ^ n12975;
  assign n13724 = n13723 ^ n13719;
  assign n13725 = n13720 & ~n13724;
  assign n13726 = n13725 ^ x109;
  assign n13727 = n13726 ^ x110;
  assign n13728 = n13287 ^ n12975;
  assign n13729 = n13721 & ~n13728;
  assign n13730 = n13729 ^ x108;
  assign n13731 = n13730 ^ x109;
  assign n13732 = n13385 & n13731;
  assign n13733 = n13732 ^ n12972;
  assign n13734 = n13733 ^ n13726;
  assign n13735 = n13727 & n13734;
  assign n13736 = n13735 ^ x110;
  assign n13737 = n13736 ^ x111;
  assign n13738 = ~n13295 & n13385;
  assign n13739 = n13738 ^ n13297;
  assign n13740 = n13739 ^ n13736;
  assign n13741 = n13737 & ~n13740;
  assign n13742 = n13741 ^ x111;
  assign n13743 = ~n13394 & n13742;
  assign n13744 = n13743 ^ n13387;
  assign n13745 = n13744 ^ n13387;
  assign n13746 = ~n13393 & ~n13745;
  assign n13747 = n13746 ^ n13387;
  assign n13748 = ~n13388 & ~n13747;
  assign n13749 = n13748 ^ x113;
  assign n13750 = n13749 ^ x114;
  assign n13751 = n13313 & n13385;
  assign n13752 = n13751 ^ n13315;
  assign n13753 = n13752 ^ n13749;
  assign n13754 = n13750 & n13753;
  assign n13755 = n13754 ^ x114;
  assign n13756 = n13755 ^ x115;
  assign n13757 = n13318 ^ x114;
  assign n13758 = n13385 & n13757;
  assign n13759 = n13758 ^ n12964;
  assign n13760 = n13759 ^ n13755;
  assign n13761 = n13756 & n13760;
  assign n13762 = n13761 ^ x115;
  assign n13763 = n13762 ^ x116;
  assign n13764 = ~n13319 & ~n13322;
  assign n13765 = n13764 ^ x115;
  assign n13766 = n13385 & n13765;
  assign n13767 = n13766 ^ n12961;
  assign n13768 = n13767 ^ n13762;
  assign n13769 = n13763 & ~n13768;
  assign n13770 = n13769 ^ x116;
  assign n13771 = n13770 ^ x117;
  assign n13772 = n13329 & n13385;
  assign n13773 = n13772 ^ n13333;
  assign n13774 = n13773 ^ n13770;
  assign n13775 = n13771 & ~n13774;
  assign n13776 = n13775 ^ x117;
  assign n13777 = n13776 ^ x118;
  assign n13778 = n13337 & n13385;
  assign n13779 = n13778 ^ n13339;
  assign n13780 = n13779 ^ n13776;
  assign n13781 = n13777 & ~n13780;
  assign n13782 = n13781 ^ x118;
  assign n13783 = n13782 ^ x119;
  assign n13784 = n13343 & n13385;
  assign n13785 = n13784 ^ n13345;
  assign n13786 = n13785 ^ n13782;
  assign n13787 = n13783 & ~n13786;
  assign n13788 = n13787 ^ x119;
  assign n13789 = n13788 ^ x120;
  assign n13790 = n13349 & n13385;
  assign n13791 = n13790 ^ n13352;
  assign n13792 = n13791 ^ n13788;
  assign n13793 = n13789 & ~n13792;
  assign n13794 = n13793 ^ x120;
  assign n13795 = n13794 ^ x121;
  assign n13796 = n13356 & n13385;
  assign n13797 = n13796 ^ n13360;
  assign n13798 = n13797 ^ n13794;
  assign n13799 = n13795 & n13798;
  assign n13800 = n13799 ^ x121;
  assign n13801 = n13800 ^ x122;
  assign n13802 = n13364 & n13385;
  assign n13803 = n13802 ^ n13368;
  assign n13804 = n13803 ^ n13800;
  assign n13805 = n13801 & ~n13804;
  assign n13806 = n13805 ^ x122;
  assign n13807 = n13806 ^ x123;
  assign n13808 = n13371 ^ x122;
  assign n13809 = n13385 & n13808;
  assign n13810 = n13809 ^ n12957;
  assign n13811 = n13810 ^ n13806;
  assign n13812 = n13807 & n13811;
  assign n13813 = n13812 ^ x123;
  assign n13814 = ~n13379 & n13813;
  assign n13815 = x124 & ~n12108;
  assign n13816 = n130 & ~n13815;
  assign n13817 = ~n13814 & n13816;
  assign n13847 = x64 & n13817;
  assign n13848 = n13427 & ~n13847;
  assign n13849 = n13419 ^ x4;
  assign n13850 = n13849 ^ n13817;
  assign n13851 = n13848 & ~n13850;
  assign n13852 = ~x66 & ~n13851;
  assign n13854 = ~x2 & ~x3;
  assign n13855 = ~n13817 & n13854;
  assign n13856 = ~x2 & x65;
  assign n13857 = ~n13855 & ~n13856;
  assign n13858 = ~n13849 & ~n13857;
  assign n13853 = x3 & n13817;
  assign n13859 = n13858 ^ n13853;
  assign n13860 = n13859 ^ n13858;
  assign n13861 = n13849 ^ x65;
  assign n13862 = x2 & ~x65;
  assign n13863 = ~n13861 & ~n13862;
  assign n13864 = n13863 ^ n13858;
  assign n13865 = n13860 & n13864;
  assign n13866 = n13865 ^ n13858;
  assign n13867 = x64 & n13866;
  assign n13868 = n13852 & ~n13867;
  assign n13869 = n13421 & ~n13817;
  assign n13870 = ~x2 & x64;
  assign n13871 = ~n13869 & n13870;
  assign n13872 = ~n13424 & n13817;
  assign n13873 = ~n13427 & n13849;
  assign n13874 = ~n13872 & n13873;
  assign n13875 = ~n13871 & n13874;
  assign n13876 = n13423 & ~n13856;
  assign n13877 = ~n13861 & n13876;
  assign n13878 = x3 & n13429;
  assign n13879 = ~n13877 & ~n13878;
  assign n13880 = n13817 & ~n13879;
  assign n13881 = ~n13875 & ~n13880;
  assign n13882 = ~n13868 & n13881;
  assign n13883 = n13882 ^ x67;
  assign n13884 = ~n13433 & n13817;
  assign n13885 = n13884 ^ n13453;
  assign n13886 = n13885 ^ n13882;
  assign n13887 = n13883 & ~n13886;
  assign n13888 = n13887 ^ x67;
  assign n13889 = n13888 ^ x68;
  assign n13818 = n13750 & n13817;
  assign n13819 = n13818 ^ n13752;
  assign n13820 = ~x115 & n13819;
  assign n13821 = n13756 & n13817;
  assign n13822 = n13821 ^ n13759;
  assign n13823 = ~x116 & n13822;
  assign n13824 = ~n13820 & ~n13823;
  assign n13825 = n13669 & n13817;
  assign n13826 = n13825 ^ n13672;
  assign n13827 = ~x102 & ~n13826;
  assign n13828 = n13676 & n13817;
  assign n13829 = n13828 ^ n13680;
  assign n13830 = ~x103 & ~n13829;
  assign n13831 = ~n13827 & ~n13830;
  assign n13832 = n13651 & n13817;
  assign n13833 = n13832 ^ n13653;
  assign n13834 = ~x99 & ~n13833;
  assign n13835 = n13657 & n13817;
  assign n13836 = n13835 ^ n13659;
  assign n13837 = ~x100 & n13836;
  assign n13838 = ~n13834 & ~n13837;
  assign n13839 = n13622 & n13817;
  assign n13840 = n13839 ^ n13628;
  assign n13841 = n13840 ^ x94;
  assign n13842 = n13615 & n13817;
  assign n13843 = n13842 ^ n13618;
  assign n13844 = x93 & ~n13843;
  assign n13845 = n13474 & n13817;
  assign n13846 = n13845 ^ n13476;
  assign n13890 = n13456 ^ x67;
  assign n13891 = n13817 & n13890;
  assign n13892 = n13891 ^ n13464;
  assign n13893 = n13892 ^ n13888;
  assign n13894 = n13889 & ~n13893;
  assign n13895 = n13894 ^ x68;
  assign n13896 = n13895 ^ x69;
  assign n13897 = n13468 & n13817;
  assign n13898 = n13897 ^ n13470;
  assign n13899 = n13898 ^ n13895;
  assign n13900 = n13896 & ~n13899;
  assign n13901 = n13900 ^ x69;
  assign n13902 = ~n13846 & n13901;
  assign n13903 = x70 & n13901;
  assign n13904 = ~n13902 & ~n13903;
  assign n13905 = n13480 & n13817;
  assign n13906 = n13905 ^ n13482;
  assign n13907 = ~n619 & n13906;
  assign n13908 = ~n13904 & ~n13907;
  assign n13909 = x71 & n13902;
  assign n13910 = n13906 ^ x71;
  assign n13911 = x70 & ~n13846;
  assign n13912 = n13911 ^ n13906;
  assign n13913 = ~n13910 & n13912;
  assign n13914 = n13913 ^ x71;
  assign n13915 = ~n13909 & ~n13914;
  assign n13916 = ~n13908 & n13915;
  assign n13917 = n13916 ^ x72;
  assign n13918 = n13486 & n13817;
  assign n13919 = n13918 ^ n13488;
  assign n13920 = n13919 ^ n13916;
  assign n13921 = ~n13917 & ~n13920;
  assign n13922 = n13921 ^ x72;
  assign n13923 = n13922 ^ x73;
  assign n13924 = n13492 & n13817;
  assign n13925 = n13924 ^ n13494;
  assign n13926 = n13925 ^ n13922;
  assign n13927 = n13923 & n13926;
  assign n13928 = n13927 ^ x73;
  assign n13929 = n13928 ^ x74;
  assign n13930 = n13498 & n13817;
  assign n13931 = n13930 ^ n13500;
  assign n13932 = n13931 ^ n13928;
  assign n13933 = n13929 & ~n13932;
  assign n13934 = n13933 ^ x74;
  assign n13935 = n13934 ^ x75;
  assign n13936 = n13503 ^ x74;
  assign n13937 = n13817 & n13936;
  assign n13938 = n13937 ^ n13411;
  assign n13939 = n13938 ^ n13934;
  assign n13940 = n13935 & n13939;
  assign n13941 = n13940 ^ x75;
  assign n13942 = n13941 ^ x76;
  assign n13943 = n13503 ^ n13411;
  assign n13944 = n13936 & n13943;
  assign n13945 = n13944 ^ x74;
  assign n13946 = n13945 ^ x75;
  assign n13947 = n13817 & n13946;
  assign n13948 = n13947 ^ n13416;
  assign n13949 = n13948 ^ n13941;
  assign n13950 = n13942 & ~n13949;
  assign n13951 = n13950 ^ x76;
  assign n13952 = n13951 ^ x77;
  assign n13953 = ~n13511 & n13817;
  assign n13954 = n13953 ^ n13513;
  assign n13955 = n13954 ^ n13951;
  assign n13956 = n13952 & n13955;
  assign n13957 = n13956 ^ x77;
  assign n13958 = n13957 ^ x78;
  assign n13959 = n13517 & n13817;
  assign n13960 = n13959 ^ n13519;
  assign n13961 = n13960 ^ n13957;
  assign n13962 = n13958 & n13961;
  assign n13963 = n13962 ^ x78;
  assign n13964 = n13963 ^ x79;
  assign n13965 = n13523 & n13817;
  assign n13966 = n13965 ^ n13525;
  assign n13967 = n13966 ^ n13963;
  assign n13968 = n13964 & ~n13967;
  assign n13969 = n13968 ^ x79;
  assign n13970 = n13969 ^ x80;
  assign n13971 = n13529 & n13817;
  assign n13972 = n13971 ^ n13531;
  assign n13973 = n13972 ^ n13969;
  assign n13974 = n13970 & n13973;
  assign n13975 = n13974 ^ x80;
  assign n13976 = n13975 ^ x81;
  assign n13977 = n13535 & n13817;
  assign n13978 = n13977 ^ n13537;
  assign n13979 = n13978 ^ n13975;
  assign n13980 = n13976 & ~n13979;
  assign n13981 = n13980 ^ x81;
  assign n13982 = n13981 ^ x82;
  assign n13983 = n13541 & n13817;
  assign n13984 = n13983 ^ n13544;
  assign n13985 = n13984 ^ n13981;
  assign n13986 = n13982 & ~n13985;
  assign n13987 = n13986 ^ x82;
  assign n13988 = n13987 ^ x83;
  assign n13989 = n13548 & n13817;
  assign n13990 = n13989 ^ n13552;
  assign n13991 = n13990 ^ n13987;
  assign n13992 = n13988 & n13991;
  assign n13993 = n13992 ^ x83;
  assign n13994 = n13993 ^ x84;
  assign n13995 = n13556 & n13817;
  assign n13996 = n13995 ^ n13559;
  assign n13997 = n13996 ^ n13993;
  assign n13998 = n13994 & n13997;
  assign n13999 = n13998 ^ x84;
  assign n14000 = n13999 ^ x85;
  assign n14001 = n13563 & n13817;
  assign n14002 = n14001 ^ n13569;
  assign n14003 = n14002 ^ n13999;
  assign n14004 = n14000 & n14003;
  assign n14005 = n14004 ^ x85;
  assign n14006 = n14005 ^ x86;
  assign n14007 = n13573 & n13817;
  assign n14008 = n14007 ^ n13576;
  assign n14009 = n14008 ^ n14005;
  assign n14010 = n14006 & ~n14009;
  assign n14011 = n14010 ^ x86;
  assign n14012 = n14011 ^ x87;
  assign n14013 = n13580 & n13817;
  assign n14014 = n14013 ^ n13586;
  assign n14015 = n14014 ^ n14011;
  assign n14016 = n14012 & n14015;
  assign n14017 = n14016 ^ x87;
  assign n14018 = n14017 ^ x88;
  assign n14019 = n13590 & n13817;
  assign n14020 = n14019 ^ n13592;
  assign n14021 = n14020 ^ n14017;
  assign n14022 = n14018 & ~n14021;
  assign n14023 = n14022 ^ x88;
  assign n14024 = n14023 ^ x89;
  assign n14025 = n13595 ^ x88;
  assign n14026 = n13817 & n14025;
  assign n14027 = n14026 ^ n13403;
  assign n14028 = n14027 ^ n14023;
  assign n14029 = n14024 & ~n14028;
  assign n14030 = n14029 ^ x89;
  assign n14031 = n14030 ^ x90;
  assign n14032 = n13595 ^ n13403;
  assign n14033 = n14025 & ~n14032;
  assign n14034 = n14033 ^ x88;
  assign n14035 = n14034 ^ x89;
  assign n14036 = n13817 & n14035;
  assign n14037 = n14036 ^ n13406;
  assign n14038 = n14037 ^ n14030;
  assign n14039 = n14031 & n14038;
  assign n14040 = n14039 ^ x90;
  assign n14041 = n14040 ^ x91;
  assign n14042 = ~n13603 & n13817;
  assign n14043 = n14042 ^ n13605;
  assign n14044 = n14043 ^ n14040;
  assign n14045 = n14041 & n14044;
  assign n14046 = n14045 ^ x91;
  assign n14047 = n14046 ^ x92;
  assign n14048 = n13609 & n13817;
  assign n14049 = n14048 ^ n13611;
  assign n14050 = n14049 ^ n14046;
  assign n14051 = n14047 & ~n14050;
  assign n14052 = n14051 ^ x92;
  assign n14053 = ~n13844 & ~n14052;
  assign n14054 = n14053 ^ n13840;
  assign n14055 = n14054 ^ n13840;
  assign n14056 = ~x93 & n13843;
  assign n14057 = n14056 ^ n13840;
  assign n14058 = n14057 ^ n13840;
  assign n14059 = ~n14055 & ~n14058;
  assign n14060 = n14059 ^ n13840;
  assign n14061 = ~n13841 & n14060;
  assign n14062 = n14061 ^ x94;
  assign n14063 = n14062 ^ x95;
  assign n14064 = n13632 & n13817;
  assign n14065 = n14064 ^ n13634;
  assign n14066 = n14065 ^ n14062;
  assign n14067 = n14063 & ~n14066;
  assign n14068 = n14067 ^ x95;
  assign n14069 = n14068 ^ x96;
  assign n14070 = n13637 ^ x95;
  assign n14071 = n13817 & n14070;
  assign n14072 = n14071 ^ n13396;
  assign n14073 = n14072 ^ n14068;
  assign n14074 = n14069 & n14073;
  assign n14075 = n14074 ^ x96;
  assign n14076 = n14075 ^ x97;
  assign n14077 = n13637 ^ n13396;
  assign n14078 = n14070 & n14077;
  assign n14079 = n14078 ^ x95;
  assign n14080 = n14079 ^ x96;
  assign n14081 = n13817 & n14080;
  assign n14082 = n14081 ^ n13399;
  assign n14083 = n14082 ^ n14075;
  assign n14084 = n14076 & n14083;
  assign n14085 = n14084 ^ x97;
  assign n14086 = n14085 ^ x98;
  assign n14087 = ~n13645 & n13817;
  assign n14088 = n14087 ^ n13647;
  assign n14089 = n14088 ^ n14085;
  assign n14090 = n14086 & n14089;
  assign n14091 = n14090 ^ x98;
  assign n14092 = n13838 & n14091;
  assign n14093 = n13836 ^ x100;
  assign n14094 = x99 & n13833;
  assign n14095 = n14094 ^ n13836;
  assign n14096 = ~n14093 & n14095;
  assign n14097 = n14096 ^ x100;
  assign n14098 = ~n14092 & ~n14097;
  assign n14099 = n14098 ^ x101;
  assign n14100 = n13663 & n13817;
  assign n14101 = n14100 ^ n13665;
  assign n14102 = n14101 ^ n14098;
  assign n14103 = ~n14099 & n14102;
  assign n14104 = n14103 ^ x101;
  assign n14105 = n13831 & n14104;
  assign n14106 = n13829 ^ x103;
  assign n14107 = x102 & n13826;
  assign n14108 = n14107 ^ n13829;
  assign n14109 = n14106 & ~n14108;
  assign n14110 = n14109 ^ x103;
  assign n14111 = ~n14105 & ~n14110;
  assign n14112 = n14111 ^ x104;
  assign n14113 = n13684 & n13817;
  assign n14114 = n14113 ^ n13686;
  assign n14115 = n14114 ^ n14111;
  assign n14116 = ~n14112 & n14115;
  assign n14117 = n14116 ^ x104;
  assign n14118 = n14117 ^ x105;
  assign n14119 = n13690 & n13817;
  assign n14120 = n14119 ^ n13692;
  assign n14121 = n14120 ^ n14117;
  assign n14122 = n14118 & ~n14121;
  assign n14123 = n14122 ^ x105;
  assign n14124 = n14123 ^ x106;
  assign n14125 = n13696 & n13817;
  assign n14126 = n14125 ^ n13698;
  assign n14127 = n14126 ^ n14123;
  assign n14128 = n14124 & ~n14127;
  assign n14129 = n14128 ^ x106;
  assign n14130 = n14129 ^ x107;
  assign n14131 = n13702 & n13817;
  assign n14132 = n14131 ^ n13704;
  assign n14133 = n14132 ^ n14129;
  assign n14134 = n14130 & ~n14133;
  assign n14135 = n14134 ^ x107;
  assign n14136 = n14135 ^ x108;
  assign n14137 = n13708 & n13817;
  assign n14138 = n14137 ^ n13710;
  assign n14139 = n14138 ^ n14135;
  assign n14140 = n14136 & ~n14139;
  assign n14141 = n14140 ^ x108;
  assign n14142 = n14141 ^ x109;
  assign n14143 = n13714 & n13817;
  assign n14144 = n14143 ^ n13716;
  assign n14145 = n14144 ^ n14141;
  assign n14146 = n14142 & n14145;
  assign n14147 = n14146 ^ x109;
  assign n14148 = n14147 ^ x110;
  assign n14149 = n13720 & n13817;
  assign n14150 = n14149 ^ n13723;
  assign n14151 = n14150 ^ n14147;
  assign n14152 = n14148 & ~n14151;
  assign n14153 = n14152 ^ x110;
  assign n14154 = n14153 ^ x111;
  assign n14155 = n13727 & n13817;
  assign n14156 = n14155 ^ n13733;
  assign n14157 = n14156 ^ n14153;
  assign n14158 = n14154 & n14157;
  assign n14159 = n14158 ^ x111;
  assign n14160 = n14159 ^ x112;
  assign n14161 = n13737 & n13817;
  assign n14162 = n14161 ^ n13739;
  assign n14163 = n14162 ^ n14159;
  assign n14164 = n14160 & ~n14163;
  assign n14165 = n14164 ^ x112;
  assign n14166 = n14165 ^ x113;
  assign n14167 = n13742 ^ x112;
  assign n14168 = n13817 & n14167;
  assign n14169 = n14168 ^ n13390;
  assign n14170 = n14169 ^ n14165;
  assign n14171 = n14166 & ~n14170;
  assign n14172 = n14171 ^ x113;
  assign n14173 = n14172 ^ x114;
  assign n14174 = ~n13391 & ~n13743;
  assign n14175 = n14174 ^ x113;
  assign n14176 = n13817 & ~n14175;
  assign n14177 = n14176 ^ n13387;
  assign n14178 = n14177 ^ n14172;
  assign n14179 = n14173 & n14178;
  assign n14180 = n14179 ^ x114;
  assign n14181 = n13824 & n14180;
  assign n14182 = n13822 ^ x116;
  assign n14183 = x115 & ~n13819;
  assign n14184 = n14183 ^ n13822;
  assign n14185 = ~n14182 & n14184;
  assign n14186 = n14185 ^ x116;
  assign n14187 = ~n14181 & ~n14186;
  assign n14188 = n14187 ^ x117;
  assign n14189 = n13763 & n13817;
  assign n14190 = n14189 ^ n13767;
  assign n14191 = n14190 ^ n14187;
  assign n14192 = ~n14188 & n14191;
  assign n14193 = n14192 ^ x117;
  assign n14194 = n14193 ^ x118;
  assign n14195 = n13771 & n13817;
  assign n14196 = n14195 ^ n13773;
  assign n14197 = n14196 ^ n14193;
  assign n14198 = n14194 & ~n14197;
  assign n14199 = n14198 ^ x118;
  assign n14200 = n14199 ^ x119;
  assign n14201 = n13777 & n13817;
  assign n14202 = n14201 ^ n13779;
  assign n14203 = n14202 ^ n14199;
  assign n14204 = n14200 & ~n14203;
  assign n14205 = n14204 ^ x119;
  assign n14206 = n14205 ^ x120;
  assign n14207 = n13783 & n13817;
  assign n14208 = n14207 ^ n13785;
  assign n14209 = n14208 ^ n14205;
  assign n14210 = n14206 & ~n14209;
  assign n14211 = n14210 ^ x120;
  assign n14212 = n14211 ^ x121;
  assign n14213 = n13789 & n13817;
  assign n14214 = n14213 ^ n13791;
  assign n14215 = n14214 ^ n14211;
  assign n14216 = n14212 & ~n14215;
  assign n14217 = n14216 ^ x121;
  assign n14218 = n14217 ^ x122;
  assign n14219 = n13795 & n13817;
  assign n14220 = n14219 ^ n13797;
  assign n14221 = n14220 ^ n14217;
  assign n14222 = n14218 & n14221;
  assign n14223 = n14222 ^ x122;
  assign n14224 = n14223 ^ x123;
  assign n14225 = n13801 & n13817;
  assign n14226 = n14225 ^ n13803;
  assign n14227 = n14226 ^ n14223;
  assign n14228 = n14224 & ~n14227;
  assign n14229 = n14228 ^ x123;
  assign n14230 = n14229 ^ x124;
  assign n14231 = n13807 & n13817;
  assign n14232 = n14231 ^ n13810;
  assign n14233 = n14232 ^ n14229;
  assign n14234 = n14230 & n14233;
  assign n14235 = n14234 ^ x124;
  assign n14236 = n14235 ^ x125;
  assign n14237 = n14235 ^ n12108;
  assign n14238 = n14237 ^ n12108;
  assign n14239 = n13813 ^ x124;
  assign n14240 = n13378 & n14239;
  assign n14241 = n130 & n14240;
  assign n14242 = n14241 ^ n13378;
  assign n14243 = n14242 ^ n12108;
  assign n14244 = n14238 & ~n14243;
  assign n14245 = n14244 ^ n12108;
  assign n14246 = n14236 & n14245;
  assign n14247 = n14246 ^ x125;
  assign n14248 = n129 & ~n14247;
  assign n14274 = n13889 & n14248;
  assign n14275 = n14274 ^ n13892;
  assign n14276 = ~x69 & ~n14275;
  assign n14277 = n13883 & n14248;
  assign n14278 = n14277 ^ n13885;
  assign n14279 = ~x68 & ~n14278;
  assign n14280 = ~n14276 & ~n14279;
  assign n14281 = x64 & n14248;
  assign n14282 = x1 & n13862;
  assign n14283 = n14282 ^ x2;
  assign n14284 = n14281 & n14283;
  assign n14285 = ~x1 & n13870;
  assign n14286 = ~n13856 & ~n14285;
  assign n14287 = ~n14248 & ~n14286;
  assign n14288 = ~x1 & x65;
  assign n14289 = n14288 ^ n13856;
  assign n14290 = x64 & n14289;
  assign n14291 = n14290 ^ n13856;
  assign n14292 = ~n14287 & ~n14291;
  assign n14293 = ~n14284 & n14292;
  assign n14294 = n14293 ^ x66;
  assign n14295 = x65 & n14248;
  assign n14296 = ~n13847 & ~n13870;
  assign n14297 = n14295 & n14296;
  assign n14298 = ~x65 & n13870;
  assign n14299 = ~n13817 & n14298;
  assign n14300 = n14248 & n14299;
  assign n14301 = x65 ^ x2;
  assign n14302 = ~n14247 & ~n14301;
  assign n14303 = n13847 & ~n14302;
  assign n14304 = ~n14300 & ~n14303;
  assign n14305 = ~n14297 & n14304;
  assign n14306 = n14305 ^ x3;
  assign n14307 = n14306 ^ n14293;
  assign n14308 = ~n14294 & n14307;
  assign n14309 = n14308 ^ x66;
  assign n14310 = n14309 ^ x67;
  assign n14313 = n13853 & ~n13862;
  assign n14314 = n13857 & ~n14313;
  assign n14315 = x64 & ~n14314;
  assign n14316 = ~n13848 & ~n14315;
  assign n14317 = n14316 ^ x66;
  assign n14318 = n14248 & ~n14317;
  assign n14311 = ~n13428 & n13872;
  assign n14312 = n14311 ^ n13849;
  assign n14319 = n14318 ^ n14312;
  assign n14320 = n14319 ^ n14309;
  assign n14321 = n14310 & n14320;
  assign n14322 = n14321 ^ x67;
  assign n14323 = n14280 & n14322;
  assign n14324 = n14275 ^ x69;
  assign n14325 = x68 & n14278;
  assign n14326 = n14325 ^ n14275;
  assign n14327 = n14324 & ~n14326;
  assign n14328 = n14327 ^ x69;
  assign n14329 = ~n14323 & ~n14328;
  assign n14330 = n14329 ^ x70;
  assign n14331 = n13896 & n14248;
  assign n14332 = n14331 ^ n13898;
  assign n14333 = n14332 ^ n14329;
  assign n14334 = ~n14330 & n14333;
  assign n14335 = n14334 ^ x70;
  assign n14336 = n14335 ^ x71;
  assign n14337 = n13901 ^ x70;
  assign n14338 = n14248 & n14337;
  assign n14339 = n14338 ^ n13846;
  assign n14340 = n14339 ^ n14335;
  assign n14341 = n14336 & n14340;
  assign n14342 = n14341 ^ x71;
  assign n14343 = n14342 ^ x72;
  assign n14344 = n13904 & ~n13911;
  assign n14345 = n14344 ^ x71;
  assign n14346 = n14248 & ~n14345;
  assign n14347 = n14346 ^ n13906;
  assign n14348 = n14347 ^ n14342;
  assign n14349 = n14343 & n14348;
  assign n14350 = n14349 ^ x72;
  assign n14351 = n14350 ^ x73;
  assign n14352 = ~n13917 & n14248;
  assign n14353 = n14352 ^ n13919;
  assign n14354 = n14353 ^ n14350;
  assign n14355 = n14351 & n14354;
  assign n14356 = n14355 ^ x73;
  assign n14357 = n14356 ^ x74;
  assign n14358 = n13923 & n14248;
  assign n14359 = n14358 ^ n13925;
  assign n14360 = n14359 ^ n14356;
  assign n14361 = n14357 & n14360;
  assign n14362 = n14361 ^ x74;
  assign n14363 = n14362 ^ x75;
  assign n14364 = n13929 & n14248;
  assign n14365 = n14364 ^ n13931;
  assign n14366 = n14365 ^ n14362;
  assign n14367 = n14363 & ~n14366;
  assign n14368 = n14367 ^ x75;
  assign n14369 = n14368 ^ x76;
  assign n14370 = n13935 & n14248;
  assign n14371 = n14370 ^ n13938;
  assign n14372 = n14371 ^ n14368;
  assign n14373 = n14369 & n14372;
  assign n14374 = n14373 ^ x76;
  assign n14375 = n14374 ^ x77;
  assign n14376 = n13942 & n14248;
  assign n14377 = n14376 ^ n13948;
  assign n14378 = n14377 ^ n14374;
  assign n14379 = n14375 & ~n14378;
  assign n14380 = n14379 ^ x77;
  assign n14381 = n14380 ^ x78;
  assign n14382 = n13952 & n14248;
  assign n14383 = n14382 ^ n13954;
  assign n14384 = n14383 ^ n14380;
  assign n14385 = n14381 & n14384;
  assign n14386 = n14385 ^ x78;
  assign n14387 = n14386 ^ x79;
  assign n14388 = n13958 & n14248;
  assign n14389 = n14388 ^ n13960;
  assign n14390 = n14389 ^ n14386;
  assign n14391 = n14387 & n14390;
  assign n14392 = n14391 ^ x79;
  assign n14393 = n14392 ^ x80;
  assign n14394 = n13964 & n14248;
  assign n14395 = n14394 ^ n13966;
  assign n14396 = n14395 ^ n14392;
  assign n14397 = n14393 & ~n14396;
  assign n14398 = n14397 ^ x80;
  assign n14399 = n14398 ^ x81;
  assign n14400 = n13970 & n14248;
  assign n14401 = n14400 ^ n13972;
  assign n14402 = n14401 ^ n14398;
  assign n14403 = n14399 & n14402;
  assign n14404 = n14403 ^ x81;
  assign n14405 = n14404 ^ x82;
  assign n14406 = n13976 & n14248;
  assign n14407 = n14406 ^ n13978;
  assign n14408 = n14407 ^ n14404;
  assign n14409 = n14405 & ~n14408;
  assign n14410 = n14409 ^ x82;
  assign n14411 = n14410 ^ x83;
  assign n14412 = n13982 & n14248;
  assign n14413 = n14412 ^ n13984;
  assign n14414 = n14413 ^ n14410;
  assign n14415 = n14411 & ~n14414;
  assign n14416 = n14415 ^ x83;
  assign n14417 = n14416 ^ x84;
  assign n14418 = n13988 & n14248;
  assign n14419 = n14418 ^ n13990;
  assign n14420 = n14419 ^ n14416;
  assign n14421 = n14417 & n14420;
  assign n14422 = n14421 ^ x84;
  assign n14423 = n14422 ^ x85;
  assign n14249 = ~n14188 & n14248;
  assign n14250 = n14249 ^ n14190;
  assign n14251 = ~x118 & ~n14250;
  assign n14252 = n14194 & n14248;
  assign n14253 = n14252 ^ n14196;
  assign n14254 = ~x119 & ~n14253;
  assign n14255 = ~n14251 & ~n14254;
  assign n14256 = n14160 & n14248;
  assign n14257 = n14256 ^ n14162;
  assign n14258 = ~x113 & ~n14257;
  assign n14259 = n14166 & n14248;
  assign n14260 = n14259 ^ n14169;
  assign n14261 = ~x114 & ~n14260;
  assign n14262 = ~n14258 & ~n14261;
  assign n14263 = n14104 ^ x102;
  assign n14264 = n14104 ^ n13826;
  assign n14265 = n14263 & ~n14264;
  assign n14266 = n14265 ^ x102;
  assign n14267 = n14266 ^ x103;
  assign n14268 = n14248 & n14267;
  assign n14269 = n14268 ^ n13829;
  assign n14270 = n14269 ^ x104;
  assign n14271 = n14248 & n14263;
  assign n14272 = n14271 ^ n13826;
  assign n14273 = ~x103 & ~n14272;
  assign n14424 = n13994 & n14248;
  assign n14425 = n14424 ^ n13996;
  assign n14426 = n14425 ^ n14422;
  assign n14427 = n14423 & n14426;
  assign n14428 = n14427 ^ x85;
  assign n14429 = n14428 ^ x86;
  assign n14430 = n14000 & n14248;
  assign n14431 = n14430 ^ n14002;
  assign n14432 = n14431 ^ n14428;
  assign n14433 = n14429 & n14432;
  assign n14434 = n14433 ^ x86;
  assign n14435 = n14434 ^ x87;
  assign n14436 = n14006 & n14248;
  assign n14437 = n14436 ^ n14008;
  assign n14438 = n14437 ^ n14434;
  assign n14439 = n14435 & ~n14438;
  assign n14440 = n14439 ^ x87;
  assign n14441 = n14440 ^ x88;
  assign n14442 = n14012 & n14248;
  assign n14443 = n14442 ^ n14014;
  assign n14444 = n14443 ^ n14440;
  assign n14445 = n14441 & n14444;
  assign n14446 = n14445 ^ x88;
  assign n14447 = n14446 ^ x89;
  assign n14448 = n14018 & n14248;
  assign n14449 = n14448 ^ n14020;
  assign n14450 = n14449 ^ n14446;
  assign n14451 = n14447 & ~n14450;
  assign n14452 = n14451 ^ x89;
  assign n14453 = n14452 ^ x90;
  assign n14454 = n14024 & n14248;
  assign n14455 = n14454 ^ n14027;
  assign n14456 = n14455 ^ n14452;
  assign n14457 = n14453 & ~n14456;
  assign n14458 = n14457 ^ x90;
  assign n14459 = n14458 ^ x91;
  assign n14460 = n14031 & n14248;
  assign n14461 = n14460 ^ n14037;
  assign n14462 = n14461 ^ n14458;
  assign n14463 = n14459 & n14462;
  assign n14464 = n14463 ^ x91;
  assign n14465 = n14464 ^ x92;
  assign n14466 = n14041 & n14248;
  assign n14467 = n14466 ^ n14043;
  assign n14468 = n14467 ^ n14464;
  assign n14469 = n14465 & n14468;
  assign n14470 = n14469 ^ x92;
  assign n14471 = n14470 ^ x93;
  assign n14472 = n14047 & n14248;
  assign n14473 = n14472 ^ n14049;
  assign n14474 = n14473 ^ n14470;
  assign n14475 = n14471 & ~n14474;
  assign n14476 = n14475 ^ x93;
  assign n14477 = n14476 ^ x94;
  assign n14478 = n14052 ^ x93;
  assign n14479 = n14248 & n14478;
  assign n14480 = n14479 ^ n13843;
  assign n14481 = n14480 ^ n14476;
  assign n14482 = n14477 & n14481;
  assign n14483 = n14482 ^ x94;
  assign n14484 = n14483 ^ x95;
  assign n14485 = ~n14053 & ~n14056;
  assign n14486 = n14485 ^ x94;
  assign n14487 = n14248 & n14486;
  assign n14488 = n14487 ^ n13840;
  assign n14489 = n14488 ^ n14483;
  assign n14490 = n14484 & n14489;
  assign n14491 = n14490 ^ x95;
  assign n14492 = n14491 ^ x96;
  assign n14493 = n14063 & n14248;
  assign n14494 = n14493 ^ n14065;
  assign n14495 = n14494 ^ n14491;
  assign n14496 = n14492 & ~n14495;
  assign n14497 = n14496 ^ x96;
  assign n14498 = n14497 ^ x97;
  assign n14499 = n14069 & n14248;
  assign n14500 = n14499 ^ n14072;
  assign n14501 = n14500 ^ n14497;
  assign n14502 = n14498 & n14501;
  assign n14503 = n14502 ^ x97;
  assign n14504 = n14503 ^ x98;
  assign n14505 = n14076 & n14248;
  assign n14506 = n14505 ^ n14082;
  assign n14507 = n14506 ^ n14503;
  assign n14508 = n14504 & n14507;
  assign n14509 = n14508 ^ x98;
  assign n14510 = n14509 ^ x99;
  assign n14511 = n14086 & n14248;
  assign n14512 = n14511 ^ n14088;
  assign n14513 = n14512 ^ n14509;
  assign n14514 = n14510 & n14513;
  assign n14515 = n14514 ^ x99;
  assign n14516 = n14515 ^ x100;
  assign n14517 = n14091 ^ x99;
  assign n14518 = n14248 & n14517;
  assign n14519 = n14518 ^ n13833;
  assign n14520 = n14519 ^ n14515;
  assign n14521 = n14516 & ~n14520;
  assign n14522 = n14521 ^ x100;
  assign n14523 = n14522 ^ x101;
  assign n14524 = n14091 ^ n13833;
  assign n14525 = n14517 & ~n14524;
  assign n14526 = n14525 ^ x99;
  assign n14527 = n14526 ^ x100;
  assign n14528 = n14248 & n14527;
  assign n14529 = n14528 ^ n13836;
  assign n14530 = n14529 ^ n14522;
  assign n14531 = n14523 & n14530;
  assign n14532 = n14531 ^ x101;
  assign n14533 = n14532 ^ x102;
  assign n14534 = ~n14099 & n14248;
  assign n14535 = n14534 ^ n14101;
  assign n14536 = n14535 ^ n14532;
  assign n14537 = n14533 & ~n14536;
  assign n14538 = n14537 ^ x102;
  assign n14539 = ~n14273 & n14538;
  assign n14540 = n14539 ^ n14269;
  assign n14541 = n14540 ^ n14269;
  assign n14542 = x103 & n14272;
  assign n14543 = n14542 ^ n14269;
  assign n14544 = n14543 ^ n14269;
  assign n14545 = ~n14541 & ~n14544;
  assign n14546 = n14545 ^ n14269;
  assign n14547 = n14270 & n14546;
  assign n14548 = n14547 ^ x104;
  assign n14549 = n14548 ^ x105;
  assign n14550 = ~n14112 & n14248;
  assign n14551 = n14550 ^ n14114;
  assign n14552 = n14551 ^ n14548;
  assign n14553 = n14549 & ~n14552;
  assign n14554 = n14553 ^ x105;
  assign n14555 = n14554 ^ x106;
  assign n14556 = n14118 & n14248;
  assign n14557 = n14556 ^ n14120;
  assign n14558 = n14557 ^ n14554;
  assign n14559 = n14555 & ~n14558;
  assign n14560 = n14559 ^ x106;
  assign n14561 = n14560 ^ x107;
  assign n14562 = n14124 & n14248;
  assign n14563 = n14562 ^ n14126;
  assign n14564 = n14563 ^ n14560;
  assign n14565 = n14561 & ~n14564;
  assign n14566 = n14565 ^ x107;
  assign n14567 = n14566 ^ x108;
  assign n14568 = n14130 & n14248;
  assign n14569 = n14568 ^ n14132;
  assign n14570 = n14569 ^ n14566;
  assign n14571 = n14567 & ~n14570;
  assign n14572 = n14571 ^ x108;
  assign n14573 = n14572 ^ x109;
  assign n14574 = n14136 & n14248;
  assign n14575 = n14574 ^ n14138;
  assign n14576 = n14575 ^ n14572;
  assign n14577 = n14573 & ~n14576;
  assign n14578 = n14577 ^ x109;
  assign n14579 = n14578 ^ x110;
  assign n14580 = n14142 & n14248;
  assign n14581 = n14580 ^ n14144;
  assign n14582 = n14581 ^ n14578;
  assign n14583 = n14579 & n14582;
  assign n14584 = n14583 ^ x110;
  assign n14585 = n14584 ^ x111;
  assign n14586 = n14148 & n14248;
  assign n14587 = n14586 ^ n14150;
  assign n14588 = n14587 ^ n14584;
  assign n14589 = n14585 & ~n14588;
  assign n14590 = n14589 ^ x111;
  assign n14591 = n14590 ^ x112;
  assign n14592 = n14154 & n14248;
  assign n14593 = n14592 ^ n14156;
  assign n14594 = n14593 ^ n14590;
  assign n14595 = n14591 & n14594;
  assign n14596 = n14595 ^ x112;
  assign n14597 = n14262 & n14596;
  assign n14598 = n14260 ^ x114;
  assign n14599 = x113 & n14257;
  assign n14600 = n14599 ^ n14260;
  assign n14601 = n14598 & ~n14600;
  assign n14602 = n14601 ^ x114;
  assign n14603 = ~n14597 & ~n14602;
  assign n14604 = n14603 ^ x115;
  assign n14605 = n14173 & n14248;
  assign n14606 = n14605 ^ n14177;
  assign n14607 = n14606 ^ n14603;
  assign n14608 = ~n14604 & ~n14607;
  assign n14609 = n14608 ^ x115;
  assign n14610 = n14609 ^ x116;
  assign n14611 = n14180 ^ x115;
  assign n14612 = n14248 & n14611;
  assign n14613 = n14612 ^ n13819;
  assign n14614 = n14613 ^ n14609;
  assign n14615 = n14610 & n14614;
  assign n14616 = n14615 ^ x116;
  assign n14617 = n14616 ^ x117;
  assign n14618 = n14180 ^ n13819;
  assign n14619 = n14611 & n14618;
  assign n14620 = n14619 ^ x115;
  assign n14621 = n14620 ^ x116;
  assign n14622 = n14248 & n14621;
  assign n14623 = n14622 ^ n13822;
  assign n14624 = n14623 ^ n14616;
  assign n14625 = n14617 & n14624;
  assign n14626 = n14625 ^ x117;
  assign n14627 = n14255 & n14626;
  assign n14628 = n14253 ^ x119;
  assign n14629 = x118 & n14250;
  assign n14630 = n14629 ^ n14253;
  assign n14631 = n14628 & ~n14630;
  assign n14632 = n14631 ^ x119;
  assign n14633 = ~n14627 & ~n14632;
  assign n14634 = n14633 ^ x120;
  assign n14635 = n14200 & n14248;
  assign n14636 = n14635 ^ n14202;
  assign n14637 = n14636 ^ n14633;
  assign n14638 = ~n14634 & n14637;
  assign n14639 = n14638 ^ x120;
  assign n14640 = n14639 ^ x121;
  assign n14641 = n14206 & n14248;
  assign n14642 = n14641 ^ n14208;
  assign n14643 = n14642 ^ n14639;
  assign n14644 = n14640 & ~n14643;
  assign n14645 = n14644 ^ x121;
  assign n14646 = n14645 ^ x122;
  assign n14647 = n14212 & n14248;
  assign n14648 = n14647 ^ n14214;
  assign n14649 = n14648 ^ n14645;
  assign n14650 = n14646 & ~n14649;
  assign n14651 = n14650 ^ x122;
  assign n14652 = n14651 ^ x123;
  assign n14653 = n14218 & n14248;
  assign n14654 = n14653 ^ n14220;
  assign n14655 = n14654 ^ n14651;
  assign n14656 = n14652 & n14655;
  assign n14657 = n14656 ^ x123;
  assign n14658 = n14657 ^ x124;
  assign n14659 = n14224 & n14248;
  assign n14660 = n14659 ^ n14226;
  assign n14661 = n14660 ^ n14657;
  assign n14662 = n14658 & ~n14661;
  assign n14663 = n14662 ^ x124;
  assign n14664 = n14663 ^ x125;
  assign n14665 = n14230 & n14248;
  assign n14666 = n14665 ^ n14232;
  assign n14667 = n14666 ^ n14663;
  assign n14668 = n14664 & n14667;
  assign n14669 = n14668 ^ x125;
  assign n14670 = n14669 ^ x126;
  assign n14671 = n14236 & n14242;
  assign n14672 = n129 & n14671;
  assign n14673 = n14672 ^ n14242;
  assign n14674 = n14673 ^ n14669;
  assign n14675 = n14670 & n14674;
  assign n14676 = n14675 ^ x126;
  assign n14677 = ~x127 & ~n14676;
  assign n14678 = n14423 & n14677;
  assign n14679 = n14678 ^ n14425;
  assign n14680 = ~x86 & n14679;
  assign n14681 = n14429 & n14677;
  assign n14682 = n14681 ^ n14431;
  assign n14683 = ~x87 & n14682;
  assign n14684 = ~n14680 & ~n14683;
  assign n14685 = n14363 & n14677;
  assign n14686 = n14685 ^ n14365;
  assign n14687 = ~x76 & ~n14686;
  assign n14688 = n14369 & n14677;
  assign n14689 = n14688 ^ n14371;
  assign n14690 = ~x77 & n14689;
  assign n14691 = ~n14687 & ~n14690;
  assign n14692 = n14336 & n14677;
  assign n14693 = n14692 ^ n14339;
  assign n14694 = n14693 ^ x72;
  assign n14695 = ~n14330 & n14677;
  assign n14696 = n14695 ^ n14332;
  assign n14697 = x71 & n14696;
  assign n14698 = x64 & n14677;
  assign n14699 = x0 & ~x65;
  assign n14700 = x1 & ~n14699;
  assign n14701 = n14698 & n14700;
  assign n14703 = x65 ^ x1;
  assign n14710 = n14703 ^ x65;
  assign n14702 = x65 ^ x0;
  assign n14704 = n14703 ^ n14702;
  assign n14705 = n14704 ^ x65;
  assign n14706 = n14702 ^ x64;
  assign n14707 = n14706 ^ n14702;
  assign n14708 = n14707 ^ n14705;
  assign n14709 = ~n14705 & ~n14708;
  assign n14711 = n14710 ^ n14709;
  assign n14712 = n14711 ^ n14705;
  assign n14713 = n14677 ^ x65;
  assign n14714 = n14713 ^ x65;
  assign n14715 = n14709 ^ n14705;
  assign n14716 = ~n14714 & ~n14715;
  assign n14717 = n14716 ^ x65;
  assign n14718 = ~n14712 & n14717;
  assign n14719 = n14718 ^ x65;
  assign n14720 = n14719 ^ x65;
  assign n14721 = n14720 ^ x65;
  assign n14722 = ~n14701 & ~n14721;
  assign n14723 = n14722 ^ x66;
  assign n14724 = x65 & ~x127;
  assign n14725 = n14724 ^ n288;
  assign n14726 = n14725 ^ n288;
  assign n14727 = n14676 ^ n288;
  assign n14728 = n14727 ^ n288;
  assign n14729 = n14726 & ~n14728;
  assign n14730 = n14729 ^ n288;
  assign n14731 = ~n14248 & n14730;
  assign n14732 = n14731 ^ n288;
  assign n14733 = x1 & n14732;
  assign n14734 = n289 & ~n14248;
  assign n14735 = n14734 ^ x65;
  assign n14736 = ~x1 & n14735;
  assign n14737 = ~n202 & ~n14736;
  assign n14738 = n14737 ^ n14281;
  assign n14739 = n14677 & ~n14738;
  assign n14740 = n14739 ^ n14281;
  assign n14741 = ~n14733 & ~n14740;
  assign n14742 = n14741 ^ x2;
  assign n14743 = n14742 ^ n14722;
  assign n14744 = ~n14723 & n14743;
  assign n14745 = n14744 ^ x66;
  assign n14746 = n14745 ^ x67;
  assign n14747 = ~n14294 & n14677;
  assign n14748 = n14747 ^ n14306;
  assign n14749 = n14748 ^ n14745;
  assign n14750 = n14746 & ~n14749;
  assign n14751 = n14750 ^ x67;
  assign n14752 = n14751 ^ x68;
  assign n14753 = n14310 & n14677;
  assign n14754 = n14753 ^ n14319;
  assign n14755 = n14754 ^ n14751;
  assign n14756 = n14752 & n14755;
  assign n14757 = n14756 ^ x68;
  assign n14758 = n14757 ^ x69;
  assign n14759 = n14322 ^ x68;
  assign n14760 = n14677 & n14759;
  assign n14761 = n14760 ^ n14278;
  assign n14762 = n14761 ^ n14757;
  assign n14763 = n14758 & ~n14762;
  assign n14764 = n14763 ^ x69;
  assign n14765 = n14764 ^ x70;
  assign n14766 = n14322 ^ n14278;
  assign n14767 = n14759 & ~n14766;
  assign n14768 = n14767 ^ x68;
  assign n14769 = n14768 ^ x69;
  assign n14770 = n14677 & n14769;
  assign n14771 = n14770 ^ n14275;
  assign n14772 = n14771 ^ n14764;
  assign n14773 = n14765 & ~n14772;
  assign n14774 = n14773 ^ x70;
  assign n14775 = ~n14697 & ~n14774;
  assign n14776 = n14775 ^ n14693;
  assign n14777 = n14776 ^ n14693;
  assign n14778 = ~x71 & ~n14696;
  assign n14779 = n14778 ^ n14693;
  assign n14780 = n14779 ^ n14693;
  assign n14781 = ~n14777 & ~n14780;
  assign n14782 = n14781 ^ n14693;
  assign n14783 = ~n14694 & n14782;
  assign n14784 = n14783 ^ x72;
  assign n14785 = n14784 ^ x73;
  assign n14786 = n14343 & n14677;
  assign n14787 = n14786 ^ n14347;
  assign n14788 = n14787 ^ n14784;
  assign n14789 = n14785 & n14788;
  assign n14790 = n14789 ^ x73;
  assign n14791 = n14790 ^ x74;
  assign n14792 = n14351 & n14677;
  assign n14793 = n14792 ^ n14353;
  assign n14794 = n14793 ^ n14790;
  assign n14795 = n14791 & n14794;
  assign n14796 = n14795 ^ x74;
  assign n14797 = n14796 ^ x75;
  assign n14798 = n14357 & n14677;
  assign n14799 = n14798 ^ n14359;
  assign n14800 = n14799 ^ n14796;
  assign n14801 = n14797 & n14800;
  assign n14802 = n14801 ^ x75;
  assign n14803 = n14691 & n14802;
  assign n14804 = n14689 ^ x77;
  assign n14805 = x76 & n14686;
  assign n14806 = n14805 ^ n14689;
  assign n14807 = ~n14804 & n14806;
  assign n14808 = n14807 ^ x77;
  assign n14809 = ~n14803 & ~n14808;
  assign n14810 = n14809 ^ x78;
  assign n14811 = n14375 & n14677;
  assign n14812 = n14811 ^ n14377;
  assign n14813 = n14812 ^ n14809;
  assign n14814 = ~n14810 & n14813;
  assign n14815 = n14814 ^ x78;
  assign n14816 = n14815 ^ x79;
  assign n14817 = n14381 & n14677;
  assign n14818 = n14817 ^ n14383;
  assign n14819 = n14818 ^ n14815;
  assign n14820 = n14816 & n14819;
  assign n14821 = n14820 ^ x79;
  assign n14822 = n14821 ^ x80;
  assign n14823 = n14387 & n14677;
  assign n14824 = n14823 ^ n14389;
  assign n14825 = n14824 ^ n14821;
  assign n14826 = n14822 & n14825;
  assign n14827 = n14826 ^ x80;
  assign n14828 = n14827 ^ x81;
  assign n14829 = n14393 & n14677;
  assign n14830 = n14829 ^ n14395;
  assign n14831 = n14830 ^ n14827;
  assign n14832 = n14828 & ~n14831;
  assign n14833 = n14832 ^ x81;
  assign n14834 = n14833 ^ x82;
  assign n14835 = n14399 & n14677;
  assign n14836 = n14835 ^ n14401;
  assign n14837 = n14836 ^ n14833;
  assign n14838 = n14834 & n14837;
  assign n14839 = n14838 ^ x82;
  assign n14840 = n14839 ^ x83;
  assign n14841 = n14405 & n14677;
  assign n14842 = n14841 ^ n14407;
  assign n14843 = n14842 ^ n14839;
  assign n14844 = n14840 & ~n14843;
  assign n14845 = n14844 ^ x83;
  assign n14846 = n14845 ^ x84;
  assign n14847 = n14411 & n14677;
  assign n14848 = n14847 ^ n14413;
  assign n14849 = n14848 ^ n14845;
  assign n14850 = n14846 & ~n14849;
  assign n14851 = n14850 ^ x84;
  assign n14852 = n14851 ^ x85;
  assign n14853 = n14417 & n14677;
  assign n14854 = n14853 ^ n14419;
  assign n14855 = n14854 ^ n14851;
  assign n14856 = n14852 & n14855;
  assign n14857 = n14856 ^ x85;
  assign n14858 = n14684 & n14857;
  assign n14859 = n14682 ^ x87;
  assign n14860 = x86 & ~n14679;
  assign n14861 = n14860 ^ n14682;
  assign n14862 = ~n14859 & n14861;
  assign n14863 = n14862 ^ x87;
  assign n14864 = ~n14858 & ~n14863;
  assign n14865 = n14864 ^ x88;
  assign n14866 = n14435 & n14677;
  assign n14867 = n14866 ^ n14437;
  assign n14868 = n14867 ^ n14864;
  assign n14869 = ~n14865 & n14868;
  assign n14870 = n14869 ^ x88;
  assign n14871 = n14870 ^ x89;
  assign n14872 = n14441 & n14677;
  assign n14873 = n14872 ^ n14443;
  assign n14874 = n14873 ^ n14870;
  assign n14875 = n14871 & n14874;
  assign n14876 = n14875 ^ x89;
  assign n14877 = n14876 ^ x90;
  assign n14878 = n14447 & n14677;
  assign n14879 = n14878 ^ n14449;
  assign n14880 = n14879 ^ n14876;
  assign n14881 = n14877 & ~n14880;
  assign n14882 = n14881 ^ x90;
  assign n14883 = n14882 ^ x91;
  assign n14884 = n14453 & n14677;
  assign n14885 = n14884 ^ n14455;
  assign n14886 = n14885 ^ n14882;
  assign n14887 = n14883 & ~n14886;
  assign n14888 = n14887 ^ x91;
  assign n14889 = n14888 ^ x92;
  assign n14890 = n14459 & n14677;
  assign n14891 = n14890 ^ n14461;
  assign n14892 = n14891 ^ n14888;
  assign n14893 = n14889 & n14892;
  assign n14894 = n14893 ^ x92;
  assign n14895 = n14894 ^ x93;
  assign n14896 = n14465 & n14677;
  assign n14897 = n14896 ^ n14467;
  assign n14898 = n14897 ^ n14894;
  assign n14899 = n14895 & n14898;
  assign n14900 = n14899 ^ x93;
  assign n14901 = n14900 ^ x94;
  assign n14902 = n14471 & n14677;
  assign n14903 = n14902 ^ n14473;
  assign n14904 = n14903 ^ n14900;
  assign n14905 = n14901 & ~n14904;
  assign n14906 = n14905 ^ x94;
  assign n14907 = n14906 ^ x95;
  assign n14908 = n14477 & n14677;
  assign n14909 = n14908 ^ n14480;
  assign n14910 = n14909 ^ n14906;
  assign n14911 = n14907 & n14910;
  assign n14912 = n14911 ^ x95;
  assign n14913 = n14912 ^ x96;
  assign n14914 = n14484 & n14677;
  assign n14915 = n14914 ^ n14488;
  assign n14916 = n14915 ^ n14912;
  assign n14917 = n14913 & n14916;
  assign n14918 = n14917 ^ x96;
  assign n14919 = n14918 ^ x97;
  assign n14920 = n14492 & n14677;
  assign n14921 = n14920 ^ n14494;
  assign n14922 = n14921 ^ n14918;
  assign n14923 = n14919 & ~n14922;
  assign n14924 = n14923 ^ x97;
  assign n14925 = n14924 ^ x98;
  assign n14926 = n14498 & n14677;
  assign n14927 = n14926 ^ n14500;
  assign n14928 = n14927 ^ n14924;
  assign n14929 = n14925 & n14928;
  assign n14930 = n14929 ^ x98;
  assign n14931 = n14930 ^ x99;
  assign n14932 = n14504 & n14677;
  assign n14933 = n14932 ^ n14506;
  assign n14934 = n14933 ^ n14930;
  assign n14935 = n14931 & n14934;
  assign n14936 = n14935 ^ x99;
  assign n14937 = n14936 ^ x100;
  assign n14938 = n14510 & n14677;
  assign n14939 = n14938 ^ n14512;
  assign n14940 = n14939 ^ n14936;
  assign n14941 = n14937 & n14940;
  assign n14942 = n14941 ^ x100;
  assign n14943 = n14942 ^ x101;
  assign n14944 = n14516 & n14677;
  assign n14945 = n14944 ^ n14519;
  assign n14946 = n14945 ^ n14942;
  assign n14947 = n14943 & ~n14946;
  assign n14948 = n14947 ^ x101;
  assign n14949 = n14948 ^ x102;
  assign n14950 = n14523 & n14677;
  assign n14951 = n14950 ^ n14529;
  assign n14952 = n14951 ^ n14948;
  assign n14953 = n14949 & n14952;
  assign n14954 = n14953 ^ x102;
  assign n14955 = n14954 ^ x103;
  assign n14956 = n14533 & n14677;
  assign n14957 = n14956 ^ n14535;
  assign n14958 = n14957 ^ n14954;
  assign n14959 = n14955 & ~n14958;
  assign n14960 = n14959 ^ x103;
  assign n14961 = n14960 ^ x104;
  assign n14962 = n14538 ^ x103;
  assign n14963 = n14677 & n14962;
  assign n14964 = n14963 ^ n14272;
  assign n14965 = n14964 ^ n14960;
  assign n14966 = n14961 & ~n14965;
  assign n14967 = n14966 ^ x104;
  assign n14968 = n14967 ^ x105;
  assign n14969 = ~n14539 & ~n14542;
  assign n14970 = n14969 ^ x104;
  assign n14971 = n14677 & ~n14970;
  assign n14972 = n14971 ^ n14269;
  assign n14973 = n14972 ^ n14967;
  assign n14974 = n14968 & ~n14973;
  assign n14975 = n14974 ^ x105;
  assign n14976 = n14975 ^ x106;
  assign n14977 = n14549 & n14677;
  assign n14978 = n14977 ^ n14551;
  assign n14979 = n14978 ^ n14975;
  assign n14980 = n14976 & ~n14979;
  assign n14981 = n14980 ^ x106;
  assign n14982 = n14981 ^ x107;
  assign n14983 = n14555 & n14677;
  assign n14984 = n14983 ^ n14557;
  assign n14985 = n14984 ^ n14981;
  assign n14986 = n14982 & ~n14985;
  assign n14987 = n14986 ^ x107;
  assign n14988 = n14987 ^ x108;
  assign n14989 = n14561 & n14677;
  assign n14990 = n14989 ^ n14563;
  assign n14991 = n14990 ^ n14987;
  assign n14992 = n14988 & ~n14991;
  assign n14993 = n14992 ^ x108;
  assign n14994 = n14993 ^ x109;
  assign n14995 = n14567 & n14677;
  assign n14996 = n14995 ^ n14569;
  assign n14997 = n14996 ^ n14993;
  assign n14998 = n14994 & ~n14997;
  assign n14999 = n14998 ^ x109;
  assign n15000 = n14999 ^ x110;
  assign n15001 = n14573 & n14677;
  assign n15002 = n15001 ^ n14575;
  assign n15003 = n15002 ^ n14999;
  assign n15004 = n15000 & ~n15003;
  assign n15005 = n15004 ^ x110;
  assign n15006 = n15005 ^ x111;
  assign n15007 = n14579 & n14677;
  assign n15008 = n15007 ^ n14581;
  assign n15009 = n15008 ^ n15005;
  assign n15010 = n15006 & n15009;
  assign n15011 = n15010 ^ x111;
  assign n15012 = n15011 ^ x112;
  assign n15013 = n14585 & n14677;
  assign n15014 = n15013 ^ n14587;
  assign n15015 = n15014 ^ n15011;
  assign n15016 = n15012 & ~n15015;
  assign n15017 = n15016 ^ x112;
  assign n15018 = n15017 ^ x113;
  assign n15019 = n14591 & n14677;
  assign n15020 = n15019 ^ n14593;
  assign n15021 = n15020 ^ n15017;
  assign n15022 = n15018 & n15021;
  assign n15023 = n15022 ^ x113;
  assign n15024 = n15023 ^ x114;
  assign n15025 = n14596 ^ x113;
  assign n15026 = n14677 & n15025;
  assign n15027 = n15026 ^ n14257;
  assign n15028 = n15027 ^ n15023;
  assign n15029 = n15024 & ~n15028;
  assign n15030 = n15029 ^ x114;
  assign n15031 = n15030 ^ x115;
  assign n15032 = n14596 ^ n14257;
  assign n15033 = n15025 & ~n15032;
  assign n15034 = n15033 ^ x113;
  assign n15035 = n15034 ^ x114;
  assign n15036 = n14677 & n15035;
  assign n15037 = n15036 ^ n14260;
  assign n15038 = n15037 ^ n15030;
  assign n15039 = n15031 & ~n15038;
  assign n15040 = n15039 ^ x115;
  assign n15041 = n15040 ^ x116;
  assign n15042 = ~n14604 & n14677;
  assign n15043 = n15042 ^ n14606;
  assign n15044 = n15043 ^ n15040;
  assign n15045 = n15041 & n15044;
  assign n15046 = n15045 ^ x116;
  assign n15047 = n15046 ^ x117;
  assign n15048 = n14610 & n14677;
  assign n15049 = n15048 ^ n14613;
  assign n15050 = n15049 ^ n15046;
  assign n15051 = n15047 & n15050;
  assign n15052 = n15051 ^ x117;
  assign n15053 = n15052 ^ x118;
  assign n15054 = n14617 & n14677;
  assign n15055 = n15054 ^ n14623;
  assign n15056 = n15055 ^ n15052;
  assign n15057 = n15053 & n15056;
  assign n15058 = n15057 ^ x118;
  assign n15059 = n15058 ^ x119;
  assign n15060 = n14626 ^ x118;
  assign n15061 = n14677 & n15060;
  assign n15062 = n15061 ^ n14250;
  assign n15063 = n15062 ^ n15058;
  assign n15064 = n15059 & ~n15063;
  assign n15065 = n15064 ^ x119;
  assign n15066 = n15065 ^ x120;
  assign n15067 = n14626 ^ n14250;
  assign n15068 = n15060 & ~n15067;
  assign n15069 = n15068 ^ x118;
  assign n15070 = n15069 ^ x119;
  assign n15071 = n14677 & n15070;
  assign n15072 = n15071 ^ n14253;
  assign n15073 = n15072 ^ n15065;
  assign n15074 = n15066 & ~n15073;
  assign n15075 = n15074 ^ x120;
  assign n15076 = n15075 ^ x121;
  assign n15077 = ~n14634 & n14677;
  assign n15078 = n15077 ^ n14636;
  assign n15079 = n15078 ^ n15075;
  assign n15080 = n15076 & ~n15079;
  assign n15081 = n15080 ^ x121;
  assign n15082 = n15081 ^ x122;
  assign n15083 = n14640 & n14677;
  assign n15084 = n15083 ^ n14642;
  assign n15085 = n15084 ^ n15081;
  assign n15086 = n15082 & ~n15085;
  assign n15087 = n15086 ^ x122;
  assign n15088 = n15087 ^ x123;
  assign n15089 = n14646 & n14677;
  assign n15090 = n15089 ^ n14648;
  assign n15091 = n15090 ^ n15087;
  assign n15092 = n15088 & ~n15091;
  assign n15093 = n15092 ^ x123;
  assign n15094 = n15093 ^ x124;
  assign n15095 = n14652 & n14677;
  assign n15096 = n15095 ^ n14654;
  assign n15097 = n15096 ^ n15093;
  assign n15098 = n15094 & n15097;
  assign n15099 = n15098 ^ x124;
  assign n15100 = n15099 ^ x125;
  assign n15101 = n14658 & n14677;
  assign n15102 = n15101 ^ n14660;
  assign n15103 = n15102 ^ n15099;
  assign n15104 = n15100 & ~n15103;
  assign n15105 = n15104 ^ x125;
  assign n15106 = n15105 ^ x126;
  assign n15107 = n14664 & n14677;
  assign n15108 = n15107 ^ n14666;
  assign n15109 = n15108 ^ n15105;
  assign n15110 = n15106 & n15109;
  assign n15111 = n15110 ^ x126;
  assign n15112 = ~n12948 & ~n15111;
  assign n15113 = ~x127 & ~n14670;
  assign n15114 = n14673 & n15113;
  assign n15115 = ~n15112 & ~n15114;
  assign n15116 = ~x62 & n227;
  assign n15117 = n15116 ^ n192;
  assign n15118 = ~x63 & x64;
  assign n15119 = ~x65 & ~x66;
  assign n15120 = ~n15118 & n15119;
  assign n15121 = n189 & n15120;
  assign n15122 = x64 & ~n15115;
  assign n15123 = n15122 ^ x0;
  assign n15124 = ~x0 & x64;
  assign n15125 = n15124 ^ n14677;
  assign n15126 = x65 ^ x64;
  assign n15127 = n15126 ^ x64;
  assign n15128 = n15124 ^ x64;
  assign n15129 = ~n15127 & n15128;
  assign n15130 = n15129 ^ x64;
  assign n15131 = n15125 & n15130;
  assign n15132 = n15131 ^ x65;
  assign n15133 = n15132 ^ n14698;
  assign n15134 = n15132 ^ n14699;
  assign n15135 = n15132 ^ n15115;
  assign n15136 = ~n15132 & n15135;
  assign n15137 = n15136 ^ n15132;
  assign n15138 = ~n15134 & ~n15137;
  assign n15139 = n15138 ^ n15136;
  assign n15140 = n15139 ^ n15132;
  assign n15141 = n15140 ^ n15115;
  assign n15142 = n15133 & n15141;
  assign n15143 = n15142 ^ n14698;
  assign n15144 = n15143 ^ x1;
  assign n15145 = ~n14723 & ~n15115;
  assign n15146 = n15145 ^ n14742;
  assign n15147 = n14746 & ~n15115;
  assign n15148 = n15147 ^ n14748;
  assign n15149 = n14752 & ~n15115;
  assign n15150 = n15149 ^ n14754;
  assign n15151 = n14758 & ~n15115;
  assign n15152 = n15151 ^ n14761;
  assign n15153 = n14765 & ~n15115;
  assign n15154 = n15153 ^ n14771;
  assign n15155 = n14774 ^ x71;
  assign n15156 = ~n15115 & n15155;
  assign n15157 = n15156 ^ n14696;
  assign n15158 = ~n14775 & ~n14778;
  assign n15159 = n15158 ^ x72;
  assign n15160 = ~n15115 & n15159;
  assign n15161 = n15160 ^ n14693;
  assign n15162 = n14785 & ~n15115;
  assign n15163 = n15162 ^ n14787;
  assign n15164 = n14791 & ~n15115;
  assign n15165 = n15164 ^ n14793;
  assign n15166 = n14797 & ~n15115;
  assign n15167 = n15166 ^ n14799;
  assign n15168 = n14802 ^ x76;
  assign n15169 = ~n15115 & n15168;
  assign n15170 = n15169 ^ n14686;
  assign n15171 = n14802 ^ n14686;
  assign n15172 = n15168 & ~n15171;
  assign n15173 = n15172 ^ x76;
  assign n15174 = n15173 ^ x77;
  assign n15175 = ~n15115 & n15174;
  assign n15176 = n15175 ^ n14689;
  assign n15177 = ~n14810 & ~n15115;
  assign n15178 = n15177 ^ n14812;
  assign n15179 = n14816 & ~n15115;
  assign n15180 = n15179 ^ n14818;
  assign n15181 = n14822 & ~n15115;
  assign n15182 = n15181 ^ n14824;
  assign n15183 = n14828 & ~n15115;
  assign n15184 = n15183 ^ n14830;
  assign n15185 = n14834 & ~n15115;
  assign n15186 = n15185 ^ n14836;
  assign n15187 = n14840 & ~n15115;
  assign n15188 = n15187 ^ n14842;
  assign n15189 = n14846 & ~n15115;
  assign n15190 = n15189 ^ n14848;
  assign n15191 = n14852 & ~n15115;
  assign n15192 = n15191 ^ n14854;
  assign n15193 = n14857 ^ x86;
  assign n15194 = ~n15115 & n15193;
  assign n15195 = n15194 ^ n14679;
  assign n15196 = n14857 ^ n14679;
  assign n15197 = n15193 & n15196;
  assign n15198 = n15197 ^ x86;
  assign n15199 = n15198 ^ x87;
  assign n15200 = ~n15115 & n15199;
  assign n15201 = n15200 ^ n14682;
  assign n15202 = ~n14865 & ~n15115;
  assign n15203 = n15202 ^ n14867;
  assign n15204 = n14871 & ~n15115;
  assign n15205 = n15204 ^ n14873;
  assign n15206 = n14877 & ~n15115;
  assign n15207 = n15206 ^ n14879;
  assign n15208 = n14883 & ~n15115;
  assign n15209 = n15208 ^ n14885;
  assign n15210 = n14889 & ~n15115;
  assign n15211 = n15210 ^ n14891;
  assign n15212 = n14895 & ~n15115;
  assign n15213 = n15212 ^ n14897;
  assign n15214 = n14901 & ~n15115;
  assign n15215 = n15214 ^ n14903;
  assign n15216 = n14907 & ~n15115;
  assign n15217 = n15216 ^ n14909;
  assign n15218 = n14913 & ~n15115;
  assign n15219 = n15218 ^ n14915;
  assign n15220 = n14919 & ~n15115;
  assign n15221 = n15220 ^ n14921;
  assign n15222 = n14925 & ~n15115;
  assign n15223 = n15222 ^ n14927;
  assign n15224 = n14931 & ~n15115;
  assign n15225 = n15224 ^ n14933;
  assign n15226 = n14937 & ~n15115;
  assign n15227 = n15226 ^ n14939;
  assign n15228 = n14943 & ~n15115;
  assign n15229 = n15228 ^ n14945;
  assign n15230 = n14949 & ~n15115;
  assign n15231 = n15230 ^ n14951;
  assign n15232 = n14955 & ~n15115;
  assign n15233 = n15232 ^ n14957;
  assign n15234 = n14961 & ~n15115;
  assign n15235 = n15234 ^ n14964;
  assign n15236 = n14968 & ~n15115;
  assign n15237 = n15236 ^ n14972;
  assign n15238 = n14976 & ~n15115;
  assign n15239 = n15238 ^ n14978;
  assign n15240 = n14982 & ~n15115;
  assign n15241 = n15240 ^ n14984;
  assign n15242 = n14988 & ~n15115;
  assign n15243 = n15242 ^ n14990;
  assign n15244 = n14994 & ~n15115;
  assign n15245 = n15244 ^ n14996;
  assign n15246 = n15000 & ~n15115;
  assign n15247 = n15246 ^ n15002;
  assign n15248 = n15006 & ~n15115;
  assign n15249 = n15248 ^ n15008;
  assign n15250 = n15012 & ~n15115;
  assign n15251 = n15250 ^ n15014;
  assign n15252 = n15018 & ~n15115;
  assign n15253 = n15252 ^ n15020;
  assign n15254 = n15024 & ~n15115;
  assign n15255 = n15254 ^ n15027;
  assign n15256 = n15031 & ~n15115;
  assign n15257 = n15256 ^ n15037;
  assign n15258 = n15041 & ~n15115;
  assign n15259 = n15258 ^ n15043;
  assign n15260 = n15047 & ~n15115;
  assign n15261 = n15260 ^ n15049;
  assign n15262 = n15053 & ~n15115;
  assign n15263 = n15262 ^ n15055;
  assign n15264 = n15059 & ~n15115;
  assign n15265 = n15264 ^ n15062;
  assign n15266 = n15066 & ~n15115;
  assign n15267 = n15266 ^ n15072;
  assign n15268 = n15076 & ~n15115;
  assign n15269 = n15268 ^ n15078;
  assign n15270 = n15082 & ~n15115;
  assign n15271 = n15270 ^ n15084;
  assign n15272 = n15088 & ~n15115;
  assign n15273 = n15272 ^ n15090;
  assign n15274 = n15094 & ~n15115;
  assign n15275 = n15274 ^ n15096;
  assign n15276 = n15100 & ~n15115;
  assign n15277 = n15276 ^ n15102;
  assign n15278 = n15106 & ~n15115;
  assign n15279 = n15278 ^ n15108;
  assign n15280 = n15111 ^ x127;
  assign n15281 = n15280 ^ x127;
  assign n15282 = n15113 ^ x127;
  assign n15283 = ~n15281 & n15282;
  assign n15284 = n15283 ^ x127;
  assign n15285 = n14673 & n15284;
  assign y0 = ~n15115;
  assign y1 = n14677;
  assign y2 = n14248;
  assign y3 = n13817;
  assign y4 = n13385;
  assign y5 = ~n12955;
  assign y6 = n12520;
  assign y7 = n12114;
  assign y8 = ~n11720;
  assign y9 = n11324;
  assign y10 = n10928;
  assign y11 = n10558;
  assign y12 = n10165;
  assign y13 = n9808;
  assign y14 = n9446;
  assign y15 = ~n9100;
  assign y16 = n8746;
  assign y17 = n8415;
  assign y18 = n8093;
  assign y19 = ~n7781;
  assign y20 = n7460;
  assign y21 = n7137;
  assign y22 = n6817;
  assign y23 = n6515;
  assign y24 = n6206;
  assign y25 = n5931;
  assign y26 = n5651;
  assign y27 = ~n5365;
  assign y28 = n5087;
  assign y29 = n4842;
  assign y30 = n4609;
  assign y31 = n4386;
  assign y32 = ~n4138;
  assign y33 = n3912;
  assign y34 = n3691;
  assign y35 = n3471;
  assign y36 = n3257;
  assign y37 = n3041;
  assign y38 = n2852;
  assign y39 = n2668;
  assign y40 = n2492;
  assign y41 = ~n2309;
  assign y42 = n2148;
  assign y43 = n1973;
  assign y44 = n1816;
  assign y45 = n1669;
  assign y46 = ~n1529;
  assign y47 = n1393;
  assign y48 = n1247;
  assign y49 = ~n1140;
  assign y50 = n1029;
  assign y51 = n921;
  assign y52 = n821;
  assign y53 = ~n728;
  assign y54 = n642;
  assign y55 = ~n562;
  assign y56 = n485;
  assign y57 = n414;
  assign y58 = n348;
  assign y59 = n302;
  assign y60 = ~n250;
  assign y61 = n215;
  assign y62 = n15117;
  assign y63 = n15121;
  assign y64 = n15123;
  assign y65 = n15144;
  assign y66 = ~n15146;
  assign y67 = ~n15148;
  assign y68 = n15150;
  assign y69 = ~n15152;
  assign y70 = ~n15154;
  assign y71 = ~n15157;
  assign y72 = n15161;
  assign y73 = n15163;
  assign y74 = n15165;
  assign y75 = n15167;
  assign y76 = ~n15170;
  assign y77 = n15176;
  assign y78 = ~n15178;
  assign y79 = n15180;
  assign y80 = n15182;
  assign y81 = ~n15184;
  assign y82 = n15186;
  assign y83 = ~n15188;
  assign y84 = ~n15190;
  assign y85 = n15192;
  assign y86 = n15195;
  assign y87 = n15201;
  assign y88 = ~n15203;
  assign y89 = n15205;
  assign y90 = ~n15207;
  assign y91 = ~n15209;
  assign y92 = n15211;
  assign y93 = n15213;
  assign y94 = ~n15215;
  assign y95 = n15217;
  assign y96 = n15219;
  assign y97 = ~n15221;
  assign y98 = n15223;
  assign y99 = n15225;
  assign y100 = n15227;
  assign y101 = ~n15229;
  assign y102 = n15231;
  assign y103 = ~n15233;
  assign y104 = ~n15235;
  assign y105 = ~n15237;
  assign y106 = ~n15239;
  assign y107 = ~n15241;
  assign y108 = ~n15243;
  assign y109 = ~n15245;
  assign y110 = ~n15247;
  assign y111 = n15249;
  assign y112 = ~n15251;
  assign y113 = n15253;
  assign y114 = ~n15255;
  assign y115 = ~n15257;
  assign y116 = n15259;
  assign y117 = n15261;
  assign y118 = n15263;
  assign y119 = ~n15265;
  assign y120 = ~n15267;
  assign y121 = ~n15269;
  assign y122 = ~n15271;
  assign y123 = ~n15273;
  assign y124 = n15275;
  assign y125 = ~n15277;
  assign y126 = n15279;
  assign y127 = n15285;
endmodule
