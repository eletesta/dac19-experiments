// Benchmark "bar" written by ABC on Mon Nov 19 13:01:30 2018

module bar ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127;
  wire n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
    n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
    n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
    n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
    n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
    n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
    n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
    n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
    n925, n926, n927, n928, n929, n931, n932, n933, n934, n935, n936, n937,
    n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
    n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
    n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
    n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
    n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
    n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
    n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
    n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
    n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
    n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
    n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
    n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
    n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
    n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
    n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1216, n1217, n1218,
    n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
    n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
    n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
    n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
    n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
    n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
    n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
    n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
    n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
    n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
    n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
    n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
    n1399, n1400, n1401, n1402, n1403, n1405, n1406, n1407, n1408, n1409,
    n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
    n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
    n1470, n1471, n1472, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
    n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
    n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
    n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
    n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
    n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
    n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1612,
    n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
    n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
    n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
    n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
    n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
    n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
    n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
    n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1750, n1751, n1752, n1753, n1754,
    n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
    n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
    n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
    n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
    n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
    n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
    n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
    n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
    n1886, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
    n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
    n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
    n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
    n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
    n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
    n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1957,
    n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
    n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
    n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
    n1998, n1999, n2000, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
    n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
    n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
    n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
    n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
    n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
    n2090, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132, n2133, n2134, n2135, n2137, n2138, n2139, n2140, n2141,
    n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2152,
    n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
    n2163, n2164, n2165, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
    n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2182, n2183, n2184,
    n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
    n2195, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2212, n2213, n2214, n2215, n2216,
    n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2227,
    n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
    n2238, n2239, n2240, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
    n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
    n2270, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
    n2281, n2282, n2283, n2284, n2285, n2287, n2288, n2289, n2290, n2291,
    n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2302,
    n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
    n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2332, n2333, n2334,
    n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
    n2345, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2362, n2363, n2364, n2365, n2366,
    n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2377,
    n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
    n2388, n2389, n2390, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
    n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
    n2420, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
    n2431, n2432, n2433, n2434, n2435, n2437, n2438, n2439, n2440, n2441,
    n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2452,
    n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
    n2463, n2464, n2465, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
    n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2482, n2483, n2484,
    n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
    n2495, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2512, n2513, n2514, n2515, n2516,
    n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2527,
    n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
    n2538, n2539, n2540, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
    n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
    n2570, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2584, n2585, n2587, n2588, n2589, n2590, n2591,
    n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2602,
    n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
    n2613, n2614, n2615, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
    n2624, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2635,
    n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2644, n2645, n2646,
    n2647, n2648, n2649, n2650, n2651, n2653, n2654, n2655, n2656, n2657,
    n2658, n2659, n2660, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
    n2669, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2680,
    n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2689, n2690, n2691,
    n2692, n2693, n2694, n2695, n2696, n2698, n2699, n2700, n2701, n2702,
    n2703, n2704, n2705, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
    n2714, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2725,
    n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2734, n2735, n2736,
    n2737, n2738, n2739, n2740, n2741, n2743, n2744, n2745, n2746, n2747,
    n2748, n2749, n2750, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
    n2759, n2761, n2762, n2764, n2765, n2767, n2768, n2770, n2771, n2773,
    n2774, n2776, n2777, n2779, n2780, n2782, n2783, n2785, n2786, n2788,
    n2789, n2791, n2792, n2794, n2795, n2797, n2798, n2800, n2801, n2803,
    n2804, n2806, n2807, n2809, n2810, n2812, n2813, n2815, n2816, n2818,
    n2819, n2821, n2822, n2824, n2825, n2827, n2828, n2830, n2831, n2833,
    n2834, n2836, n2837, n2839, n2840, n2842, n2843, n2845, n2846, n2848,
    n2849, n2851, n2852, n2854, n2855, n2857, n2858, n2860, n2861, n2863,
    n2864, n2866, n2867, n2869, n2870, n2872, n2873, n2875, n2876, n2878,
    n2879, n2881, n2882, n2884, n2885, n2887, n2888, n2890, n2891, n2893,
    n2894, n2896, n2897, n2899, n2900, n2902, n2903, n2905, n2906, n2908,
    n2909, n2911, n2912, n2914, n2915, n2917, n2918, n2920, n2921, n2923,
    n2924, n2926, n2927, n2929, n2930, n2932, n2933, n2935, n2936, n2938,
    n2939, n2941, n2942, n2944, n2945, n2947, n2948, n2950, n2951;
  assign n265 = pi062 & pi129;
  assign n266 = pi064 & ~pi129;
  assign n267 = ~n265 & ~n266;
  assign n268 = n267 & ~pi128;
  assign n269 = pi061 & pi129;
  assign n270 = pi063 & ~pi129;
  assign n271 = ~n269 & ~n270;
  assign n272 = n271 & pi128;
  assign n273 = ~n268 & ~n272;
  assign n274 = n273 & ~pi131;
  assign n275 = pi054 & pi129;
  assign n276 = pi056 & ~pi129;
  assign n277 = ~n275 & ~n276;
  assign n278 = n277 & ~pi128;
  assign n279 = pi053 & pi129;
  assign n280 = pi055 & ~pi129;
  assign n281 = ~n279 & ~n280;
  assign n282 = n281 & pi128;
  assign n283 = ~n278 & ~n282;
  assign n284 = n283 & pi131;
  assign n285 = ~n274 & ~n284;
  assign n286 = n285 & ~pi130;
  assign n287 = pi058 & pi129;
  assign n288 = pi060 & ~pi129;
  assign n289 = ~n287 & ~n288;
  assign n290 = n289 & ~pi128;
  assign n291 = pi057 & pi129;
  assign n292 = pi059 & ~pi129;
  assign n293 = ~n291 & ~n292;
  assign n294 = n293 & pi128;
  assign n295 = ~n290 & ~n294;
  assign n296 = n295 & ~pi131;
  assign n297 = pi050 & pi129;
  assign n298 = pi052 & ~pi129;
  assign n299 = ~n297 & ~n298;
  assign n300 = n299 & ~pi128;
  assign n301 = pi049 & pi129;
  assign n302 = pi051 & ~pi129;
  assign n303 = ~n301 & ~n302;
  assign n304 = n303 & pi128;
  assign n305 = ~n300 & ~n304;
  assign n306 = n305 & pi131;
  assign n307 = ~n296 & ~n306;
  assign n308 = n307 & pi130;
  assign n309 = ~n286 & ~n308;
  assign n310 = n309 & ~pi133;
  assign n311 = pi030 & pi129;
  assign n312 = pi032 & ~pi129;
  assign n313 = ~n311 & ~n312;
  assign n314 = n313 & ~pi128;
  assign n315 = pi029 & pi129;
  assign n316 = pi031 & ~pi129;
  assign n317 = ~n315 & ~n316;
  assign n318 = n317 & pi128;
  assign n319 = ~n314 & ~n318;
  assign n320 = n319 & ~pi131;
  assign n321 = pi022 & pi129;
  assign n322 = pi024 & ~pi129;
  assign n323 = ~n321 & ~n322;
  assign n324 = n323 & ~pi128;
  assign n325 = pi021 & pi129;
  assign n326 = pi023 & ~pi129;
  assign n327 = ~n325 & ~n326;
  assign n328 = n327 & pi128;
  assign n329 = ~n324 & ~n328;
  assign n330 = n329 & pi131;
  assign n331 = ~n320 & ~n330;
  assign n332 = n331 & ~pi130;
  assign n333 = pi026 & pi129;
  assign n334 = pi028 & ~pi129;
  assign n335 = ~n333 & ~n334;
  assign n336 = n335 & ~pi128;
  assign n337 = pi025 & pi129;
  assign n338 = pi027 & ~pi129;
  assign n339 = ~n337 & ~n338;
  assign n340 = n339 & pi128;
  assign n341 = ~n336 & ~n340;
  assign n342 = n341 & ~pi131;
  assign n343 = pi018 & pi129;
  assign n344 = pi020 & ~pi129;
  assign n345 = ~n343 & ~n344;
  assign n346 = n345 & ~pi128;
  assign n347 = pi017 & pi129;
  assign n348 = pi019 & ~pi129;
  assign n349 = ~n347 & ~n348;
  assign n350 = n349 & pi128;
  assign n351 = ~n346 & ~n350;
  assign n352 = n351 & pi131;
  assign n353 = ~n342 & ~n352;
  assign n354 = n353 & pi130;
  assign n355 = ~n332 & ~n354;
  assign n356 = n355 & pi133;
  assign n357 = ~n310 & ~n356;
  assign n358 = n357 & ~pi132;
  assign n359 = pi046 & pi129;
  assign n360 = pi048 & ~pi129;
  assign n361 = ~n359 & ~n360;
  assign n362 = n361 & ~pi128;
  assign n363 = pi045 & pi129;
  assign n364 = pi047 & ~pi129;
  assign n365 = ~n363 & ~n364;
  assign n366 = n365 & pi128;
  assign n367 = ~n362 & ~n366;
  assign n368 = ~n367 & ~pi131;
  assign n369 = pi038 & pi129;
  assign n370 = pi040 & ~pi129;
  assign n371 = ~n369 & ~n370;
  assign n372 = n371 & ~pi128;
  assign n373 = pi037 & pi129;
  assign n374 = pi039 & ~pi129;
  assign n375 = ~n373 & ~n374;
  assign n376 = n375 & pi128;
  assign n377 = ~n372 & ~n376;
  assign n378 = ~n377 & pi131;
  assign n379 = ~n368 & ~n378;
  assign n380 = ~n379 & ~pi130;
  assign n381 = pi042 & pi129;
  assign n382 = pi044 & ~pi129;
  assign n383 = ~n381 & ~n382;
  assign n384 = n383 & ~pi128;
  assign n385 = pi041 & pi129;
  assign n386 = pi043 & ~pi129;
  assign n387 = ~n385 & ~n386;
  assign n388 = n387 & pi128;
  assign n389 = ~n384 & ~n388;
  assign n390 = n389 & ~pi131;
  assign n391 = pi034 & pi129;
  assign n392 = pi036 & ~pi129;
  assign n393 = ~n391 & ~n392;
  assign n394 = n393 & ~pi128;
  assign n395 = pi033 & pi129;
  assign n396 = pi035 & ~pi129;
  assign n397 = ~n395 & ~n396;
  assign n398 = n397 & pi128;
  assign n399 = ~n394 & ~n398;
  assign n400 = n399 & pi131;
  assign n401 = ~n390 & ~n400;
  assign n402 = n401 & pi130;
  assign n403 = ~n380 & ~n402;
  assign n404 = n403 & ~pi133;
  assign n405 = pi014 & pi129;
  assign n406 = pi016 & ~pi129;
  assign n407 = ~n405 & ~n406;
  assign n408 = n407 & ~pi128;
  assign n409 = pi013 & pi129;
  assign n410 = pi015 & ~pi129;
  assign n411 = ~n409 & ~n410;
  assign n412 = n411 & pi128;
  assign n413 = ~n408 & ~n412;
  assign n414 = n413 & ~pi131;
  assign n415 = pi006 & pi129;
  assign n416 = pi008 & ~pi129;
  assign n417 = ~n415 & ~n416;
  assign n418 = n417 & ~pi128;
  assign n419 = pi005 & pi129;
  assign n420 = pi007 & ~pi129;
  assign n421 = ~n419 & ~n420;
  assign n422 = n421 & pi128;
  assign n423 = ~n418 & ~n422;
  assign n424 = n423 & pi131;
  assign n425 = ~n414 & ~n424;
  assign n426 = n425 & ~pi130;
  assign n427 = pi010 & pi129;
  assign n428 = pi012 & ~pi129;
  assign n429 = ~n427 & ~n428;
  assign n430 = n429 & ~pi128;
  assign n431 = pi009 & pi129;
  assign n432 = pi011 & ~pi129;
  assign n433 = ~n431 & ~n432;
  assign n434 = n433 & pi128;
  assign n435 = ~n430 & ~n434;
  assign n436 = n435 & ~pi131;
  assign n437 = pi002 & pi129;
  assign n438 = pi004 & ~pi129;
  assign n439 = ~n437 & ~n438;
  assign n440 = n439 & ~pi128;
  assign n441 = pi001 & pi129;
  assign n442 = pi003 & ~pi129;
  assign n443 = ~n441 & ~n442;
  assign n444 = n443 & pi128;
  assign n445 = ~n440 & ~n444;
  assign n446 = n445 & pi131;
  assign n447 = ~n436 & ~n446;
  assign n448 = n447 & pi130;
  assign n449 = ~n426 & ~n448;
  assign n450 = n449 & pi133;
  assign n451 = ~n404 & ~n450;
  assign n452 = n451 & pi132;
  assign n453 = ~n358 & ~n452;
  assign n454 = n453 & pi134;
  assign n455 = pi126 & pi129;
  assign n456 = pi000 & ~pi129;
  assign n457 = ~n455 & ~n456;
  assign n458 = n457 & ~pi128;
  assign n459 = pi125 & pi129;
  assign n460 = pi127 & ~pi129;
  assign n461 = ~n459 & ~n460;
  assign n462 = n461 & pi128;
  assign n463 = ~n458 & ~n462;
  assign n464 = n463 & ~pi131;
  assign n465 = pi118 & pi129;
  assign n466 = pi120 & ~pi129;
  assign n467 = ~n465 & ~n466;
  assign n468 = n467 & ~pi128;
  assign n469 = pi117 & pi129;
  assign n470 = pi119 & ~pi129;
  assign n471 = ~n469 & ~n470;
  assign n472 = n471 & pi128;
  assign n473 = ~n468 & ~n472;
  assign n474 = n473 & pi131;
  assign n475 = ~n464 & ~n474;
  assign n476 = n475 & ~pi130;
  assign n477 = pi122 & pi129;
  assign n478 = pi124 & ~pi129;
  assign n479 = ~n477 & ~n478;
  assign n480 = n479 & ~pi128;
  assign n481 = pi121 & pi129;
  assign n482 = pi123 & ~pi129;
  assign n483 = ~n481 & ~n482;
  assign n484 = n483 & pi128;
  assign n485 = ~n480 & ~n484;
  assign n486 = n485 & ~pi131;
  assign n487 = pi114 & pi129;
  assign n488 = pi116 & ~pi129;
  assign n489 = ~n487 & ~n488;
  assign n490 = n489 & ~pi128;
  assign n491 = pi113 & pi129;
  assign n492 = pi115 & ~pi129;
  assign n493 = ~n491 & ~n492;
  assign n494 = n493 & pi128;
  assign n495 = ~n490 & ~n494;
  assign n496 = n495 & pi131;
  assign n497 = ~n486 & ~n496;
  assign n498 = n497 & pi130;
  assign n499 = ~n476 & ~n498;
  assign n500 = n499 & ~pi133;
  assign n501 = pi094 & pi129;
  assign n502 = pi096 & ~pi129;
  assign n503 = ~n501 & ~n502;
  assign n504 = n503 & ~pi128;
  assign n505 = pi093 & pi129;
  assign n506 = pi095 & ~pi129;
  assign n507 = ~n505 & ~n506;
  assign n508 = n507 & pi128;
  assign n509 = ~n504 & ~n508;
  assign n510 = n509 & ~pi131;
  assign n511 = pi086 & pi129;
  assign n512 = pi088 & ~pi129;
  assign n513 = ~n511 & ~n512;
  assign n514 = n513 & ~pi128;
  assign n515 = pi085 & pi129;
  assign n516 = pi087 & ~pi129;
  assign n517 = ~n515 & ~n516;
  assign n518 = n517 & pi128;
  assign n519 = ~n514 & ~n518;
  assign n520 = n519 & pi131;
  assign n521 = ~n510 & ~n520;
  assign n522 = n521 & ~pi130;
  assign n523 = pi090 & pi129;
  assign n524 = pi092 & ~pi129;
  assign n525 = ~n523 & ~n524;
  assign n526 = n525 & ~pi128;
  assign n527 = pi089 & pi129;
  assign n528 = pi091 & ~pi129;
  assign n529 = ~n527 & ~n528;
  assign n530 = n529 & pi128;
  assign n531 = ~n526 & ~n530;
  assign n532 = n531 & ~pi131;
  assign n533 = pi082 & pi129;
  assign n534 = pi084 & ~pi129;
  assign n535 = ~n533 & ~n534;
  assign n536 = n535 & ~pi128;
  assign n537 = pi081 & pi129;
  assign n538 = pi083 & ~pi129;
  assign n539 = ~n537 & ~n538;
  assign n540 = n539 & pi128;
  assign n541 = ~n536 & ~n540;
  assign n542 = n541 & pi131;
  assign n543 = ~n532 & ~n542;
  assign n544 = n543 & pi130;
  assign n545 = ~n522 & ~n544;
  assign n546 = n545 & pi133;
  assign n547 = ~n500 & ~n546;
  assign n548 = n547 & ~pi132;
  assign n549 = pi110 & pi129;
  assign n550 = pi112 & ~pi129;
  assign n551 = ~n549 & ~n550;
  assign n552 = n551 & ~pi128;
  assign n553 = pi109 & pi129;
  assign n554 = pi111 & ~pi129;
  assign n555 = ~n553 & ~n554;
  assign n556 = n555 & pi128;
  assign n557 = ~n552 & ~n556;
  assign n558 = n557 & ~pi131;
  assign n559 = pi102 & pi129;
  assign n560 = pi104 & ~pi129;
  assign n561 = ~n559 & ~n560;
  assign n562 = n561 & ~pi128;
  assign n563 = pi101 & pi129;
  assign n564 = pi103 & ~pi129;
  assign n565 = ~n563 & ~n564;
  assign n566 = n565 & pi128;
  assign n567 = ~n562 & ~n566;
  assign n568 = n567 & pi131;
  assign n569 = ~n558 & ~n568;
  assign n570 = n569 & ~pi130;
  assign n571 = pi106 & pi129;
  assign n572 = pi108 & ~pi129;
  assign n573 = ~n571 & ~n572;
  assign n574 = n573 & ~pi128;
  assign n575 = pi105 & pi129;
  assign n576 = pi107 & ~pi129;
  assign n577 = ~n575 & ~n576;
  assign n578 = n577 & pi128;
  assign n579 = ~n574 & ~n578;
  assign n580 = n579 & ~pi131;
  assign n581 = pi098 & pi129;
  assign n582 = pi100 & ~pi129;
  assign n583 = ~n581 & ~n582;
  assign n584 = n583 & ~pi128;
  assign n585 = pi097 & pi129;
  assign n586 = pi099 & ~pi129;
  assign n587 = ~n585 & ~n586;
  assign n588 = n587 & pi128;
  assign n589 = ~n584 & ~n588;
  assign n590 = n589 & pi131;
  assign n591 = ~n580 & ~n590;
  assign n592 = n591 & pi130;
  assign n593 = ~n570 & ~n592;
  assign n594 = n593 & ~pi133;
  assign n595 = pi078 & pi129;
  assign n596 = pi080 & ~pi129;
  assign n597 = ~n595 & ~n596;
  assign n598 = n597 & ~pi128;
  assign n599 = pi077 & pi129;
  assign n600 = pi079 & ~pi129;
  assign n601 = ~n599 & ~n600;
  assign n602 = n601 & pi128;
  assign n603 = ~n598 & ~n602;
  assign n604 = n603 & ~pi131;
  assign n605 = pi070 & pi129;
  assign n606 = pi072 & ~pi129;
  assign n607 = ~n605 & ~n606;
  assign n608 = n607 & ~pi128;
  assign n609 = pi069 & pi129;
  assign n610 = pi071 & ~pi129;
  assign n611 = ~n609 & ~n610;
  assign n612 = n611 & pi128;
  assign n613 = ~n608 & ~n612;
  assign n614 = n613 & pi131;
  assign n615 = ~n604 & ~n614;
  assign n616 = n615 & ~pi130;
  assign n617 = pi074 & pi129;
  assign n618 = pi076 & ~pi129;
  assign n619 = ~n617 & ~n618;
  assign n620 = n619 & ~pi128;
  assign n621 = pi073 & pi129;
  assign n622 = pi075 & ~pi129;
  assign n623 = ~n621 & ~n622;
  assign n624 = n623 & pi128;
  assign n625 = ~n620 & ~n624;
  assign n626 = n625 & ~pi131;
  assign n627 = pi066 & pi129;
  assign n628 = pi068 & ~pi129;
  assign n629 = ~n627 & ~n628;
  assign n630 = n629 & ~pi128;
  assign n631 = pi065 & pi129;
  assign n632 = pi067 & ~pi129;
  assign n633 = ~n631 & ~n632;
  assign n634 = n633 & pi128;
  assign n635 = ~n630 & ~n634;
  assign n636 = n635 & pi131;
  assign n637 = ~n626 & ~n636;
  assign n638 = n637 & pi130;
  assign n639 = ~n616 & ~n638;
  assign n640 = n639 & pi133;
  assign n641 = ~n594 & ~n640;
  assign n642 = n641 & pi132;
  assign n643 = ~n548 & ~n642;
  assign n644 = n643 & ~pi134;
  assign po000 = n454 | n644;
  assign n646 = pi063 & pi129;
  assign n647 = pi065 & ~pi129;
  assign n648 = ~n646 & ~n647;
  assign n649 = n648 & ~pi128;
  assign n650 = n267 & pi128;
  assign n651 = ~n649 & ~n650;
  assign n652 = ~n651 & ~pi131;
  assign n653 = pi055 & pi129;
  assign n654 = pi057 & ~pi129;
  assign n655 = ~n653 & ~n654;
  assign n656 = n655 & ~pi128;
  assign n657 = n277 & pi128;
  assign n658 = ~n656 & ~n657;
  assign n659 = ~n658 & pi131;
  assign n660 = ~n652 & ~n659;
  assign n661 = ~n660 & ~pi130;
  assign n662 = pi059 & pi129;
  assign n663 = pi061 & ~pi129;
  assign n664 = ~n662 & ~n663;
  assign n665 = n664 & ~pi128;
  assign n666 = n289 & pi128;
  assign n667 = ~n665 & ~n666;
  assign n668 = ~n667 & ~pi131;
  assign n669 = pi051 & pi129;
  assign n670 = pi053 & ~pi129;
  assign n671 = ~n669 & ~n670;
  assign n672 = n671 & ~pi128;
  assign n673 = n299 & pi128;
  assign n674 = ~n672 & ~n673;
  assign n675 = ~n674 & pi131;
  assign n676 = ~n668 & ~n675;
  assign n677 = ~n676 & pi130;
  assign n678 = ~n661 & ~n677;
  assign n679 = n678 & ~pi133;
  assign n680 = pi031 & pi129;
  assign n681 = pi033 & ~pi129;
  assign n682 = ~n680 & ~n681;
  assign n683 = n682 & ~pi128;
  assign n684 = n313 & pi128;
  assign n685 = ~n683 & ~n684;
  assign n686 = ~n685 & ~pi131;
  assign n687 = pi023 & pi129;
  assign n688 = pi025 & ~pi129;
  assign n689 = ~n687 & ~n688;
  assign n690 = n689 & ~pi128;
  assign n691 = n323 & pi128;
  assign n692 = ~n690 & ~n691;
  assign n693 = ~n692 & pi131;
  assign n694 = ~n686 & ~n693;
  assign n695 = ~n694 & ~pi130;
  assign n696 = pi027 & pi129;
  assign n697 = pi029 & ~pi129;
  assign n698 = ~n696 & ~n697;
  assign n699 = n698 & ~pi128;
  assign n700 = n335 & pi128;
  assign n701 = ~n699 & ~n700;
  assign n702 = ~n701 & ~pi131;
  assign n703 = pi019 & pi129;
  assign n704 = pi021 & ~pi129;
  assign n705 = ~n703 & ~n704;
  assign n706 = n705 & ~pi128;
  assign n707 = n345 & pi128;
  assign n708 = ~n706 & ~n707;
  assign n709 = ~n708 & pi131;
  assign n710 = ~n702 & ~n709;
  assign n711 = ~n710 & pi130;
  assign n712 = ~n695 & ~n711;
  assign n713 = n712 & pi133;
  assign n714 = ~n679 & ~n713;
  assign n715 = n714 & ~pi132;
  assign n716 = pi047 & pi129;
  assign n717 = pi049 & ~pi129;
  assign n718 = ~n716 & ~n717;
  assign n719 = n718 & ~pi128;
  assign n720 = n361 & pi128;
  assign n721 = ~n719 & ~n720;
  assign n722 = ~n721 & ~pi131;
  assign n723 = pi039 & pi129;
  assign n724 = pi041 & ~pi129;
  assign n725 = ~n723 & ~n724;
  assign n726 = n725 & ~pi128;
  assign n727 = n371 & pi128;
  assign n728 = ~n726 & ~n727;
  assign n729 = ~n728 & pi131;
  assign n730 = ~n722 & ~n729;
  assign n731 = ~n730 & ~pi130;
  assign n732 = pi043 & pi129;
  assign n733 = pi045 & ~pi129;
  assign n734 = ~n732 & ~n733;
  assign n735 = n734 & ~pi128;
  assign n736 = n383 & pi128;
  assign n737 = ~n735 & ~n736;
  assign n738 = ~n737 & ~pi131;
  assign n739 = pi035 & pi129;
  assign n740 = pi037 & ~pi129;
  assign n741 = ~n739 & ~n740;
  assign n742 = n741 & ~pi128;
  assign n743 = n393 & pi128;
  assign n744 = ~n742 & ~n743;
  assign n745 = ~n744 & pi131;
  assign n746 = ~n738 & ~n745;
  assign n747 = ~n746 & pi130;
  assign n748 = ~n731 & ~n747;
  assign n749 = n748 & ~pi133;
  assign n750 = pi015 & pi129;
  assign n751 = pi017 & ~pi129;
  assign n752 = ~n750 & ~n751;
  assign n753 = n752 & ~pi128;
  assign n754 = n407 & pi128;
  assign n755 = ~n753 & ~n754;
  assign n756 = ~n755 & ~pi131;
  assign n757 = pi007 & pi129;
  assign n758 = pi009 & ~pi129;
  assign n759 = ~n757 & ~n758;
  assign n760 = n759 & ~pi128;
  assign n761 = n417 & pi128;
  assign n762 = ~n760 & ~n761;
  assign n763 = ~n762 & pi131;
  assign n764 = ~n756 & ~n763;
  assign n765 = ~n764 & ~pi130;
  assign n766 = pi011 & pi129;
  assign n767 = pi013 & ~pi129;
  assign n768 = ~n766 & ~n767;
  assign n769 = n768 & ~pi128;
  assign n770 = n429 & pi128;
  assign n771 = ~n769 & ~n770;
  assign n772 = ~n771 & ~pi131;
  assign n773 = pi003 & pi129;
  assign n774 = pi005 & ~pi129;
  assign n775 = ~n773 & ~n774;
  assign n776 = n775 & ~pi128;
  assign n777 = n439 & pi128;
  assign n778 = ~n776 & ~n777;
  assign n779 = ~n778 & pi131;
  assign n780 = ~n772 & ~n779;
  assign n781 = ~n780 & pi130;
  assign n782 = ~n765 & ~n781;
  assign n783 = n782 & pi133;
  assign n784 = ~n749 & ~n783;
  assign n785 = n784 & pi132;
  assign n786 = ~n715 & ~n785;
  assign n787 = n786 & pi134;
  assign n788 = pi127 & pi129;
  assign n789 = pi001 & ~pi129;
  assign n790 = ~n788 & ~n789;
  assign n791 = n790 & ~pi128;
  assign n792 = n457 & pi128;
  assign n793 = ~n791 & ~n792;
  assign n794 = ~n793 & ~pi131;
  assign n795 = pi119 & pi129;
  assign n796 = pi121 & ~pi129;
  assign n797 = ~n795 & ~n796;
  assign n798 = n797 & ~pi128;
  assign n799 = n467 & pi128;
  assign n800 = ~n798 & ~n799;
  assign n801 = ~n800 & pi131;
  assign n802 = ~n794 & ~n801;
  assign n803 = ~n802 & ~pi130;
  assign n804 = pi123 & pi129;
  assign n805 = pi125 & ~pi129;
  assign n806 = ~n804 & ~n805;
  assign n807 = n806 & ~pi128;
  assign n808 = n479 & pi128;
  assign n809 = ~n807 & ~n808;
  assign n810 = ~n809 & ~pi131;
  assign n811 = pi115 & pi129;
  assign n812 = pi117 & ~pi129;
  assign n813 = ~n811 & ~n812;
  assign n814 = n813 & ~pi128;
  assign n815 = n489 & pi128;
  assign n816 = ~n814 & ~n815;
  assign n817 = ~n816 & pi131;
  assign n818 = ~n810 & ~n817;
  assign n819 = ~n818 & pi130;
  assign n820 = ~n803 & ~n819;
  assign n821 = n820 & ~pi133;
  assign n822 = pi095 & pi129;
  assign n823 = pi097 & ~pi129;
  assign n824 = ~n822 & ~n823;
  assign n825 = n824 & ~pi128;
  assign n826 = n503 & pi128;
  assign n827 = ~n825 & ~n826;
  assign n828 = ~n827 & ~pi131;
  assign n829 = pi087 & pi129;
  assign n830 = pi089 & ~pi129;
  assign n831 = ~n829 & ~n830;
  assign n832 = n831 & ~pi128;
  assign n833 = n513 & pi128;
  assign n834 = ~n832 & ~n833;
  assign n835 = ~n834 & pi131;
  assign n836 = ~n828 & ~n835;
  assign n837 = ~n836 & ~pi130;
  assign n838 = pi091 & pi129;
  assign n839 = pi093 & ~pi129;
  assign n840 = ~n838 & ~n839;
  assign n841 = n840 & ~pi128;
  assign n842 = n525 & pi128;
  assign n843 = ~n841 & ~n842;
  assign n844 = ~n843 & ~pi131;
  assign n845 = pi083 & pi129;
  assign n846 = pi085 & ~pi129;
  assign n847 = ~n845 & ~n846;
  assign n848 = n847 & ~pi128;
  assign n849 = n535 & pi128;
  assign n850 = ~n848 & ~n849;
  assign n851 = ~n850 & pi131;
  assign n852 = ~n844 & ~n851;
  assign n853 = ~n852 & pi130;
  assign n854 = ~n837 & ~n853;
  assign n855 = n854 & pi133;
  assign n856 = ~n821 & ~n855;
  assign n857 = n856 & ~pi132;
  assign n858 = pi111 & pi129;
  assign n859 = pi113 & ~pi129;
  assign n860 = ~n858 & ~n859;
  assign n861 = n860 & ~pi128;
  assign n862 = n551 & pi128;
  assign n863 = ~n861 & ~n862;
  assign n864 = ~n863 & ~pi131;
  assign n865 = pi103 & pi129;
  assign n866 = pi105 & ~pi129;
  assign n867 = ~n865 & ~n866;
  assign n868 = n867 & ~pi128;
  assign n869 = n561 & pi128;
  assign n870 = ~n868 & ~n869;
  assign n871 = ~n870 & pi131;
  assign n872 = ~n864 & ~n871;
  assign n873 = ~n872 & ~pi130;
  assign n874 = pi107 & pi129;
  assign n875 = pi109 & ~pi129;
  assign n876 = ~n874 & ~n875;
  assign n877 = n876 & ~pi128;
  assign n878 = n573 & pi128;
  assign n879 = ~n877 & ~n878;
  assign n880 = ~n879 & ~pi131;
  assign n881 = pi099 & pi129;
  assign n882 = pi101 & ~pi129;
  assign n883 = ~n881 & ~n882;
  assign n884 = n883 & ~pi128;
  assign n885 = n583 & pi128;
  assign n886 = ~n884 & ~n885;
  assign n887 = ~n886 & pi131;
  assign n888 = ~n880 & ~n887;
  assign n889 = ~n888 & pi130;
  assign n890 = ~n873 & ~n889;
  assign n891 = n890 & ~pi133;
  assign n892 = pi079 & pi129;
  assign n893 = pi081 & ~pi129;
  assign n894 = ~n892 & ~n893;
  assign n895 = n894 & ~pi128;
  assign n896 = n597 & pi128;
  assign n897 = ~n895 & ~n896;
  assign n898 = ~n897 & ~pi131;
  assign n899 = pi071 & pi129;
  assign n900 = pi073 & ~pi129;
  assign n901 = ~n899 & ~n900;
  assign n902 = n901 & ~pi128;
  assign n903 = n607 & pi128;
  assign n904 = ~n902 & ~n903;
  assign n905 = ~n904 & pi131;
  assign n906 = ~n898 & ~n905;
  assign n907 = ~n906 & ~pi130;
  assign n908 = pi075 & pi129;
  assign n909 = pi077 & ~pi129;
  assign n910 = ~n908 & ~n909;
  assign n911 = n910 & ~pi128;
  assign n912 = n619 & pi128;
  assign n913 = ~n911 & ~n912;
  assign n914 = ~n913 & ~pi131;
  assign n915 = pi067 & pi129;
  assign n916 = pi069 & ~pi129;
  assign n917 = ~n915 & ~n916;
  assign n918 = n917 & ~pi128;
  assign n919 = n629 & pi128;
  assign n920 = ~n918 & ~n919;
  assign n921 = ~n920 & pi131;
  assign n922 = ~n914 & ~n921;
  assign n923 = ~n922 & pi130;
  assign n924 = ~n907 & ~n923;
  assign n925 = n924 & pi133;
  assign n926 = ~n891 & ~n925;
  assign n927 = n926 & pi132;
  assign n928 = ~n857 & ~n927;
  assign n929 = n928 & ~pi134;
  assign po001 = n787 | n929;
  assign n931 = pi064 & pi129;
  assign n932 = pi066 & ~pi129;
  assign n933 = ~n931 & ~n932;
  assign n934 = n933 & ~pi128;
  assign n935 = n648 & pi128;
  assign n936 = ~n934 & ~n935;
  assign n937 = ~n936 & ~pi131;
  assign n938 = pi056 & pi129;
  assign n939 = pi058 & ~pi129;
  assign n940 = ~n938 & ~n939;
  assign n941 = n940 & ~pi128;
  assign n942 = n655 & pi128;
  assign n943 = ~n941 & ~n942;
  assign n944 = ~n943 & pi131;
  assign n945 = ~n937 & ~n944;
  assign n946 = ~n945 & ~pi130;
  assign n947 = pi060 & pi129;
  assign n948 = pi062 & ~pi129;
  assign n949 = ~n947 & ~n948;
  assign n950 = n949 & ~pi128;
  assign n951 = n664 & pi128;
  assign n952 = ~n950 & ~n951;
  assign n953 = ~n952 & ~pi131;
  assign n954 = pi052 & pi129;
  assign n955 = pi054 & ~pi129;
  assign n956 = ~n954 & ~n955;
  assign n957 = n956 & ~pi128;
  assign n958 = n671 & pi128;
  assign n959 = ~n957 & ~n958;
  assign n960 = ~n959 & pi131;
  assign n961 = ~n953 & ~n960;
  assign n962 = ~n961 & pi130;
  assign n963 = ~n946 & ~n962;
  assign n964 = n963 & ~pi133;
  assign n965 = pi032 & pi129;
  assign n966 = pi034 & ~pi129;
  assign n967 = ~n965 & ~n966;
  assign n968 = n967 & ~pi128;
  assign n969 = n682 & pi128;
  assign n970 = ~n968 & ~n969;
  assign n971 = ~n970 & ~pi131;
  assign n972 = pi024 & pi129;
  assign n973 = pi026 & ~pi129;
  assign n974 = ~n972 & ~n973;
  assign n975 = n974 & ~pi128;
  assign n976 = n689 & pi128;
  assign n977 = ~n975 & ~n976;
  assign n978 = ~n977 & pi131;
  assign n979 = ~n971 & ~n978;
  assign n980 = ~n979 & ~pi130;
  assign n981 = pi028 & pi129;
  assign n982 = pi030 & ~pi129;
  assign n983 = ~n981 & ~n982;
  assign n984 = n983 & ~pi128;
  assign n985 = n698 & pi128;
  assign n986 = ~n984 & ~n985;
  assign n987 = ~n986 & ~pi131;
  assign n988 = pi020 & pi129;
  assign n989 = pi022 & ~pi129;
  assign n990 = ~n988 & ~n989;
  assign n991 = n990 & ~pi128;
  assign n992 = n705 & pi128;
  assign n993 = ~n991 & ~n992;
  assign n994 = ~n993 & pi131;
  assign n995 = ~n987 & ~n994;
  assign n996 = ~n995 & pi130;
  assign n997 = ~n980 & ~n996;
  assign n998 = n997 & pi133;
  assign n999 = ~n964 & ~n998;
  assign n1000 = n999 & ~pi132;
  assign n1001 = pi048 & pi129;
  assign n1002 = pi050 & ~pi129;
  assign n1003 = ~n1001 & ~n1002;
  assign n1004 = n1003 & ~pi128;
  assign n1005 = n718 & pi128;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = ~n1006 & ~pi131;
  assign n1008 = pi040 & pi129;
  assign n1009 = pi042 & ~pi129;
  assign n1010 = ~n1008 & ~n1009;
  assign n1011 = n1010 & ~pi128;
  assign n1012 = n725 & pi128;
  assign n1013 = ~n1011 & ~n1012;
  assign n1014 = ~n1013 & pi131;
  assign n1015 = ~n1007 & ~n1014;
  assign n1016 = ~n1015 & ~pi130;
  assign n1017 = pi044 & pi129;
  assign n1018 = pi046 & ~pi129;
  assign n1019 = ~n1017 & ~n1018;
  assign n1020 = n1019 & ~pi128;
  assign n1021 = n734 & pi128;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = ~n1022 & ~pi131;
  assign n1024 = pi036 & pi129;
  assign n1025 = pi038 & ~pi129;
  assign n1026 = ~n1024 & ~n1025;
  assign n1027 = n1026 & ~pi128;
  assign n1028 = n741 & pi128;
  assign n1029 = ~n1027 & ~n1028;
  assign n1030 = ~n1029 & pi131;
  assign n1031 = ~n1023 & ~n1030;
  assign n1032 = ~n1031 & pi130;
  assign n1033 = ~n1016 & ~n1032;
  assign n1034 = n1033 & ~pi133;
  assign n1035 = pi016 & pi129;
  assign n1036 = pi018 & ~pi129;
  assign n1037 = ~n1035 & ~n1036;
  assign n1038 = n1037 & ~pi128;
  assign n1039 = n752 & pi128;
  assign n1040 = ~n1038 & ~n1039;
  assign n1041 = ~n1040 & ~pi131;
  assign n1042 = pi008 & pi129;
  assign n1043 = pi010 & ~pi129;
  assign n1044 = ~n1042 & ~n1043;
  assign n1045 = n1044 & ~pi128;
  assign n1046 = n759 & pi128;
  assign n1047 = ~n1045 & ~n1046;
  assign n1048 = ~n1047 & pi131;
  assign n1049 = ~n1041 & ~n1048;
  assign n1050 = ~n1049 & ~pi130;
  assign n1051 = pi012 & pi129;
  assign n1052 = pi014 & ~pi129;
  assign n1053 = ~n1051 & ~n1052;
  assign n1054 = n1053 & ~pi128;
  assign n1055 = n768 & pi128;
  assign n1056 = ~n1054 & ~n1055;
  assign n1057 = ~n1056 & ~pi131;
  assign n1058 = pi004 & pi129;
  assign n1059 = pi006 & ~pi129;
  assign n1060 = ~n1058 & ~n1059;
  assign n1061 = n1060 & ~pi128;
  assign n1062 = n775 & pi128;
  assign n1063 = ~n1061 & ~n1062;
  assign n1064 = ~n1063 & pi131;
  assign n1065 = ~n1057 & ~n1064;
  assign n1066 = ~n1065 & pi130;
  assign n1067 = ~n1050 & ~n1066;
  assign n1068 = n1067 & pi133;
  assign n1069 = ~n1034 & ~n1068;
  assign n1070 = n1069 & pi132;
  assign n1071 = ~n1000 & ~n1070;
  assign n1072 = n1071 & pi134;
  assign n1073 = pi000 & pi129;
  assign n1074 = pi002 & ~pi129;
  assign n1075 = ~n1073 & ~n1074;
  assign n1076 = n1075 & ~pi128;
  assign n1077 = n790 & pi128;
  assign n1078 = ~n1076 & ~n1077;
  assign n1079 = ~n1078 & ~pi131;
  assign n1080 = pi120 & pi129;
  assign n1081 = pi122 & ~pi129;
  assign n1082 = ~n1080 & ~n1081;
  assign n1083 = n1082 & ~pi128;
  assign n1084 = n797 & pi128;
  assign n1085 = ~n1083 & ~n1084;
  assign n1086 = ~n1085 & pi131;
  assign n1087 = ~n1079 & ~n1086;
  assign n1088 = ~n1087 & ~pi130;
  assign n1089 = pi124 & pi129;
  assign n1090 = pi126 & ~pi129;
  assign n1091 = ~n1089 & ~n1090;
  assign n1092 = n1091 & ~pi128;
  assign n1093 = n806 & pi128;
  assign n1094 = ~n1092 & ~n1093;
  assign n1095 = ~n1094 & ~pi131;
  assign n1096 = pi116 & pi129;
  assign n1097 = pi118 & ~pi129;
  assign n1098 = ~n1096 & ~n1097;
  assign n1099 = n1098 & ~pi128;
  assign n1100 = n813 & pi128;
  assign n1101 = ~n1099 & ~n1100;
  assign n1102 = ~n1101 & pi131;
  assign n1103 = ~n1095 & ~n1102;
  assign n1104 = ~n1103 & pi130;
  assign n1105 = ~n1088 & ~n1104;
  assign n1106 = n1105 & ~pi133;
  assign n1107 = pi096 & pi129;
  assign n1108 = pi098 & ~pi129;
  assign n1109 = ~n1107 & ~n1108;
  assign n1110 = n1109 & ~pi128;
  assign n1111 = n824 & pi128;
  assign n1112 = ~n1110 & ~n1111;
  assign n1113 = ~n1112 & ~pi131;
  assign n1114 = pi088 & pi129;
  assign n1115 = pi090 & ~pi129;
  assign n1116 = ~n1114 & ~n1115;
  assign n1117 = n1116 & ~pi128;
  assign n1118 = n831 & pi128;
  assign n1119 = ~n1117 & ~n1118;
  assign n1120 = ~n1119 & pi131;
  assign n1121 = ~n1113 & ~n1120;
  assign n1122 = ~n1121 & ~pi130;
  assign n1123 = pi092 & pi129;
  assign n1124 = pi094 & ~pi129;
  assign n1125 = ~n1123 & ~n1124;
  assign n1126 = n1125 & ~pi128;
  assign n1127 = n840 & pi128;
  assign n1128 = ~n1126 & ~n1127;
  assign n1129 = ~n1128 & ~pi131;
  assign n1130 = pi084 & pi129;
  assign n1131 = pi086 & ~pi129;
  assign n1132 = ~n1130 & ~n1131;
  assign n1133 = n1132 & ~pi128;
  assign n1134 = n847 & pi128;
  assign n1135 = ~n1133 & ~n1134;
  assign n1136 = ~n1135 & pi131;
  assign n1137 = ~n1129 & ~n1136;
  assign n1138 = ~n1137 & pi130;
  assign n1139 = ~n1122 & ~n1138;
  assign n1140 = n1139 & pi133;
  assign n1141 = ~n1106 & ~n1140;
  assign n1142 = n1141 & ~pi132;
  assign n1143 = pi112 & pi129;
  assign n1144 = pi114 & ~pi129;
  assign n1145 = ~n1143 & ~n1144;
  assign n1146 = n1145 & ~pi128;
  assign n1147 = n860 & pi128;
  assign n1148 = ~n1146 & ~n1147;
  assign n1149 = ~n1148 & ~pi131;
  assign n1150 = pi104 & pi129;
  assign n1151 = pi106 & ~pi129;
  assign n1152 = ~n1150 & ~n1151;
  assign n1153 = n1152 & ~pi128;
  assign n1154 = n867 & pi128;
  assign n1155 = ~n1153 & ~n1154;
  assign n1156 = ~n1155 & pi131;
  assign n1157 = ~n1149 & ~n1156;
  assign n1158 = ~n1157 & ~pi130;
  assign n1159 = pi108 & pi129;
  assign n1160 = pi110 & ~pi129;
  assign n1161 = ~n1159 & ~n1160;
  assign n1162 = n1161 & ~pi128;
  assign n1163 = n876 & pi128;
  assign n1164 = ~n1162 & ~n1163;
  assign n1165 = ~n1164 & ~pi131;
  assign n1166 = pi100 & pi129;
  assign n1167 = pi102 & ~pi129;
  assign n1168 = ~n1166 & ~n1167;
  assign n1169 = n1168 & ~pi128;
  assign n1170 = n883 & pi128;
  assign n1171 = ~n1169 & ~n1170;
  assign n1172 = ~n1171 & pi131;
  assign n1173 = ~n1165 & ~n1172;
  assign n1174 = ~n1173 & pi130;
  assign n1175 = ~n1158 & ~n1174;
  assign n1176 = n1175 & ~pi133;
  assign n1177 = pi080 & pi129;
  assign n1178 = pi082 & ~pi129;
  assign n1179 = ~n1177 & ~n1178;
  assign n1180 = n1179 & ~pi128;
  assign n1181 = n894 & pi128;
  assign n1182 = ~n1180 & ~n1181;
  assign n1183 = ~n1182 & ~pi131;
  assign n1184 = pi072 & pi129;
  assign n1185 = pi074 & ~pi129;
  assign n1186 = ~n1184 & ~n1185;
  assign n1187 = n1186 & ~pi128;
  assign n1188 = n901 & pi128;
  assign n1189 = ~n1187 & ~n1188;
  assign n1190 = ~n1189 & pi131;
  assign n1191 = ~n1183 & ~n1190;
  assign n1192 = ~n1191 & ~pi130;
  assign n1193 = pi076 & pi129;
  assign n1194 = pi078 & ~pi129;
  assign n1195 = ~n1193 & ~n1194;
  assign n1196 = n1195 & ~pi128;
  assign n1197 = n910 & pi128;
  assign n1198 = ~n1196 & ~n1197;
  assign n1199 = ~n1198 & ~pi131;
  assign n1200 = pi068 & pi129;
  assign n1201 = pi070 & ~pi129;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = n1202 & ~pi128;
  assign n1204 = n917 & pi128;
  assign n1205 = ~n1203 & ~n1204;
  assign n1206 = ~n1205 & pi131;
  assign n1207 = ~n1199 & ~n1206;
  assign n1208 = ~n1207 & pi130;
  assign n1209 = ~n1192 & ~n1208;
  assign n1210 = n1209 & pi133;
  assign n1211 = ~n1176 & ~n1210;
  assign n1212 = n1211 & pi132;
  assign n1213 = ~n1142 & ~n1212;
  assign n1214 = n1213 & ~pi134;
  assign po002 = n1072 | n1214;
  assign n1216 = n933 & pi128;
  assign n1217 = n633 & ~pi128;
  assign n1218 = ~n1216 & ~n1217;
  assign n1219 = ~n1218 & ~pi131;
  assign n1220 = n940 & pi128;
  assign n1221 = n293 & ~pi128;
  assign n1222 = ~n1220 & ~n1221;
  assign n1223 = ~n1222 & pi131;
  assign n1224 = ~n1219 & ~n1223;
  assign n1225 = ~n1224 & ~pi130;
  assign n1226 = n949 & pi128;
  assign n1227 = n271 & ~pi128;
  assign n1228 = ~n1226 & ~n1227;
  assign n1229 = n1228 & ~pi131;
  assign n1230 = n956 & pi128;
  assign n1231 = n281 & ~pi128;
  assign n1232 = ~n1230 & ~n1231;
  assign n1233 = n1232 & pi131;
  assign n1234 = ~n1229 & ~n1233;
  assign n1235 = n1234 & pi130;
  assign n1236 = ~n1225 & ~n1235;
  assign n1237 = n1236 & ~pi133;
  assign n1238 = n967 & pi128;
  assign n1239 = n397 & ~pi128;
  assign n1240 = ~n1238 & ~n1239;
  assign n1241 = ~n1240 & ~pi131;
  assign n1242 = n974 & pi128;
  assign n1243 = n339 & ~pi128;
  assign n1244 = ~n1242 & ~n1243;
  assign n1245 = ~n1244 & pi131;
  assign n1246 = ~n1241 & ~n1245;
  assign n1247 = ~n1246 & ~pi130;
  assign n1248 = n983 & pi128;
  assign n1249 = n317 & ~pi128;
  assign n1250 = ~n1248 & ~n1249;
  assign n1251 = n1250 & ~pi131;
  assign n1252 = n990 & pi128;
  assign n1253 = n327 & ~pi128;
  assign n1254 = ~n1252 & ~n1253;
  assign n1255 = n1254 & pi131;
  assign n1256 = ~n1251 & ~n1255;
  assign n1257 = n1256 & pi130;
  assign n1258 = ~n1247 & ~n1257;
  assign n1259 = n1258 & pi133;
  assign n1260 = ~n1237 & ~n1259;
  assign n1261 = n1260 & ~pi132;
  assign n1262 = n1003 & pi128;
  assign n1263 = n303 & ~pi128;
  assign n1264 = ~n1262 & ~n1263;
  assign n1265 = n1264 & ~pi131;
  assign n1266 = n1010 & pi128;
  assign n1267 = n387 & ~pi128;
  assign n1268 = ~n1266 & ~n1267;
  assign n1269 = n1268 & pi131;
  assign n1270 = ~n1265 & ~n1269;
  assign n1271 = n1270 & ~pi130;
  assign n1272 = n1019 & pi128;
  assign n1273 = n365 & ~pi128;
  assign n1274 = ~n1272 & ~n1273;
  assign n1275 = ~n1274 & ~pi131;
  assign n1276 = n1026 & pi128;
  assign n1277 = n375 & ~pi128;
  assign n1278 = ~n1276 & ~n1277;
  assign n1279 = ~n1278 & pi131;
  assign n1280 = ~n1275 & ~n1279;
  assign n1281 = ~n1280 & pi130;
  assign n1282 = ~n1271 & ~n1281;
  assign n1283 = n1282 & ~pi133;
  assign n1284 = n1037 & pi128;
  assign n1285 = n349 & ~pi128;
  assign n1286 = ~n1284 & ~n1285;
  assign n1287 = n1286 & ~pi131;
  assign n1288 = n1044 & pi128;
  assign n1289 = n433 & ~pi128;
  assign n1290 = ~n1288 & ~n1289;
  assign n1291 = n1290 & pi131;
  assign n1292 = ~n1287 & ~n1291;
  assign n1293 = n1292 & ~pi130;
  assign n1294 = n1053 & pi128;
  assign n1295 = n411 & ~pi128;
  assign n1296 = ~n1294 & ~n1295;
  assign n1297 = n1296 & ~pi131;
  assign n1298 = n1060 & pi128;
  assign n1299 = n421 & ~pi128;
  assign n1300 = ~n1298 & ~n1299;
  assign n1301 = n1300 & pi131;
  assign n1302 = ~n1297 & ~n1301;
  assign n1303 = n1302 & pi130;
  assign n1304 = ~n1293 & ~n1303;
  assign n1305 = n1304 & pi133;
  assign n1306 = ~n1283 & ~n1305;
  assign n1307 = n1306 & pi132;
  assign n1308 = ~n1261 & ~n1307;
  assign n1309 = n1308 & pi134;
  assign n1310 = n1075 & pi128;
  assign n1311 = n443 & ~pi128;
  assign n1312 = ~n1310 & ~n1311;
  assign n1313 = n1312 & ~pi131;
  assign n1314 = n1082 & pi128;
  assign n1315 = n483 & ~pi128;
  assign n1316 = ~n1314 & ~n1315;
  assign n1317 = n1316 & pi131;
  assign n1318 = ~n1313 & ~n1317;
  assign n1319 = n1318 & ~pi130;
  assign n1320 = n1091 & pi128;
  assign n1321 = n461 & ~pi128;
  assign n1322 = ~n1320 & ~n1321;
  assign n1323 = n1322 & ~pi131;
  assign n1324 = n1098 & pi128;
  assign n1325 = n471 & ~pi128;
  assign n1326 = ~n1324 & ~n1325;
  assign n1327 = n1326 & pi131;
  assign n1328 = ~n1323 & ~n1327;
  assign n1329 = n1328 & pi130;
  assign n1330 = ~n1319 & ~n1329;
  assign n1331 = n1330 & ~pi133;
  assign n1332 = n1109 & pi128;
  assign n1333 = n587 & ~pi128;
  assign n1334 = ~n1332 & ~n1333;
  assign n1335 = ~n1334 & ~pi131;
  assign n1336 = n1116 & pi128;
  assign n1337 = n529 & ~pi128;
  assign n1338 = ~n1336 & ~n1337;
  assign n1339 = ~n1338 & pi131;
  assign n1340 = ~n1335 & ~n1339;
  assign n1341 = ~n1340 & ~pi130;
  assign n1342 = n1125 & pi128;
  assign n1343 = n507 & ~pi128;
  assign n1344 = ~n1342 & ~n1343;
  assign n1345 = n1344 & ~pi131;
  assign n1346 = n1132 & pi128;
  assign n1347 = n517 & ~pi128;
  assign n1348 = ~n1346 & ~n1347;
  assign n1349 = n1348 & pi131;
  assign n1350 = ~n1345 & ~n1349;
  assign n1351 = n1350 & pi130;
  assign n1352 = ~n1341 & ~n1351;
  assign n1353 = n1352 & pi133;
  assign n1354 = ~n1331 & ~n1353;
  assign n1355 = n1354 & ~pi132;
  assign n1356 = n1145 & pi128;
  assign n1357 = n493 & ~pi128;
  assign n1358 = ~n1356 & ~n1357;
  assign n1359 = n1358 & ~pi131;
  assign n1360 = n1152 & pi128;
  assign n1361 = n577 & ~pi128;
  assign n1362 = ~n1360 & ~n1361;
  assign n1363 = n1362 & pi131;
  assign n1364 = ~n1359 & ~n1363;
  assign n1365 = n1364 & ~pi130;
  assign n1366 = n1161 & pi128;
  assign n1367 = n555 & ~pi128;
  assign n1368 = ~n1366 & ~n1367;
  assign n1369 = n1368 & ~pi131;
  assign n1370 = n1168 & pi128;
  assign n1371 = n565 & ~pi128;
  assign n1372 = ~n1370 & ~n1371;
  assign n1373 = n1372 & pi131;
  assign n1374 = ~n1369 & ~n1373;
  assign n1375 = n1374 & pi130;
  assign n1376 = ~n1365 & ~n1375;
  assign n1377 = n1376 & ~pi133;
  assign n1378 = n1179 & pi128;
  assign n1379 = n539 & ~pi128;
  assign n1380 = ~n1378 & ~n1379;
  assign n1381 = n1380 & ~pi131;
  assign n1382 = n1186 & pi128;
  assign n1383 = n623 & ~pi128;
  assign n1384 = ~n1382 & ~n1383;
  assign n1385 = n1384 & pi131;
  assign n1386 = ~n1381 & ~n1385;
  assign n1387 = n1386 & ~pi130;
  assign n1388 = n1195 & pi128;
  assign n1389 = n601 & ~pi128;
  assign n1390 = ~n1388 & ~n1389;
  assign n1391 = n1390 & ~pi131;
  assign n1392 = n1202 & pi128;
  assign n1393 = n611 & ~pi128;
  assign n1394 = ~n1392 & ~n1393;
  assign n1395 = n1394 & pi131;
  assign n1396 = ~n1391 & ~n1395;
  assign n1397 = n1396 & pi130;
  assign n1398 = ~n1387 & ~n1397;
  assign n1399 = n1398 & pi133;
  assign n1400 = ~n1377 & ~n1399;
  assign n1401 = n1400 & pi132;
  assign n1402 = ~n1355 & ~n1401;
  assign n1403 = n1402 & ~pi134;
  assign po003 = n1309 | n1403;
  assign n1405 = ~n635 & ~pi131;
  assign n1406 = ~n295 & pi131;
  assign n1407 = ~n1405 & ~n1406;
  assign n1408 = ~n1407 & ~pi130;
  assign n1409 = n285 & pi130;
  assign n1410 = ~n1408 & ~n1409;
  assign n1411 = ~n1410 & ~pi133;
  assign n1412 = ~n399 & ~pi131;
  assign n1413 = ~n341 & pi131;
  assign n1414 = ~n1412 & ~n1413;
  assign n1415 = ~n1414 & ~pi130;
  assign n1416 = n331 & pi130;
  assign n1417 = ~n1415 & ~n1416;
  assign n1418 = ~n1417 & pi133;
  assign n1419 = ~n1411 & ~n1418;
  assign n1420 = ~n1419 & ~pi132;
  assign n1421 = n305 & ~pi131;
  assign n1422 = n389 & pi131;
  assign n1423 = ~n1421 & ~n1422;
  assign n1424 = n1423 & ~pi130;
  assign n1425 = ~n379 & pi130;
  assign n1426 = ~n1424 & ~n1425;
  assign n1427 = ~n1426 & ~pi133;
  assign n1428 = n351 & ~pi131;
  assign n1429 = n435 & pi131;
  assign n1430 = ~n1428 & ~n1429;
  assign n1431 = n1430 & ~pi130;
  assign n1432 = n425 & pi130;
  assign n1433 = ~n1431 & ~n1432;
  assign n1434 = ~n1433 & pi133;
  assign n1435 = ~n1427 & ~n1434;
  assign n1436 = ~n1435 & pi132;
  assign n1437 = ~n1420 & ~n1436;
  assign n1438 = n1437 & pi134;
  assign n1439 = n445 & ~pi131;
  assign n1440 = n485 & pi131;
  assign n1441 = ~n1439 & ~n1440;
  assign n1442 = n1441 & ~pi130;
  assign n1443 = n475 & pi130;
  assign n1444 = ~n1442 & ~n1443;
  assign n1445 = ~n1444 & ~pi133;
  assign n1446 = ~n589 & ~pi131;
  assign n1447 = ~n531 & pi131;
  assign n1448 = ~n1446 & ~n1447;
  assign n1449 = ~n1448 & ~pi130;
  assign n1450 = n521 & pi130;
  assign n1451 = ~n1449 & ~n1450;
  assign n1452 = ~n1451 & pi133;
  assign n1453 = ~n1445 & ~n1452;
  assign n1454 = ~n1453 & ~pi132;
  assign n1455 = n495 & ~pi131;
  assign n1456 = n579 & pi131;
  assign n1457 = ~n1455 & ~n1456;
  assign n1458 = n1457 & ~pi130;
  assign n1459 = n569 & pi130;
  assign n1460 = ~n1458 & ~n1459;
  assign n1461 = ~n1460 & ~pi133;
  assign n1462 = n541 & ~pi131;
  assign n1463 = n625 & pi131;
  assign n1464 = ~n1462 & ~n1463;
  assign n1465 = n1464 & ~pi130;
  assign n1466 = n615 & pi130;
  assign n1467 = ~n1465 & ~n1466;
  assign n1468 = ~n1467 & pi133;
  assign n1469 = ~n1461 & ~n1468;
  assign n1470 = ~n1469 & pi132;
  assign n1471 = ~n1454 & ~n1470;
  assign n1472 = n1471 & ~pi134;
  assign po004 = n1438 | n1472;
  assign n1474 = ~n920 & ~pi131;
  assign n1475 = ~n667 & pi131;
  assign n1476 = ~n1474 & ~n1475;
  assign n1477 = ~n1476 & ~pi130;
  assign n1478 = ~n660 & pi130;
  assign n1479 = ~n1477 & ~n1478;
  assign n1480 = ~n1479 & ~pi133;
  assign n1481 = ~n744 & ~pi131;
  assign n1482 = ~n701 & pi131;
  assign n1483 = ~n1481 & ~n1482;
  assign n1484 = ~n1483 & ~pi130;
  assign n1485 = ~n694 & pi130;
  assign n1486 = ~n1484 & ~n1485;
  assign n1487 = ~n1486 & pi133;
  assign n1488 = ~n1480 & ~n1487;
  assign n1489 = ~n1488 & ~pi132;
  assign n1490 = ~n674 & ~pi131;
  assign n1491 = ~n737 & pi131;
  assign n1492 = ~n1490 & ~n1491;
  assign n1493 = ~n1492 & ~pi130;
  assign n1494 = ~n730 & pi130;
  assign n1495 = ~n1493 & ~n1494;
  assign n1496 = ~n1495 & ~pi133;
  assign n1497 = ~n708 & ~pi131;
  assign n1498 = ~n771 & pi131;
  assign n1499 = ~n1497 & ~n1498;
  assign n1500 = ~n1499 & ~pi130;
  assign n1501 = ~n764 & pi130;
  assign n1502 = ~n1500 & ~n1501;
  assign n1503 = ~n1502 & pi133;
  assign n1504 = ~n1496 & ~n1503;
  assign n1505 = ~n1504 & pi132;
  assign n1506 = ~n1489 & ~n1505;
  assign n1507 = n1506 & pi134;
  assign n1508 = ~n778 & ~pi131;
  assign n1509 = ~n809 & pi131;
  assign n1510 = ~n1508 & ~n1509;
  assign n1511 = ~n1510 & ~pi130;
  assign n1512 = ~n802 & pi130;
  assign n1513 = ~n1511 & ~n1512;
  assign n1514 = ~n1513 & ~pi133;
  assign n1515 = ~n886 & ~pi131;
  assign n1516 = ~n843 & pi131;
  assign n1517 = ~n1515 & ~n1516;
  assign n1518 = ~n1517 & ~pi130;
  assign n1519 = ~n836 & pi130;
  assign n1520 = ~n1518 & ~n1519;
  assign n1521 = ~n1520 & pi133;
  assign n1522 = ~n1514 & ~n1521;
  assign n1523 = ~n1522 & ~pi132;
  assign n1524 = ~n816 & ~pi131;
  assign n1525 = ~n879 & pi131;
  assign n1526 = ~n1524 & ~n1525;
  assign n1527 = ~n1526 & ~pi130;
  assign n1528 = ~n872 & pi130;
  assign n1529 = ~n1527 & ~n1528;
  assign n1530 = ~n1529 & ~pi133;
  assign n1531 = ~n850 & ~pi131;
  assign n1532 = ~n913 & pi131;
  assign n1533 = ~n1531 & ~n1532;
  assign n1534 = ~n1533 & ~pi130;
  assign n1535 = ~n906 & pi130;
  assign n1536 = ~n1534 & ~n1535;
  assign n1537 = ~n1536 & pi133;
  assign n1538 = ~n1530 & ~n1537;
  assign n1539 = ~n1538 & pi132;
  assign n1540 = ~n1523 & ~n1539;
  assign n1541 = n1540 & ~pi134;
  assign po005 = n1507 | n1541;
  assign n1543 = ~n1205 & ~pi131;
  assign n1544 = ~n952 & pi131;
  assign n1545 = ~n1543 & ~n1544;
  assign n1546 = ~n1545 & ~pi130;
  assign n1547 = ~n945 & pi130;
  assign n1548 = ~n1546 & ~n1547;
  assign n1549 = ~n1548 & ~pi133;
  assign n1550 = ~n1029 & ~pi131;
  assign n1551 = ~n986 & pi131;
  assign n1552 = ~n1550 & ~n1551;
  assign n1553 = ~n1552 & ~pi130;
  assign n1554 = ~n979 & pi130;
  assign n1555 = ~n1553 & ~n1554;
  assign n1556 = ~n1555 & pi133;
  assign n1557 = ~n1549 & ~n1556;
  assign n1558 = ~n1557 & ~pi132;
  assign n1559 = ~n959 & ~pi131;
  assign n1560 = ~n1022 & pi131;
  assign n1561 = ~n1559 & ~n1560;
  assign n1562 = ~n1561 & ~pi130;
  assign n1563 = ~n1015 & pi130;
  assign n1564 = ~n1562 & ~n1563;
  assign n1565 = ~n1564 & ~pi133;
  assign n1566 = ~n993 & ~pi131;
  assign n1567 = ~n1056 & pi131;
  assign n1568 = ~n1566 & ~n1567;
  assign n1569 = ~n1568 & ~pi130;
  assign n1570 = ~n1049 & pi130;
  assign n1571 = ~n1569 & ~n1570;
  assign n1572 = ~n1571 & pi133;
  assign n1573 = ~n1565 & ~n1572;
  assign n1574 = ~n1573 & pi132;
  assign n1575 = ~n1558 & ~n1574;
  assign n1576 = n1575 & pi134;
  assign n1577 = ~n1063 & ~pi131;
  assign n1578 = ~n1094 & pi131;
  assign n1579 = ~n1577 & ~n1578;
  assign n1580 = ~n1579 & ~pi130;
  assign n1581 = ~n1087 & pi130;
  assign n1582 = ~n1580 & ~n1581;
  assign n1583 = ~n1582 & ~pi133;
  assign n1584 = ~n1171 & ~pi131;
  assign n1585 = ~n1128 & pi131;
  assign n1586 = ~n1584 & ~n1585;
  assign n1587 = ~n1586 & ~pi130;
  assign n1588 = ~n1121 & pi130;
  assign n1589 = ~n1587 & ~n1588;
  assign n1590 = ~n1589 & pi133;
  assign n1591 = ~n1583 & ~n1590;
  assign n1592 = ~n1591 & ~pi132;
  assign n1593 = ~n1101 & ~pi131;
  assign n1594 = ~n1164 & pi131;
  assign n1595 = ~n1593 & ~n1594;
  assign n1596 = ~n1595 & ~pi130;
  assign n1597 = ~n1157 & pi130;
  assign n1598 = ~n1596 & ~n1597;
  assign n1599 = ~n1598 & ~pi133;
  assign n1600 = ~n1135 & ~pi131;
  assign n1601 = ~n1198 & pi131;
  assign n1602 = ~n1600 & ~n1601;
  assign n1603 = ~n1602 & ~pi130;
  assign n1604 = ~n1191 & pi130;
  assign n1605 = ~n1603 & ~n1604;
  assign n1606 = ~n1605 & pi133;
  assign n1607 = ~n1599 & ~n1606;
  assign n1608 = ~n1607 & pi132;
  assign n1609 = ~n1592 & ~n1608;
  assign n1610 = n1609 & ~pi134;
  assign po006 = n1576 | n1610;
  assign n1612 = ~n1394 & ~pi131;
  assign n1613 = ~n1228 & pi131;
  assign n1614 = ~n1612 & ~n1613;
  assign n1615 = ~n1614 & ~pi130;
  assign n1616 = ~n1224 & pi130;
  assign n1617 = ~n1615 & ~n1616;
  assign n1618 = ~n1617 & ~pi133;
  assign n1619 = ~n1278 & ~pi131;
  assign n1620 = ~n1250 & pi131;
  assign n1621 = ~n1619 & ~n1620;
  assign n1622 = ~n1621 & ~pi130;
  assign n1623 = ~n1246 & pi130;
  assign n1624 = ~n1622 & ~n1623;
  assign n1625 = ~n1624 & pi133;
  assign n1626 = ~n1618 & ~n1625;
  assign n1627 = ~n1626 & ~pi132;
  assign n1628 = n1232 & ~pi131;
  assign n1629 = n1274 & pi131;
  assign n1630 = ~n1628 & ~n1629;
  assign n1631 = n1630 & ~pi130;
  assign n1632 = n1270 & pi130;
  assign n1633 = ~n1631 & ~n1632;
  assign n1634 = ~n1633 & ~pi133;
  assign n1635 = n1254 & ~pi131;
  assign n1636 = n1296 & pi131;
  assign n1637 = ~n1635 & ~n1636;
  assign n1638 = n1637 & ~pi130;
  assign n1639 = n1292 & pi130;
  assign n1640 = ~n1638 & ~n1639;
  assign n1641 = ~n1640 & pi133;
  assign n1642 = ~n1634 & ~n1641;
  assign n1643 = ~n1642 & pi132;
  assign n1644 = ~n1627 & ~n1643;
  assign n1645 = n1644 & pi134;
  assign n1646 = n1300 & ~pi131;
  assign n1647 = n1322 & pi131;
  assign n1648 = ~n1646 & ~n1647;
  assign n1649 = n1648 & ~pi130;
  assign n1650 = n1318 & pi130;
  assign n1651 = ~n1649 & ~n1650;
  assign n1652 = ~n1651 & ~pi133;
  assign n1653 = ~n1372 & ~pi131;
  assign n1654 = ~n1344 & pi131;
  assign n1655 = ~n1653 & ~n1654;
  assign n1656 = ~n1655 & ~pi130;
  assign n1657 = ~n1340 & pi130;
  assign n1658 = ~n1656 & ~n1657;
  assign n1659 = ~n1658 & pi133;
  assign n1660 = ~n1652 & ~n1659;
  assign n1661 = ~n1660 & ~pi132;
  assign n1662 = n1326 & ~pi131;
  assign n1663 = n1368 & pi131;
  assign n1664 = ~n1662 & ~n1663;
  assign n1665 = n1664 & ~pi130;
  assign n1666 = n1364 & pi130;
  assign n1667 = ~n1665 & ~n1666;
  assign n1668 = ~n1667 & ~pi133;
  assign n1669 = n1348 & ~pi131;
  assign n1670 = n1390 & pi131;
  assign n1671 = ~n1669 & ~n1670;
  assign n1672 = n1671 & ~pi130;
  assign n1673 = n1386 & pi130;
  assign n1674 = ~n1672 & ~n1673;
  assign n1675 = ~n1674 & pi133;
  assign n1676 = ~n1668 & ~n1675;
  assign n1677 = ~n1676 & pi132;
  assign n1678 = ~n1661 & ~n1677;
  assign n1679 = n1678 & ~pi134;
  assign po007 = n1645 | n1679;
  assign n1681 = ~n613 & ~pi131;
  assign n1682 = ~n273 & pi131;
  assign n1683 = ~n1681 & ~n1682;
  assign n1684 = ~n1683 & ~pi130;
  assign n1685 = ~n1407 & pi130;
  assign n1686 = ~n1684 & ~n1685;
  assign n1687 = ~n1686 & ~pi133;
  assign n1688 = ~n377 & ~pi131;
  assign n1689 = ~n319 & pi131;
  assign n1690 = ~n1688 & ~n1689;
  assign n1691 = ~n1690 & ~pi130;
  assign n1692 = ~n1414 & pi130;
  assign n1693 = ~n1691 & ~n1692;
  assign n1694 = ~n1693 & pi133;
  assign n1695 = ~n1687 & ~n1694;
  assign n1696 = ~n1695 & ~pi132;
  assign n1697 = n283 & ~pi131;
  assign n1698 = n367 & pi131;
  assign n1699 = ~n1697 & ~n1698;
  assign n1700 = n1699 & ~pi130;
  assign n1701 = n1423 & pi130;
  assign n1702 = ~n1700 & ~n1701;
  assign n1703 = ~n1702 & ~pi133;
  assign n1704 = n329 & ~pi131;
  assign n1705 = n413 & pi131;
  assign n1706 = ~n1704 & ~n1705;
  assign n1707 = n1706 & ~pi130;
  assign n1708 = n1430 & pi130;
  assign n1709 = ~n1707 & ~n1708;
  assign n1710 = ~n1709 & pi133;
  assign n1711 = ~n1703 & ~n1710;
  assign n1712 = ~n1711 & pi132;
  assign n1713 = ~n1696 & ~n1712;
  assign n1714 = n1713 & pi134;
  assign n1715 = n423 & ~pi131;
  assign n1716 = n463 & pi131;
  assign n1717 = ~n1715 & ~n1716;
  assign n1718 = n1717 & ~pi130;
  assign n1719 = n1441 & pi130;
  assign n1720 = ~n1718 & ~n1719;
  assign n1721 = ~n1720 & ~pi133;
  assign n1722 = ~n567 & ~pi131;
  assign n1723 = ~n509 & pi131;
  assign n1724 = ~n1722 & ~n1723;
  assign n1725 = ~n1724 & ~pi130;
  assign n1726 = ~n1448 & pi130;
  assign n1727 = ~n1725 & ~n1726;
  assign n1728 = ~n1727 & pi133;
  assign n1729 = ~n1721 & ~n1728;
  assign n1730 = ~n1729 & ~pi132;
  assign n1731 = n473 & ~pi131;
  assign n1732 = n557 & pi131;
  assign n1733 = ~n1731 & ~n1732;
  assign n1734 = n1733 & ~pi130;
  assign n1735 = n1457 & pi130;
  assign n1736 = ~n1734 & ~n1735;
  assign n1737 = ~n1736 & ~pi133;
  assign n1738 = n519 & ~pi131;
  assign n1739 = n603 & pi131;
  assign n1740 = ~n1738 & ~n1739;
  assign n1741 = n1740 & ~pi130;
  assign n1742 = n1464 & pi130;
  assign n1743 = ~n1741 & ~n1742;
  assign n1744 = ~n1743 & pi133;
  assign n1745 = ~n1737 & ~n1744;
  assign n1746 = ~n1745 & pi132;
  assign n1747 = ~n1730 & ~n1746;
  assign n1748 = n1747 & ~pi134;
  assign po008 = n1714 | n1748;
  assign n1750 = ~n904 & ~pi131;
  assign n1751 = ~n651 & pi131;
  assign n1752 = ~n1750 & ~n1751;
  assign n1753 = ~n1752 & ~pi130;
  assign n1754 = ~n1476 & pi130;
  assign n1755 = ~n1753 & ~n1754;
  assign n1756 = ~n1755 & ~pi133;
  assign n1757 = ~n728 & ~pi131;
  assign n1758 = ~n685 & pi131;
  assign n1759 = ~n1757 & ~n1758;
  assign n1760 = ~n1759 & ~pi130;
  assign n1761 = ~n1483 & pi130;
  assign n1762 = ~n1760 & ~n1761;
  assign n1763 = ~n1762 & pi133;
  assign n1764 = ~n1756 & ~n1763;
  assign n1765 = ~n1764 & ~pi132;
  assign n1766 = ~n658 & ~pi131;
  assign n1767 = ~n721 & pi131;
  assign n1768 = ~n1766 & ~n1767;
  assign n1769 = ~n1768 & ~pi130;
  assign n1770 = ~n1492 & pi130;
  assign n1771 = ~n1769 & ~n1770;
  assign n1772 = ~n1771 & ~pi133;
  assign n1773 = ~n692 & ~pi131;
  assign n1774 = ~n755 & pi131;
  assign n1775 = ~n1773 & ~n1774;
  assign n1776 = ~n1775 & ~pi130;
  assign n1777 = ~n1499 & pi130;
  assign n1778 = ~n1776 & ~n1777;
  assign n1779 = ~n1778 & pi133;
  assign n1780 = ~n1772 & ~n1779;
  assign n1781 = ~n1780 & pi132;
  assign n1782 = ~n1765 & ~n1781;
  assign n1783 = n1782 & pi134;
  assign n1784 = ~n762 & ~pi131;
  assign n1785 = ~n793 & pi131;
  assign n1786 = ~n1784 & ~n1785;
  assign n1787 = ~n1786 & ~pi130;
  assign n1788 = ~n1510 & pi130;
  assign n1789 = ~n1787 & ~n1788;
  assign n1790 = ~n1789 & ~pi133;
  assign n1791 = ~n870 & ~pi131;
  assign n1792 = ~n827 & pi131;
  assign n1793 = ~n1791 & ~n1792;
  assign n1794 = ~n1793 & ~pi130;
  assign n1795 = ~n1517 & pi130;
  assign n1796 = ~n1794 & ~n1795;
  assign n1797 = ~n1796 & pi133;
  assign n1798 = ~n1790 & ~n1797;
  assign n1799 = ~n1798 & ~pi132;
  assign n1800 = ~n800 & ~pi131;
  assign n1801 = ~n863 & pi131;
  assign n1802 = ~n1800 & ~n1801;
  assign n1803 = ~n1802 & ~pi130;
  assign n1804 = ~n1526 & pi130;
  assign n1805 = ~n1803 & ~n1804;
  assign n1806 = ~n1805 & ~pi133;
  assign n1807 = ~n834 & ~pi131;
  assign n1808 = ~n897 & pi131;
  assign n1809 = ~n1807 & ~n1808;
  assign n1810 = ~n1809 & ~pi130;
  assign n1811 = ~n1533 & pi130;
  assign n1812 = ~n1810 & ~n1811;
  assign n1813 = ~n1812 & pi133;
  assign n1814 = ~n1806 & ~n1813;
  assign n1815 = ~n1814 & pi132;
  assign n1816 = ~n1799 & ~n1815;
  assign n1817 = n1816 & ~pi134;
  assign po009 = n1783 | n1817;
  assign n1819 = ~n1189 & ~pi131;
  assign n1820 = ~n936 & pi131;
  assign n1821 = ~n1819 & ~n1820;
  assign n1822 = ~n1821 & ~pi130;
  assign n1823 = ~n1545 & pi130;
  assign n1824 = ~n1822 & ~n1823;
  assign n1825 = ~n1824 & ~pi133;
  assign n1826 = ~n1013 & ~pi131;
  assign n1827 = ~n970 & pi131;
  assign n1828 = ~n1826 & ~n1827;
  assign n1829 = ~n1828 & ~pi130;
  assign n1830 = ~n1552 & pi130;
  assign n1831 = ~n1829 & ~n1830;
  assign n1832 = ~n1831 & pi133;
  assign n1833 = ~n1825 & ~n1832;
  assign n1834 = ~n1833 & ~pi132;
  assign n1835 = ~n943 & ~pi131;
  assign n1836 = ~n1006 & pi131;
  assign n1837 = ~n1835 & ~n1836;
  assign n1838 = ~n1837 & ~pi130;
  assign n1839 = ~n1561 & pi130;
  assign n1840 = ~n1838 & ~n1839;
  assign n1841 = ~n1840 & ~pi133;
  assign n1842 = ~n977 & ~pi131;
  assign n1843 = ~n1040 & pi131;
  assign n1844 = ~n1842 & ~n1843;
  assign n1845 = ~n1844 & ~pi130;
  assign n1846 = ~n1568 & pi130;
  assign n1847 = ~n1845 & ~n1846;
  assign n1848 = ~n1847 & pi133;
  assign n1849 = ~n1841 & ~n1848;
  assign n1850 = ~n1849 & pi132;
  assign n1851 = ~n1834 & ~n1850;
  assign n1852 = n1851 & pi134;
  assign n1853 = ~n1047 & ~pi131;
  assign n1854 = ~n1078 & pi131;
  assign n1855 = ~n1853 & ~n1854;
  assign n1856 = ~n1855 & ~pi130;
  assign n1857 = ~n1579 & pi130;
  assign n1858 = ~n1856 & ~n1857;
  assign n1859 = ~n1858 & ~pi133;
  assign n1860 = ~n1155 & ~pi131;
  assign n1861 = ~n1112 & pi131;
  assign n1862 = ~n1860 & ~n1861;
  assign n1863 = ~n1862 & ~pi130;
  assign n1864 = ~n1586 & pi130;
  assign n1865 = ~n1863 & ~n1864;
  assign n1866 = ~n1865 & pi133;
  assign n1867 = ~n1859 & ~n1866;
  assign n1868 = ~n1867 & ~pi132;
  assign n1869 = ~n1085 & ~pi131;
  assign n1870 = ~n1148 & pi131;
  assign n1871 = ~n1869 & ~n1870;
  assign n1872 = ~n1871 & ~pi130;
  assign n1873 = ~n1595 & pi130;
  assign n1874 = ~n1872 & ~n1873;
  assign n1875 = ~n1874 & ~pi133;
  assign n1876 = ~n1119 & ~pi131;
  assign n1877 = ~n1182 & pi131;
  assign n1878 = ~n1876 & ~n1877;
  assign n1879 = ~n1878 & ~pi130;
  assign n1880 = ~n1602 & pi130;
  assign n1881 = ~n1879 & ~n1880;
  assign n1882 = ~n1881 & pi133;
  assign n1883 = ~n1875 & ~n1882;
  assign n1884 = ~n1883 & pi132;
  assign n1885 = ~n1868 & ~n1884;
  assign n1886 = n1885 & ~pi134;
  assign po010 = n1852 | n1886;
  assign n1888 = n1218 & pi131;
  assign n1889 = n1384 & ~pi131;
  assign n1890 = ~n1888 & ~n1889;
  assign n1891 = n1890 & ~pi130;
  assign n1892 = ~n1614 & pi130;
  assign n1893 = ~n1891 & ~n1892;
  assign n1894 = ~n1893 & ~pi133;
  assign n1895 = n1240 & pi131;
  assign n1896 = n1268 & ~pi131;
  assign n1897 = ~n1895 & ~n1896;
  assign n1898 = n1897 & ~pi130;
  assign n1899 = ~n1621 & pi130;
  assign n1900 = ~n1898 & ~n1899;
  assign n1901 = ~n1900 & pi133;
  assign n1902 = ~n1894 & ~n1901;
  assign n1903 = ~n1902 & ~pi132;
  assign n1904 = n1222 & ~pi131;
  assign n1905 = n1264 & pi131;
  assign n1906 = ~n1904 & ~n1905;
  assign n1907 = n1906 & ~pi130;
  assign n1908 = n1630 & pi130;
  assign n1909 = ~n1907 & ~n1908;
  assign n1910 = ~n1909 & ~pi133;
  assign n1911 = n1244 & ~pi131;
  assign n1912 = n1286 & pi131;
  assign n1913 = ~n1911 & ~n1912;
  assign n1914 = n1913 & ~pi130;
  assign n1915 = n1637 & pi130;
  assign n1916 = ~n1914 & ~n1915;
  assign n1917 = ~n1916 & pi133;
  assign n1918 = ~n1910 & ~n1917;
  assign n1919 = ~n1918 & pi132;
  assign n1920 = ~n1903 & ~n1919;
  assign n1921 = n1920 & pi134;
  assign n1922 = n1290 & ~pi131;
  assign n1923 = n1312 & pi131;
  assign n1924 = ~n1922 & ~n1923;
  assign n1925 = n1924 & ~pi130;
  assign n1926 = n1648 & pi130;
  assign n1927 = ~n1925 & ~n1926;
  assign n1928 = ~n1927 & ~pi133;
  assign n1929 = n1334 & pi131;
  assign n1930 = n1362 & ~pi131;
  assign n1931 = ~n1929 & ~n1930;
  assign n1932 = n1931 & ~pi130;
  assign n1933 = ~n1655 & pi130;
  assign n1934 = ~n1932 & ~n1933;
  assign n1935 = ~n1934 & pi133;
  assign n1936 = ~n1928 & ~n1935;
  assign n1937 = ~n1936 & ~pi132;
  assign n1938 = n1316 & ~pi131;
  assign n1939 = n1358 & pi131;
  assign n1940 = ~n1938 & ~n1939;
  assign n1941 = n1940 & ~pi130;
  assign n1942 = n1664 & pi130;
  assign n1943 = ~n1941 & ~n1942;
  assign n1944 = ~n1943 & ~pi133;
  assign n1945 = n1338 & ~pi131;
  assign n1946 = n1380 & pi131;
  assign n1947 = ~n1945 & ~n1946;
  assign n1948 = n1947 & ~pi130;
  assign n1949 = n1671 & pi130;
  assign n1950 = ~n1948 & ~n1949;
  assign n1951 = ~n1950 & pi133;
  assign n1952 = ~n1944 & ~n1951;
  assign n1953 = ~n1952 & pi132;
  assign n1954 = ~n1937 & ~n1953;
  assign n1955 = n1954 & ~pi134;
  assign po011 = n1921 | n1955;
  assign n1957 = ~n1683 & pi130;
  assign n1958 = n637 & ~pi130;
  assign n1959 = ~n1957 & ~n1958;
  assign n1960 = ~n1959 & ~pi133;
  assign n1961 = ~n1690 & pi130;
  assign n1962 = n401 & ~pi130;
  assign n1963 = ~n1961 & ~n1962;
  assign n1964 = ~n1963 & pi133;
  assign n1965 = ~n1960 & ~n1964;
  assign n1966 = ~n1965 & ~pi132;
  assign n1967 = n1699 & pi130;
  assign n1968 = n307 & ~pi130;
  assign n1969 = ~n1967 & ~n1968;
  assign n1970 = n1969 & ~pi133;
  assign n1971 = n1706 & pi130;
  assign n1972 = n353 & ~pi130;
  assign n1973 = ~n1971 & ~n1972;
  assign n1974 = n1973 & pi133;
  assign n1975 = ~n1970 & ~n1974;
  assign n1976 = n1975 & pi132;
  assign n1977 = ~n1966 & ~n1976;
  assign n1978 = n1977 & pi134;
  assign n1979 = n1717 & pi130;
  assign n1980 = n447 & ~pi130;
  assign n1981 = ~n1979 & ~n1980;
  assign n1982 = n1981 & ~pi133;
  assign n1983 = ~n1724 & pi130;
  assign n1984 = n591 & ~pi130;
  assign n1985 = ~n1983 & ~n1984;
  assign n1986 = n1985 & pi133;
  assign n1987 = ~n1982 & ~n1986;
  assign n1988 = n1987 & ~pi132;
  assign n1989 = n1733 & pi130;
  assign n1990 = n497 & ~pi130;
  assign n1991 = ~n1989 & ~n1990;
  assign n1992 = n1991 & ~pi133;
  assign n1993 = n1740 & pi130;
  assign n1994 = n543 & ~pi130;
  assign n1995 = ~n1993 & ~n1994;
  assign n1996 = n1995 & pi133;
  assign n1997 = ~n1992 & ~n1996;
  assign n1998 = n1997 & pi132;
  assign n1999 = ~n1988 & ~n1998;
  assign n2000 = n1999 & ~pi134;
  assign po012 = n1978 | n2000;
  assign n2002 = ~n1752 & pi130;
  assign n2003 = ~n922 & ~pi130;
  assign n2004 = ~n2002 & ~n2003;
  assign n2005 = ~n2004 & ~pi133;
  assign n2006 = ~n1759 & pi130;
  assign n2007 = ~n746 & ~pi130;
  assign n2008 = ~n2006 & ~n2007;
  assign n2009 = ~n2008 & pi133;
  assign n2010 = ~n2005 & ~n2009;
  assign n2011 = ~n2010 & ~pi132;
  assign n2012 = ~n1768 & pi130;
  assign n2013 = ~n676 & ~pi130;
  assign n2014 = ~n2012 & ~n2013;
  assign n2015 = n2014 & ~pi133;
  assign n2016 = ~n1775 & pi130;
  assign n2017 = ~n710 & ~pi130;
  assign n2018 = ~n2016 & ~n2017;
  assign n2019 = n2018 & pi133;
  assign n2020 = ~n2015 & ~n2019;
  assign n2021 = n2020 & pi132;
  assign n2022 = ~n2011 & ~n2021;
  assign n2023 = n2022 & pi134;
  assign n2024 = ~n1786 & pi130;
  assign n2025 = ~n780 & ~pi130;
  assign n2026 = ~n2024 & ~n2025;
  assign n2027 = n2026 & ~pi133;
  assign n2028 = ~n1793 & pi130;
  assign n2029 = ~n888 & ~pi130;
  assign n2030 = ~n2028 & ~n2029;
  assign n2031 = n2030 & pi133;
  assign n2032 = ~n2027 & ~n2031;
  assign n2033 = n2032 & ~pi132;
  assign n2034 = ~n1802 & pi130;
  assign n2035 = ~n818 & ~pi130;
  assign n2036 = ~n2034 & ~n2035;
  assign n2037 = n2036 & ~pi133;
  assign n2038 = ~n1809 & pi130;
  assign n2039 = ~n852 & ~pi130;
  assign n2040 = ~n2038 & ~n2039;
  assign n2041 = n2040 & pi133;
  assign n2042 = ~n2037 & ~n2041;
  assign n2043 = n2042 & pi132;
  assign n2044 = ~n2033 & ~n2043;
  assign n2045 = n2044 & ~pi134;
  assign po013 = n2023 | n2045;
  assign n2047 = ~n1821 & pi130;
  assign n2048 = ~n1207 & ~pi130;
  assign n2049 = ~n2047 & ~n2048;
  assign n2050 = ~n2049 & ~pi133;
  assign n2051 = ~n1828 & pi130;
  assign n2052 = ~n1031 & ~pi130;
  assign n2053 = ~n2051 & ~n2052;
  assign n2054 = ~n2053 & pi133;
  assign n2055 = ~n2050 & ~n2054;
  assign n2056 = ~n2055 & ~pi132;
  assign n2057 = ~n1837 & pi130;
  assign n2058 = ~n961 & ~pi130;
  assign n2059 = ~n2057 & ~n2058;
  assign n2060 = n2059 & ~pi133;
  assign n2061 = ~n1844 & pi130;
  assign n2062 = ~n995 & ~pi130;
  assign n2063 = ~n2061 & ~n2062;
  assign n2064 = n2063 & pi133;
  assign n2065 = ~n2060 & ~n2064;
  assign n2066 = n2065 & pi132;
  assign n2067 = ~n2056 & ~n2066;
  assign n2068 = n2067 & pi134;
  assign n2069 = ~n1855 & pi130;
  assign n2070 = ~n1065 & ~pi130;
  assign n2071 = ~n2069 & ~n2070;
  assign n2072 = n2071 & ~pi133;
  assign n2073 = ~n1862 & pi130;
  assign n2074 = ~n1173 & ~pi130;
  assign n2075 = ~n2073 & ~n2074;
  assign n2076 = n2075 & pi133;
  assign n2077 = ~n2072 & ~n2076;
  assign n2078 = n2077 & ~pi132;
  assign n2079 = ~n1871 & pi130;
  assign n2080 = ~n1103 & ~pi130;
  assign n2081 = ~n2079 & ~n2080;
  assign n2082 = n2081 & ~pi133;
  assign n2083 = ~n1878 & pi130;
  assign n2084 = ~n1137 & ~pi130;
  assign n2085 = ~n2083 & ~n2084;
  assign n2086 = n2085 & pi133;
  assign n2087 = ~n2082 & ~n2086;
  assign n2088 = n2087 & pi132;
  assign n2089 = ~n2078 & ~n2088;
  assign n2090 = n2089 & ~pi134;
  assign po014 = n2068 | n2090;
  assign n2092 = n1890 & pi130;
  assign n2093 = n1396 & ~pi130;
  assign n2094 = ~n2092 & ~n2093;
  assign n2095 = ~n2094 & ~pi133;
  assign n2096 = n1897 & pi130;
  assign n2097 = ~n1280 & ~pi130;
  assign n2098 = ~n2096 & ~n2097;
  assign n2099 = ~n2098 & pi133;
  assign n2100 = ~n2095 & ~n2099;
  assign n2101 = ~n2100 & ~pi132;
  assign n2102 = n1906 & pi130;
  assign n2103 = n1234 & ~pi130;
  assign n2104 = ~n2102 & ~n2103;
  assign n2105 = n2104 & ~pi133;
  assign n2106 = n1913 & pi130;
  assign n2107 = n1256 & ~pi130;
  assign n2108 = ~n2106 & ~n2107;
  assign n2109 = n2108 & pi133;
  assign n2110 = ~n2105 & ~n2109;
  assign n2111 = n2110 & pi132;
  assign n2112 = ~n2101 & ~n2111;
  assign n2113 = n2112 & pi134;
  assign n2114 = n1924 & pi130;
  assign n2115 = n1302 & ~pi130;
  assign n2116 = ~n2114 & ~n2115;
  assign n2117 = n2116 & ~pi133;
  assign n2118 = n1931 & pi130;
  assign n2119 = n1374 & ~pi130;
  assign n2120 = ~n2118 & ~n2119;
  assign n2121 = n2120 & pi133;
  assign n2122 = ~n2117 & ~n2121;
  assign n2123 = n2122 & ~pi132;
  assign n2124 = n1940 & pi130;
  assign n2125 = n1328 & ~pi130;
  assign n2126 = ~n2124 & ~n2125;
  assign n2127 = n2126 & ~pi133;
  assign n2128 = n1947 & pi130;
  assign n2129 = n1350 & ~pi130;
  assign n2130 = ~n2128 & ~n2129;
  assign n2131 = n2130 & pi133;
  assign n2132 = ~n2127 & ~n2131;
  assign n2133 = n2132 & pi132;
  assign n2134 = ~n2123 & ~n2133;
  assign n2135 = n2134 & ~pi134;
  assign po015 = n2113 | n2135;
  assign n2137 = ~n639 & ~pi133;
  assign n2138 = ~n403 & pi133;
  assign n2139 = ~n2137 & ~n2138;
  assign n2140 = ~n2139 & ~pi132;
  assign n2141 = n357 & pi132;
  assign n2142 = ~n2140 & ~n2141;
  assign n2143 = n2142 & pi134;
  assign n2144 = n449 & ~pi133;
  assign n2145 = n593 & pi133;
  assign n2146 = ~n2144 & ~n2145;
  assign n2147 = n2146 & ~pi132;
  assign n2148 = n547 & pi132;
  assign n2149 = ~n2147 & ~n2148;
  assign n2150 = n2149 & ~pi134;
  assign po016 = n2143 | n2150;
  assign n2152 = ~n924 & ~pi133;
  assign n2153 = ~n748 & pi133;
  assign n2154 = ~n2152 & ~n2153;
  assign n2155 = ~n2154 & ~pi132;
  assign n2156 = n714 & pi132;
  assign n2157 = ~n2155 & ~n2156;
  assign n2158 = n2157 & pi134;
  assign n2159 = n782 & ~pi133;
  assign n2160 = n890 & pi133;
  assign n2161 = ~n2159 & ~n2160;
  assign n2162 = n2161 & ~pi132;
  assign n2163 = n856 & pi132;
  assign n2164 = ~n2162 & ~n2163;
  assign n2165 = n2164 & ~pi134;
  assign po017 = n2158 | n2165;
  assign n2167 = ~n1209 & ~pi133;
  assign n2168 = ~n1033 & pi133;
  assign n2169 = ~n2167 & ~n2168;
  assign n2170 = ~n2169 & ~pi132;
  assign n2171 = n999 & pi132;
  assign n2172 = ~n2170 & ~n2171;
  assign n2173 = n2172 & pi134;
  assign n2174 = n1067 & ~pi133;
  assign n2175 = n1175 & pi133;
  assign n2176 = ~n2174 & ~n2175;
  assign n2177 = n2176 & ~pi132;
  assign n2178 = n1141 & pi132;
  assign n2179 = ~n2177 & ~n2178;
  assign n2180 = n2179 & ~pi134;
  assign po018 = n2173 | n2180;
  assign n2182 = ~n1398 & ~pi133;
  assign n2183 = ~n1282 & pi133;
  assign n2184 = ~n2182 & ~n2183;
  assign n2185 = ~n2184 & ~pi132;
  assign n2186 = n1260 & pi132;
  assign n2187 = ~n2185 & ~n2186;
  assign n2188 = n2187 & pi134;
  assign n2189 = n1304 & ~pi133;
  assign n2190 = n1376 & pi133;
  assign n2191 = ~n2189 & ~n2190;
  assign n2192 = n2191 & ~pi132;
  assign n2193 = n1354 & pi132;
  assign n2194 = ~n2192 & ~n2193;
  assign n2195 = n2194 & ~pi134;
  assign po019 = n2188 | n2195;
  assign n2197 = ~n1467 & ~pi133;
  assign n2198 = ~n1426 & pi133;
  assign n2199 = ~n2197 & ~n2198;
  assign n2200 = ~n2199 & ~pi132;
  assign n2201 = ~n1419 & pi132;
  assign n2202 = ~n2200 & ~n2201;
  assign n2203 = n2202 & pi134;
  assign n2204 = ~n1433 & ~pi133;
  assign n2205 = ~n1460 & pi133;
  assign n2206 = ~n2204 & ~n2205;
  assign n2207 = ~n2206 & ~pi132;
  assign n2208 = ~n1453 & pi132;
  assign n2209 = ~n2207 & ~n2208;
  assign n2210 = n2209 & ~pi134;
  assign po020 = n2203 | n2210;
  assign n2212 = ~n1536 & ~pi133;
  assign n2213 = ~n1495 & pi133;
  assign n2214 = ~n2212 & ~n2213;
  assign n2215 = ~n2214 & ~pi132;
  assign n2216 = ~n1488 & pi132;
  assign n2217 = ~n2215 & ~n2216;
  assign n2218 = n2217 & pi134;
  assign n2219 = ~n1502 & ~pi133;
  assign n2220 = ~n1529 & pi133;
  assign n2221 = ~n2219 & ~n2220;
  assign n2222 = ~n2221 & ~pi132;
  assign n2223 = ~n1522 & pi132;
  assign n2224 = ~n2222 & ~n2223;
  assign n2225 = n2224 & ~pi134;
  assign po021 = n2218 | n2225;
  assign n2227 = ~n1605 & ~pi133;
  assign n2228 = ~n1564 & pi133;
  assign n2229 = ~n2227 & ~n2228;
  assign n2230 = ~n2229 & ~pi132;
  assign n2231 = ~n1557 & pi132;
  assign n2232 = ~n2230 & ~n2231;
  assign n2233 = n2232 & pi134;
  assign n2234 = ~n1571 & ~pi133;
  assign n2235 = ~n1598 & pi133;
  assign n2236 = ~n2234 & ~n2235;
  assign n2237 = ~n2236 & ~pi132;
  assign n2238 = ~n1591 & pi132;
  assign n2239 = ~n2237 & ~n2238;
  assign n2240 = n2239 & ~pi134;
  assign po022 = n2233 | n2240;
  assign n2242 = ~n1674 & ~pi133;
  assign n2243 = ~n1633 & pi133;
  assign n2244 = ~n2242 & ~n2243;
  assign n2245 = ~n2244 & ~pi132;
  assign n2246 = ~n1626 & pi132;
  assign n2247 = ~n2245 & ~n2246;
  assign n2248 = n2247 & pi134;
  assign n2249 = ~n1640 & ~pi133;
  assign n2250 = ~n1667 & pi133;
  assign n2251 = ~n2249 & ~n2250;
  assign n2252 = ~n2251 & ~pi132;
  assign n2253 = ~n1660 & pi132;
  assign n2254 = ~n2252 & ~n2253;
  assign n2255 = n2254 & ~pi134;
  assign po023 = n2248 | n2255;
  assign n2257 = ~n1743 & ~pi133;
  assign n2258 = ~n1702 & pi133;
  assign n2259 = ~n2257 & ~n2258;
  assign n2260 = ~n2259 & ~pi132;
  assign n2261 = ~n1695 & pi132;
  assign n2262 = ~n2260 & ~n2261;
  assign n2263 = n2262 & pi134;
  assign n2264 = ~n1709 & ~pi133;
  assign n2265 = ~n1736 & pi133;
  assign n2266 = ~n2264 & ~n2265;
  assign n2267 = ~n2266 & ~pi132;
  assign n2268 = ~n1729 & pi132;
  assign n2269 = ~n2267 & ~n2268;
  assign n2270 = n2269 & ~pi134;
  assign po024 = n2263 | n2270;
  assign n2272 = ~n1812 & ~pi133;
  assign n2273 = ~n1771 & pi133;
  assign n2274 = ~n2272 & ~n2273;
  assign n2275 = ~n2274 & ~pi132;
  assign n2276 = ~n1764 & pi132;
  assign n2277 = ~n2275 & ~n2276;
  assign n2278 = n2277 & pi134;
  assign n2279 = ~n1778 & ~pi133;
  assign n2280 = ~n1805 & pi133;
  assign n2281 = ~n2279 & ~n2280;
  assign n2282 = ~n2281 & ~pi132;
  assign n2283 = ~n1798 & pi132;
  assign n2284 = ~n2282 & ~n2283;
  assign n2285 = n2284 & ~pi134;
  assign po025 = n2278 | n2285;
  assign n2287 = ~n1881 & ~pi133;
  assign n2288 = ~n1840 & pi133;
  assign n2289 = ~n2287 & ~n2288;
  assign n2290 = ~n2289 & ~pi132;
  assign n2291 = ~n1833 & pi132;
  assign n2292 = ~n2290 & ~n2291;
  assign n2293 = n2292 & pi134;
  assign n2294 = ~n1847 & ~pi133;
  assign n2295 = ~n1874 & pi133;
  assign n2296 = ~n2294 & ~n2295;
  assign n2297 = ~n2296 & ~pi132;
  assign n2298 = ~n1867 & pi132;
  assign n2299 = ~n2297 & ~n2298;
  assign n2300 = n2299 & ~pi134;
  assign po026 = n2293 | n2300;
  assign n2302 = ~n1950 & ~pi133;
  assign n2303 = ~n1909 & pi133;
  assign n2304 = ~n2302 & ~n2303;
  assign n2305 = ~n2304 & ~pi132;
  assign n2306 = ~n1902 & pi132;
  assign n2307 = ~n2305 & ~n2306;
  assign n2308 = n2307 & pi134;
  assign n2309 = ~n1916 & ~pi133;
  assign n2310 = ~n1943 & pi133;
  assign n2311 = ~n2309 & ~n2310;
  assign n2312 = ~n2311 & ~pi132;
  assign n2313 = ~n1936 & pi132;
  assign n2314 = ~n2312 & ~n2313;
  assign n2315 = n2314 & ~pi134;
  assign po027 = n2308 | n2315;
  assign n2317 = ~n1995 & ~pi133;
  assign n2318 = ~n1969 & pi133;
  assign n2319 = ~n2317 & ~n2318;
  assign n2320 = ~n2319 & ~pi132;
  assign n2321 = ~n1965 & pi132;
  assign n2322 = ~n2320 & ~n2321;
  assign n2323 = n2322 & pi134;
  assign n2324 = n1973 & ~pi133;
  assign n2325 = n1991 & pi133;
  assign n2326 = ~n2324 & ~n2325;
  assign n2327 = n2326 & ~pi132;
  assign n2328 = n1987 & pi132;
  assign n2329 = ~n2327 & ~n2328;
  assign n2330 = n2329 & ~pi134;
  assign po028 = n2323 | n2330;
  assign n2332 = ~n2040 & ~pi133;
  assign n2333 = ~n2014 & pi133;
  assign n2334 = ~n2332 & ~n2333;
  assign n2335 = ~n2334 & ~pi132;
  assign n2336 = ~n2010 & pi132;
  assign n2337 = ~n2335 & ~n2336;
  assign n2338 = n2337 & pi134;
  assign n2339 = n2018 & ~pi133;
  assign n2340 = n2036 & pi133;
  assign n2341 = ~n2339 & ~n2340;
  assign n2342 = n2341 & ~pi132;
  assign n2343 = n2032 & pi132;
  assign n2344 = ~n2342 & ~n2343;
  assign n2345 = n2344 & ~pi134;
  assign po029 = n2338 | n2345;
  assign n2347 = ~n2085 & ~pi133;
  assign n2348 = ~n2059 & pi133;
  assign n2349 = ~n2347 & ~n2348;
  assign n2350 = ~n2349 & ~pi132;
  assign n2351 = ~n2055 & pi132;
  assign n2352 = ~n2350 & ~n2351;
  assign n2353 = n2352 & pi134;
  assign n2354 = n2063 & ~pi133;
  assign n2355 = n2081 & pi133;
  assign n2356 = ~n2354 & ~n2355;
  assign n2357 = n2356 & ~pi132;
  assign n2358 = n2077 & pi132;
  assign n2359 = ~n2357 & ~n2358;
  assign n2360 = n2359 & ~pi134;
  assign po030 = n2353 | n2360;
  assign n2362 = ~n2130 & ~pi133;
  assign n2363 = ~n2104 & pi133;
  assign n2364 = ~n2362 & ~n2363;
  assign n2365 = ~n2364 & ~pi132;
  assign n2366 = ~n2100 & pi132;
  assign n2367 = ~n2365 & ~n2366;
  assign n2368 = n2367 & pi134;
  assign n2369 = n2108 & ~pi133;
  assign n2370 = n2126 & pi133;
  assign n2371 = ~n2369 & ~n2370;
  assign n2372 = n2371 & ~pi132;
  assign n2373 = n2122 & pi132;
  assign n2374 = ~n2372 & ~n2373;
  assign n2375 = n2374 & ~pi134;
  assign po031 = n2368 | n2375;
  assign n2377 = ~n545 & ~pi133;
  assign n2378 = ~n309 & pi133;
  assign n2379 = ~n2377 & ~n2378;
  assign n2380 = ~n2379 & ~pi132;
  assign n2381 = ~n2139 & pi132;
  assign n2382 = ~n2380 & ~n2381;
  assign n2383 = n2382 & pi134;
  assign n2384 = n355 & ~pi133;
  assign n2385 = n499 & pi133;
  assign n2386 = ~n2384 & ~n2385;
  assign n2387 = n2386 & ~pi132;
  assign n2388 = n2146 & pi132;
  assign n2389 = ~n2387 & ~n2388;
  assign n2390 = n2389 & ~pi134;
  assign po032 = n2383 | n2390;
  assign n2392 = ~n854 & ~pi133;
  assign n2393 = ~n678 & pi133;
  assign n2394 = ~n2392 & ~n2393;
  assign n2395 = ~n2394 & ~pi132;
  assign n2396 = ~n2154 & pi132;
  assign n2397 = ~n2395 & ~n2396;
  assign n2398 = n2397 & pi134;
  assign n2399 = n712 & ~pi133;
  assign n2400 = n820 & pi133;
  assign n2401 = ~n2399 & ~n2400;
  assign n2402 = n2401 & ~pi132;
  assign n2403 = n2161 & pi132;
  assign n2404 = ~n2402 & ~n2403;
  assign n2405 = n2404 & ~pi134;
  assign po033 = n2398 | n2405;
  assign n2407 = ~n1139 & ~pi133;
  assign n2408 = ~n963 & pi133;
  assign n2409 = ~n2407 & ~n2408;
  assign n2410 = ~n2409 & ~pi132;
  assign n2411 = ~n2169 & pi132;
  assign n2412 = ~n2410 & ~n2411;
  assign n2413 = n2412 & pi134;
  assign n2414 = n997 & ~pi133;
  assign n2415 = n1105 & pi133;
  assign n2416 = ~n2414 & ~n2415;
  assign n2417 = n2416 & ~pi132;
  assign n2418 = n2176 & pi132;
  assign n2419 = ~n2417 & ~n2418;
  assign n2420 = n2419 & ~pi134;
  assign po034 = n2413 | n2420;
  assign n2422 = ~n1352 & ~pi133;
  assign n2423 = ~n1236 & pi133;
  assign n2424 = ~n2422 & ~n2423;
  assign n2425 = ~n2424 & ~pi132;
  assign n2426 = ~n2184 & pi132;
  assign n2427 = ~n2425 & ~n2426;
  assign n2428 = n2427 & pi134;
  assign n2429 = n1258 & ~pi133;
  assign n2430 = n1330 & pi133;
  assign n2431 = ~n2429 & ~n2430;
  assign n2432 = n2431 & ~pi132;
  assign n2433 = n2191 & pi132;
  assign n2434 = ~n2432 & ~n2433;
  assign n2435 = n2434 & ~pi134;
  assign po035 = n2428 | n2435;
  assign n2437 = ~n1451 & ~pi133;
  assign n2438 = ~n1410 & pi133;
  assign n2439 = ~n2437 & ~n2438;
  assign n2440 = ~n2439 & ~pi132;
  assign n2441 = ~n2199 & pi132;
  assign n2442 = ~n2440 & ~n2441;
  assign n2443 = n2442 & pi134;
  assign n2444 = ~n1417 & ~pi133;
  assign n2445 = ~n1444 & pi133;
  assign n2446 = ~n2444 & ~n2445;
  assign n2447 = ~n2446 & ~pi132;
  assign n2448 = ~n2206 & pi132;
  assign n2449 = ~n2447 & ~n2448;
  assign n2450 = n2449 & ~pi134;
  assign po036 = n2443 | n2450;
  assign n2452 = ~n1520 & ~pi133;
  assign n2453 = ~n1479 & pi133;
  assign n2454 = ~n2452 & ~n2453;
  assign n2455 = ~n2454 & ~pi132;
  assign n2456 = ~n2214 & pi132;
  assign n2457 = ~n2455 & ~n2456;
  assign n2458 = n2457 & pi134;
  assign n2459 = ~n1486 & ~pi133;
  assign n2460 = ~n1513 & pi133;
  assign n2461 = ~n2459 & ~n2460;
  assign n2462 = ~n2461 & ~pi132;
  assign n2463 = ~n2221 & pi132;
  assign n2464 = ~n2462 & ~n2463;
  assign n2465 = n2464 & ~pi134;
  assign po037 = n2458 | n2465;
  assign n2467 = ~n1589 & ~pi133;
  assign n2468 = ~n1548 & pi133;
  assign n2469 = ~n2467 & ~n2468;
  assign n2470 = ~n2469 & ~pi132;
  assign n2471 = ~n2229 & pi132;
  assign n2472 = ~n2470 & ~n2471;
  assign n2473 = n2472 & pi134;
  assign n2474 = ~n1555 & ~pi133;
  assign n2475 = ~n1582 & pi133;
  assign n2476 = ~n2474 & ~n2475;
  assign n2477 = ~n2476 & ~pi132;
  assign n2478 = ~n2236 & pi132;
  assign n2479 = ~n2477 & ~n2478;
  assign n2480 = n2479 & ~pi134;
  assign po038 = n2473 | n2480;
  assign n2482 = ~n1658 & ~pi133;
  assign n2483 = ~n1617 & pi133;
  assign n2484 = ~n2482 & ~n2483;
  assign n2485 = ~n2484 & ~pi132;
  assign n2486 = ~n2244 & pi132;
  assign n2487 = ~n2485 & ~n2486;
  assign n2488 = n2487 & pi134;
  assign n2489 = ~n1624 & ~pi133;
  assign n2490 = ~n1651 & pi133;
  assign n2491 = ~n2489 & ~n2490;
  assign n2492 = ~n2491 & ~pi132;
  assign n2493 = ~n2251 & pi132;
  assign n2494 = ~n2492 & ~n2493;
  assign n2495 = n2494 & ~pi134;
  assign po039 = n2488 | n2495;
  assign n2497 = ~n1727 & ~pi133;
  assign n2498 = ~n1686 & pi133;
  assign n2499 = ~n2497 & ~n2498;
  assign n2500 = ~n2499 & ~pi132;
  assign n2501 = ~n2259 & pi132;
  assign n2502 = ~n2500 & ~n2501;
  assign n2503 = n2502 & pi134;
  assign n2504 = ~n1693 & ~pi133;
  assign n2505 = ~n1720 & pi133;
  assign n2506 = ~n2504 & ~n2505;
  assign n2507 = ~n2506 & ~pi132;
  assign n2508 = ~n2266 & pi132;
  assign n2509 = ~n2507 & ~n2508;
  assign n2510 = n2509 & ~pi134;
  assign po040 = n2503 | n2510;
  assign n2512 = ~n1796 & ~pi133;
  assign n2513 = ~n1755 & pi133;
  assign n2514 = ~n2512 & ~n2513;
  assign n2515 = ~n2514 & ~pi132;
  assign n2516 = ~n2274 & pi132;
  assign n2517 = ~n2515 & ~n2516;
  assign n2518 = n2517 & pi134;
  assign n2519 = ~n1762 & ~pi133;
  assign n2520 = ~n1789 & pi133;
  assign n2521 = ~n2519 & ~n2520;
  assign n2522 = ~n2521 & ~pi132;
  assign n2523 = ~n2281 & pi132;
  assign n2524 = ~n2522 & ~n2523;
  assign n2525 = n2524 & ~pi134;
  assign po041 = n2518 | n2525;
  assign n2527 = ~n1865 & ~pi133;
  assign n2528 = ~n1824 & pi133;
  assign n2529 = ~n2527 & ~n2528;
  assign n2530 = ~n2529 & ~pi132;
  assign n2531 = ~n2289 & pi132;
  assign n2532 = ~n2530 & ~n2531;
  assign n2533 = n2532 & pi134;
  assign n2534 = ~n1831 & ~pi133;
  assign n2535 = ~n1858 & pi133;
  assign n2536 = ~n2534 & ~n2535;
  assign n2537 = ~n2536 & ~pi132;
  assign n2538 = ~n2296 & pi132;
  assign n2539 = ~n2537 & ~n2538;
  assign n2540 = n2539 & ~pi134;
  assign po042 = n2533 | n2540;
  assign n2542 = ~n1934 & ~pi133;
  assign n2543 = ~n1893 & pi133;
  assign n2544 = ~n2542 & ~n2543;
  assign n2545 = ~n2544 & ~pi132;
  assign n2546 = ~n2304 & pi132;
  assign n2547 = ~n2545 & ~n2546;
  assign n2548 = n2547 & pi134;
  assign n2549 = ~n1900 & ~pi133;
  assign n2550 = ~n1927 & pi133;
  assign n2551 = ~n2549 & ~n2550;
  assign n2552 = ~n2551 & ~pi132;
  assign n2553 = ~n2311 & pi132;
  assign n2554 = ~n2552 & ~n2553;
  assign n2555 = n2554 & ~pi134;
  assign po043 = n2548 | n2555;
  assign n2557 = n1959 & pi133;
  assign n2558 = n1985 & ~pi133;
  assign n2559 = ~n2557 & ~n2558;
  assign n2560 = n2559 & ~pi132;
  assign n2561 = ~n2319 & pi132;
  assign n2562 = ~n2560 & ~n2561;
  assign n2563 = n2562 & pi134;
  assign n2564 = n1963 & ~pi133;
  assign n2565 = n1981 & pi133;
  assign n2566 = ~n2564 & ~n2565;
  assign n2567 = n2566 & ~pi132;
  assign n2568 = n2326 & pi132;
  assign n2569 = ~n2567 & ~n2568;
  assign n2570 = n2569 & ~pi134;
  assign po044 = n2563 | n2570;
  assign n2572 = n2004 & pi133;
  assign n2573 = n2030 & ~pi133;
  assign n2574 = ~n2572 & ~n2573;
  assign n2575 = n2574 & ~pi132;
  assign n2576 = ~n2334 & pi132;
  assign n2577 = ~n2575 & ~n2576;
  assign n2578 = n2577 & pi134;
  assign n2579 = n2008 & ~pi133;
  assign n2580 = n2026 & pi133;
  assign n2581 = ~n2579 & ~n2580;
  assign n2582 = n2581 & ~pi132;
  assign n2583 = n2341 & pi132;
  assign n2584 = ~n2582 & ~n2583;
  assign n2585 = n2584 & ~pi134;
  assign po045 = n2578 | n2585;
  assign n2587 = n2049 & pi133;
  assign n2588 = n2075 & ~pi133;
  assign n2589 = ~n2587 & ~n2588;
  assign n2590 = n2589 & ~pi132;
  assign n2591 = ~n2349 & pi132;
  assign n2592 = ~n2590 & ~n2591;
  assign n2593 = n2592 & pi134;
  assign n2594 = n2053 & ~pi133;
  assign n2595 = n2071 & pi133;
  assign n2596 = ~n2594 & ~n2595;
  assign n2597 = n2596 & ~pi132;
  assign n2598 = n2356 & pi132;
  assign n2599 = ~n2597 & ~n2598;
  assign n2600 = n2599 & ~pi134;
  assign po046 = n2593 | n2600;
  assign n2602 = n2094 & pi133;
  assign n2603 = n2120 & ~pi133;
  assign n2604 = ~n2602 & ~n2603;
  assign n2605 = n2604 & ~pi132;
  assign n2606 = ~n2364 & pi132;
  assign n2607 = ~n2605 & ~n2606;
  assign n2608 = n2607 & pi134;
  assign n2609 = n2098 & ~pi133;
  assign n2610 = n2116 & pi133;
  assign n2611 = ~n2609 & ~n2610;
  assign n2612 = n2611 & ~pi132;
  assign n2613 = n2371 & pi132;
  assign n2614 = ~n2612 & ~n2613;
  assign n2615 = n2614 & ~pi134;
  assign po047 = n2608 | n2615;
  assign n2617 = ~n2379 & pi132;
  assign n2618 = n641 & ~pi132;
  assign n2619 = ~n2617 & ~n2618;
  assign n2620 = n2619 & pi134;
  assign n2621 = n2386 & pi132;
  assign n2622 = n451 & ~pi132;
  assign n2623 = ~n2621 & ~n2622;
  assign n2624 = n2623 & ~pi134;
  assign po048 = n2620 | n2624;
  assign n2626 = ~n2394 & pi132;
  assign n2627 = n926 & ~pi132;
  assign n2628 = ~n2626 & ~n2627;
  assign n2629 = n2628 & pi134;
  assign n2630 = n2401 & pi132;
  assign n2631 = n784 & ~pi132;
  assign n2632 = ~n2630 & ~n2631;
  assign n2633 = n2632 & ~pi134;
  assign po049 = n2629 | n2633;
  assign n2635 = ~n2409 & pi132;
  assign n2636 = n1211 & ~pi132;
  assign n2637 = ~n2635 & ~n2636;
  assign n2638 = n2637 & pi134;
  assign n2639 = n2416 & pi132;
  assign n2640 = n1069 & ~pi132;
  assign n2641 = ~n2639 & ~n2640;
  assign n2642 = n2641 & ~pi134;
  assign po050 = n2638 | n2642;
  assign n2644 = ~n2424 & pi132;
  assign n2645 = n1400 & ~pi132;
  assign n2646 = ~n2644 & ~n2645;
  assign n2647 = n2646 & pi134;
  assign n2648 = n2431 & pi132;
  assign n2649 = n1306 & ~pi132;
  assign n2650 = ~n2648 & ~n2649;
  assign n2651 = n2650 & ~pi134;
  assign po051 = n2647 | n2651;
  assign n2653 = ~n2439 & pi132;
  assign n2654 = ~n1469 & ~pi132;
  assign n2655 = ~n2653 & ~n2654;
  assign n2656 = n2655 & pi134;
  assign n2657 = ~n2446 & pi132;
  assign n2658 = ~n1435 & ~pi132;
  assign n2659 = ~n2657 & ~n2658;
  assign n2660 = n2659 & ~pi134;
  assign po052 = n2656 | n2660;
  assign n2662 = ~n2454 & pi132;
  assign n2663 = ~n1538 & ~pi132;
  assign n2664 = ~n2662 & ~n2663;
  assign n2665 = n2664 & pi134;
  assign n2666 = ~n2461 & pi132;
  assign n2667 = ~n1504 & ~pi132;
  assign n2668 = ~n2666 & ~n2667;
  assign n2669 = n2668 & ~pi134;
  assign po053 = n2665 | n2669;
  assign n2671 = ~n2469 & pi132;
  assign n2672 = ~n1607 & ~pi132;
  assign n2673 = ~n2671 & ~n2672;
  assign n2674 = n2673 & pi134;
  assign n2675 = ~n2476 & pi132;
  assign n2676 = ~n1573 & ~pi132;
  assign n2677 = ~n2675 & ~n2676;
  assign n2678 = n2677 & ~pi134;
  assign po054 = n2674 | n2678;
  assign n2680 = ~n2484 & pi132;
  assign n2681 = ~n1676 & ~pi132;
  assign n2682 = ~n2680 & ~n2681;
  assign n2683 = n2682 & pi134;
  assign n2684 = ~n2491 & pi132;
  assign n2685 = ~n1642 & ~pi132;
  assign n2686 = ~n2684 & ~n2685;
  assign n2687 = n2686 & ~pi134;
  assign po055 = n2683 | n2687;
  assign n2689 = ~n2499 & pi132;
  assign n2690 = ~n1745 & ~pi132;
  assign n2691 = ~n2689 & ~n2690;
  assign n2692 = n2691 & pi134;
  assign n2693 = ~n2506 & pi132;
  assign n2694 = ~n1711 & ~pi132;
  assign n2695 = ~n2693 & ~n2694;
  assign n2696 = n2695 & ~pi134;
  assign po056 = n2692 | n2696;
  assign n2698 = ~n2514 & pi132;
  assign n2699 = ~n1814 & ~pi132;
  assign n2700 = ~n2698 & ~n2699;
  assign n2701 = n2700 & pi134;
  assign n2702 = ~n2521 & pi132;
  assign n2703 = ~n1780 & ~pi132;
  assign n2704 = ~n2702 & ~n2703;
  assign n2705 = n2704 & ~pi134;
  assign po057 = n2701 | n2705;
  assign n2707 = ~n2529 & pi132;
  assign n2708 = ~n1883 & ~pi132;
  assign n2709 = ~n2707 & ~n2708;
  assign n2710 = n2709 & pi134;
  assign n2711 = ~n2536 & pi132;
  assign n2712 = ~n1849 & ~pi132;
  assign n2713 = ~n2711 & ~n2712;
  assign n2714 = n2713 & ~pi134;
  assign po058 = n2710 | n2714;
  assign n2716 = ~n2544 & pi132;
  assign n2717 = ~n1952 & ~pi132;
  assign n2718 = ~n2716 & ~n2717;
  assign n2719 = n2718 & pi134;
  assign n2720 = ~n2551 & pi132;
  assign n2721 = ~n1918 & ~pi132;
  assign n2722 = ~n2720 & ~n2721;
  assign n2723 = n2722 & ~pi134;
  assign po059 = n2719 | n2723;
  assign n2725 = n2559 & pi132;
  assign n2726 = n1997 & ~pi132;
  assign n2727 = ~n2725 & ~n2726;
  assign n2728 = n2727 & pi134;
  assign n2729 = n2566 & pi132;
  assign n2730 = n1975 & ~pi132;
  assign n2731 = ~n2729 & ~n2730;
  assign n2732 = n2731 & ~pi134;
  assign po060 = n2728 | n2732;
  assign n2734 = n2574 & pi132;
  assign n2735 = n2042 & ~pi132;
  assign n2736 = ~n2734 & ~n2735;
  assign n2737 = n2736 & pi134;
  assign n2738 = n2581 & pi132;
  assign n2739 = n2020 & ~pi132;
  assign n2740 = ~n2738 & ~n2739;
  assign n2741 = n2740 & ~pi134;
  assign po061 = n2737 | n2741;
  assign n2743 = n2589 & pi132;
  assign n2744 = n2087 & ~pi132;
  assign n2745 = ~n2743 & ~n2744;
  assign n2746 = n2745 & pi134;
  assign n2747 = n2596 & pi132;
  assign n2748 = n2065 & ~pi132;
  assign n2749 = ~n2747 & ~n2748;
  assign n2750 = n2749 & ~pi134;
  assign po062 = n2746 | n2750;
  assign n2752 = n2604 & pi132;
  assign n2753 = n2132 & ~pi132;
  assign n2754 = ~n2752 & ~n2753;
  assign n2755 = n2754 & pi134;
  assign n2756 = n2611 & pi132;
  assign n2757 = n2110 & ~pi132;
  assign n2758 = ~n2756 & ~n2757;
  assign n2759 = n2758 & ~pi134;
  assign po063 = n2755 | n2759;
  assign n2761 = n453 & ~pi134;
  assign n2762 = n643 & pi134;
  assign po064 = n2761 | n2762;
  assign n2764 = n786 & ~pi134;
  assign n2765 = n928 & pi134;
  assign po065 = n2764 | n2765;
  assign n2767 = n1071 & ~pi134;
  assign n2768 = n1213 & pi134;
  assign po066 = n2767 | n2768;
  assign n2770 = n1308 & ~pi134;
  assign n2771 = n1402 & pi134;
  assign po067 = n2770 | n2771;
  assign n2773 = n1437 & ~pi134;
  assign n2774 = n1471 & pi134;
  assign po068 = n2773 | n2774;
  assign n2776 = n1506 & ~pi134;
  assign n2777 = n1540 & pi134;
  assign po069 = n2776 | n2777;
  assign n2779 = n1575 & ~pi134;
  assign n2780 = n1609 & pi134;
  assign po070 = n2779 | n2780;
  assign n2782 = n1644 & ~pi134;
  assign n2783 = n1678 & pi134;
  assign po071 = n2782 | n2783;
  assign n2785 = n1713 & ~pi134;
  assign n2786 = n1747 & pi134;
  assign po072 = n2785 | n2786;
  assign n2788 = n1782 & ~pi134;
  assign n2789 = n1816 & pi134;
  assign po073 = n2788 | n2789;
  assign n2791 = n1851 & ~pi134;
  assign n2792 = n1885 & pi134;
  assign po074 = n2791 | n2792;
  assign n2794 = n1920 & ~pi134;
  assign n2795 = n1954 & pi134;
  assign po075 = n2794 | n2795;
  assign n2797 = n1977 & ~pi134;
  assign n2798 = n1999 & pi134;
  assign po076 = n2797 | n2798;
  assign n2800 = n2022 & ~pi134;
  assign n2801 = n2044 & pi134;
  assign po077 = n2800 | n2801;
  assign n2803 = n2067 & ~pi134;
  assign n2804 = n2089 & pi134;
  assign po078 = n2803 | n2804;
  assign n2806 = n2112 & ~pi134;
  assign n2807 = n2134 & pi134;
  assign po079 = n2806 | n2807;
  assign n2809 = n2142 & ~pi134;
  assign n2810 = n2149 & pi134;
  assign po080 = n2809 | n2810;
  assign n2812 = n2157 & ~pi134;
  assign n2813 = n2164 & pi134;
  assign po081 = n2812 | n2813;
  assign n2815 = n2172 & ~pi134;
  assign n2816 = n2179 & pi134;
  assign po082 = n2815 | n2816;
  assign n2818 = n2187 & ~pi134;
  assign n2819 = n2194 & pi134;
  assign po083 = n2818 | n2819;
  assign n2821 = n2202 & ~pi134;
  assign n2822 = n2209 & pi134;
  assign po084 = n2821 | n2822;
  assign n2824 = n2217 & ~pi134;
  assign n2825 = n2224 & pi134;
  assign po085 = n2824 | n2825;
  assign n2827 = n2232 & ~pi134;
  assign n2828 = n2239 & pi134;
  assign po086 = n2827 | n2828;
  assign n2830 = n2247 & ~pi134;
  assign n2831 = n2254 & pi134;
  assign po087 = n2830 | n2831;
  assign n2833 = n2262 & ~pi134;
  assign n2834 = n2269 & pi134;
  assign po088 = n2833 | n2834;
  assign n2836 = n2277 & ~pi134;
  assign n2837 = n2284 & pi134;
  assign po089 = n2836 | n2837;
  assign n2839 = n2292 & ~pi134;
  assign n2840 = n2299 & pi134;
  assign po090 = n2839 | n2840;
  assign n2842 = n2307 & ~pi134;
  assign n2843 = n2314 & pi134;
  assign po091 = n2842 | n2843;
  assign n2845 = n2322 & ~pi134;
  assign n2846 = n2329 & pi134;
  assign po092 = n2845 | n2846;
  assign n2848 = n2337 & ~pi134;
  assign n2849 = n2344 & pi134;
  assign po093 = n2848 | n2849;
  assign n2851 = n2352 & ~pi134;
  assign n2852 = n2359 & pi134;
  assign po094 = n2851 | n2852;
  assign n2854 = n2367 & ~pi134;
  assign n2855 = n2374 & pi134;
  assign po095 = n2854 | n2855;
  assign n2857 = n2382 & ~pi134;
  assign n2858 = n2389 & pi134;
  assign po096 = n2857 | n2858;
  assign n2860 = n2397 & ~pi134;
  assign n2861 = n2404 & pi134;
  assign po097 = n2860 | n2861;
  assign n2863 = n2412 & ~pi134;
  assign n2864 = n2419 & pi134;
  assign po098 = n2863 | n2864;
  assign n2866 = n2427 & ~pi134;
  assign n2867 = n2434 & pi134;
  assign po099 = n2866 | n2867;
  assign n2869 = n2442 & ~pi134;
  assign n2870 = n2449 & pi134;
  assign po100 = n2869 | n2870;
  assign n2872 = n2457 & ~pi134;
  assign n2873 = n2464 & pi134;
  assign po101 = n2872 | n2873;
  assign n2875 = n2472 & ~pi134;
  assign n2876 = n2479 & pi134;
  assign po102 = n2875 | n2876;
  assign n2878 = n2487 & ~pi134;
  assign n2879 = n2494 & pi134;
  assign po103 = n2878 | n2879;
  assign n2881 = n2502 & ~pi134;
  assign n2882 = n2509 & pi134;
  assign po104 = n2881 | n2882;
  assign n2884 = n2517 & ~pi134;
  assign n2885 = n2524 & pi134;
  assign po105 = n2884 | n2885;
  assign n2887 = n2532 & ~pi134;
  assign n2888 = n2539 & pi134;
  assign po106 = n2887 | n2888;
  assign n2890 = n2547 & ~pi134;
  assign n2891 = n2554 & pi134;
  assign po107 = n2890 | n2891;
  assign n2893 = n2562 & ~pi134;
  assign n2894 = n2569 & pi134;
  assign po108 = n2893 | n2894;
  assign n2896 = n2577 & ~pi134;
  assign n2897 = n2584 & pi134;
  assign po109 = n2896 | n2897;
  assign n2899 = n2592 & ~pi134;
  assign n2900 = n2599 & pi134;
  assign po110 = n2899 | n2900;
  assign n2902 = n2607 & ~pi134;
  assign n2903 = n2614 & pi134;
  assign po111 = n2902 | n2903;
  assign n2905 = n2619 & ~pi134;
  assign n2906 = n2623 & pi134;
  assign po112 = n2905 | n2906;
  assign n2908 = n2628 & ~pi134;
  assign n2909 = n2632 & pi134;
  assign po113 = n2908 | n2909;
  assign n2911 = n2637 & ~pi134;
  assign n2912 = n2641 & pi134;
  assign po114 = n2911 | n2912;
  assign n2914 = n2646 & ~pi134;
  assign n2915 = n2650 & pi134;
  assign po115 = n2914 | n2915;
  assign n2917 = n2655 & ~pi134;
  assign n2918 = n2659 & pi134;
  assign po116 = n2917 | n2918;
  assign n2920 = n2664 & ~pi134;
  assign n2921 = n2668 & pi134;
  assign po117 = n2920 | n2921;
  assign n2923 = n2673 & ~pi134;
  assign n2924 = n2677 & pi134;
  assign po118 = n2923 | n2924;
  assign n2926 = n2682 & ~pi134;
  assign n2927 = n2686 & pi134;
  assign po119 = n2926 | n2927;
  assign n2929 = n2691 & ~pi134;
  assign n2930 = n2695 & pi134;
  assign po120 = n2929 | n2930;
  assign n2932 = n2700 & ~pi134;
  assign n2933 = n2704 & pi134;
  assign po121 = n2932 | n2933;
  assign n2935 = n2709 & ~pi134;
  assign n2936 = n2713 & pi134;
  assign po122 = n2935 | n2936;
  assign n2938 = n2718 & ~pi134;
  assign n2939 = n2722 & pi134;
  assign po123 = n2938 | n2939;
  assign n2941 = n2727 & ~pi134;
  assign n2942 = n2731 & pi134;
  assign po124 = n2941 | n2942;
  assign n2944 = n2736 & ~pi134;
  assign n2945 = n2740 & pi134;
  assign po125 = n2944 | n2945;
  assign n2947 = n2745 & ~pi134;
  assign n2948 = n2749 & pi134;
  assign po126 = n2947 | n2948;
  assign n2950 = n2754 & ~pi134;
  assign n2951 = n2758 & pi134;
  assign po127 = n2950 | n2951;
endmodule


