module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127;
  wire n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833;
  assign n129 = x0 & x64;
  assign n131 = x0 & x65;
  assign n130 = x1 & x64;
  assign n132 = n131 ^ n130;
  assign n133 = x66 ^ x2;
  assign n134 = n129 & ~n133;
  assign n140 = x2 & x64;
  assign n139 = ~x64 & x66;
  assign n141 = n140 ^ n139;
  assign n142 = ~x0 & n141;
  assign n143 = n142 ^ n139;
  assign n135 = x1 & x65;
  assign n136 = x64 & ~n135;
  assign n137 = x0 & n136;
  assign n138 = n137 ^ n135;
  assign n144 = n143 ^ n138;
  assign n145 = ~n134 & n144;
  assign n159 = x64 & x65;
  assign n160 = ~x66 & ~n159;
  assign n161 = x65 & x66;
  assign n162 = ~n160 & ~n161;
  assign n163 = x2 ^ x1;
  assign n164 = ~n162 & n163;
  assign n165 = n164 ^ x1;
  assign n166 = n165 ^ x67;
  assign n155 = x1 & n133;
  assign n156 = ~x1 & x2;
  assign n157 = ~x65 & n156;
  assign n158 = ~n155 & ~n157;
  assign n167 = n166 ^ n158;
  assign n168 = ~x0 & ~n167;
  assign n169 = n168 ^ n166;
  assign n146 = x3 & x64;
  assign n147 = n146 ^ x2;
  assign n148 = ~x0 & ~n135;
  assign n149 = ~x64 & x65;
  assign n150 = ~n139 & ~n149;
  assign n151 = ~n148 & ~n150;
  assign n152 = ~n146 & n151;
  assign n153 = n147 & n152;
  assign n154 = n153 ^ n147;
  assign n170 = n169 ^ n154;
  assign n180 = x67 & ~n160;
  assign n181 = ~x67 & ~n161;
  assign n182 = ~n180 & ~n181;
  assign n183 = n163 & ~n182;
  assign n184 = n183 ^ x1;
  assign n185 = n184 ^ x68;
  assign n186 = x0 & ~n185;
  assign n187 = ~x66 & n156;
  assign n188 = ~x0 & ~n187;
  assign n189 = x67 ^ x2;
  assign n190 = x1 & n189;
  assign n191 = n188 & ~n190;
  assign n192 = ~n186 & ~n191;
  assign n172 = x3 ^ x2;
  assign n173 = x65 ^ x3;
  assign n174 = n172 & ~n173;
  assign n175 = n174 ^ x2;
  assign n176 = n175 ^ x4;
  assign n177 = x64 & n176;
  assign n178 = n149 & n172;
  assign n179 = ~n177 & ~n178;
  assign n193 = n192 ^ n179;
  assign n171 = n154 & n169;
  assign n194 = n193 ^ n171;
  assign n227 = ~x68 & ~n180;
  assign n228 = x68 & ~n181;
  assign n229 = ~n227 & ~n228;
  assign n230 = n163 & ~n229;
  assign n231 = n230 ^ x1;
  assign n232 = n231 ^ x69;
  assign n233 = x0 & n232;
  assign n234 = ~x1 & x67;
  assign n235 = ~x0 & ~n234;
  assign n236 = x1 & x68;
  assign n237 = n236 ^ x2;
  assign n238 = n235 & n237;
  assign n239 = ~n233 & ~n238;
  assign n208 = ~x64 & ~x66;
  assign n209 = x5 ^ x4;
  assign n210 = n172 & n209;
  assign n211 = n208 & n210;
  assign n203 = x2 & x3;
  assign n198 = ~x2 & ~x3;
  assign n212 = n203 ^ n198;
  assign n213 = x4 & n212;
  assign n214 = n213 ^ n203;
  assign n215 = ~n211 & ~n214;
  assign n216 = x65 & ~n215;
  assign n217 = x4 ^ x3;
  assign n218 = n209 & ~n217;
  assign n219 = ~n172 & n218;
  assign n220 = x64 & n219;
  assign n221 = n149 & n209;
  assign n222 = x66 & n172;
  assign n223 = ~n221 & n222;
  assign n224 = ~n220 & ~n223;
  assign n225 = ~n216 & n224;
  assign n199 = x4 & x64;
  assign n200 = n198 & ~n199;
  assign n201 = ~x64 & ~x65;
  assign n202 = ~n200 & ~n201;
  assign n204 = ~x4 & x64;
  assign n205 = n203 & ~n204;
  assign n206 = n202 & ~n205;
  assign n207 = x5 & n206;
  assign n226 = n225 ^ n207;
  assign n240 = n239 ^ n226;
  assign n195 = n179 ^ n171;
  assign n196 = ~n193 & n195;
  assign n197 = n196 ^ n192;
  assign n241 = n240 ^ n197;
  assign n258 = x66 & n214;
  assign n259 = n172 & ~n209;
  assign n260 = x67 & n259;
  assign n261 = ~n258 & ~n260;
  assign n262 = x65 & n219;
  assign n263 = n261 & ~n262;
  assign n264 = n162 ^ x67;
  assign n265 = n210 & n264;
  assign n266 = n263 & ~n265;
  assign n267 = n266 ^ x5;
  assign n268 = x6 ^ x5;
  assign n269 = n267 & n268;
  assign n270 = x5 & ~n206;
  assign n271 = n225 & n270;
  assign n272 = ~x6 & n271;
  assign n273 = ~n269 & ~n272;
  assign n274 = x64 & ~n273;
  assign n275 = x64 & n268;
  assign n276 = ~n271 & ~n275;
  assign n277 = n276 ^ n271;
  assign n278 = ~n267 & n277;
  assign n279 = n278 ^ n271;
  assign n280 = ~n274 & ~n279;
  assign n245 = x69 & ~n227;
  assign n246 = ~x69 & ~n228;
  assign n247 = ~n245 & ~n246;
  assign n248 = n163 & ~n247;
  assign n249 = n248 ^ x1;
  assign n250 = n249 ^ x70;
  assign n251 = x0 & ~n250;
  assign n252 = x69 ^ x2;
  assign n253 = x1 & n252;
  assign n254 = ~x0 & ~n253;
  assign n255 = ~x68 & n156;
  assign n256 = n254 & ~n255;
  assign n257 = ~n251 & ~n256;
  assign n281 = n280 ^ n257;
  assign n242 = n239 ^ n197;
  assign n243 = ~n240 & ~n242;
  assign n244 = n243 ^ n197;
  assign n282 = n281 ^ n244;
  assign n337 = ~n267 & ~n276;
  assign n300 = n182 ^ x68;
  assign n301 = n210 & n300;
  assign n302 = x67 & n214;
  assign n303 = x66 & n219;
  assign n304 = ~n302 & ~n303;
  assign n305 = x68 & n259;
  assign n306 = n304 & ~n305;
  assign n307 = ~n301 & n306;
  assign n308 = ~x5 & ~n307;
  assign n310 = ~x5 & ~x6;
  assign n311 = x65 & ~n310;
  assign n309 = x7 & x64;
  assign n312 = n311 ^ n309;
  assign n313 = n308 & n312;
  assign n314 = x5 & x6;
  assign n315 = ~x7 & n314;
  assign n316 = x5 & ~x6;
  assign n317 = x7 & ~x65;
  assign n318 = n316 & n317;
  assign n319 = ~n315 & ~n318;
  assign n320 = n307 & ~n319;
  assign n321 = ~n313 & ~n320;
  assign n322 = x64 & ~n321;
  assign n323 = x6 & n307;
  assign n324 = x65 & ~n309;
  assign n325 = ~n323 & n324;
  assign n326 = ~x5 & x6;
  assign n327 = ~n307 & ~n326;
  assign n328 = n325 & ~n327;
  assign n329 = ~n322 & ~n328;
  assign n330 = n307 ^ x5;
  assign n331 = ~x7 & x64;
  assign n332 = n331 ^ n312;
  assign n333 = n314 & n332;
  assign n334 = n333 ^ n312;
  assign n335 = n330 & ~n334;
  assign n336 = n329 & ~n335;
  assign n338 = n337 ^ n336;
  assign n291 = ~x70 & ~n245;
  assign n292 = x70 & ~n246;
  assign n293 = ~n291 & ~n292;
  assign n294 = n163 & ~n293;
  assign n295 = n294 ^ x1;
  assign n296 = n295 ^ x71;
  assign n287 = x2 & ~x69;
  assign n286 = x70 ^ x2;
  assign n288 = n287 ^ n286;
  assign n289 = x1 & n288;
  assign n290 = n289 ^ n287;
  assign n297 = n296 ^ n290;
  assign n298 = ~x0 & n297;
  assign n299 = n298 ^ n296;
  assign n339 = n338 ^ n299;
  assign n283 = n280 ^ n244;
  assign n284 = n281 & ~n283;
  assign n285 = n284 ^ n244;
  assign n340 = n339 ^ n285;
  assign n371 = x8 ^ x7;
  assign n372 = n268 & n371;
  assign n373 = n208 & n372;
  assign n374 = n314 ^ n310;
  assign n375 = ~x7 & n374;
  assign n376 = n375 ^ n310;
  assign n377 = ~n373 & ~n376;
  assign n378 = x65 & ~n377;
  assign n379 = n149 & n371;
  assign n380 = x66 & n268;
  assign n381 = ~n379 & n380;
  assign n382 = ~n378 & ~n381;
  assign n383 = n310 & n331;
  assign n384 = n382 & ~n383;
  assign n367 = n314 & ~n331;
  assign n368 = ~n309 & n310;
  assign n369 = ~n201 & ~n368;
  assign n370 = ~n367 & n369;
  assign n385 = n384 ^ n370;
  assign n386 = x8 & n385;
  assign n387 = n309 & n314;
  assign n388 = ~x8 & ~n387;
  assign n389 = n382 & n388;
  assign n390 = ~n386 & ~n389;
  assign n358 = n229 ^ x69;
  assign n359 = n210 & n358;
  assign n360 = x68 & n214;
  assign n361 = x67 & n219;
  assign n362 = ~n360 & ~n361;
  assign n363 = x69 & n259;
  assign n364 = n362 & ~n363;
  assign n365 = ~n359 & n364;
  assign n366 = n365 ^ x5;
  assign n391 = n390 ^ n366;
  assign n356 = n336 & ~n337;
  assign n357 = n356 ^ n335;
  assign n392 = n391 ^ n357;
  assign n344 = x71 ^ x70;
  assign n345 = ~n293 & n344;
  assign n346 = n163 & ~n345;
  assign n347 = n346 ^ x1;
  assign n348 = n347 ^ x72;
  assign n349 = x0 & n348;
  assign n350 = x70 & n156;
  assign n351 = ~x0 & ~n350;
  assign n352 = x1 & x71;
  assign n353 = n352 ^ x2;
  assign n354 = n351 & n353;
  assign n355 = ~n349 & ~n354;
  assign n393 = n392 ^ n355;
  assign n341 = n338 ^ n285;
  assign n342 = ~n339 & n341;
  assign n343 = n342 ^ n285;
  assign n394 = n393 ^ n343;
  assign n440 = n384 & n386;
  assign n427 = x66 & n376;
  assign n428 = n268 & ~n371;
  assign n429 = x67 & n428;
  assign n430 = ~n427 & ~n429;
  assign n431 = x7 ^ x6;
  assign n432 = n371 & ~n431;
  assign n433 = ~n268 & n432;
  assign n434 = x65 & n433;
  assign n435 = n430 & ~n434;
  assign n436 = n264 & n372;
  assign n437 = n435 & ~n436;
  assign n438 = n437 ^ x8;
  assign n425 = x9 ^ x8;
  assign n426 = x64 & n425;
  assign n439 = n438 ^ n426;
  assign n441 = n440 ^ n439;
  assign n416 = n247 ^ x70;
  assign n417 = n210 & n416;
  assign n418 = x69 & n214;
  assign n419 = x70 & n259;
  assign n420 = ~n418 & ~n419;
  assign n421 = x68 & n219;
  assign n422 = n420 & ~n421;
  assign n423 = ~n417 & n422;
  assign n424 = n423 ^ x5;
  assign n442 = n441 ^ n424;
  assign n413 = n390 ^ n357;
  assign n414 = n391 & ~n413;
  assign n415 = n414 ^ n357;
  assign n443 = n442 ^ n415;
  assign n402 = x71 & ~x72;
  assign n403 = ~n291 & n402;
  assign n404 = ~x71 & x72;
  assign n405 = ~n292 & n404;
  assign n406 = ~n403 & ~n405;
  assign n407 = n163 & n406;
  assign n408 = n407 ^ x1;
  assign n409 = n408 ^ x73;
  assign n398 = ~x71 & n156;
  assign n399 = x72 ^ x2;
  assign n400 = x1 & n399;
  assign n401 = ~n398 & ~n400;
  assign n410 = n409 ^ n401;
  assign n411 = ~x0 & ~n410;
  assign n412 = n411 ^ n409;
  assign n444 = n443 ^ n412;
  assign n395 = n392 ^ n343;
  assign n396 = n393 & n395;
  assign n397 = n396 ^ n343;
  assign n445 = n444 ^ n397;
  assign n491 = ~n426 & ~n440;
  assign n492 = ~n438 & ~n491;
  assign n484 = x65 ^ x9;
  assign n485 = n425 & ~n484;
  assign n486 = n485 ^ x8;
  assign n487 = n486 ^ x10;
  assign n488 = x64 & n487;
  assign n489 = n149 & n425;
  assign n490 = ~n488 & ~n489;
  assign n493 = n492 ^ n490;
  assign n476 = n300 & n372;
  assign n477 = x67 & n376;
  assign n478 = x66 & n433;
  assign n479 = ~n477 & ~n478;
  assign n480 = x68 & n428;
  assign n481 = n479 & ~n480;
  assign n482 = ~n476 & n481;
  assign n483 = n482 ^ x8;
  assign n494 = n493 ^ n483;
  assign n467 = n293 ^ x71;
  assign n468 = n210 & n467;
  assign n469 = x70 & n214;
  assign n470 = x69 & n219;
  assign n471 = ~n469 & ~n470;
  assign n472 = x71 & n259;
  assign n473 = n471 & ~n472;
  assign n474 = ~n468 & n473;
  assign n475 = n474 ^ x5;
  assign n495 = n494 ^ n475;
  assign n464 = n441 ^ n415;
  assign n465 = ~n442 & n464;
  assign n466 = n465 ^ n415;
  assign n496 = n495 ^ n466;
  assign n453 = ~x72 & ~n403;
  assign n454 = x73 & n453;
  assign n455 = x72 & ~x73;
  assign n456 = ~n405 & n455;
  assign n457 = ~n454 & ~n456;
  assign n458 = n163 & n457;
  assign n459 = n458 ^ x1;
  assign n460 = n459 ^ x74;
  assign n449 = x1 & x73;
  assign n450 = n449 ^ x2;
  assign n451 = ~x1 & x72;
  assign n452 = n450 & ~n451;
  assign n461 = n460 ^ n452;
  assign n462 = ~x0 & n461;
  assign n463 = n462 ^ n460;
  assign n497 = n496 ^ n463;
  assign n446 = n443 ^ n397;
  assign n447 = n444 & ~n446;
  assign n448 = n447 ^ n397;
  assign n498 = n497 ^ n448;
  assign n544 = ~x8 & ~x9;
  assign n554 = x10 & x64;
  assign n563 = n544 & ~n554;
  assign n564 = ~n201 & ~n563;
  assign n543 = x8 & x9;
  assign n557 = ~x10 & x64;
  assign n565 = n543 & ~n557;
  assign n566 = n564 & ~n565;
  assign n567 = x11 & ~n566;
  assign n540 = x11 ^ x10;
  assign n541 = n425 & n540;
  assign n542 = n208 & n541;
  assign n545 = n544 ^ n543;
  assign n546 = x10 & n545;
  assign n547 = n546 ^ n543;
  assign n548 = ~n542 & ~n547;
  assign n549 = x65 & ~n548;
  assign n550 = n149 & n540;
  assign n551 = x66 & n425;
  assign n552 = ~n550 & n551;
  assign n553 = ~n549 & ~n552;
  assign n558 = n544 & n557;
  assign n559 = n553 & ~n558;
  assign n555 = n543 & n554;
  assign n556 = n553 & ~n555;
  assign n560 = n559 ^ n556;
  assign n561 = ~x11 & ~n560;
  assign n562 = n561 ^ n559;
  assign n568 = n567 ^ n562;
  assign n532 = n358 & n372;
  assign n533 = x68 & n376;
  assign n534 = x67 & n433;
  assign n535 = ~n533 & ~n534;
  assign n536 = x69 & n428;
  assign n537 = n535 & ~n536;
  assign n538 = ~n532 & n537;
  assign n539 = n538 ^ x8;
  assign n569 = n568 ^ n539;
  assign n529 = n490 ^ n483;
  assign n530 = ~n493 & ~n529;
  assign n531 = n530 ^ n492;
  assign n570 = n569 ^ n531;
  assign n520 = n345 ^ x72;
  assign n521 = n210 & n520;
  assign n522 = x71 & n214;
  assign n523 = x70 & n219;
  assign n524 = ~n522 & ~n523;
  assign n525 = x72 & n259;
  assign n526 = n524 & ~n525;
  assign n527 = ~n521 & n526;
  assign n528 = n527 ^ x5;
  assign n571 = n570 ^ n528;
  assign n517 = n494 ^ n466;
  assign n518 = n495 & ~n517;
  assign n519 = n518 ^ n466;
  assign n572 = n571 ^ n519;
  assign n502 = x73 & ~n453;
  assign n503 = ~x74 & ~n502;
  assign n504 = ~x73 & ~n456;
  assign n505 = x74 & ~n504;
  assign n506 = ~n503 & ~n505;
  assign n507 = n163 & ~n506;
  assign n508 = n507 ^ x1;
  assign n509 = n508 ^ x75;
  assign n510 = x0 & ~n509;
  assign n511 = x74 ^ x2;
  assign n512 = x1 & n511;
  assign n513 = ~x0 & ~n512;
  assign n514 = ~x73 & n156;
  assign n515 = n513 & ~n514;
  assign n516 = ~n510 & ~n515;
  assign n573 = n572 ^ n516;
  assign n499 = n496 ^ n448;
  assign n500 = ~n497 & n499;
  assign n501 = n500 ^ n448;
  assign n574 = n573 ^ n501;
  assign n623 = n372 & n416;
  assign n624 = x68 & n433;
  assign n625 = x70 & n428;
  assign n626 = ~n624 & ~n625;
  assign n627 = x69 & n376;
  assign n628 = n626 & ~n627;
  assign n629 = ~n623 & n628;
  assign n630 = n629 ^ x8;
  assign n609 = x66 & n547;
  assign n610 = x10 ^ x9;
  assign n611 = n540 & ~n610;
  assign n612 = ~n425 & n611;
  assign n613 = x65 & n612;
  assign n614 = ~n609 & ~n613;
  assign n615 = n425 & ~n540;
  assign n616 = x67 & n615;
  assign n617 = n614 & ~n616;
  assign n618 = n264 & n541;
  assign n619 = n617 & ~n618;
  assign n620 = n619 ^ x11;
  assign n607 = x12 ^ x11;
  assign n608 = x64 & n607;
  assign n621 = n620 ^ n608;
  assign n606 = n559 & n567;
  assign n622 = n621 ^ n606;
  assign n631 = n630 ^ n622;
  assign n603 = n568 ^ n531;
  assign n604 = n569 & n603;
  assign n605 = n604 ^ n531;
  assign n632 = n631 ^ n605;
  assign n594 = n406 ^ x73;
  assign n595 = n210 & ~n594;
  assign n596 = x72 & n214;
  assign n597 = x71 & n219;
  assign n598 = ~n596 & ~n597;
  assign n599 = x73 & n259;
  assign n600 = n598 & ~n599;
  assign n601 = ~n595 & n600;
  assign n602 = n601 ^ x5;
  assign n633 = n632 ^ n602;
  assign n591 = n570 ^ n519;
  assign n592 = ~n571 & n591;
  assign n593 = n592 ^ n519;
  assign n634 = n633 ^ n593;
  assign n582 = x75 & ~n503;
  assign n583 = ~x75 & ~n505;
  assign n584 = ~n582 & ~n583;
  assign n585 = n163 & ~n584;
  assign n586 = n585 ^ x1;
  assign n587 = n586 ^ x76;
  assign n578 = x1 & x75;
  assign n579 = n578 ^ x2;
  assign n580 = ~x1 & x74;
  assign n581 = n579 & ~n580;
  assign n588 = n587 ^ n581;
  assign n589 = ~x0 & n588;
  assign n590 = n589 ^ n587;
  assign n635 = n634 ^ n590;
  assign n575 = n572 ^ n501;
  assign n576 = n573 & ~n575;
  assign n577 = n576 ^ n501;
  assign n636 = n635 ^ n577;
  assign n691 = ~n606 & ~n608;
  assign n692 = ~n620 & ~n691;
  assign n684 = x65 ^ x12;
  assign n685 = n607 & ~n684;
  assign n686 = n685 ^ x11;
  assign n687 = n686 ^ x13;
  assign n688 = x64 & n687;
  assign n689 = n149 & n607;
  assign n690 = ~n688 & ~n689;
  assign n693 = n692 ^ n690;
  assign n676 = n300 & n541;
  assign n677 = x66 & n612;
  assign n678 = x67 & n547;
  assign n679 = ~n677 & ~n678;
  assign n680 = x68 & n615;
  assign n681 = n679 & ~n680;
  assign n682 = ~n676 & n681;
  assign n683 = n682 ^ x11;
  assign n694 = n693 ^ n683;
  assign n668 = n372 & n467;
  assign n669 = x69 & n433;
  assign n670 = x70 & n376;
  assign n671 = ~n669 & ~n670;
  assign n672 = x71 & n428;
  assign n673 = n671 & ~n672;
  assign n674 = ~n668 & n673;
  assign n675 = n674 ^ x8;
  assign n695 = n694 ^ n675;
  assign n665 = n630 ^ n605;
  assign n666 = ~n631 & ~n665;
  assign n667 = n666 ^ n605;
  assign n696 = n695 ^ n667;
  assign n656 = n457 ^ x74;
  assign n657 = n210 & ~n656;
  assign n658 = x73 & n214;
  assign n659 = x74 & n259;
  assign n660 = ~n658 & ~n659;
  assign n661 = x72 & n219;
  assign n662 = n660 & ~n661;
  assign n663 = ~n657 & n662;
  assign n664 = n663 ^ x5;
  assign n697 = n696 ^ n664;
  assign n653 = n632 ^ n593;
  assign n654 = n633 & ~n653;
  assign n655 = n654 ^ n593;
  assign n698 = n697 ^ n655;
  assign n640 = ~x76 & ~n582;
  assign n641 = x76 & ~n583;
  assign n642 = ~n640 & ~n641;
  assign n643 = n163 & ~n642;
  assign n644 = n643 ^ x1;
  assign n645 = n644 ^ x77;
  assign n646 = x0 & ~n645;
  assign n647 = ~x75 & n156;
  assign n648 = ~x0 & ~n647;
  assign n649 = x76 ^ x2;
  assign n650 = x1 & n649;
  assign n651 = n648 & ~n650;
  assign n652 = ~n646 & ~n651;
  assign n699 = n698 ^ n652;
  assign n637 = n634 ^ n577;
  assign n638 = ~n635 & n637;
  assign n639 = n638 ^ n577;
  assign n700 = n699 ^ n639;
  assign n765 = n358 & n541;
  assign n766 = x67 & n612;
  assign n767 = x68 & n547;
  assign n768 = ~n766 & ~n767;
  assign n769 = x69 & n615;
  assign n770 = n768 & ~n769;
  assign n771 = ~n765 & n770;
  assign n772 = n771 ^ x11;
  assign n751 = x14 ^ x13;
  assign n752 = n607 & n751;
  assign n753 = n208 & n752;
  assign n754 = ~x11 & ~x12;
  assign n744 = x11 & x12;
  assign n755 = n754 ^ n744;
  assign n756 = x13 & n755;
  assign n757 = n756 ^ n744;
  assign n758 = ~n753 & ~n757;
  assign n759 = x65 & ~n758;
  assign n760 = n149 & n751;
  assign n761 = x66 & n607;
  assign n762 = ~n760 & n761;
  assign n763 = ~n759 & ~n762;
  assign n743 = ~x64 & ~n689;
  assign n745 = x13 & x64;
  assign n746 = n744 & n745;
  assign n747 = ~n743 & ~n746;
  assign n748 = n747 ^ n746;
  assign n749 = x14 & n748;
  assign n750 = n749 ^ n746;
  assign n764 = n763 ^ n750;
  assign n773 = n772 ^ n764;
  assign n740 = n690 ^ n683;
  assign n741 = ~n693 & ~n740;
  assign n742 = n741 ^ n692;
  assign n774 = n773 ^ n742;
  assign n732 = n372 & n520;
  assign n733 = x71 & n376;
  assign n734 = x70 & n433;
  assign n735 = ~n733 & ~n734;
  assign n736 = x72 & n428;
  assign n737 = n735 & ~n736;
  assign n738 = ~n732 & n737;
  assign n739 = n738 ^ x8;
  assign n775 = n774 ^ n739;
  assign n729 = n694 ^ n667;
  assign n730 = n695 & n729;
  assign n731 = n730 ^ n667;
  assign n776 = n775 ^ n731;
  assign n720 = n506 ^ x75;
  assign n721 = n210 & n720;
  assign n722 = x73 & n219;
  assign n723 = x74 & n214;
  assign n724 = ~n722 & ~n723;
  assign n725 = x75 & n259;
  assign n726 = n724 & ~n725;
  assign n727 = ~n721 & n726;
  assign n728 = n727 ^ x5;
  assign n777 = n776 ^ n728;
  assign n717 = n696 ^ n655;
  assign n718 = ~n697 & n717;
  assign n719 = n718 ^ n655;
  assign n778 = n777 ^ n719;
  assign n704 = x77 & ~n640;
  assign n705 = ~x77 & ~n641;
  assign n706 = ~n704 & ~n705;
  assign n707 = n163 & ~n706;
  assign n708 = n707 ^ x1;
  assign n709 = n708 ^ x78;
  assign n710 = x0 & ~n709;
  assign n711 = x77 ^ x2;
  assign n712 = x1 & n711;
  assign n713 = ~x0 & ~n712;
  assign n714 = ~x76 & n156;
  assign n715 = n713 & ~n714;
  assign n716 = ~n710 & ~n715;
  assign n779 = n778 ^ n716;
  assign n701 = n698 ^ n639;
  assign n702 = n699 & ~n701;
  assign n703 = n702 ^ n639;
  assign n780 = n779 ^ n703;
  assign n840 = n416 & n541;
  assign n841 = x69 & n547;
  assign n842 = x68 & n612;
  assign n843 = ~n841 & ~n842;
  assign n844 = x70 & n615;
  assign n845 = n843 & ~n844;
  assign n846 = ~n840 & n845;
  assign n847 = n846 ^ x11;
  assign n836 = x14 & ~n747;
  assign n837 = n763 & n836;
  assign n834 = x15 ^ x14;
  assign n835 = x64 & n834;
  assign n838 = n837 ^ n835;
  assign n822 = x66 & n757;
  assign n823 = x13 ^ x12;
  assign n824 = n751 & ~n823;
  assign n825 = ~n607 & n824;
  assign n826 = x65 & n825;
  assign n827 = ~n822 & ~n826;
  assign n828 = n607 & ~n751;
  assign n829 = x67 & n828;
  assign n830 = n827 & ~n829;
  assign n831 = n264 & n752;
  assign n832 = n830 & ~n831;
  assign n833 = n832 ^ x14;
  assign n839 = n838 ^ n833;
  assign n848 = n847 ^ n839;
  assign n819 = n772 ^ n742;
  assign n820 = ~n773 & ~n819;
  assign n821 = n820 ^ n742;
  assign n849 = n848 ^ n821;
  assign n811 = n372 & ~n594;
  assign n812 = x72 & n376;
  assign n813 = x71 & n433;
  assign n814 = ~n812 & ~n813;
  assign n815 = x73 & n428;
  assign n816 = n814 & ~n815;
  assign n817 = ~n811 & n816;
  assign n818 = n817 ^ x8;
  assign n850 = n849 ^ n818;
  assign n808 = n774 ^ n731;
  assign n809 = n775 & n808;
  assign n810 = n809 ^ n731;
  assign n851 = n850 ^ n810;
  assign n799 = n584 ^ x76;
  assign n800 = n210 & n799;
  assign n801 = x74 & n219;
  assign n802 = x75 & n214;
  assign n803 = ~n801 & ~n802;
  assign n804 = x76 & n259;
  assign n805 = n803 & ~n804;
  assign n806 = ~n800 & n805;
  assign n807 = n806 ^ x5;
  assign n852 = n851 ^ n807;
  assign n796 = n776 ^ n719;
  assign n797 = ~n777 & n796;
  assign n798 = n797 ^ n719;
  assign n853 = n852 ^ n798;
  assign n788 = x78 ^ x77;
  assign n789 = ~n706 & n788;
  assign n790 = n163 & ~n789;
  assign n791 = n790 ^ x1;
  assign n792 = n791 ^ x79;
  assign n784 = ~x77 & n156;
  assign n785 = x78 ^ x2;
  assign n786 = x1 & n785;
  assign n787 = ~n784 & ~n786;
  assign n793 = n792 ^ n787;
  assign n794 = ~x0 & ~n793;
  assign n795 = n794 ^ n792;
  assign n854 = n853 ^ n795;
  assign n781 = n778 ^ n703;
  assign n782 = n779 & ~n781;
  assign n783 = n782 ^ n703;
  assign n855 = n854 ^ n783;
  assign n923 = ~n835 & ~n837;
  assign n924 = ~n833 & ~n923;
  assign n916 = x65 ^ x15;
  assign n917 = n834 & ~n916;
  assign n918 = n917 ^ x14;
  assign n919 = n918 ^ x16;
  assign n920 = x64 & n919;
  assign n921 = n149 & n834;
  assign n922 = ~n920 & ~n921;
  assign n925 = n924 ^ n922;
  assign n908 = n300 & n752;
  assign n909 = x67 & n757;
  assign n910 = x66 & n825;
  assign n911 = ~n909 & ~n910;
  assign n912 = x68 & n828;
  assign n913 = n911 & ~n912;
  assign n914 = ~n908 & n913;
  assign n915 = n914 ^ x14;
  assign n926 = n925 ^ n915;
  assign n900 = n467 & n541;
  assign n901 = x69 & n612;
  assign n902 = x70 & n547;
  assign n903 = ~n901 & ~n902;
  assign n904 = x71 & n615;
  assign n905 = n903 & ~n904;
  assign n906 = ~n900 & n905;
  assign n907 = n906 ^ x11;
  assign n927 = n926 ^ n907;
  assign n897 = n847 ^ n821;
  assign n898 = ~n848 & ~n897;
  assign n899 = n898 ^ n821;
  assign n928 = n927 ^ n899;
  assign n889 = n372 & ~n656;
  assign n890 = x73 & n376;
  assign n891 = x72 & n433;
  assign n892 = ~n890 & ~n891;
  assign n893 = x74 & n428;
  assign n894 = n892 & ~n893;
  assign n895 = ~n889 & n894;
  assign n896 = n895 ^ x8;
  assign n929 = n928 ^ n896;
  assign n886 = n849 ^ n810;
  assign n887 = n850 & n886;
  assign n888 = n887 ^ n810;
  assign n930 = n929 ^ n888;
  assign n877 = n642 ^ x77;
  assign n878 = n210 & n877;
  assign n879 = x75 & n219;
  assign n880 = x76 & n214;
  assign n881 = ~n879 & ~n880;
  assign n882 = x77 & n259;
  assign n883 = n881 & ~n882;
  assign n884 = ~n878 & n883;
  assign n885 = n884 ^ x5;
  assign n931 = n930 ^ n885;
  assign n874 = n851 ^ n798;
  assign n875 = ~n852 & n874;
  assign n876 = n875 ^ n798;
  assign n932 = n931 ^ n876;
  assign n859 = ~x78 & x79;
  assign n860 = ~n704 & n859;
  assign n861 = x78 & ~x79;
  assign n862 = ~n705 & n861;
  assign n863 = ~n860 & ~n862;
  assign n864 = n163 & n863;
  assign n865 = n864 ^ x1;
  assign n866 = n865 ^ x80;
  assign n867 = x0 & ~n866;
  assign n868 = ~x78 & n156;
  assign n869 = ~x0 & ~n868;
  assign n870 = x79 ^ x2;
  assign n871 = x1 & n870;
  assign n872 = n869 & ~n871;
  assign n873 = ~n867 & ~n872;
  assign n933 = n932 ^ n873;
  assign n856 = n853 ^ n783;
  assign n857 = n854 & ~n856;
  assign n858 = n857 ^ n783;
  assign n934 = n933 ^ n858;
  assign n996 = ~x14 & ~x15;
  assign n1004 = ~x16 & x17;
  assign n1005 = n996 & n1004;
  assign n1006 = x64 & n1005;
  assign n1007 = x17 ^ x16;
  assign n1008 = n834 & n1007;
  assign n1009 = n208 & n1008;
  assign n999 = x14 & x15;
  assign n1010 = n999 ^ n996;
  assign n1011 = x16 & n1010;
  assign n1012 = n1011 ^ n999;
  assign n1013 = ~n1009 & ~n1012;
  assign n1014 = x65 & ~n1013;
  assign n1015 = n149 & n1007;
  assign n1016 = x66 & n834;
  assign n1017 = ~n1015 & n1016;
  assign n1018 = ~n1014 & ~n1017;
  assign n1019 = n1018 ^ x17;
  assign n995 = x16 & x64;
  assign n1020 = n995 & n999;
  assign n1021 = n1018 & n1020;
  assign n1022 = n1019 & n1021;
  assign n1023 = n1022 ^ n1019;
  assign n1024 = ~n1006 & ~n1023;
  assign n997 = ~n201 & ~n996;
  assign n998 = ~n995 & ~n997;
  assign n1000 = ~x16 & x64;
  assign n1001 = n999 & ~n1000;
  assign n1002 = ~n998 & ~n1001;
  assign n1003 = x17 & ~n1002;
  assign n1025 = n1024 ^ n1003;
  assign n987 = n358 & n752;
  assign n988 = x68 & n757;
  assign n989 = x67 & n825;
  assign n990 = ~n988 & ~n989;
  assign n991 = x69 & n828;
  assign n992 = n990 & ~n991;
  assign n993 = ~n987 & n992;
  assign n994 = n993 ^ x14;
  assign n1026 = n1025 ^ n994;
  assign n984 = n922 ^ n915;
  assign n985 = ~n925 & ~n984;
  assign n986 = n985 ^ n924;
  assign n1027 = n1026 ^ n986;
  assign n976 = n520 & n541;
  assign n977 = x71 & n547;
  assign n978 = x70 & n612;
  assign n979 = ~n977 & ~n978;
  assign n980 = x72 & n615;
  assign n981 = n979 & ~n980;
  assign n982 = ~n976 & n981;
  assign n983 = n982 ^ x11;
  assign n1028 = n1027 ^ n983;
  assign n973 = n926 ^ n899;
  assign n974 = n927 & n973;
  assign n975 = n974 ^ n899;
  assign n1029 = n1028 ^ n975;
  assign n965 = n372 & n720;
  assign n966 = x74 & n376;
  assign n967 = x73 & n433;
  assign n968 = ~n966 & ~n967;
  assign n969 = x75 & n428;
  assign n970 = n968 & ~n969;
  assign n971 = ~n965 & n970;
  assign n972 = n971 ^ x8;
  assign n1030 = n1029 ^ n972;
  assign n962 = n928 ^ n888;
  assign n963 = ~n929 & ~n962;
  assign n964 = n963 ^ n888;
  assign n1031 = n1030 ^ n964;
  assign n953 = n706 ^ x78;
  assign n954 = n210 & n953;
  assign n955 = x76 & n219;
  assign n956 = x78 & n259;
  assign n957 = ~n955 & ~n956;
  assign n958 = x77 & n214;
  assign n959 = n957 & ~n958;
  assign n960 = ~n954 & n959;
  assign n961 = n960 ^ x5;
  assign n1032 = n1031 ^ n961;
  assign n950 = n930 ^ n876;
  assign n951 = n931 & ~n950;
  assign n952 = n951 ^ n876;
  assign n1033 = n1032 ^ n952;
  assign n938 = x80 ^ x79;
  assign n939 = n863 & n938;
  assign n940 = n163 & ~n939;
  assign n941 = n940 ^ x1;
  assign n942 = n941 ^ x81;
  assign n943 = x0 & n942;
  assign n944 = ~x1 & x79;
  assign n945 = ~x0 & ~n944;
  assign n946 = x1 & x80;
  assign n947 = n946 ^ x2;
  assign n948 = n945 & n947;
  assign n949 = ~n943 & ~n948;
  assign n1034 = n1033 ^ n949;
  assign n935 = n932 ^ n858;
  assign n936 = ~n933 & n935;
  assign n937 = n936 ^ n858;
  assign n1035 = n1034 ^ n937;
  assign n1111 = n1003 & n1024;
  assign n1098 = x66 & n1012;
  assign n1099 = x16 ^ x15;
  assign n1100 = n1007 & ~n1099;
  assign n1101 = ~n834 & n1100;
  assign n1102 = x65 & n1101;
  assign n1103 = ~n1098 & ~n1102;
  assign n1104 = n834 & ~n1007;
  assign n1105 = x67 & n1104;
  assign n1106 = n1103 & ~n1105;
  assign n1107 = n264 & n1008;
  assign n1108 = n1106 & ~n1107;
  assign n1109 = n1108 ^ x17;
  assign n1096 = x18 ^ x17;
  assign n1097 = x64 & n1096;
  assign n1110 = n1109 ^ n1097;
  assign n1112 = n1111 ^ n1110;
  assign n1088 = n416 & n752;
  assign n1089 = x69 & n757;
  assign n1090 = x68 & n825;
  assign n1091 = ~n1089 & ~n1090;
  assign n1092 = x70 & n828;
  assign n1093 = n1091 & ~n1092;
  assign n1094 = ~n1088 & n1093;
  assign n1095 = n1094 ^ x14;
  assign n1113 = n1112 ^ n1095;
  assign n1085 = n1025 ^ n986;
  assign n1086 = n1026 & n1085;
  assign n1087 = n1086 ^ n986;
  assign n1114 = n1113 ^ n1087;
  assign n1077 = n541 & ~n594;
  assign n1078 = x71 & n612;
  assign n1079 = x73 & n615;
  assign n1080 = ~n1078 & ~n1079;
  assign n1081 = x72 & n547;
  assign n1082 = n1080 & ~n1081;
  assign n1083 = ~n1077 & n1082;
  assign n1084 = n1083 ^ x11;
  assign n1115 = n1114 ^ n1084;
  assign n1074 = n1027 ^ n975;
  assign n1075 = ~n1028 & ~n1074;
  assign n1076 = n1075 ^ n975;
  assign n1116 = n1115 ^ n1076;
  assign n1066 = n372 & n799;
  assign n1067 = x74 & n433;
  assign n1068 = x75 & n376;
  assign n1069 = ~n1067 & ~n1068;
  assign n1070 = x76 & n428;
  assign n1071 = n1069 & ~n1070;
  assign n1072 = ~n1066 & n1071;
  assign n1073 = n1072 ^ x8;
  assign n1117 = n1116 ^ n1073;
  assign n1063 = n1029 ^ n964;
  assign n1064 = n1030 & n1063;
  assign n1065 = n1064 ^ n964;
  assign n1118 = n1117 ^ n1065;
  assign n1054 = n789 ^ x79;
  assign n1055 = n210 & n1054;
  assign n1056 = x77 & n219;
  assign n1057 = x79 & n259;
  assign n1058 = ~n1056 & ~n1057;
  assign n1059 = x78 & n214;
  assign n1060 = n1058 & ~n1059;
  assign n1061 = ~n1055 & n1060;
  assign n1062 = n1061 ^ x5;
  assign n1119 = n1118 ^ n1062;
  assign n1051 = n1031 ^ n952;
  assign n1052 = ~n1032 & n1051;
  assign n1053 = n1052 ^ n952;
  assign n1120 = n1119 ^ n1053;
  assign n1043 = x81 ^ x80;
  assign n1044 = ~n939 & n1043;
  assign n1045 = n163 & ~n1044;
  assign n1046 = n1045 ^ x1;
  assign n1047 = n1046 ^ x82;
  assign n1039 = ~x80 & n156;
  assign n1040 = x81 ^ x2;
  assign n1041 = x1 & n1040;
  assign n1042 = ~n1039 & ~n1041;
  assign n1048 = n1047 ^ n1042;
  assign n1049 = ~x0 & ~n1048;
  assign n1050 = n1049 ^ n1047;
  assign n1121 = n1120 ^ n1050;
  assign n1036 = n1033 ^ n937;
  assign n1037 = ~n1034 & ~n1036;
  assign n1038 = n1037 ^ n937;
  assign n1122 = n1121 ^ n1038;
  assign n1199 = ~n1097 & ~n1111;
  assign n1200 = ~n1109 & ~n1199;
  assign n1190 = n300 & n1008;
  assign n1191 = x67 & n1012;
  assign n1192 = x66 & n1101;
  assign n1193 = ~n1191 & ~n1192;
  assign n1194 = x68 & n1104;
  assign n1195 = n1193 & ~n1194;
  assign n1196 = ~n1190 & n1195;
  assign n1197 = n1196 ^ x17;
  assign n1183 = x65 ^ x18;
  assign n1184 = n1096 & ~n1183;
  assign n1185 = n1184 ^ x17;
  assign n1186 = n1185 ^ x19;
  assign n1187 = x64 & n1186;
  assign n1188 = n149 & n1096;
  assign n1189 = ~n1187 & ~n1188;
  assign n1198 = n1197 ^ n1189;
  assign n1201 = n1200 ^ n1198;
  assign n1175 = n467 & n752;
  assign n1176 = x70 & n757;
  assign n1177 = x69 & n825;
  assign n1178 = ~n1176 & ~n1177;
  assign n1179 = x71 & n828;
  assign n1180 = n1178 & ~n1179;
  assign n1181 = ~n1175 & n1180;
  assign n1182 = n1181 ^ x14;
  assign n1202 = n1201 ^ n1182;
  assign n1172 = n1112 ^ n1087;
  assign n1173 = ~n1113 & ~n1172;
  assign n1174 = n1173 ^ n1087;
  assign n1203 = n1202 ^ n1174;
  assign n1164 = n541 & ~n656;
  assign n1165 = x73 & n547;
  assign n1166 = x72 & n612;
  assign n1167 = ~n1165 & ~n1166;
  assign n1168 = x74 & n615;
  assign n1169 = n1167 & ~n1168;
  assign n1170 = ~n1164 & n1169;
  assign n1171 = n1170 ^ x11;
  assign n1204 = n1203 ^ n1171;
  assign n1161 = n1114 ^ n1076;
  assign n1162 = n1115 & n1161;
  assign n1163 = n1162 ^ n1076;
  assign n1205 = n1204 ^ n1163;
  assign n1153 = n372 & n877;
  assign n1154 = x75 & n433;
  assign n1155 = x76 & n376;
  assign n1156 = ~n1154 & ~n1155;
  assign n1157 = x77 & n428;
  assign n1158 = n1156 & ~n1157;
  assign n1159 = ~n1153 & n1158;
  assign n1160 = n1159 ^ x8;
  assign n1206 = n1205 ^ n1160;
  assign n1150 = n1116 ^ n1065;
  assign n1151 = ~n1117 & ~n1150;
  assign n1152 = n1151 ^ n1065;
  assign n1207 = n1206 ^ n1152;
  assign n1141 = n863 ^ x80;
  assign n1142 = n210 & ~n1141;
  assign n1143 = x79 & n214;
  assign n1144 = x80 & n259;
  assign n1145 = ~n1143 & ~n1144;
  assign n1146 = x78 & n219;
  assign n1147 = n1145 & ~n1146;
  assign n1148 = ~n1142 & n1147;
  assign n1149 = n1148 ^ x5;
  assign n1208 = n1207 ^ n1149;
  assign n1138 = n1118 ^ n1053;
  assign n1139 = n1119 & ~n1138;
  assign n1140 = n1139 ^ n1053;
  assign n1209 = n1208 ^ n1140;
  assign n1126 = x82 ^ x81;
  assign n1127 = ~n1044 & n1126;
  assign n1128 = n163 & ~n1127;
  assign n1129 = n1128 ^ x1;
  assign n1130 = n1129 ^ x83;
  assign n1131 = x0 & ~n1130;
  assign n1132 = ~x81 & n156;
  assign n1133 = ~x0 & ~n1132;
  assign n1134 = x82 ^ x2;
  assign n1135 = x1 & n1134;
  assign n1136 = n1133 & ~n1135;
  assign n1137 = ~n1131 & ~n1136;
  assign n1210 = n1209 ^ n1137;
  assign n1123 = n1120 ^ n1038;
  assign n1124 = ~n1121 & n1123;
  assign n1125 = n1124 ^ n1038;
  assign n1211 = n1210 ^ n1125;
  assign n1283 = ~x17 & ~x18;
  assign n1292 = ~x19 & x20;
  assign n1293 = n1283 & n1292;
  assign n1294 = x64 & n1293;
  assign n1295 = x20 ^ x19;
  assign n1296 = n1096 & n1295;
  assign n1297 = n208 & n1296;
  assign n1287 = x17 & x18;
  assign n1298 = n1287 ^ n1283;
  assign n1299 = x19 & n1298;
  assign n1300 = n1299 ^ n1287;
  assign n1301 = ~n1297 & ~n1300;
  assign n1302 = x65 & ~n1301;
  assign n1303 = n149 & n1295;
  assign n1304 = x66 & n1096;
  assign n1305 = ~n1303 & n1304;
  assign n1306 = ~n1302 & ~n1305;
  assign n1307 = n1306 ^ x20;
  assign n1284 = x19 & x64;
  assign n1308 = n1284 & n1287;
  assign n1309 = n1306 & n1308;
  assign n1310 = n1307 & n1309;
  assign n1311 = n1310 ^ n1307;
  assign n1312 = ~n1294 & ~n1311;
  assign n1285 = n1283 & ~n1284;
  assign n1286 = ~n201 & ~n1285;
  assign n1288 = ~x19 & x64;
  assign n1289 = n1287 & ~n1288;
  assign n1290 = n1286 & ~n1289;
  assign n1291 = x20 & ~n1290;
  assign n1313 = n1312 ^ n1291;
  assign n1275 = n358 & n1008;
  assign n1276 = x67 & n1101;
  assign n1277 = x69 & n1104;
  assign n1278 = ~n1276 & ~n1277;
  assign n1279 = x68 & n1012;
  assign n1280 = n1278 & ~n1279;
  assign n1281 = ~n1275 & n1280;
  assign n1282 = n1281 ^ x17;
  assign n1314 = n1313 ^ n1282;
  assign n1272 = n1200 ^ n1197;
  assign n1273 = ~n1198 & ~n1272;
  assign n1274 = n1273 ^ n1200;
  assign n1315 = n1314 ^ n1274;
  assign n1264 = n520 & n752;
  assign n1265 = x71 & n757;
  assign n1266 = x70 & n825;
  assign n1267 = ~n1265 & ~n1266;
  assign n1268 = x72 & n828;
  assign n1269 = n1267 & ~n1268;
  assign n1270 = ~n1264 & n1269;
  assign n1271 = n1270 ^ x14;
  assign n1316 = n1315 ^ n1271;
  assign n1261 = n1201 ^ n1174;
  assign n1262 = n1202 & n1261;
  assign n1263 = n1262 ^ n1174;
  assign n1317 = n1316 ^ n1263;
  assign n1253 = n541 & n720;
  assign n1254 = x73 & n612;
  assign n1255 = x75 & n615;
  assign n1256 = ~n1254 & ~n1255;
  assign n1257 = x74 & n547;
  assign n1258 = n1256 & ~n1257;
  assign n1259 = ~n1253 & n1258;
  assign n1260 = n1259 ^ x11;
  assign n1318 = n1317 ^ n1260;
  assign n1250 = n1203 ^ n1163;
  assign n1251 = ~n1204 & ~n1250;
  assign n1252 = n1251 ^ n1163;
  assign n1319 = n1318 ^ n1252;
  assign n1242 = n372 & n953;
  assign n1243 = x76 & n433;
  assign n1244 = x78 & n428;
  assign n1245 = ~n1243 & ~n1244;
  assign n1246 = x77 & n376;
  assign n1247 = n1245 & ~n1246;
  assign n1248 = ~n1242 & n1247;
  assign n1249 = n1248 ^ x8;
  assign n1320 = n1319 ^ n1249;
  assign n1239 = n1205 ^ n1152;
  assign n1240 = n1206 & n1239;
  assign n1241 = n1240 ^ n1152;
  assign n1321 = n1320 ^ n1241;
  assign n1230 = n939 ^ x81;
  assign n1231 = n210 & n1230;
  assign n1232 = x79 & n219;
  assign n1233 = x80 & n214;
  assign n1234 = ~n1232 & ~n1233;
  assign n1235 = x81 & n259;
  assign n1236 = n1234 & ~n1235;
  assign n1237 = ~n1231 & n1236;
  assign n1238 = n1237 ^ x5;
  assign n1322 = n1321 ^ n1238;
  assign n1227 = n1207 ^ n1140;
  assign n1228 = ~n1208 & n1227;
  assign n1229 = n1228 ^ n1140;
  assign n1323 = n1322 ^ n1229;
  assign n1215 = x83 ^ x82;
  assign n1216 = ~n1127 & n1215;
  assign n1217 = n163 & ~n1216;
  assign n1218 = n1217 ^ x1;
  assign n1219 = n1218 ^ x84;
  assign n1220 = x0 & n1219;
  assign n1221 = x1 & x83;
  assign n1222 = n1221 ^ x2;
  assign n1223 = ~x1 & x82;
  assign n1224 = ~x0 & ~n1223;
  assign n1225 = n1222 & n1224;
  assign n1226 = ~n1220 & ~n1225;
  assign n1324 = n1323 ^ n1226;
  assign n1212 = n1209 ^ n1125;
  assign n1213 = n1210 & ~n1212;
  assign n1214 = n1213 ^ n1125;
  assign n1325 = n1324 ^ n1214;
  assign n1413 = n1291 & n1312;
  assign n1400 = x66 & n1300;
  assign n1401 = x19 ^ x18;
  assign n1402 = n1295 & ~n1401;
  assign n1403 = ~n1096 & n1402;
  assign n1404 = x65 & n1403;
  assign n1405 = ~n1400 & ~n1404;
  assign n1406 = n1096 & ~n1295;
  assign n1407 = x67 & n1406;
  assign n1408 = n1405 & ~n1407;
  assign n1409 = n264 & n1296;
  assign n1410 = n1408 & ~n1409;
  assign n1411 = n1410 ^ x20;
  assign n1398 = x21 ^ x20;
  assign n1399 = x64 & n1398;
  assign n1412 = n1411 ^ n1399;
  assign n1414 = n1413 ^ n1412;
  assign n1390 = n416 & n1008;
  assign n1391 = x68 & n1101;
  assign n1392 = x70 & n1104;
  assign n1393 = ~n1391 & ~n1392;
  assign n1394 = x69 & n1012;
  assign n1395 = n1393 & ~n1394;
  assign n1396 = ~n1390 & n1395;
  assign n1397 = n1396 ^ x17;
  assign n1415 = n1414 ^ n1397;
  assign n1387 = n1313 ^ n1274;
  assign n1388 = n1314 & n1387;
  assign n1389 = n1388 ^ n1274;
  assign n1416 = n1415 ^ n1389;
  assign n1379 = ~n594 & n752;
  assign n1380 = x71 & n825;
  assign n1381 = x73 & n828;
  assign n1382 = ~n1380 & ~n1381;
  assign n1383 = x72 & n757;
  assign n1384 = n1382 & ~n1383;
  assign n1385 = ~n1379 & n1384;
  assign n1386 = n1385 ^ x14;
  assign n1417 = n1416 ^ n1386;
  assign n1376 = n1315 ^ n1263;
  assign n1377 = ~n1316 & ~n1376;
  assign n1378 = n1377 ^ n1263;
  assign n1418 = n1417 ^ n1378;
  assign n1368 = n541 & n799;
  assign n1369 = x75 & n547;
  assign n1370 = x76 & n615;
  assign n1371 = ~n1369 & ~n1370;
  assign n1372 = x74 & n612;
  assign n1373 = n1371 & ~n1372;
  assign n1374 = ~n1368 & n1373;
  assign n1375 = n1374 ^ x11;
  assign n1419 = n1418 ^ n1375;
  assign n1365 = n1317 ^ n1252;
  assign n1366 = n1318 & n1365;
  assign n1367 = n1366 ^ n1252;
  assign n1420 = n1419 ^ n1367;
  assign n1357 = n372 & n1054;
  assign n1358 = x77 & n433;
  assign n1359 = x78 & n376;
  assign n1360 = ~n1358 & ~n1359;
  assign n1361 = x79 & n428;
  assign n1362 = n1360 & ~n1361;
  assign n1363 = ~n1357 & n1362;
  assign n1364 = n1363 ^ x8;
  assign n1421 = n1420 ^ n1364;
  assign n1354 = n1319 ^ n1241;
  assign n1355 = ~n1320 & ~n1354;
  assign n1356 = n1355 ^ n1241;
  assign n1422 = n1421 ^ n1356;
  assign n1345 = n1044 ^ x82;
  assign n1346 = n210 & n1345;
  assign n1347 = x80 & n219;
  assign n1348 = x81 & n214;
  assign n1349 = ~n1347 & ~n1348;
  assign n1350 = x82 & n259;
  assign n1351 = n1349 & ~n1350;
  assign n1352 = ~n1346 & n1351;
  assign n1353 = n1352 ^ x5;
  assign n1423 = n1422 ^ n1353;
  assign n1342 = n1321 ^ n1229;
  assign n1343 = n1322 & ~n1342;
  assign n1344 = n1343 ^ n1229;
  assign n1424 = n1423 ^ n1344;
  assign n1334 = x84 ^ x83;
  assign n1335 = ~n1216 & n1334;
  assign n1336 = n163 & ~n1335;
  assign n1337 = n1336 ^ x1;
  assign n1338 = n1337 ^ x85;
  assign n1330 = x2 & ~x83;
  assign n1329 = x84 ^ x2;
  assign n1331 = n1330 ^ n1329;
  assign n1332 = x1 & n1331;
  assign n1333 = n1332 ^ n1330;
  assign n1339 = n1338 ^ n1333;
  assign n1340 = ~x0 & n1339;
  assign n1341 = n1340 ^ n1338;
  assign n1425 = n1424 ^ n1341;
  assign n1326 = n1323 ^ n1214;
  assign n1327 = n1324 & n1326;
  assign n1328 = n1327 ^ n1214;
  assign n1426 = n1425 ^ n1328;
  assign n1514 = ~n1399 & ~n1413;
  assign n1515 = ~n1411 & ~n1514;
  assign n1505 = n300 & n1296;
  assign n1506 = x66 & n1403;
  assign n1507 = x68 & n1406;
  assign n1508 = ~n1506 & ~n1507;
  assign n1509 = x67 & n1300;
  assign n1510 = n1508 & ~n1509;
  assign n1511 = ~n1505 & n1510;
  assign n1512 = n1511 ^ x20;
  assign n1498 = x65 ^ x21;
  assign n1499 = n1398 & ~n1498;
  assign n1500 = n1499 ^ x20;
  assign n1501 = n1500 ^ x22;
  assign n1502 = x64 & n1501;
  assign n1503 = n149 & n1398;
  assign n1504 = ~n1502 & ~n1503;
  assign n1513 = n1512 ^ n1504;
  assign n1516 = n1515 ^ n1513;
  assign n1490 = n467 & n1008;
  assign n1491 = x69 & n1101;
  assign n1492 = x71 & n1104;
  assign n1493 = ~n1491 & ~n1492;
  assign n1494 = x70 & n1012;
  assign n1495 = n1493 & ~n1494;
  assign n1496 = ~n1490 & n1495;
  assign n1497 = n1496 ^ x17;
  assign n1517 = n1516 ^ n1497;
  assign n1487 = n1414 ^ n1389;
  assign n1488 = ~n1415 & ~n1487;
  assign n1489 = n1488 ^ n1389;
  assign n1518 = n1517 ^ n1489;
  assign n1479 = ~n656 & n752;
  assign n1480 = x73 & n757;
  assign n1481 = x72 & n825;
  assign n1482 = ~n1480 & ~n1481;
  assign n1483 = x74 & n828;
  assign n1484 = n1482 & ~n1483;
  assign n1485 = ~n1479 & n1484;
  assign n1486 = n1485 ^ x14;
  assign n1519 = n1518 ^ n1486;
  assign n1476 = n1416 ^ n1378;
  assign n1477 = n1417 & n1476;
  assign n1478 = n1477 ^ n1378;
  assign n1520 = n1519 ^ n1478;
  assign n1468 = n541 & n877;
  assign n1469 = x75 & n612;
  assign n1470 = x76 & n547;
  assign n1471 = ~n1469 & ~n1470;
  assign n1472 = x77 & n615;
  assign n1473 = n1471 & ~n1472;
  assign n1474 = ~n1468 & n1473;
  assign n1475 = n1474 ^ x11;
  assign n1521 = n1520 ^ n1475;
  assign n1465 = n1418 ^ n1367;
  assign n1466 = ~n1419 & ~n1465;
  assign n1467 = n1466 ^ n1367;
  assign n1522 = n1521 ^ n1467;
  assign n1457 = n372 & ~n1141;
  assign n1458 = x79 & n376;
  assign n1459 = x78 & n433;
  assign n1460 = ~n1458 & ~n1459;
  assign n1461 = x80 & n428;
  assign n1462 = n1460 & ~n1461;
  assign n1463 = ~n1457 & n1462;
  assign n1464 = n1463 ^ x8;
  assign n1523 = n1522 ^ n1464;
  assign n1454 = n1420 ^ n1356;
  assign n1455 = n1421 & n1454;
  assign n1456 = n1455 ^ n1356;
  assign n1524 = n1523 ^ n1456;
  assign n1445 = n1127 ^ x83;
  assign n1446 = n210 & n1445;
  assign n1447 = x81 & n219;
  assign n1448 = x83 & n259;
  assign n1449 = ~n1447 & ~n1448;
  assign n1450 = x82 & n214;
  assign n1451 = n1449 & ~n1450;
  assign n1452 = ~n1446 & n1451;
  assign n1453 = n1452 ^ x5;
  assign n1525 = n1524 ^ n1453;
  assign n1442 = n1422 ^ n1344;
  assign n1443 = ~n1423 & n1442;
  assign n1444 = n1443 ^ n1344;
  assign n1526 = n1525 ^ n1444;
  assign n1434 = x85 ^ x84;
  assign n1435 = ~n1335 & n1434;
  assign n1436 = n163 & ~n1435;
  assign n1437 = n1436 ^ x1;
  assign n1438 = n1437 ^ x86;
  assign n1430 = ~x84 & n156;
  assign n1431 = x85 ^ x2;
  assign n1432 = x1 & n1431;
  assign n1433 = ~n1430 & ~n1432;
  assign n1439 = n1438 ^ n1433;
  assign n1440 = ~x0 & ~n1439;
  assign n1441 = n1440 ^ n1438;
  assign n1527 = n1526 ^ n1441;
  assign n1427 = n1424 ^ n1328;
  assign n1428 = n1425 & ~n1427;
  assign n1429 = n1428 ^ n1328;
  assign n1528 = n1527 ^ n1429;
  assign n1612 = ~x20 & ~x21;
  assign n1620 = ~x22 & x23;
  assign n1621 = n1612 & n1620;
  assign n1622 = x64 & n1621;
  assign n1623 = x23 ^ x22;
  assign n1624 = n1398 & n1623;
  assign n1625 = n208 & n1624;
  assign n1615 = x20 & x21;
  assign n1626 = n1615 ^ n1612;
  assign n1627 = x22 & n1626;
  assign n1628 = n1627 ^ n1615;
  assign n1629 = ~n1625 & ~n1628;
  assign n1630 = x65 & ~n1629;
  assign n1631 = n149 & n1623;
  assign n1632 = x66 & n1398;
  assign n1633 = ~n1631 & n1632;
  assign n1634 = ~n1630 & ~n1633;
  assign n1635 = n1634 ^ x23;
  assign n1611 = x22 & x64;
  assign n1636 = n1611 & n1615;
  assign n1637 = n1634 & n1636;
  assign n1638 = n1635 & n1637;
  assign n1639 = n1638 ^ n1635;
  assign n1640 = ~n1622 & ~n1639;
  assign n1613 = ~n201 & ~n1612;
  assign n1614 = ~n1611 & ~n1613;
  assign n1616 = ~x22 & x64;
  assign n1617 = n1615 & ~n1616;
  assign n1618 = ~n1614 & ~n1617;
  assign n1619 = x23 & ~n1618;
  assign n1641 = n1640 ^ n1619;
  assign n1603 = n358 & n1296;
  assign n1604 = x67 & n1403;
  assign n1605 = x69 & n1406;
  assign n1606 = ~n1604 & ~n1605;
  assign n1607 = x68 & n1300;
  assign n1608 = n1606 & ~n1607;
  assign n1609 = ~n1603 & n1608;
  assign n1610 = n1609 ^ x20;
  assign n1642 = n1641 ^ n1610;
  assign n1600 = n1515 ^ n1512;
  assign n1601 = ~n1513 & ~n1600;
  assign n1602 = n1601 ^ n1515;
  assign n1643 = n1642 ^ n1602;
  assign n1592 = n520 & n1008;
  assign n1593 = x70 & n1101;
  assign n1594 = x72 & n1104;
  assign n1595 = ~n1593 & ~n1594;
  assign n1596 = x71 & n1012;
  assign n1597 = n1595 & ~n1596;
  assign n1598 = ~n1592 & n1597;
  assign n1599 = n1598 ^ x17;
  assign n1644 = n1643 ^ n1599;
  assign n1589 = n1516 ^ n1489;
  assign n1590 = n1517 & n1589;
  assign n1591 = n1590 ^ n1489;
  assign n1645 = n1644 ^ n1591;
  assign n1581 = n720 & n752;
  assign n1582 = x73 & n825;
  assign n1583 = x75 & n828;
  assign n1584 = ~n1582 & ~n1583;
  assign n1585 = x74 & n757;
  assign n1586 = n1584 & ~n1585;
  assign n1587 = ~n1581 & n1586;
  assign n1588 = n1587 ^ x14;
  assign n1646 = n1645 ^ n1588;
  assign n1578 = n1518 ^ n1478;
  assign n1579 = ~n1519 & ~n1578;
  assign n1580 = n1579 ^ n1478;
  assign n1647 = n1646 ^ n1580;
  assign n1570 = n541 & n953;
  assign n1571 = x76 & n612;
  assign n1572 = x77 & n547;
  assign n1573 = ~n1571 & ~n1572;
  assign n1574 = x78 & n615;
  assign n1575 = n1573 & ~n1574;
  assign n1576 = ~n1570 & n1575;
  assign n1577 = n1576 ^ x11;
  assign n1648 = n1647 ^ n1577;
  assign n1567 = n1520 ^ n1467;
  assign n1568 = n1521 & n1567;
  assign n1569 = n1568 ^ n1467;
  assign n1649 = n1648 ^ n1569;
  assign n1559 = n372 & n1230;
  assign n1560 = x79 & n433;
  assign n1561 = x81 & n428;
  assign n1562 = ~n1560 & ~n1561;
  assign n1563 = x80 & n376;
  assign n1564 = n1562 & ~n1563;
  assign n1565 = ~n1559 & n1564;
  assign n1566 = n1565 ^ x8;
  assign n1650 = n1649 ^ n1566;
  assign n1556 = n1522 ^ n1456;
  assign n1557 = ~n1523 & ~n1556;
  assign n1558 = n1557 ^ n1456;
  assign n1651 = n1650 ^ n1558;
  assign n1547 = n1216 ^ x84;
  assign n1548 = n210 & n1547;
  assign n1549 = x82 & n219;
  assign n1550 = x84 & n259;
  assign n1551 = ~n1549 & ~n1550;
  assign n1552 = x83 & n214;
  assign n1553 = n1551 & ~n1552;
  assign n1554 = ~n1548 & n1553;
  assign n1555 = n1554 ^ x5;
  assign n1652 = n1651 ^ n1555;
  assign n1544 = n1524 ^ n1444;
  assign n1545 = n1525 & ~n1544;
  assign n1546 = n1545 ^ n1444;
  assign n1653 = n1652 ^ n1546;
  assign n1536 = x86 ^ x85;
  assign n1537 = ~n1435 & n1536;
  assign n1538 = n163 & ~n1537;
  assign n1539 = n1538 ^ x1;
  assign n1540 = n1539 ^ x87;
  assign n1532 = ~x85 & n156;
  assign n1533 = x86 ^ x2;
  assign n1534 = x1 & n1533;
  assign n1535 = ~n1532 & ~n1534;
  assign n1541 = n1540 ^ n1535;
  assign n1542 = ~x0 & ~n1541;
  assign n1543 = n1542 ^ n1540;
  assign n1654 = n1653 ^ n1543;
  assign n1529 = n1526 ^ n1429;
  assign n1530 = ~n1527 & n1529;
  assign n1531 = n1530 ^ n1429;
  assign n1655 = n1654 ^ n1531;
  assign n1753 = n1619 & n1640;
  assign n1740 = x22 ^ x21;
  assign n1741 = n1623 & ~n1740;
  assign n1742 = ~n1398 & n1741;
  assign n1743 = x65 & n1742;
  assign n1744 = n1398 & ~n1623;
  assign n1745 = x67 & n1744;
  assign n1746 = ~n1743 & ~n1745;
  assign n1747 = x66 & n1628;
  assign n1748 = n1746 & ~n1747;
  assign n1749 = n264 & n1624;
  assign n1750 = n1748 & ~n1749;
  assign n1751 = n1750 ^ x23;
  assign n1738 = x24 ^ x23;
  assign n1739 = x64 & n1738;
  assign n1752 = n1751 ^ n1739;
  assign n1754 = n1753 ^ n1752;
  assign n1730 = n416 & n1296;
  assign n1731 = x68 & n1403;
  assign n1732 = x69 & n1300;
  assign n1733 = ~n1731 & ~n1732;
  assign n1734 = x70 & n1406;
  assign n1735 = n1733 & ~n1734;
  assign n1736 = ~n1730 & n1735;
  assign n1737 = n1736 ^ x20;
  assign n1755 = n1754 ^ n1737;
  assign n1727 = n1641 ^ n1602;
  assign n1728 = n1642 & n1727;
  assign n1729 = n1728 ^ n1602;
  assign n1756 = n1755 ^ n1729;
  assign n1719 = ~n594 & n1008;
  assign n1720 = x71 & n1101;
  assign n1721 = x73 & n1104;
  assign n1722 = ~n1720 & ~n1721;
  assign n1723 = x72 & n1012;
  assign n1724 = n1722 & ~n1723;
  assign n1725 = ~n1719 & n1724;
  assign n1726 = n1725 ^ x17;
  assign n1757 = n1756 ^ n1726;
  assign n1716 = n1643 ^ n1591;
  assign n1717 = ~n1644 & ~n1716;
  assign n1718 = n1717 ^ n1591;
  assign n1758 = n1757 ^ n1718;
  assign n1708 = n752 & n799;
  assign n1709 = x74 & n825;
  assign n1710 = x75 & n757;
  assign n1711 = ~n1709 & ~n1710;
  assign n1712 = x76 & n828;
  assign n1713 = n1711 & ~n1712;
  assign n1714 = ~n1708 & n1713;
  assign n1715 = n1714 ^ x14;
  assign n1759 = n1758 ^ n1715;
  assign n1705 = n1645 ^ n1580;
  assign n1706 = n1646 & n1705;
  assign n1707 = n1706 ^ n1580;
  assign n1760 = n1759 ^ n1707;
  assign n1697 = n541 & n1054;
  assign n1698 = x77 & n612;
  assign n1699 = x79 & n615;
  assign n1700 = ~n1698 & ~n1699;
  assign n1701 = x78 & n547;
  assign n1702 = n1700 & ~n1701;
  assign n1703 = ~n1697 & n1702;
  assign n1704 = n1703 ^ x11;
  assign n1761 = n1760 ^ n1704;
  assign n1694 = n1647 ^ n1569;
  assign n1695 = ~n1648 & ~n1694;
  assign n1696 = n1695 ^ n1569;
  assign n1762 = n1761 ^ n1696;
  assign n1686 = n372 & n1345;
  assign n1687 = x80 & n433;
  assign n1688 = x81 & n376;
  assign n1689 = ~n1687 & ~n1688;
  assign n1690 = x82 & n428;
  assign n1691 = n1689 & ~n1690;
  assign n1692 = ~n1686 & n1691;
  assign n1693 = n1692 ^ x8;
  assign n1763 = n1762 ^ n1693;
  assign n1683 = n1649 ^ n1558;
  assign n1684 = n1650 & n1683;
  assign n1685 = n1684 ^ n1558;
  assign n1764 = n1763 ^ n1685;
  assign n1674 = n1335 ^ x85;
  assign n1675 = n210 & n1674;
  assign n1676 = x83 & n219;
  assign n1677 = x84 & n214;
  assign n1678 = ~n1676 & ~n1677;
  assign n1679 = x85 & n259;
  assign n1680 = n1678 & ~n1679;
  assign n1681 = ~n1675 & n1680;
  assign n1682 = n1681 ^ x5;
  assign n1765 = n1764 ^ n1682;
  assign n1671 = n1651 ^ n1546;
  assign n1672 = ~n1652 & n1671;
  assign n1673 = n1672 ^ n1546;
  assign n1766 = n1765 ^ n1673;
  assign n1663 = x87 ^ x86;
  assign n1664 = ~n1537 & n1663;
  assign n1665 = n163 & ~n1664;
  assign n1666 = n1665 ^ x1;
  assign n1667 = n1666 ^ x88;
  assign n1659 = x1 & x87;
  assign n1660 = n1659 ^ x2;
  assign n1661 = ~x1 & x86;
  assign n1662 = n1660 & ~n1661;
  assign n1668 = n1667 ^ n1662;
  assign n1669 = ~x0 & n1668;
  assign n1670 = n1669 ^ n1667;
  assign n1767 = n1766 ^ n1670;
  assign n1656 = n1653 ^ n1531;
  assign n1657 = n1654 & ~n1656;
  assign n1658 = n1657 ^ n1531;
  assign n1768 = n1767 ^ n1658;
  assign n1867 = ~n1739 & ~n1753;
  assign n1868 = ~n1751 & ~n1867;
  assign n1858 = n300 & n1624;
  assign n1859 = x66 & n1742;
  assign n1860 = x68 & n1744;
  assign n1861 = ~n1859 & ~n1860;
  assign n1862 = x67 & n1628;
  assign n1863 = n1861 & ~n1862;
  assign n1864 = ~n1858 & n1863;
  assign n1865 = n1864 ^ x23;
  assign n1851 = x65 ^ x24;
  assign n1852 = n1738 & ~n1851;
  assign n1853 = n1852 ^ x23;
  assign n1854 = n1853 ^ x25;
  assign n1855 = x64 & n1854;
  assign n1856 = n149 & n1738;
  assign n1857 = ~n1855 & ~n1856;
  assign n1866 = n1865 ^ n1857;
  assign n1869 = n1868 ^ n1866;
  assign n1843 = n467 & n1296;
  assign n1844 = x69 & n1403;
  assign n1845 = x70 & n1300;
  assign n1846 = ~n1844 & ~n1845;
  assign n1847 = x71 & n1406;
  assign n1848 = n1846 & ~n1847;
  assign n1849 = ~n1843 & n1848;
  assign n1850 = n1849 ^ x20;
  assign n1870 = n1869 ^ n1850;
  assign n1840 = n1754 ^ n1729;
  assign n1841 = ~n1755 & ~n1840;
  assign n1842 = n1841 ^ n1729;
  assign n1871 = n1870 ^ n1842;
  assign n1832 = ~n656 & n1008;
  assign n1833 = x73 & n1012;
  assign n1834 = x72 & n1101;
  assign n1835 = ~n1833 & ~n1834;
  assign n1836 = x74 & n1104;
  assign n1837 = n1835 & ~n1836;
  assign n1838 = ~n1832 & n1837;
  assign n1839 = n1838 ^ x17;
  assign n1872 = n1871 ^ n1839;
  assign n1829 = n1756 ^ n1718;
  assign n1830 = n1757 & n1829;
  assign n1831 = n1830 ^ n1718;
  assign n1873 = n1872 ^ n1831;
  assign n1821 = n752 & n877;
  assign n1822 = x75 & n825;
  assign n1823 = x76 & n757;
  assign n1824 = ~n1822 & ~n1823;
  assign n1825 = x77 & n828;
  assign n1826 = n1824 & ~n1825;
  assign n1827 = ~n1821 & n1826;
  assign n1828 = n1827 ^ x14;
  assign n1874 = n1873 ^ n1828;
  assign n1818 = n1758 ^ n1707;
  assign n1819 = ~n1759 & ~n1818;
  assign n1820 = n1819 ^ n1707;
  assign n1875 = n1874 ^ n1820;
  assign n1810 = n541 & ~n1141;
  assign n1811 = x78 & n612;
  assign n1812 = x79 & n547;
  assign n1813 = ~n1811 & ~n1812;
  assign n1814 = x80 & n615;
  assign n1815 = n1813 & ~n1814;
  assign n1816 = ~n1810 & n1815;
  assign n1817 = n1816 ^ x11;
  assign n1876 = n1875 ^ n1817;
  assign n1807 = n1760 ^ n1696;
  assign n1808 = n1761 & n1807;
  assign n1809 = n1808 ^ n1696;
  assign n1877 = n1876 ^ n1809;
  assign n1799 = n372 & n1445;
  assign n1800 = x81 & n433;
  assign n1801 = x82 & n376;
  assign n1802 = ~n1800 & ~n1801;
  assign n1803 = x83 & n428;
  assign n1804 = n1802 & ~n1803;
  assign n1805 = ~n1799 & n1804;
  assign n1806 = n1805 ^ x8;
  assign n1878 = n1877 ^ n1806;
  assign n1796 = n1762 ^ n1685;
  assign n1797 = ~n1763 & ~n1796;
  assign n1798 = n1797 ^ n1685;
  assign n1879 = n1878 ^ n1798;
  assign n1787 = n1435 ^ x86;
  assign n1788 = n210 & n1787;
  assign n1789 = x84 & n219;
  assign n1790 = x86 & n259;
  assign n1791 = ~n1789 & ~n1790;
  assign n1792 = x85 & n214;
  assign n1793 = n1791 & ~n1792;
  assign n1794 = ~n1788 & n1793;
  assign n1795 = n1794 ^ x5;
  assign n1880 = n1879 ^ n1795;
  assign n1784 = n1764 ^ n1673;
  assign n1785 = n1765 & ~n1784;
  assign n1786 = n1785 ^ n1673;
  assign n1881 = n1880 ^ n1786;
  assign n1776 = x88 ^ x87;
  assign n1777 = ~n1664 & n1776;
  assign n1778 = n163 & ~n1777;
  assign n1779 = n1778 ^ x1;
  assign n1780 = n1779 ^ x89;
  assign n1772 = ~x87 & n156;
  assign n1773 = x88 ^ x2;
  assign n1774 = x1 & n1773;
  assign n1775 = ~n1772 & ~n1774;
  assign n1781 = n1780 ^ n1775;
  assign n1782 = ~x0 & ~n1781;
  assign n1783 = n1782 ^ n1780;
  assign n1882 = n1881 ^ n1783;
  assign n1769 = n1766 ^ n1658;
  assign n1770 = ~n1767 & n1769;
  assign n1771 = n1770 ^ n1658;
  assign n1883 = n1882 ^ n1771;
  assign n2001 = n720 & n1008;
  assign n2002 = x74 & n1012;
  assign n2003 = x73 & n1101;
  assign n2004 = ~n2002 & ~n2003;
  assign n2005 = x75 & n1104;
  assign n2006 = n2004 & ~n2005;
  assign n2007 = ~n2001 & n2006;
  assign n2008 = n2007 ^ x17;
  assign n1998 = n1871 ^ n1831;
  assign n1999 = ~n1872 & ~n1998;
  assign n2000 = n1999 ^ n1831;
  assign n2009 = n2008 ^ n2000;
  assign n1986 = n358 & n1624;
  assign n1987 = x67 & n1742;
  assign n1988 = x69 & n1744;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = x68 & n1628;
  assign n1991 = n1989 & ~n1990;
  assign n1992 = ~n1986 & n1991;
  assign n1993 = n1992 ^ x23;
  assign n1968 = x26 ^ x25;
  assign n1969 = n1738 & n1968;
  assign n1970 = n208 & n1969;
  assign n1963 = x23 & x24;
  assign n1959 = ~x23 & ~x24;
  assign n1971 = n1963 ^ n1959;
  assign n1972 = x25 & n1971;
  assign n1973 = n1972 ^ n1963;
  assign n1974 = ~n1970 & ~n1973;
  assign n1975 = x65 & ~n1974;
  assign n1976 = x25 ^ x24;
  assign n1977 = n1968 & ~n1976;
  assign n1978 = ~n1738 & n1977;
  assign n1979 = x64 & n1978;
  assign n1980 = n149 & n1968;
  assign n1981 = x66 & n1738;
  assign n1982 = ~n1980 & n1981;
  assign n1983 = ~n1979 & ~n1982;
  assign n1984 = ~n1975 & n1983;
  assign n1960 = x25 & x64;
  assign n1961 = n1959 & ~n1960;
  assign n1962 = ~n201 & ~n1961;
  assign n1964 = ~x25 & x64;
  assign n1965 = n1963 & ~n1964;
  assign n1966 = n1962 & ~n1965;
  assign n1967 = x26 & n1966;
  assign n1985 = n1984 ^ n1967;
  assign n1994 = n1993 ^ n1985;
  assign n1956 = n1868 ^ n1865;
  assign n1957 = ~n1866 & ~n1956;
  assign n1958 = n1957 ^ n1868;
  assign n1995 = n1994 ^ n1958;
  assign n1948 = n520 & n1296;
  assign n1949 = x70 & n1403;
  assign n1950 = x72 & n1406;
  assign n1951 = ~n1949 & ~n1950;
  assign n1952 = x71 & n1300;
  assign n1953 = n1951 & ~n1952;
  assign n1954 = ~n1948 & n1953;
  assign n1955 = n1954 ^ x20;
  assign n1996 = n1995 ^ n1955;
  assign n1945 = n1869 ^ n1842;
  assign n1946 = n1870 & n1945;
  assign n1947 = n1946 ^ n1842;
  assign n1997 = n1996 ^ n1947;
  assign n2010 = n2009 ^ n1997;
  assign n1937 = n752 & n953;
  assign n1938 = x76 & n825;
  assign n1939 = x77 & n757;
  assign n1940 = ~n1938 & ~n1939;
  assign n1941 = x78 & n828;
  assign n1942 = n1940 & ~n1941;
  assign n1943 = ~n1937 & n1942;
  assign n1944 = n1943 ^ x14;
  assign n2011 = n2010 ^ n1944;
  assign n1934 = n1873 ^ n1820;
  assign n1935 = n1874 & n1934;
  assign n1936 = n1935 ^ n1820;
  assign n2012 = n2011 ^ n1936;
  assign n1926 = n541 & n1230;
  assign n1927 = x79 & n612;
  assign n1928 = x81 & n615;
  assign n1929 = ~n1927 & ~n1928;
  assign n1930 = x80 & n547;
  assign n1931 = n1929 & ~n1930;
  assign n1932 = ~n1926 & n1931;
  assign n1933 = n1932 ^ x11;
  assign n2013 = n2012 ^ n1933;
  assign n1923 = n1875 ^ n1809;
  assign n1924 = ~n1876 & ~n1923;
  assign n1925 = n1924 ^ n1809;
  assign n2014 = n2013 ^ n1925;
  assign n1915 = n372 & n1547;
  assign n1916 = x82 & n433;
  assign n1917 = x84 & n428;
  assign n1918 = ~n1916 & ~n1917;
  assign n1919 = x83 & n376;
  assign n1920 = n1918 & ~n1919;
  assign n1921 = ~n1915 & n1920;
  assign n1922 = n1921 ^ x8;
  assign n2015 = n2014 ^ n1922;
  assign n1912 = n1877 ^ n1798;
  assign n1913 = n1878 & n1912;
  assign n1914 = n1913 ^ n1798;
  assign n2016 = n2015 ^ n1914;
  assign n1903 = n1537 ^ x87;
  assign n1904 = n210 & n1903;
  assign n1905 = x85 & n219;
  assign n1906 = x87 & n259;
  assign n1907 = ~n1905 & ~n1906;
  assign n1908 = x86 & n214;
  assign n1909 = n1907 & ~n1908;
  assign n1910 = ~n1904 & n1909;
  assign n1911 = n1910 ^ x5;
  assign n2017 = n2016 ^ n1911;
  assign n1900 = n1879 ^ n1786;
  assign n1901 = ~n1880 & n1900;
  assign n1902 = n1901 ^ n1786;
  assign n2018 = n2017 ^ n1902;
  assign n1887 = x89 ^ x88;
  assign n1888 = ~n1777 & n1887;
  assign n1889 = n163 & ~n1888;
  assign n1890 = n1889 ^ x1;
  assign n1891 = n1890 ^ x90;
  assign n1892 = x0 & ~n1891;
  assign n1893 = x2 & ~x88;
  assign n1894 = ~x1 & n1893;
  assign n1895 = ~x0 & ~n1894;
  assign n1896 = x89 ^ x2;
  assign n1897 = x1 & n1896;
  assign n1898 = n1895 & ~n1897;
  assign n1899 = ~n1892 & ~n1898;
  assign n2019 = n2018 ^ n1899;
  assign n1884 = n1881 ^ n1771;
  assign n1885 = n1882 & ~n1884;
  assign n1886 = n1885 ^ n1771;
  assign n2020 = n2019 ^ n1886;
  assign n2122 = n416 & n1624;
  assign n2123 = x68 & n1742;
  assign n2124 = x70 & n1744;
  assign n2125 = ~n2123 & ~n2124;
  assign n2126 = x69 & n1628;
  assign n2127 = n2125 & ~n2126;
  assign n2128 = ~n2122 & n2127;
  assign n2129 = n2128 ^ x23;
  assign n2118 = x26 & ~n1966;
  assign n2119 = n1984 & n2118;
  assign n2116 = x27 ^ x26;
  assign n2117 = x64 & n2116;
  assign n2120 = n2119 ^ n2117;
  assign n2107 = n264 & n1969;
  assign n2108 = n1738 & ~n1968;
  assign n2109 = x67 & n2108;
  assign n2110 = ~n2107 & ~n2109;
  assign n2111 = x65 & n1978;
  assign n2112 = x66 & n1973;
  assign n2113 = ~n2111 & ~n2112;
  assign n2114 = n2110 & n2113;
  assign n2115 = n2114 ^ x26;
  assign n2121 = n2120 ^ n2115;
  assign n2130 = n2129 ^ n2121;
  assign n2104 = n1993 ^ n1958;
  assign n2105 = ~n1994 & ~n2104;
  assign n2106 = n2105 ^ n1958;
  assign n2131 = n2130 ^ n2106;
  assign n2096 = ~n594 & n1296;
  assign n2097 = x71 & n1403;
  assign n2098 = x73 & n1406;
  assign n2099 = ~n2097 & ~n2098;
  assign n2100 = x72 & n1300;
  assign n2101 = n2099 & ~n2100;
  assign n2102 = ~n2096 & n2101;
  assign n2103 = n2102 ^ x20;
  assign n2132 = n2131 ^ n2103;
  assign n2093 = n1995 ^ n1947;
  assign n2094 = n1996 & n2093;
  assign n2095 = n2094 ^ n1947;
  assign n2133 = n2132 ^ n2095;
  assign n2085 = n799 & n1008;
  assign n2086 = x74 & n1101;
  assign n2087 = x76 & n1104;
  assign n2088 = ~n2086 & ~n2087;
  assign n2089 = x75 & n1012;
  assign n2090 = n2088 & ~n2089;
  assign n2091 = ~n2085 & n2090;
  assign n2092 = n2091 ^ x17;
  assign n2134 = n2133 ^ n2092;
  assign n2082 = n2008 ^ n1997;
  assign n2083 = ~n2009 & ~n2082;
  assign n2084 = n2083 ^ n2000;
  assign n2135 = n2134 ^ n2084;
  assign n2074 = n752 & n1054;
  assign n2075 = x77 & n825;
  assign n2076 = x79 & n828;
  assign n2077 = ~n2075 & ~n2076;
  assign n2078 = x78 & n757;
  assign n2079 = n2077 & ~n2078;
  assign n2080 = ~n2074 & n2079;
  assign n2081 = n2080 ^ x14;
  assign n2136 = n2135 ^ n2081;
  assign n2071 = n2010 ^ n1936;
  assign n2072 = n2011 & n2071;
  assign n2073 = n2072 ^ n1936;
  assign n2137 = n2136 ^ n2073;
  assign n2063 = n541 & n1345;
  assign n2064 = x80 & n612;
  assign n2065 = x81 & n547;
  assign n2066 = ~n2064 & ~n2065;
  assign n2067 = x82 & n615;
  assign n2068 = n2066 & ~n2067;
  assign n2069 = ~n2063 & n2068;
  assign n2070 = n2069 ^ x11;
  assign n2138 = n2137 ^ n2070;
  assign n2060 = n2012 ^ n1925;
  assign n2061 = ~n2013 & ~n2060;
  assign n2062 = n2061 ^ n1925;
  assign n2139 = n2138 ^ n2062;
  assign n2052 = n372 & n1674;
  assign n2053 = x83 & n433;
  assign n2054 = x84 & n376;
  assign n2055 = ~n2053 & ~n2054;
  assign n2056 = x85 & n428;
  assign n2057 = n2055 & ~n2056;
  assign n2058 = ~n2052 & n2057;
  assign n2059 = n2058 ^ x8;
  assign n2140 = n2139 ^ n2059;
  assign n2049 = n2014 ^ n1914;
  assign n2050 = n2015 & n2049;
  assign n2051 = n2050 ^ n1914;
  assign n2141 = n2140 ^ n2051;
  assign n2040 = n1664 ^ x88;
  assign n2041 = n210 & n2040;
  assign n2042 = x86 & n219;
  assign n2043 = x87 & n214;
  assign n2044 = ~n2042 & ~n2043;
  assign n2045 = x88 & n259;
  assign n2046 = n2044 & ~n2045;
  assign n2047 = ~n2041 & n2046;
  assign n2048 = n2047 ^ x5;
  assign n2142 = n2141 ^ n2048;
  assign n2037 = n2016 ^ n1902;
  assign n2038 = ~n2017 & n2037;
  assign n2039 = n2038 ^ n1902;
  assign n2143 = n2142 ^ n2039;
  assign n2024 = x90 ^ x89;
  assign n2025 = ~n1888 & n2024;
  assign n2026 = n163 & ~n2025;
  assign n2027 = n2026 ^ x1;
  assign n2028 = n2027 ^ x91;
  assign n2029 = x0 & ~n2028;
  assign n2030 = x2 & ~x89;
  assign n2031 = ~x1 & n2030;
  assign n2032 = ~x0 & ~n2031;
  assign n2033 = x90 ^ x2;
  assign n2034 = x1 & n2033;
  assign n2035 = n2032 & ~n2034;
  assign n2036 = ~n2029 & ~n2035;
  assign n2144 = n2143 ^ n2036;
  assign n2021 = n2018 ^ n1886;
  assign n2022 = n2019 & ~n2021;
  assign n2023 = n2022 ^ n1886;
  assign n2145 = n2144 ^ n2023;
  assign n2250 = n467 & n1624;
  assign n2251 = x70 & n1628;
  assign n2252 = x69 & n1742;
  assign n2253 = ~n2251 & ~n2252;
  assign n2254 = x71 & n1744;
  assign n2255 = n2253 & ~n2254;
  assign n2256 = ~n2250 & n2255;
  assign n2257 = n2256 ^ x23;
  assign n2247 = ~n2117 & ~n2119;
  assign n2248 = ~n2115 & ~n2247;
  assign n2238 = n300 & n1969;
  assign n2239 = x66 & n1978;
  assign n2240 = x67 & n1973;
  assign n2241 = ~n2239 & ~n2240;
  assign n2242 = x68 & n2108;
  assign n2243 = n2241 & ~n2242;
  assign n2244 = ~n2238 & n2243;
  assign n2245 = n2244 ^ x26;
  assign n2231 = x65 ^ x27;
  assign n2232 = n2116 & ~n2231;
  assign n2233 = n2232 ^ x26;
  assign n2234 = n2233 ^ x28;
  assign n2235 = x64 & n2234;
  assign n2236 = n149 & n2116;
  assign n2237 = ~n2235 & ~n2236;
  assign n2246 = n2245 ^ n2237;
  assign n2249 = n2248 ^ n2246;
  assign n2258 = n2257 ^ n2249;
  assign n2228 = n2129 ^ n2106;
  assign n2229 = ~n2130 & ~n2228;
  assign n2230 = n2229 ^ n2106;
  assign n2259 = n2258 ^ n2230;
  assign n2220 = ~n656 & n1296;
  assign n2221 = x73 & n1300;
  assign n2222 = x74 & n1406;
  assign n2223 = ~n2221 & ~n2222;
  assign n2224 = x72 & n1403;
  assign n2225 = n2223 & ~n2224;
  assign n2226 = ~n2220 & n2225;
  assign n2227 = n2226 ^ x20;
  assign n2260 = n2259 ^ n2227;
  assign n2217 = n2131 ^ n2095;
  assign n2218 = n2132 & n2217;
  assign n2219 = n2218 ^ n2095;
  assign n2261 = n2260 ^ n2219;
  assign n2209 = n877 & n1008;
  assign n2210 = x75 & n1101;
  assign n2211 = x76 & n1012;
  assign n2212 = ~n2210 & ~n2211;
  assign n2213 = x77 & n1104;
  assign n2214 = n2212 & ~n2213;
  assign n2215 = ~n2209 & n2214;
  assign n2216 = n2215 ^ x17;
  assign n2262 = n2261 ^ n2216;
  assign n2206 = n2133 ^ n2084;
  assign n2207 = ~n2134 & ~n2206;
  assign n2208 = n2207 ^ n2084;
  assign n2263 = n2262 ^ n2208;
  assign n2198 = n752 & ~n1141;
  assign n2199 = x78 & n825;
  assign n2200 = x80 & n828;
  assign n2201 = ~n2199 & ~n2200;
  assign n2202 = x79 & n757;
  assign n2203 = n2201 & ~n2202;
  assign n2204 = ~n2198 & n2203;
  assign n2205 = n2204 ^ x14;
  assign n2264 = n2263 ^ n2205;
  assign n2195 = n2135 ^ n2073;
  assign n2196 = n2136 & n2195;
  assign n2197 = n2196 ^ n2073;
  assign n2265 = n2264 ^ n2197;
  assign n2187 = n541 & n1445;
  assign n2188 = x81 & n612;
  assign n2189 = x82 & n547;
  assign n2190 = ~n2188 & ~n2189;
  assign n2191 = x83 & n615;
  assign n2192 = n2190 & ~n2191;
  assign n2193 = ~n2187 & n2192;
  assign n2194 = n2193 ^ x11;
  assign n2266 = n2265 ^ n2194;
  assign n2184 = n2137 ^ n2062;
  assign n2185 = ~n2138 & ~n2184;
  assign n2186 = n2185 ^ n2062;
  assign n2267 = n2266 ^ n2186;
  assign n2176 = n372 & n1787;
  assign n2177 = x84 & n433;
  assign n2178 = x86 & n428;
  assign n2179 = ~n2177 & ~n2178;
  assign n2180 = x85 & n376;
  assign n2181 = n2179 & ~n2180;
  assign n2182 = ~n2176 & n2181;
  assign n2183 = n2182 ^ x8;
  assign n2268 = n2267 ^ n2183;
  assign n2173 = n2139 ^ n2051;
  assign n2174 = n2140 & n2173;
  assign n2175 = n2174 ^ n2051;
  assign n2269 = n2268 ^ n2175;
  assign n2164 = n1777 ^ x89;
  assign n2165 = n210 & n2164;
  assign n2166 = x87 & n219;
  assign n2167 = x88 & n214;
  assign n2168 = ~n2166 & ~n2167;
  assign n2169 = x89 & n259;
  assign n2170 = n2168 & ~n2169;
  assign n2171 = ~n2165 & n2170;
  assign n2172 = n2171 ^ x5;
  assign n2270 = n2269 ^ n2172;
  assign n2161 = n2141 ^ n2039;
  assign n2162 = ~n2142 & n2161;
  assign n2163 = n2162 ^ n2039;
  assign n2271 = n2270 ^ n2163;
  assign n2149 = x91 ^ x90;
  assign n2150 = ~n2025 & n2149;
  assign n2151 = n163 & ~n2150;
  assign n2152 = n2151 ^ x1;
  assign n2153 = n2152 ^ x92;
  assign n2154 = x0 & n2153;
  assign n2155 = ~x1 & x90;
  assign n2156 = ~x0 & ~n2155;
  assign n2157 = x1 & x91;
  assign n2158 = n2157 ^ x2;
  assign n2159 = n2156 & n2158;
  assign n2160 = ~n2154 & ~n2159;
  assign n2272 = n2271 ^ n2160;
  assign n2146 = n2143 ^ n2023;
  assign n2147 = n2144 & ~n2146;
  assign n2148 = n2147 ^ n2023;
  assign n2273 = n2272 ^ n2148;
  assign n2402 = n520 & n1624;
  assign n2403 = x70 & n1742;
  assign n2404 = x72 & n1744;
  assign n2405 = ~n2403 & ~n2404;
  assign n2406 = x71 & n1628;
  assign n2407 = n2405 & ~n2406;
  assign n2408 = ~n2402 & n2407;
  assign n2409 = n2408 ^ x23;
  assign n2370 = x29 ^ x28;
  assign n2371 = n2116 & n2370;
  assign n2372 = n208 & n2371;
  assign n2374 = x26 & x27;
  assign n2373 = ~x26 & ~x27;
  assign n2375 = n2374 ^ n2373;
  assign n2376 = x28 & n2375;
  assign n2377 = n2376 ^ n2374;
  assign n2378 = ~n2372 & ~n2377;
  assign n2379 = x65 & ~n2378;
  assign n2380 = n149 & n2370;
  assign n2381 = x66 & n2116;
  assign n2382 = ~n2380 & n2381;
  assign n2383 = ~n2379 & ~n2382;
  assign n2384 = x28 & x64;
  assign n2385 = n2373 & ~n2384;
  assign n2386 = ~n201 & ~n2385;
  assign n2387 = ~x28 & x64;
  assign n2388 = n2374 & ~n2387;
  assign n2389 = n2386 & ~n2388;
  assign n2390 = x29 & ~n2387;
  assign n2391 = ~n2389 & n2390;
  assign n2392 = n2383 & n2391;
  assign n2395 = x29 & n2389;
  assign n2393 = n2374 & n2384;
  assign n2394 = ~x29 & ~n2393;
  assign n2396 = n2395 ^ n2394;
  assign n2397 = n2383 & n2396;
  assign n2398 = n2397 ^ n2395;
  assign n2399 = ~n2392 & ~n2398;
  assign n2362 = n358 & n1969;
  assign n2363 = x68 & n1973;
  assign n2364 = x67 & n1978;
  assign n2365 = ~n2363 & ~n2364;
  assign n2366 = x69 & n2108;
  assign n2367 = n2365 & ~n2366;
  assign n2368 = ~n2362 & n2367;
  assign n2369 = n2368 ^ x26;
  assign n2400 = n2399 ^ n2369;
  assign n2359 = n2248 ^ n2245;
  assign n2360 = ~n2246 & ~n2359;
  assign n2361 = n2360 ^ n2248;
  assign n2401 = n2400 ^ n2361;
  assign n2410 = n2409 ^ n2401;
  assign n2356 = n2257 ^ n2230;
  assign n2357 = n2258 & ~n2356;
  assign n2358 = n2357 ^ n2230;
  assign n2411 = n2410 ^ n2358;
  assign n2348 = n720 & n1296;
  assign n2349 = x74 & n1300;
  assign n2350 = x75 & n1406;
  assign n2351 = ~n2349 & ~n2350;
  assign n2352 = x73 & n1403;
  assign n2353 = n2351 & ~n2352;
  assign n2354 = ~n2348 & n2353;
  assign n2355 = n2354 ^ x20;
  assign n2412 = n2411 ^ n2355;
  assign n2345 = n2259 ^ n2219;
  assign n2346 = ~n2260 & ~n2345;
  assign n2347 = n2346 ^ n2219;
  assign n2413 = n2412 ^ n2347;
  assign n2337 = n953 & n1008;
  assign n2338 = x76 & n1101;
  assign n2339 = x77 & n1012;
  assign n2340 = ~n2338 & ~n2339;
  assign n2341 = x78 & n1104;
  assign n2342 = n2340 & ~n2341;
  assign n2343 = ~n2337 & n2342;
  assign n2344 = n2343 ^ x17;
  assign n2414 = n2413 ^ n2344;
  assign n2334 = n2261 ^ n2208;
  assign n2335 = n2262 & n2334;
  assign n2336 = n2335 ^ n2208;
  assign n2415 = n2414 ^ n2336;
  assign n2326 = n752 & n1230;
  assign n2327 = x79 & n825;
  assign n2328 = x81 & n828;
  assign n2329 = ~n2327 & ~n2328;
  assign n2330 = x80 & n757;
  assign n2331 = n2329 & ~n2330;
  assign n2332 = ~n2326 & n2331;
  assign n2333 = n2332 ^ x14;
  assign n2416 = n2415 ^ n2333;
  assign n2323 = n2263 ^ n2197;
  assign n2324 = ~n2264 & ~n2323;
  assign n2325 = n2324 ^ n2197;
  assign n2417 = n2416 ^ n2325;
  assign n2315 = n541 & n1547;
  assign n2316 = x82 & n612;
  assign n2317 = x83 & n547;
  assign n2318 = ~n2316 & ~n2317;
  assign n2319 = x84 & n615;
  assign n2320 = n2318 & ~n2319;
  assign n2321 = ~n2315 & n2320;
  assign n2322 = n2321 ^ x11;
  assign n2418 = n2417 ^ n2322;
  assign n2312 = n2265 ^ n2186;
  assign n2313 = n2266 & n2312;
  assign n2314 = n2313 ^ n2186;
  assign n2419 = n2418 ^ n2314;
  assign n2304 = n372 & n1903;
  assign n2305 = x85 & n433;
  assign n2306 = x86 & n376;
  assign n2307 = ~n2305 & ~n2306;
  assign n2308 = x87 & n428;
  assign n2309 = n2307 & ~n2308;
  assign n2310 = ~n2304 & n2309;
  assign n2311 = n2310 ^ x8;
  assign n2420 = n2419 ^ n2311;
  assign n2301 = n2267 ^ n2175;
  assign n2302 = ~n2268 & ~n2301;
  assign n2303 = n2302 ^ n2175;
  assign n2421 = n2420 ^ n2303;
  assign n2292 = n1888 ^ x90;
  assign n2293 = n210 & n2292;
  assign n2294 = x88 & n219;
  assign n2295 = x89 & n214;
  assign n2296 = ~n2294 & ~n2295;
  assign n2297 = x90 & n259;
  assign n2298 = n2296 & ~n2297;
  assign n2299 = ~n2293 & n2298;
  assign n2300 = n2299 ^ x5;
  assign n2422 = n2421 ^ n2300;
  assign n2289 = n2269 ^ n2163;
  assign n2290 = n2270 & ~n2289;
  assign n2291 = n2290 ^ n2163;
  assign n2423 = n2422 ^ n2291;
  assign n2277 = x92 ^ x91;
  assign n2278 = ~n2150 & n2277;
  assign n2279 = n163 & ~n2278;
  assign n2280 = n2279 ^ x1;
  assign n2281 = n2280 ^ x93;
  assign n2282 = x0 & n2281;
  assign n2283 = ~x1 & x91;
  assign n2284 = ~x0 & ~n2283;
  assign n2285 = x1 & x92;
  assign n2286 = n2285 ^ x2;
  assign n2287 = n2284 & n2286;
  assign n2288 = ~n2282 & ~n2287;
  assign n2424 = n2423 ^ n2288;
  assign n2274 = n2271 ^ n2148;
  assign n2275 = n2272 & n2274;
  assign n2276 = n2275 ^ n2148;
  assign n2425 = n2424 ^ n2276;
  assign n2541 = n416 & n1969;
  assign n2542 = x68 & n1978;
  assign n2543 = x69 & n1973;
  assign n2544 = ~n2542 & ~n2543;
  assign n2545 = x70 & n2108;
  assign n2546 = n2544 & ~n2545;
  assign n2547 = ~n2541 & n2546;
  assign n2548 = n2547 ^ x26;
  assign n2537 = x30 ^ x29;
  assign n2538 = x64 & n2537;
  assign n2539 = n2538 ^ n2392;
  assign n2525 = x66 & n2377;
  assign n2526 = x28 ^ x27;
  assign n2527 = n2370 & ~n2526;
  assign n2528 = ~n2116 & n2527;
  assign n2529 = x65 & n2528;
  assign n2530 = ~n2525 & ~n2529;
  assign n2531 = n2116 & ~n2370;
  assign n2532 = x67 & n2531;
  assign n2533 = n2530 & ~n2532;
  assign n2534 = n264 & n2371;
  assign n2535 = n2533 & ~n2534;
  assign n2536 = n2535 ^ x29;
  assign n2540 = n2539 ^ n2536;
  assign n2549 = n2548 ^ n2540;
  assign n2522 = n2399 ^ n2361;
  assign n2523 = n2400 & n2522;
  assign n2524 = n2523 ^ n2361;
  assign n2550 = n2549 ^ n2524;
  assign n2514 = ~n594 & n1624;
  assign n2515 = x71 & n1742;
  assign n2516 = x73 & n1744;
  assign n2517 = ~n2515 & ~n2516;
  assign n2518 = x72 & n1628;
  assign n2519 = n2517 & ~n2518;
  assign n2520 = ~n2514 & n2519;
  assign n2521 = n2520 ^ x23;
  assign n2551 = n2550 ^ n2521;
  assign n2511 = n2409 ^ n2358;
  assign n2512 = ~n2410 & ~n2511;
  assign n2513 = n2512 ^ n2358;
  assign n2552 = n2551 ^ n2513;
  assign n2503 = n799 & n1296;
  assign n2504 = x75 & n1300;
  assign n2505 = x74 & n1403;
  assign n2506 = ~n2504 & ~n2505;
  assign n2507 = x76 & n1406;
  assign n2508 = n2506 & ~n2507;
  assign n2509 = ~n2503 & n2508;
  assign n2510 = n2509 ^ x20;
  assign n2553 = n2552 ^ n2510;
  assign n2500 = n2411 ^ n2347;
  assign n2501 = n2412 & n2500;
  assign n2502 = n2501 ^ n2347;
  assign n2554 = n2553 ^ n2502;
  assign n2492 = n1008 & n1054;
  assign n2493 = x77 & n1101;
  assign n2494 = x78 & n1012;
  assign n2495 = ~n2493 & ~n2494;
  assign n2496 = x79 & n1104;
  assign n2497 = n2495 & ~n2496;
  assign n2498 = ~n2492 & n2497;
  assign n2499 = n2498 ^ x17;
  assign n2555 = n2554 ^ n2499;
  assign n2489 = n2413 ^ n2336;
  assign n2490 = ~n2414 & ~n2489;
  assign n2491 = n2490 ^ n2336;
  assign n2556 = n2555 ^ n2491;
  assign n2481 = n752 & n1345;
  assign n2482 = x80 & n825;
  assign n2483 = x81 & n757;
  assign n2484 = ~n2482 & ~n2483;
  assign n2485 = x82 & n828;
  assign n2486 = n2484 & ~n2485;
  assign n2487 = ~n2481 & n2486;
  assign n2488 = n2487 ^ x14;
  assign n2557 = n2556 ^ n2488;
  assign n2478 = n2415 ^ n2325;
  assign n2479 = n2416 & n2478;
  assign n2480 = n2479 ^ n2325;
  assign n2558 = n2557 ^ n2480;
  assign n2470 = n541 & n1674;
  assign n2471 = x83 & n612;
  assign n2472 = x85 & n615;
  assign n2473 = ~n2471 & ~n2472;
  assign n2474 = x84 & n547;
  assign n2475 = n2473 & ~n2474;
  assign n2476 = ~n2470 & n2475;
  assign n2477 = n2476 ^ x11;
  assign n2559 = n2558 ^ n2477;
  assign n2467 = n2417 ^ n2314;
  assign n2468 = ~n2418 & ~n2467;
  assign n2469 = n2468 ^ n2314;
  assign n2560 = n2559 ^ n2469;
  assign n2459 = n372 & n2040;
  assign n2460 = x86 & n433;
  assign n2461 = x87 & n376;
  assign n2462 = ~n2460 & ~n2461;
  assign n2463 = x88 & n428;
  assign n2464 = n2462 & ~n2463;
  assign n2465 = ~n2459 & n2464;
  assign n2466 = n2465 ^ x8;
  assign n2561 = n2560 ^ n2466;
  assign n2456 = n2419 ^ n2303;
  assign n2457 = n2420 & n2456;
  assign n2458 = n2457 ^ n2303;
  assign n2562 = n2561 ^ n2458;
  assign n2447 = n2025 ^ x91;
  assign n2448 = n210 & n2447;
  assign n2449 = x89 & n219;
  assign n2450 = x91 & n259;
  assign n2451 = ~n2449 & ~n2450;
  assign n2452 = x90 & n214;
  assign n2453 = n2451 & ~n2452;
  assign n2454 = ~n2448 & n2453;
  assign n2455 = n2454 ^ x5;
  assign n2563 = n2562 ^ n2455;
  assign n2444 = n2421 ^ n2291;
  assign n2445 = ~n2422 & n2444;
  assign n2446 = n2445 ^ n2291;
  assign n2564 = n2563 ^ n2446;
  assign n2433 = x93 ^ x92;
  assign n2434 = x93 ^ x91;
  assign n2435 = ~n2150 & ~n2434;
  assign n2436 = n2433 & n2435;
  assign n2437 = n2436 ^ n2433;
  assign n2438 = n163 & ~n2437;
  assign n2439 = n2438 ^ x1;
  assign n2440 = n2439 ^ x94;
  assign n2429 = ~x92 & n156;
  assign n2430 = x93 ^ x2;
  assign n2431 = x1 & n2430;
  assign n2432 = ~n2429 & ~n2431;
  assign n2441 = n2440 ^ n2432;
  assign n2442 = ~x0 & ~n2441;
  assign n2443 = n2442 ^ n2440;
  assign n2565 = n2564 ^ n2443;
  assign n2426 = n2423 ^ n2276;
  assign n2427 = ~n2424 & ~n2426;
  assign n2428 = n2427 ^ n2276;
  assign n2566 = n2565 ^ n2428;
  assign n2682 = n467 & n1969;
  assign n2683 = x70 & n1973;
  assign n2684 = x69 & n1978;
  assign n2685 = ~n2683 & ~n2684;
  assign n2686 = x71 & n2108;
  assign n2687 = n2685 & ~n2686;
  assign n2688 = ~n2682 & n2687;
  assign n2689 = n2688 ^ x26;
  assign n2679 = n2548 ^ n2524;
  assign n2680 = ~n2549 & ~n2679;
  assign n2681 = n2680 ^ n2524;
  assign n2690 = n2689 ^ n2681;
  assign n2676 = ~n2392 & ~n2538;
  assign n2677 = ~n2536 & ~n2676;
  assign n2667 = n300 & n2371;
  assign n2668 = x66 & n2528;
  assign n2669 = x68 & n2531;
  assign n2670 = ~n2668 & ~n2669;
  assign n2671 = x67 & n2377;
  assign n2672 = n2670 & ~n2671;
  assign n2673 = ~n2667 & n2672;
  assign n2674 = n2673 ^ x29;
  assign n2660 = x65 ^ x30;
  assign n2661 = n2537 & ~n2660;
  assign n2662 = n2661 ^ x29;
  assign n2663 = n2662 ^ x31;
  assign n2664 = x64 & n2663;
  assign n2665 = n149 & n2537;
  assign n2666 = ~n2664 & ~n2665;
  assign n2675 = n2674 ^ n2666;
  assign n2678 = n2677 ^ n2675;
  assign n2691 = n2690 ^ n2678;
  assign n2652 = ~n656 & n1624;
  assign n2653 = x73 & n1628;
  assign n2654 = x72 & n1742;
  assign n2655 = ~n2653 & ~n2654;
  assign n2656 = x74 & n1744;
  assign n2657 = n2655 & ~n2656;
  assign n2658 = ~n2652 & n2657;
  assign n2659 = n2658 ^ x23;
  assign n2692 = n2691 ^ n2659;
  assign n2649 = n2550 ^ n2513;
  assign n2650 = n2551 & n2649;
  assign n2651 = n2650 ^ n2513;
  assign n2693 = n2692 ^ n2651;
  assign n2641 = n877 & n1296;
  assign n2642 = x75 & n1403;
  assign n2643 = x76 & n1300;
  assign n2644 = ~n2642 & ~n2643;
  assign n2645 = x77 & n1406;
  assign n2646 = n2644 & ~n2645;
  assign n2647 = ~n2641 & n2646;
  assign n2648 = n2647 ^ x20;
  assign n2694 = n2693 ^ n2648;
  assign n2638 = n2552 ^ n2502;
  assign n2639 = ~n2553 & ~n2638;
  assign n2640 = n2639 ^ n2502;
  assign n2695 = n2694 ^ n2640;
  assign n2630 = n1008 & ~n1141;
  assign n2631 = x78 & n1101;
  assign n2632 = x79 & n1012;
  assign n2633 = ~n2631 & ~n2632;
  assign n2634 = x80 & n1104;
  assign n2635 = n2633 & ~n2634;
  assign n2636 = ~n2630 & n2635;
  assign n2637 = n2636 ^ x17;
  assign n2696 = n2695 ^ n2637;
  assign n2627 = n2554 ^ n2491;
  assign n2628 = n2555 & n2627;
  assign n2629 = n2628 ^ n2491;
  assign n2697 = n2696 ^ n2629;
  assign n2619 = n752 & n1445;
  assign n2620 = x81 & n825;
  assign n2621 = x82 & n757;
  assign n2622 = ~n2620 & ~n2621;
  assign n2623 = x83 & n828;
  assign n2624 = n2622 & ~n2623;
  assign n2625 = ~n2619 & n2624;
  assign n2626 = n2625 ^ x14;
  assign n2698 = n2697 ^ n2626;
  assign n2616 = n2556 ^ n2480;
  assign n2617 = ~n2557 & ~n2616;
  assign n2618 = n2617 ^ n2480;
  assign n2699 = n2698 ^ n2618;
  assign n2608 = n541 & n1787;
  assign n2609 = x84 & n612;
  assign n2610 = x85 & n547;
  assign n2611 = ~n2609 & ~n2610;
  assign n2612 = x86 & n615;
  assign n2613 = n2611 & ~n2612;
  assign n2614 = ~n2608 & n2613;
  assign n2615 = n2614 ^ x11;
  assign n2700 = n2699 ^ n2615;
  assign n2605 = n2558 ^ n2469;
  assign n2606 = n2559 & n2605;
  assign n2607 = n2606 ^ n2469;
  assign n2701 = n2700 ^ n2607;
  assign n2597 = n372 & n2164;
  assign n2598 = x87 & n433;
  assign n2599 = x88 & n376;
  assign n2600 = ~n2598 & ~n2599;
  assign n2601 = x89 & n428;
  assign n2602 = n2600 & ~n2601;
  assign n2603 = ~n2597 & n2602;
  assign n2604 = n2603 ^ x8;
  assign n2702 = n2701 ^ n2604;
  assign n2594 = n2560 ^ n2458;
  assign n2595 = ~n2561 & ~n2594;
  assign n2596 = n2595 ^ n2458;
  assign n2703 = n2702 ^ n2596;
  assign n2585 = n2150 ^ x92;
  assign n2586 = n210 & n2585;
  assign n2587 = x90 & n219;
  assign n2588 = x91 & n214;
  assign n2589 = ~n2587 & ~n2588;
  assign n2590 = x92 & n259;
  assign n2591 = n2589 & ~n2590;
  assign n2592 = ~n2586 & n2591;
  assign n2593 = n2592 ^ x5;
  assign n2704 = n2703 ^ n2593;
  assign n2582 = n2562 ^ n2446;
  assign n2583 = n2563 & ~n2582;
  assign n2584 = n2583 ^ n2446;
  assign n2705 = n2704 ^ n2584;
  assign n2570 = x94 ^ x93;
  assign n2571 = ~n2437 & n2570;
  assign n2572 = n163 & ~n2571;
  assign n2573 = n2572 ^ x1;
  assign n2574 = n2573 ^ x95;
  assign n2575 = x0 & n2574;
  assign n2576 = ~x1 & x93;
  assign n2577 = ~x0 & ~n2576;
  assign n2578 = x1 & x94;
  assign n2579 = n2578 ^ x2;
  assign n2580 = n2577 & n2579;
  assign n2581 = ~n2575 & ~n2580;
  assign n2706 = n2705 ^ n2581;
  assign n2567 = n2564 ^ n2428;
  assign n2568 = ~n2565 & n2567;
  assign n2569 = n2568 ^ n2428;
  assign n2707 = n2706 ^ n2569;
  assign n2823 = ~x29 & ~x30;
  assign n2832 = ~x31 & x32;
  assign n2833 = n2823 & n2832;
  assign n2834 = x64 & n2833;
  assign n2835 = x32 ^ x31;
  assign n2836 = n2537 & n2835;
  assign n2837 = n208 & n2836;
  assign n2827 = x29 & x30;
  assign n2838 = n2827 ^ n2823;
  assign n2839 = ~x31 & n2838;
  assign n2840 = n2839 ^ n2823;
  assign n2841 = ~n2837 & ~n2840;
  assign n2842 = x65 & ~n2841;
  assign n2843 = n149 & n2835;
  assign n2844 = x66 & n2537;
  assign n2845 = ~n2843 & n2844;
  assign n2846 = ~n2842 & ~n2845;
  assign n2847 = n2846 ^ x32;
  assign n2824 = x31 & x64;
  assign n2848 = n2824 & n2827;
  assign n2849 = n2846 & n2848;
  assign n2850 = n2847 & n2849;
  assign n2851 = n2850 ^ n2847;
  assign n2852 = ~n2834 & ~n2851;
  assign n2825 = n2823 & ~n2824;
  assign n2826 = ~n201 & ~n2825;
  assign n2828 = ~x31 & x64;
  assign n2829 = n2827 & ~n2828;
  assign n2830 = n2826 & ~n2829;
  assign n2831 = x32 & ~n2830;
  assign n2853 = n2852 ^ n2831;
  assign n2815 = n358 & n2371;
  assign n2816 = x67 & n2528;
  assign n2817 = x69 & n2531;
  assign n2818 = ~n2816 & ~n2817;
  assign n2819 = x68 & n2377;
  assign n2820 = n2818 & ~n2819;
  assign n2821 = ~n2815 & n2820;
  assign n2822 = n2821 ^ x29;
  assign n2854 = n2853 ^ n2822;
  assign n2812 = n2677 ^ n2674;
  assign n2813 = ~n2675 & ~n2812;
  assign n2814 = n2813 ^ n2677;
  assign n2855 = n2854 ^ n2814;
  assign n2804 = n520 & n1969;
  assign n2805 = x71 & n1973;
  assign n2806 = x70 & n1978;
  assign n2807 = ~n2805 & ~n2806;
  assign n2808 = x72 & n2108;
  assign n2809 = n2807 & ~n2808;
  assign n2810 = ~n2804 & n2809;
  assign n2811 = n2810 ^ x26;
  assign n2856 = n2855 ^ n2811;
  assign n2801 = n2689 ^ n2678;
  assign n2802 = ~n2690 & n2801;
  assign n2803 = n2802 ^ n2681;
  assign n2857 = n2856 ^ n2803;
  assign n2793 = n720 & n1624;
  assign n2794 = x73 & n1742;
  assign n2795 = x74 & n1628;
  assign n2796 = ~n2794 & ~n2795;
  assign n2797 = x75 & n1744;
  assign n2798 = n2796 & ~n2797;
  assign n2799 = ~n2793 & n2798;
  assign n2800 = n2799 ^ x23;
  assign n2858 = n2857 ^ n2800;
  assign n2790 = n2691 ^ n2651;
  assign n2791 = ~n2692 & ~n2790;
  assign n2792 = n2791 ^ n2651;
  assign n2859 = n2858 ^ n2792;
  assign n2782 = n953 & n1296;
  assign n2783 = x76 & n1403;
  assign n2784 = x77 & n1300;
  assign n2785 = ~n2783 & ~n2784;
  assign n2786 = x78 & n1406;
  assign n2787 = n2785 & ~n2786;
  assign n2788 = ~n2782 & n2787;
  assign n2789 = n2788 ^ x20;
  assign n2860 = n2859 ^ n2789;
  assign n2779 = n2693 ^ n2640;
  assign n2780 = n2694 & n2779;
  assign n2781 = n2780 ^ n2640;
  assign n2861 = n2860 ^ n2781;
  assign n2771 = n1008 & n1230;
  assign n2772 = x79 & n1101;
  assign n2773 = x80 & n1012;
  assign n2774 = ~n2772 & ~n2773;
  assign n2775 = x81 & n1104;
  assign n2776 = n2774 & ~n2775;
  assign n2777 = ~n2771 & n2776;
  assign n2778 = n2777 ^ x17;
  assign n2862 = n2861 ^ n2778;
  assign n2768 = n2695 ^ n2629;
  assign n2769 = ~n2696 & ~n2768;
  assign n2770 = n2769 ^ n2629;
  assign n2863 = n2862 ^ n2770;
  assign n2760 = n752 & n1547;
  assign n2761 = x82 & n825;
  assign n2762 = x84 & n828;
  assign n2763 = ~n2761 & ~n2762;
  assign n2764 = x83 & n757;
  assign n2765 = n2763 & ~n2764;
  assign n2766 = ~n2760 & n2765;
  assign n2767 = n2766 ^ x14;
  assign n2864 = n2863 ^ n2767;
  assign n2757 = n2697 ^ n2618;
  assign n2758 = n2698 & n2757;
  assign n2759 = n2758 ^ n2618;
  assign n2865 = n2864 ^ n2759;
  assign n2749 = n541 & n1903;
  assign n2750 = x85 & n612;
  assign n2751 = x87 & n615;
  assign n2752 = ~n2750 & ~n2751;
  assign n2753 = x86 & n547;
  assign n2754 = n2752 & ~n2753;
  assign n2755 = ~n2749 & n2754;
  assign n2756 = n2755 ^ x11;
  assign n2866 = n2865 ^ n2756;
  assign n2746 = n2699 ^ n2607;
  assign n2747 = ~n2700 & ~n2746;
  assign n2748 = n2747 ^ n2607;
  assign n2867 = n2866 ^ n2748;
  assign n2738 = n372 & n2292;
  assign n2739 = x89 & n376;
  assign n2740 = x88 & n433;
  assign n2741 = ~n2739 & ~n2740;
  assign n2742 = x90 & n428;
  assign n2743 = n2741 & ~n2742;
  assign n2744 = ~n2738 & n2743;
  assign n2745 = n2744 ^ x8;
  assign n2868 = n2867 ^ n2745;
  assign n2735 = n2701 ^ n2596;
  assign n2736 = n2702 & n2735;
  assign n2737 = n2736 ^ n2596;
  assign n2869 = n2868 ^ n2737;
  assign n2726 = n2278 ^ x93;
  assign n2727 = n210 & n2726;
  assign n2728 = x91 & n219;
  assign n2729 = x92 & n214;
  assign n2730 = ~n2728 & ~n2729;
  assign n2731 = x93 & n259;
  assign n2732 = n2730 & ~n2731;
  assign n2733 = ~n2727 & n2732;
  assign n2734 = n2733 ^ x5;
  assign n2870 = n2869 ^ n2734;
  assign n2723 = n2703 ^ n2584;
  assign n2724 = ~n2704 & n2723;
  assign n2725 = n2724 ^ n2584;
  assign n2871 = n2870 ^ n2725;
  assign n2715 = x95 ^ x94;
  assign n2716 = ~n2571 & n2715;
  assign n2717 = n163 & ~n2716;
  assign n2718 = n2717 ^ x1;
  assign n2719 = n2718 ^ x96;
  assign n2711 = x1 & x95;
  assign n2712 = n2711 ^ x2;
  assign n2713 = ~x1 & x94;
  assign n2714 = n2712 & ~n2713;
  assign n2720 = n2719 ^ n2714;
  assign n2721 = ~x0 & n2720;
  assign n2722 = n2721 ^ n2719;
  assign n2872 = n2871 ^ n2722;
  assign n2708 = n2705 ^ n2569;
  assign n2709 = ~n2706 & ~n2708;
  assign n2710 = n2709 ^ n2569;
  assign n2873 = n2872 ^ n2710;
  assign n3007 = n2831 & n2852;
  assign n2994 = x31 ^ x30;
  assign n2995 = n2835 & ~n2994;
  assign n2996 = ~n2537 & n2995;
  assign n2997 = x65 & n2996;
  assign n2998 = n2537 & ~n2835;
  assign n2999 = x67 & n2998;
  assign n3000 = ~n2997 & ~n2999;
  assign n3001 = x66 & n2840;
  assign n3002 = n3000 & ~n3001;
  assign n3003 = n264 & n2836;
  assign n3004 = n3002 & ~n3003;
  assign n3005 = n3004 ^ x32;
  assign n2992 = x33 ^ x32;
  assign n2993 = x64 & n2992;
  assign n3006 = n3005 ^ n2993;
  assign n3008 = n3007 ^ n3006;
  assign n2984 = n416 & n2371;
  assign n2985 = x69 & n2377;
  assign n2986 = x68 & n2528;
  assign n2987 = ~n2985 & ~n2986;
  assign n2988 = x70 & n2531;
  assign n2989 = n2987 & ~n2988;
  assign n2990 = ~n2984 & n2989;
  assign n2991 = n2990 ^ x29;
  assign n3009 = n3008 ^ n2991;
  assign n2981 = n2853 ^ n2814;
  assign n2982 = n2854 & n2981;
  assign n2983 = n2982 ^ n2814;
  assign n3010 = n3009 ^ n2983;
  assign n2973 = ~n594 & n1969;
  assign n2974 = x72 & n1973;
  assign n2975 = x71 & n1978;
  assign n2976 = ~n2974 & ~n2975;
  assign n2977 = x73 & n2108;
  assign n2978 = n2976 & ~n2977;
  assign n2979 = ~n2973 & n2978;
  assign n2980 = n2979 ^ x26;
  assign n3011 = n3010 ^ n2980;
  assign n2970 = n2855 ^ n2803;
  assign n2971 = ~n2856 & ~n2970;
  assign n2972 = n2971 ^ n2803;
  assign n3012 = n3011 ^ n2972;
  assign n2962 = n799 & n1624;
  assign n2963 = x74 & n1742;
  assign n2964 = x76 & n1744;
  assign n2965 = ~n2963 & ~n2964;
  assign n2966 = x75 & n1628;
  assign n2967 = n2965 & ~n2966;
  assign n2968 = ~n2962 & n2967;
  assign n2969 = n2968 ^ x23;
  assign n3013 = n3012 ^ n2969;
  assign n2959 = n2857 ^ n2792;
  assign n2960 = n2858 & n2959;
  assign n2961 = n2960 ^ n2792;
  assign n3014 = n3013 ^ n2961;
  assign n2951 = n1054 & n1296;
  assign n2952 = x77 & n1403;
  assign n2953 = x78 & n1300;
  assign n2954 = ~n2952 & ~n2953;
  assign n2955 = x79 & n1406;
  assign n2956 = n2954 & ~n2955;
  assign n2957 = ~n2951 & n2956;
  assign n2958 = n2957 ^ x20;
  assign n3015 = n3014 ^ n2958;
  assign n2948 = n2859 ^ n2781;
  assign n2949 = ~n2860 & ~n2948;
  assign n2950 = n2949 ^ n2781;
  assign n3016 = n3015 ^ n2950;
  assign n2940 = n1008 & n1345;
  assign n2941 = x80 & n1101;
  assign n2942 = x81 & n1012;
  assign n2943 = ~n2941 & ~n2942;
  assign n2944 = x82 & n1104;
  assign n2945 = n2943 & ~n2944;
  assign n2946 = ~n2940 & n2945;
  assign n2947 = n2946 ^ x17;
  assign n3017 = n3016 ^ n2947;
  assign n2937 = n2861 ^ n2770;
  assign n2938 = n2862 & n2937;
  assign n2939 = n2938 ^ n2770;
  assign n3018 = n3017 ^ n2939;
  assign n2929 = n752 & n1674;
  assign n2930 = x83 & n825;
  assign n2931 = x85 & n828;
  assign n2932 = ~n2930 & ~n2931;
  assign n2933 = x84 & n757;
  assign n2934 = n2932 & ~n2933;
  assign n2935 = ~n2929 & n2934;
  assign n2936 = n2935 ^ x14;
  assign n3019 = n3018 ^ n2936;
  assign n2926 = n2863 ^ n2759;
  assign n2927 = ~n2864 & ~n2926;
  assign n2928 = n2927 ^ n2759;
  assign n3020 = n3019 ^ n2928;
  assign n2918 = n541 & n2040;
  assign n2919 = x86 & n612;
  assign n2920 = x87 & n547;
  assign n2921 = ~n2919 & ~n2920;
  assign n2922 = x88 & n615;
  assign n2923 = n2921 & ~n2922;
  assign n2924 = ~n2918 & n2923;
  assign n2925 = n2924 ^ x11;
  assign n3021 = n3020 ^ n2925;
  assign n2915 = n2865 ^ n2748;
  assign n2916 = n2866 & n2915;
  assign n2917 = n2916 ^ n2748;
  assign n3022 = n3021 ^ n2917;
  assign n2907 = n372 & n2447;
  assign n2908 = x89 & n433;
  assign n2909 = x91 & n428;
  assign n2910 = ~n2908 & ~n2909;
  assign n2911 = x90 & n376;
  assign n2912 = n2910 & ~n2911;
  assign n2913 = ~n2907 & n2912;
  assign n2914 = n2913 ^ x8;
  assign n3023 = n3022 ^ n2914;
  assign n2904 = n2867 ^ n2737;
  assign n2905 = ~n2868 & ~n2904;
  assign n2906 = n2905 ^ n2737;
  assign n3024 = n3023 ^ n2906;
  assign n2895 = n2437 ^ x94;
  assign n2896 = n210 & n2895;
  assign n2897 = x92 & n219;
  assign n2898 = x94 & n259;
  assign n2899 = ~n2897 & ~n2898;
  assign n2900 = x93 & n214;
  assign n2901 = n2899 & ~n2900;
  assign n2902 = ~n2896 & n2901;
  assign n2903 = n2902 ^ x5;
  assign n3025 = n3024 ^ n2903;
  assign n2892 = n2869 ^ n2725;
  assign n2893 = n2870 & ~n2892;
  assign n2894 = n2893 ^ n2725;
  assign n3026 = n3025 ^ n2894;
  assign n2881 = x96 ^ x95;
  assign n2882 = x96 ^ x94;
  assign n2883 = ~n2571 & ~n2882;
  assign n2884 = n2881 & n2883;
  assign n2885 = n2884 ^ n2881;
  assign n2886 = n163 & ~n2885;
  assign n2887 = n2886 ^ x1;
  assign n2888 = n2887 ^ x97;
  assign n2877 = ~x95 & n156;
  assign n2878 = x96 ^ x2;
  assign n2879 = x1 & n2878;
  assign n2880 = ~n2877 & ~n2879;
  assign n2889 = n2888 ^ n2880;
  assign n2890 = ~x0 & ~n2889;
  assign n2891 = n2890 ^ n2888;
  assign n3027 = n3026 ^ n2891;
  assign n2874 = n2871 ^ n2710;
  assign n2875 = ~n2872 & n2874;
  assign n2876 = n2875 ^ n2710;
  assign n3028 = n3027 ^ n2876;
  assign n3167 = ~n2993 & ~n3007;
  assign n3168 = ~n3005 & ~n3167;
  assign n3158 = n300 & n2836;
  assign n3159 = x67 & n2840;
  assign n3160 = x66 & n2996;
  assign n3161 = ~n3159 & ~n3160;
  assign n3162 = x68 & n2998;
  assign n3163 = n3161 & ~n3162;
  assign n3164 = ~n3158 & n3163;
  assign n3165 = n3164 ^ x32;
  assign n3151 = x65 ^ x33;
  assign n3152 = n2992 & ~n3151;
  assign n3153 = n3152 ^ x32;
  assign n3154 = n3153 ^ x34;
  assign n3155 = x64 & n3154;
  assign n3156 = n149 & n2992;
  assign n3157 = ~n3155 & ~n3156;
  assign n3166 = n3165 ^ n3157;
  assign n3169 = n3168 ^ n3166;
  assign n3143 = n467 & n2371;
  assign n3144 = x69 & n2528;
  assign n3145 = x71 & n2531;
  assign n3146 = ~n3144 & ~n3145;
  assign n3147 = x70 & n2377;
  assign n3148 = n3146 & ~n3147;
  assign n3149 = ~n3143 & n3148;
  assign n3150 = n3149 ^ x29;
  assign n3170 = n3169 ^ n3150;
  assign n3140 = n3008 ^ n2983;
  assign n3141 = ~n3009 & ~n3140;
  assign n3142 = n3141 ^ n2983;
  assign n3171 = n3170 ^ n3142;
  assign n3132 = ~n656 & n1969;
  assign n3133 = x73 & n1973;
  assign n3134 = x72 & n1978;
  assign n3135 = ~n3133 & ~n3134;
  assign n3136 = x74 & n2108;
  assign n3137 = n3135 & ~n3136;
  assign n3138 = ~n3132 & n3137;
  assign n3139 = n3138 ^ x26;
  assign n3172 = n3171 ^ n3139;
  assign n3129 = n3010 ^ n2972;
  assign n3130 = n3011 & n3129;
  assign n3131 = n3130 ^ n2972;
  assign n3173 = n3172 ^ n3131;
  assign n3121 = n877 & n1624;
  assign n3122 = x75 & n1742;
  assign n3123 = x76 & n1628;
  assign n3124 = ~n3122 & ~n3123;
  assign n3125 = x77 & n1744;
  assign n3126 = n3124 & ~n3125;
  assign n3127 = ~n3121 & n3126;
  assign n3128 = n3127 ^ x23;
  assign n3174 = n3173 ^ n3128;
  assign n3118 = n3012 ^ n2961;
  assign n3119 = ~n3013 & ~n3118;
  assign n3120 = n3119 ^ n2961;
  assign n3175 = n3174 ^ n3120;
  assign n3110 = ~n1141 & n1296;
  assign n3111 = x78 & n1403;
  assign n3112 = x79 & n1300;
  assign n3113 = ~n3111 & ~n3112;
  assign n3114 = x80 & n1406;
  assign n3115 = n3113 & ~n3114;
  assign n3116 = ~n3110 & n3115;
  assign n3117 = n3116 ^ x20;
  assign n3176 = n3175 ^ n3117;
  assign n3107 = n3014 ^ n2950;
  assign n3108 = n3015 & n3107;
  assign n3109 = n3108 ^ n2950;
  assign n3177 = n3176 ^ n3109;
  assign n3099 = n1008 & n1445;
  assign n3100 = x82 & n1012;
  assign n3101 = x81 & n1101;
  assign n3102 = ~n3100 & ~n3101;
  assign n3103 = x83 & n1104;
  assign n3104 = n3102 & ~n3103;
  assign n3105 = ~n3099 & n3104;
  assign n3106 = n3105 ^ x17;
  assign n3178 = n3177 ^ n3106;
  assign n3096 = n3016 ^ n2939;
  assign n3097 = ~n3017 & ~n3096;
  assign n3098 = n3097 ^ n2939;
  assign n3179 = n3178 ^ n3098;
  assign n3088 = n752 & n1787;
  assign n3089 = x84 & n825;
  assign n3090 = x85 & n757;
  assign n3091 = ~n3089 & ~n3090;
  assign n3092 = x86 & n828;
  assign n3093 = n3091 & ~n3092;
  assign n3094 = ~n3088 & n3093;
  assign n3095 = n3094 ^ x14;
  assign n3180 = n3179 ^ n3095;
  assign n3085 = n3018 ^ n2928;
  assign n3086 = n3019 & n3085;
  assign n3087 = n3086 ^ n2928;
  assign n3181 = n3180 ^ n3087;
  assign n3077 = n541 & n2164;
  assign n3078 = x87 & n612;
  assign n3079 = x89 & n615;
  assign n3080 = ~n3078 & ~n3079;
  assign n3081 = x88 & n547;
  assign n3082 = n3080 & ~n3081;
  assign n3083 = ~n3077 & n3082;
  assign n3084 = n3083 ^ x11;
  assign n3182 = n3181 ^ n3084;
  assign n3074 = n3020 ^ n2917;
  assign n3075 = ~n3021 & ~n3074;
  assign n3076 = n3075 ^ n2917;
  assign n3183 = n3182 ^ n3076;
  assign n3066 = n372 & n2585;
  assign n3067 = x90 & n433;
  assign n3068 = x91 & n376;
  assign n3069 = ~n3067 & ~n3068;
  assign n3070 = x92 & n428;
  assign n3071 = n3069 & ~n3070;
  assign n3072 = ~n3066 & n3071;
  assign n3073 = n3072 ^ x8;
  assign n3184 = n3183 ^ n3073;
  assign n3063 = n3022 ^ n2906;
  assign n3064 = n3023 & n3063;
  assign n3065 = n3064 ^ n2906;
  assign n3185 = n3184 ^ n3065;
  assign n3054 = n2571 ^ x95;
  assign n3055 = n210 & n3054;
  assign n3056 = x93 & n219;
  assign n3057 = x94 & n214;
  assign n3058 = ~n3056 & ~n3057;
  assign n3059 = x95 & n259;
  assign n3060 = n3058 & ~n3059;
  assign n3061 = ~n3055 & n3060;
  assign n3062 = n3061 ^ x5;
  assign n3186 = n3185 ^ n3062;
  assign n3051 = n3024 ^ n2894;
  assign n3052 = ~n3025 & n3051;
  assign n3053 = n3052 ^ n2894;
  assign n3187 = n3186 ^ n3053;
  assign n3032 = ~x94 & ~n2571;
  assign n3033 = x95 & x97;
  assign n3034 = ~n3032 & n3033;
  assign n3035 = ~x96 & ~n3034;
  assign n3036 = x94 & ~n2571;
  assign n3037 = ~x95 & ~x97;
  assign n3038 = ~n3036 & n3037;
  assign n3039 = ~n3035 & ~n3038;
  assign n3040 = n3039 ^ x97;
  assign n3041 = n163 & ~n3040;
  assign n3042 = n3041 ^ x1;
  assign n3043 = n3042 ^ x98;
  assign n3044 = x0 & ~n3043;
  assign n3045 = x97 ^ x2;
  assign n3046 = x1 & n3045;
  assign n3047 = ~x0 & ~n3046;
  assign n3048 = ~x96 & n156;
  assign n3049 = n3047 & ~n3048;
  assign n3050 = ~n3044 & ~n3049;
  assign n3188 = n3187 ^ n3050;
  assign n3029 = n3026 ^ n2876;
  assign n3030 = n3027 & ~n3029;
  assign n3031 = n3030 ^ n2876;
  assign n3189 = n3188 ^ n3031;
  assign n3317 = ~x32 & ~x33;
  assign n3326 = ~x34 & x35;
  assign n3327 = n3317 & n3326;
  assign n3328 = x64 & n3327;
  assign n3329 = x35 ^ x34;
  assign n3330 = n2992 & n3329;
  assign n3331 = n208 & n3330;
  assign n3321 = x32 & x33;
  assign n3332 = n3321 ^ n3317;
  assign n3333 = x34 & n3332;
  assign n3334 = n3333 ^ n3321;
  assign n3335 = ~n3331 & ~n3334;
  assign n3336 = x65 & ~n3335;
  assign n3337 = n149 & n3329;
  assign n3338 = x66 & n2992;
  assign n3339 = ~n3337 & n3338;
  assign n3340 = ~n3336 & ~n3339;
  assign n3341 = n3340 ^ x35;
  assign n3318 = x34 & x64;
  assign n3342 = n3318 & n3321;
  assign n3343 = n3340 & n3342;
  assign n3344 = n3341 & n3343;
  assign n3345 = n3344 ^ n3341;
  assign n3346 = ~n3328 & ~n3345;
  assign n3319 = n3317 & ~n3318;
  assign n3320 = ~n201 & ~n3319;
  assign n3322 = ~x34 & x64;
  assign n3323 = n3321 & ~n3322;
  assign n3324 = n3320 & ~n3323;
  assign n3325 = x35 & ~n3324;
  assign n3347 = n3346 ^ n3325;
  assign n3309 = n358 & n2836;
  assign n3310 = x68 & n2840;
  assign n3311 = x67 & n2996;
  assign n3312 = ~n3310 & ~n3311;
  assign n3313 = x69 & n2998;
  assign n3314 = n3312 & ~n3313;
  assign n3315 = ~n3309 & n3314;
  assign n3316 = n3315 ^ x32;
  assign n3348 = n3347 ^ n3316;
  assign n3306 = n3168 ^ n3165;
  assign n3307 = ~n3166 & ~n3306;
  assign n3308 = n3307 ^ n3168;
  assign n3349 = n3348 ^ n3308;
  assign n3298 = n520 & n2371;
  assign n3299 = x70 & n2528;
  assign n3300 = x72 & n2531;
  assign n3301 = ~n3299 & ~n3300;
  assign n3302 = x71 & n2377;
  assign n3303 = n3301 & ~n3302;
  assign n3304 = ~n3298 & n3303;
  assign n3305 = n3304 ^ x29;
  assign n3350 = n3349 ^ n3305;
  assign n3295 = n3169 ^ n3142;
  assign n3296 = n3170 & n3295;
  assign n3297 = n3296 ^ n3142;
  assign n3351 = n3350 ^ n3297;
  assign n3287 = n720 & n1969;
  assign n3288 = x73 & n1978;
  assign n3289 = x74 & n1973;
  assign n3290 = ~n3288 & ~n3289;
  assign n3291 = x75 & n2108;
  assign n3292 = n3290 & ~n3291;
  assign n3293 = ~n3287 & n3292;
  assign n3294 = n3293 ^ x26;
  assign n3352 = n3351 ^ n3294;
  assign n3284 = n3171 ^ n3131;
  assign n3285 = ~n3172 & ~n3284;
  assign n3286 = n3285 ^ n3131;
  assign n3353 = n3352 ^ n3286;
  assign n3276 = n953 & n1624;
  assign n3277 = x76 & n1742;
  assign n3278 = x78 & n1744;
  assign n3279 = ~n3277 & ~n3278;
  assign n3280 = x77 & n1628;
  assign n3281 = n3279 & ~n3280;
  assign n3282 = ~n3276 & n3281;
  assign n3283 = n3282 ^ x23;
  assign n3354 = n3353 ^ n3283;
  assign n3273 = n3173 ^ n3120;
  assign n3274 = n3174 & n3273;
  assign n3275 = n3274 ^ n3120;
  assign n3355 = n3354 ^ n3275;
  assign n3265 = n1230 & n1296;
  assign n3266 = x79 & n1403;
  assign n3267 = x81 & n1406;
  assign n3268 = ~n3266 & ~n3267;
  assign n3269 = x80 & n1300;
  assign n3270 = n3268 & ~n3269;
  assign n3271 = ~n3265 & n3270;
  assign n3272 = n3271 ^ x20;
  assign n3356 = n3355 ^ n3272;
  assign n3262 = n3175 ^ n3109;
  assign n3263 = ~n3176 & ~n3262;
  assign n3264 = n3263 ^ n3109;
  assign n3357 = n3356 ^ n3264;
  assign n3254 = n1008 & n1547;
  assign n3255 = x83 & n1012;
  assign n3256 = x82 & n1101;
  assign n3257 = ~n3255 & ~n3256;
  assign n3258 = x84 & n1104;
  assign n3259 = n3257 & ~n3258;
  assign n3260 = ~n3254 & n3259;
  assign n3261 = n3260 ^ x17;
  assign n3358 = n3357 ^ n3261;
  assign n3251 = n3177 ^ n3098;
  assign n3252 = n3178 & n3251;
  assign n3253 = n3252 ^ n3098;
  assign n3359 = n3358 ^ n3253;
  assign n3243 = n752 & n1903;
  assign n3244 = x85 & n825;
  assign n3245 = x86 & n757;
  assign n3246 = ~n3244 & ~n3245;
  assign n3247 = x87 & n828;
  assign n3248 = n3246 & ~n3247;
  assign n3249 = ~n3243 & n3248;
  assign n3250 = n3249 ^ x14;
  assign n3360 = n3359 ^ n3250;
  assign n3240 = n3179 ^ n3087;
  assign n3241 = ~n3180 & ~n3240;
  assign n3242 = n3241 ^ n3087;
  assign n3361 = n3360 ^ n3242;
  assign n3232 = n541 & n2292;
  assign n3233 = x88 & n612;
  assign n3234 = x90 & n615;
  assign n3235 = ~n3233 & ~n3234;
  assign n3236 = x89 & n547;
  assign n3237 = n3235 & ~n3236;
  assign n3238 = ~n3232 & n3237;
  assign n3239 = n3238 ^ x11;
  assign n3362 = n3361 ^ n3239;
  assign n3229 = n3181 ^ n3076;
  assign n3230 = n3182 & n3229;
  assign n3231 = n3230 ^ n3076;
  assign n3363 = n3362 ^ n3231;
  assign n3221 = n372 & n2726;
  assign n3222 = x91 & n433;
  assign n3223 = x93 & n428;
  assign n3224 = ~n3222 & ~n3223;
  assign n3225 = x92 & n376;
  assign n3226 = n3224 & ~n3225;
  assign n3227 = ~n3221 & n3226;
  assign n3228 = n3227 ^ x8;
  assign n3364 = n3363 ^ n3228;
  assign n3218 = n3183 ^ n3065;
  assign n3219 = ~n3184 & ~n3218;
  assign n3220 = n3219 ^ n3065;
  assign n3365 = n3364 ^ n3220;
  assign n3209 = n2716 ^ x96;
  assign n3210 = n210 & n3209;
  assign n3211 = x94 & n219;
  assign n3212 = x95 & n214;
  assign n3213 = ~n3211 & ~n3212;
  assign n3214 = x96 & n259;
  assign n3215 = n3213 & ~n3214;
  assign n3216 = ~n3210 & n3215;
  assign n3217 = n3216 ^ x5;
  assign n3366 = n3365 ^ n3217;
  assign n3206 = n3185 ^ n3053;
  assign n3207 = n3186 & ~n3206;
  assign n3208 = n3207 ^ n3053;
  assign n3367 = n3366 ^ n3208;
  assign n3198 = x98 ^ x97;
  assign n3199 = ~n3040 & n3198;
  assign n3200 = n163 & ~n3199;
  assign n3201 = n3200 ^ x1;
  assign n3202 = n3201 ^ x99;
  assign n3194 = x2 & ~x97;
  assign n3193 = x98 ^ x2;
  assign n3195 = n3194 ^ n3193;
  assign n3196 = x1 & n3195;
  assign n3197 = n3196 ^ n3194;
  assign n3203 = n3202 ^ n3197;
  assign n3204 = ~x0 & n3203;
  assign n3205 = n3204 ^ n3202;
  assign n3368 = n3367 ^ n3205;
  assign n3190 = n3187 ^ n3031;
  assign n3191 = ~n3188 & n3190;
  assign n3192 = n3191 ^ n3031;
  assign n3369 = n3368 ^ n3192;
  assign n3511 = n3325 & n3346;
  assign n3498 = x34 ^ x33;
  assign n3499 = n3329 & ~n3498;
  assign n3500 = ~n2992 & n3499;
  assign n3501 = x65 & n3500;
  assign n3502 = n2992 & ~n3329;
  assign n3503 = x67 & n3502;
  assign n3504 = ~n3501 & ~n3503;
  assign n3505 = x66 & n3334;
  assign n3506 = n3504 & ~n3505;
  assign n3507 = n264 & n3330;
  assign n3508 = n3506 & ~n3507;
  assign n3509 = n3508 ^ x35;
  assign n3496 = x36 ^ x35;
  assign n3497 = x64 & n3496;
  assign n3510 = n3509 ^ n3497;
  assign n3512 = n3511 ^ n3510;
  assign n3488 = n416 & n2836;
  assign n3489 = x68 & n2996;
  assign n3490 = x70 & n2998;
  assign n3491 = ~n3489 & ~n3490;
  assign n3492 = x69 & n2840;
  assign n3493 = n3491 & ~n3492;
  assign n3494 = ~n3488 & n3493;
  assign n3495 = n3494 ^ x32;
  assign n3513 = n3512 ^ n3495;
  assign n3485 = n3347 ^ n3308;
  assign n3486 = n3348 & n3485;
  assign n3487 = n3486 ^ n3308;
  assign n3514 = n3513 ^ n3487;
  assign n3477 = ~n594 & n2371;
  assign n3478 = x71 & n2528;
  assign n3479 = x73 & n2531;
  assign n3480 = ~n3478 & ~n3479;
  assign n3481 = x72 & n2377;
  assign n3482 = n3480 & ~n3481;
  assign n3483 = ~n3477 & n3482;
  assign n3484 = n3483 ^ x29;
  assign n3515 = n3514 ^ n3484;
  assign n3474 = n3349 ^ n3297;
  assign n3475 = ~n3350 & ~n3474;
  assign n3476 = n3475 ^ n3297;
  assign n3516 = n3515 ^ n3476;
  assign n3466 = n799 & n1969;
  assign n3467 = x74 & n1978;
  assign n3468 = x76 & n2108;
  assign n3469 = ~n3467 & ~n3468;
  assign n3470 = x75 & n1973;
  assign n3471 = n3469 & ~n3470;
  assign n3472 = ~n3466 & n3471;
  assign n3473 = n3472 ^ x26;
  assign n3517 = n3516 ^ n3473;
  assign n3463 = n3351 ^ n3286;
  assign n3464 = n3352 & n3463;
  assign n3465 = n3464 ^ n3286;
  assign n3518 = n3517 ^ n3465;
  assign n3455 = n1054 & n1624;
  assign n3456 = x77 & n1742;
  assign n3457 = x78 & n1628;
  assign n3458 = ~n3456 & ~n3457;
  assign n3459 = x79 & n1744;
  assign n3460 = n3458 & ~n3459;
  assign n3461 = ~n3455 & n3460;
  assign n3462 = n3461 ^ x23;
  assign n3519 = n3518 ^ n3462;
  assign n3452 = n3353 ^ n3275;
  assign n3453 = ~n3354 & ~n3452;
  assign n3454 = n3453 ^ n3275;
  assign n3520 = n3519 ^ n3454;
  assign n3444 = n1296 & n1345;
  assign n3445 = x80 & n1403;
  assign n3446 = x81 & n1300;
  assign n3447 = ~n3445 & ~n3446;
  assign n3448 = x82 & n1406;
  assign n3449 = n3447 & ~n3448;
  assign n3450 = ~n3444 & n3449;
  assign n3451 = n3450 ^ x20;
  assign n3521 = n3520 ^ n3451;
  assign n3441 = n3355 ^ n3264;
  assign n3442 = n3356 & n3441;
  assign n3443 = n3442 ^ n3264;
  assign n3522 = n3521 ^ n3443;
  assign n3433 = n1008 & n1674;
  assign n3434 = x84 & n1012;
  assign n3435 = x83 & n1101;
  assign n3436 = ~n3434 & ~n3435;
  assign n3437 = x85 & n1104;
  assign n3438 = n3436 & ~n3437;
  assign n3439 = ~n3433 & n3438;
  assign n3440 = n3439 ^ x17;
  assign n3523 = n3522 ^ n3440;
  assign n3430 = n3357 ^ n3253;
  assign n3431 = ~n3358 & ~n3430;
  assign n3432 = n3431 ^ n3253;
  assign n3524 = n3523 ^ n3432;
  assign n3422 = n752 & n2040;
  assign n3423 = x86 & n825;
  assign n3424 = x87 & n757;
  assign n3425 = ~n3423 & ~n3424;
  assign n3426 = x88 & n828;
  assign n3427 = n3425 & ~n3426;
  assign n3428 = ~n3422 & n3427;
  assign n3429 = n3428 ^ x14;
  assign n3525 = n3524 ^ n3429;
  assign n3419 = n3359 ^ n3242;
  assign n3420 = n3360 & n3419;
  assign n3421 = n3420 ^ n3242;
  assign n3526 = n3525 ^ n3421;
  assign n3411 = n541 & n2447;
  assign n3412 = x89 & n612;
  assign n3413 = x90 & n547;
  assign n3414 = ~n3412 & ~n3413;
  assign n3415 = x91 & n615;
  assign n3416 = n3414 & ~n3415;
  assign n3417 = ~n3411 & n3416;
  assign n3418 = n3417 ^ x11;
  assign n3527 = n3526 ^ n3418;
  assign n3408 = n3361 ^ n3231;
  assign n3409 = ~n3362 & ~n3408;
  assign n3410 = n3409 ^ n3231;
  assign n3528 = n3527 ^ n3410;
  assign n3400 = n372 & n2895;
  assign n3401 = x92 & n433;
  assign n3402 = x93 & n376;
  assign n3403 = ~n3401 & ~n3402;
  assign n3404 = x94 & n428;
  assign n3405 = n3403 & ~n3404;
  assign n3406 = ~n3400 & n3405;
  assign n3407 = n3406 ^ x8;
  assign n3529 = n3528 ^ n3407;
  assign n3397 = n3363 ^ n3220;
  assign n3398 = n3364 & n3397;
  assign n3399 = n3398 ^ n3220;
  assign n3530 = n3529 ^ n3399;
  assign n3388 = n2885 ^ x97;
  assign n3389 = n210 & n3388;
  assign n3390 = x95 & n219;
  assign n3391 = x97 & n259;
  assign n3392 = ~n3390 & ~n3391;
  assign n3393 = x96 & n214;
  assign n3394 = n3392 & ~n3393;
  assign n3395 = ~n3389 & n3394;
  assign n3396 = n3395 ^ x5;
  assign n3531 = n3530 ^ n3396;
  assign n3385 = n3365 ^ n3208;
  assign n3386 = ~n3366 & n3385;
  assign n3387 = n3386 ^ n3208;
  assign n3532 = n3531 ^ n3387;
  assign n3373 = x99 ^ x98;
  assign n3374 = ~n3199 & n3373;
  assign n3375 = n163 & ~n3374;
  assign n3376 = n3375 ^ x1;
  assign n3377 = n3376 ^ x100;
  assign n3378 = x0 & ~n3377;
  assign n3379 = ~x98 & n156;
  assign n3380 = ~x0 & ~n3379;
  assign n3381 = x99 ^ x2;
  assign n3382 = x1 & n3381;
  assign n3383 = n3380 & ~n3382;
  assign n3384 = ~n3378 & ~n3383;
  assign n3533 = n3532 ^ n3384;
  assign n3370 = n3367 ^ n3192;
  assign n3371 = n3368 & ~n3370;
  assign n3372 = n3371 ^ n3192;
  assign n3534 = n3533 ^ n3372;
  assign n3679 = ~n3497 & ~n3511;
  assign n3680 = ~n3509 & ~n3679;
  assign n3672 = x65 ^ x36;
  assign n3673 = n3496 & ~n3672;
  assign n3674 = n3673 ^ x35;
  assign n3675 = n3674 ^ x37;
  assign n3676 = x64 & n3675;
  assign n3677 = n149 & n3496;
  assign n3678 = ~n3676 & ~n3677;
  assign n3681 = n3680 ^ n3678;
  assign n3664 = n300 & n3330;
  assign n3665 = x66 & n3500;
  assign n3666 = x68 & n3502;
  assign n3667 = ~n3665 & ~n3666;
  assign n3668 = x67 & n3334;
  assign n3669 = n3667 & ~n3668;
  assign n3670 = ~n3664 & n3669;
  assign n3671 = n3670 ^ x35;
  assign n3682 = n3681 ^ n3671;
  assign n3656 = n467 & n2836;
  assign n3657 = x70 & n2840;
  assign n3658 = x69 & n2996;
  assign n3659 = ~n3657 & ~n3658;
  assign n3660 = x71 & n2998;
  assign n3661 = n3659 & ~n3660;
  assign n3662 = ~n3656 & n3661;
  assign n3663 = n3662 ^ x32;
  assign n3683 = n3682 ^ n3663;
  assign n3653 = n3512 ^ n3487;
  assign n3654 = ~n3513 & ~n3653;
  assign n3655 = n3654 ^ n3487;
  assign n3684 = n3683 ^ n3655;
  assign n3645 = ~n656 & n2371;
  assign n3646 = x72 & n2528;
  assign n3647 = x74 & n2531;
  assign n3648 = ~n3646 & ~n3647;
  assign n3649 = x73 & n2377;
  assign n3650 = n3648 & ~n3649;
  assign n3651 = ~n3645 & n3650;
  assign n3652 = n3651 ^ x29;
  assign n3685 = n3684 ^ n3652;
  assign n3642 = n3484 ^ n3476;
  assign n3643 = ~n3515 & n3642;
  assign n3644 = n3643 ^ n3514;
  assign n3686 = n3685 ^ n3644;
  assign n3634 = n877 & n1969;
  assign n3635 = x75 & n1978;
  assign n3636 = x77 & n2108;
  assign n3637 = ~n3635 & ~n3636;
  assign n3638 = x76 & n1973;
  assign n3639 = n3637 & ~n3638;
  assign n3640 = ~n3634 & n3639;
  assign n3641 = n3640 ^ x26;
  assign n3687 = n3686 ^ n3641;
  assign n3631 = n3516 ^ n3465;
  assign n3632 = ~n3517 & ~n3631;
  assign n3633 = n3632 ^ n3465;
  assign n3688 = n3687 ^ n3633;
  assign n3623 = ~n1141 & n1624;
  assign n3624 = x78 & n1742;
  assign n3625 = x79 & n1628;
  assign n3626 = ~n3624 & ~n3625;
  assign n3627 = x80 & n1744;
  assign n3628 = n3626 & ~n3627;
  assign n3629 = ~n3623 & n3628;
  assign n3630 = n3629 ^ x23;
  assign n3689 = n3688 ^ n3630;
  assign n3620 = n3518 ^ n3454;
  assign n3621 = n3519 & n3620;
  assign n3622 = n3621 ^ n3454;
  assign n3690 = n3689 ^ n3622;
  assign n3612 = n1296 & n1445;
  assign n3613 = x81 & n1403;
  assign n3614 = x82 & n1300;
  assign n3615 = ~n3613 & ~n3614;
  assign n3616 = x83 & n1406;
  assign n3617 = n3615 & ~n3616;
  assign n3618 = ~n3612 & n3617;
  assign n3619 = n3618 ^ x20;
  assign n3691 = n3690 ^ n3619;
  assign n3609 = n3520 ^ n3443;
  assign n3610 = ~n3521 & ~n3609;
  assign n3611 = n3610 ^ n3443;
  assign n3692 = n3691 ^ n3611;
  assign n3601 = n1008 & n1787;
  assign n3602 = x85 & n1012;
  assign n3603 = x84 & n1101;
  assign n3604 = ~n3602 & ~n3603;
  assign n3605 = x86 & n1104;
  assign n3606 = n3604 & ~n3605;
  assign n3607 = ~n3601 & n3606;
  assign n3608 = n3607 ^ x17;
  assign n3693 = n3692 ^ n3608;
  assign n3598 = n3522 ^ n3432;
  assign n3599 = n3523 & n3598;
  assign n3600 = n3599 ^ n3432;
  assign n3694 = n3693 ^ n3600;
  assign n3590 = n752 & n2164;
  assign n3591 = x87 & n825;
  assign n3592 = x89 & n828;
  assign n3593 = ~n3591 & ~n3592;
  assign n3594 = x88 & n757;
  assign n3595 = n3593 & ~n3594;
  assign n3596 = ~n3590 & n3595;
  assign n3597 = n3596 ^ x14;
  assign n3695 = n3694 ^ n3597;
  assign n3587 = n3524 ^ n3421;
  assign n3588 = ~n3525 & ~n3587;
  assign n3589 = n3588 ^ n3421;
  assign n3696 = n3695 ^ n3589;
  assign n3579 = n541 & n2585;
  assign n3580 = x90 & n612;
  assign n3581 = x92 & n615;
  assign n3582 = ~n3580 & ~n3581;
  assign n3583 = x91 & n547;
  assign n3584 = n3582 & ~n3583;
  assign n3585 = ~n3579 & n3584;
  assign n3586 = n3585 ^ x11;
  assign n3697 = n3696 ^ n3586;
  assign n3576 = n3526 ^ n3410;
  assign n3577 = n3527 & n3576;
  assign n3578 = n3577 ^ n3410;
  assign n3698 = n3697 ^ n3578;
  assign n3568 = n372 & n3054;
  assign n3569 = x93 & n433;
  assign n3570 = x94 & n376;
  assign n3571 = ~n3569 & ~n3570;
  assign n3572 = x95 & n428;
  assign n3573 = n3571 & ~n3572;
  assign n3574 = ~n3568 & n3573;
  assign n3575 = n3574 ^ x8;
  assign n3699 = n3698 ^ n3575;
  assign n3565 = n3528 ^ n3399;
  assign n3566 = ~n3529 & ~n3565;
  assign n3567 = n3566 ^ n3399;
  assign n3700 = n3699 ^ n3567;
  assign n3556 = n3198 ^ n3039;
  assign n3557 = n210 & n3556;
  assign n3558 = x96 & n219;
  assign n3559 = x98 & n259;
  assign n3560 = ~n3558 & ~n3559;
  assign n3561 = x97 & n214;
  assign n3562 = n3560 & ~n3561;
  assign n3563 = ~n3557 & n3562;
  assign n3564 = n3563 ^ x5;
  assign n3701 = n3700 ^ n3564;
  assign n3553 = n3530 ^ n3387;
  assign n3554 = n3531 & ~n3553;
  assign n3555 = n3554 ^ n3387;
  assign n3702 = n3701 ^ n3555;
  assign n3538 = x100 ^ x99;
  assign n3539 = x100 ^ x98;
  assign n3540 = ~n3199 & ~n3539;
  assign n3541 = n3538 & n3540;
  assign n3542 = n3541 ^ n3538;
  assign n3543 = n163 & ~n3542;
  assign n3544 = n3543 ^ x1;
  assign n3545 = n3544 ^ x101;
  assign n3546 = x0 & n3545;
  assign n3547 = ~x1 & x99;
  assign n3548 = ~x0 & ~n3547;
  assign n3549 = x1 & x100;
  assign n3550 = n3549 ^ x2;
  assign n3551 = n3548 & n3550;
  assign n3552 = ~n3546 & ~n3551;
  assign n3703 = n3702 ^ n3552;
  assign n3535 = n3532 ^ n3372;
  assign n3536 = ~n3533 & n3535;
  assign n3537 = n3536 ^ n3372;
  assign n3704 = n3703 ^ n3537;
  assign n3880 = n1230 & n1624;
  assign n3881 = x80 & n1628;
  assign n3882 = x79 & n1742;
  assign n3883 = ~n3881 & ~n3882;
  assign n3884 = x81 & n1744;
  assign n3885 = n3883 & ~n3884;
  assign n3886 = ~n3880 & n3885;
  assign n3887 = n3886 ^ x23;
  assign n3877 = n3688 ^ n3622;
  assign n3878 = ~n3689 & ~n3877;
  assign n3879 = n3878 ^ n3622;
  assign n3888 = n3887 ^ n3879;
  assign n3867 = n953 & n1969;
  assign n3868 = x76 & n1978;
  assign n3869 = x77 & n1973;
  assign n3870 = ~n3868 & ~n3869;
  assign n3871 = x78 & n2108;
  assign n3872 = n3870 & ~n3871;
  assign n3873 = ~n3867 & n3872;
  assign n3874 = n3873 ^ x26;
  assign n3864 = n3686 ^ n3633;
  assign n3865 = n3687 & n3864;
  assign n3866 = n3865 ^ n3633;
  assign n3875 = n3874 ^ n3866;
  assign n3854 = n720 & n2371;
  assign n3855 = x74 & n2377;
  assign n3856 = x73 & n2528;
  assign n3857 = ~n3855 & ~n3856;
  assign n3858 = x75 & n2531;
  assign n3859 = n3857 & ~n3858;
  assign n3860 = ~n3854 & n3859;
  assign n3861 = n3860 ^ x29;
  assign n3851 = n3684 ^ n3644;
  assign n3852 = ~n3685 & ~n3851;
  assign n3853 = n3852 ^ n3644;
  assign n3862 = n3861 ^ n3853;
  assign n3816 = ~x35 & ~x36;
  assign n3825 = ~x37 & x38;
  assign n3826 = n3816 & n3825;
  assign n3827 = x64 & n3826;
  assign n3828 = x38 ^ x37;
  assign n3829 = n3496 & n3828;
  assign n3830 = n208 & n3829;
  assign n3820 = x35 & x36;
  assign n3831 = n3820 ^ n3816;
  assign n3832 = x37 & n3831;
  assign n3833 = n3832 ^ n3820;
  assign n3834 = ~n3830 & ~n3833;
  assign n3835 = x65 & ~n3834;
  assign n3836 = n149 & n3828;
  assign n3837 = x66 & n3496;
  assign n3838 = ~n3836 & n3837;
  assign n3839 = ~n3835 & ~n3838;
  assign n3840 = n3839 ^ x38;
  assign n3817 = x37 & x64;
  assign n3841 = n3817 & n3820;
  assign n3842 = n3839 & n3841;
  assign n3843 = n3840 & n3842;
  assign n3844 = n3843 ^ n3840;
  assign n3845 = ~n3827 & ~n3844;
  assign n3818 = n3816 & ~n3817;
  assign n3819 = ~n201 & ~n3818;
  assign n3821 = ~x37 & x64;
  assign n3822 = n3820 & ~n3821;
  assign n3823 = n3819 & ~n3822;
  assign n3824 = x38 & ~n3823;
  assign n3846 = n3845 ^ n3824;
  assign n3808 = n358 & n3330;
  assign n3809 = x68 & n3334;
  assign n3810 = x67 & n3500;
  assign n3811 = ~n3809 & ~n3810;
  assign n3812 = x69 & n3502;
  assign n3813 = n3811 & ~n3812;
  assign n3814 = ~n3808 & n3813;
  assign n3815 = n3814 ^ x35;
  assign n3847 = n3846 ^ n3815;
  assign n3805 = n3678 ^ n3671;
  assign n3806 = ~n3681 & ~n3805;
  assign n3807 = n3806 ^ n3680;
  assign n3848 = n3847 ^ n3807;
  assign n3797 = n520 & n2836;
  assign n3798 = x70 & n2996;
  assign n3799 = x72 & n2998;
  assign n3800 = ~n3798 & ~n3799;
  assign n3801 = x71 & n2840;
  assign n3802 = n3800 & ~n3801;
  assign n3803 = ~n3797 & n3802;
  assign n3804 = n3803 ^ x32;
  assign n3849 = n3848 ^ n3804;
  assign n3794 = n3682 ^ n3655;
  assign n3795 = n3683 & n3794;
  assign n3796 = n3795 ^ n3655;
  assign n3850 = n3849 ^ n3796;
  assign n3863 = n3862 ^ n3850;
  assign n3876 = n3875 ^ n3863;
  assign n3889 = n3888 ^ n3876;
  assign n3786 = n1296 & n1547;
  assign n3787 = x82 & n1403;
  assign n3788 = x83 & n1300;
  assign n3789 = ~n3787 & ~n3788;
  assign n3790 = x84 & n1406;
  assign n3791 = n3789 & ~n3790;
  assign n3792 = ~n3786 & n3791;
  assign n3793 = n3792 ^ x20;
  assign n3890 = n3889 ^ n3793;
  assign n3783 = n3690 ^ n3611;
  assign n3784 = n3691 & n3783;
  assign n3785 = n3784 ^ n3611;
  assign n3891 = n3890 ^ n3785;
  assign n3775 = n1008 & n1903;
  assign n3776 = x86 & n1012;
  assign n3777 = x85 & n1101;
  assign n3778 = ~n3776 & ~n3777;
  assign n3779 = x87 & n1104;
  assign n3780 = n3778 & ~n3779;
  assign n3781 = ~n3775 & n3780;
  assign n3782 = n3781 ^ x17;
  assign n3892 = n3891 ^ n3782;
  assign n3772 = n3692 ^ n3600;
  assign n3773 = ~n3693 & ~n3772;
  assign n3774 = n3773 ^ n3600;
  assign n3893 = n3892 ^ n3774;
  assign n3764 = n752 & n2292;
  assign n3765 = x88 & n825;
  assign n3766 = x90 & n828;
  assign n3767 = ~n3765 & ~n3766;
  assign n3768 = x89 & n757;
  assign n3769 = n3767 & ~n3768;
  assign n3770 = ~n3764 & n3769;
  assign n3771 = n3770 ^ x14;
  assign n3894 = n3893 ^ n3771;
  assign n3761 = n3694 ^ n3589;
  assign n3762 = n3695 & n3761;
  assign n3763 = n3762 ^ n3589;
  assign n3895 = n3894 ^ n3763;
  assign n3753 = n541 & n2726;
  assign n3754 = x91 & n612;
  assign n3755 = x92 & n547;
  assign n3756 = ~n3754 & ~n3755;
  assign n3757 = x93 & n615;
  assign n3758 = n3756 & ~n3757;
  assign n3759 = ~n3753 & n3758;
  assign n3760 = n3759 ^ x11;
  assign n3896 = n3895 ^ n3760;
  assign n3750 = n3696 ^ n3578;
  assign n3751 = ~n3697 & ~n3750;
  assign n3752 = n3751 ^ n3578;
  assign n3897 = n3896 ^ n3752;
  assign n3742 = n372 & n3209;
  assign n3743 = x94 & n433;
  assign n3744 = x95 & n376;
  assign n3745 = ~n3743 & ~n3744;
  assign n3746 = x96 & n428;
  assign n3747 = n3745 & ~n3746;
  assign n3748 = ~n3742 & n3747;
  assign n3749 = n3748 ^ x8;
  assign n3898 = n3897 ^ n3749;
  assign n3739 = n3698 ^ n3567;
  assign n3740 = n3699 & n3739;
  assign n3741 = n3740 ^ n3567;
  assign n3899 = n3898 ^ n3741;
  assign n3730 = n3199 ^ x99;
  assign n3731 = n210 & n3730;
  assign n3732 = x98 & n214;
  assign n3733 = x97 & n219;
  assign n3734 = ~n3732 & ~n3733;
  assign n3735 = x99 & n259;
  assign n3736 = n3734 & ~n3735;
  assign n3737 = ~n3731 & n3736;
  assign n3738 = n3737 ^ x5;
  assign n3900 = n3899 ^ n3738;
  assign n3727 = n3700 ^ n3555;
  assign n3728 = ~n3701 & n3727;
  assign n3729 = n3728 ^ n3555;
  assign n3901 = n3900 ^ n3729;
  assign n3712 = ~x98 & ~n3199;
  assign n3713 = x99 & x101;
  assign n3714 = ~n3712 & n3713;
  assign n3715 = ~x100 & ~n3714;
  assign n3716 = x98 & ~n3199;
  assign n3717 = ~x99 & ~x101;
  assign n3718 = ~n3716 & n3717;
  assign n3719 = ~n3715 & ~n3718;
  assign n3720 = n3719 ^ x101;
  assign n3721 = n163 & ~n3720;
  assign n3722 = n3721 ^ x1;
  assign n3723 = n3722 ^ x102;
  assign n3708 = x100 & n156;
  assign n3709 = x1 & x101;
  assign n3710 = ~n3708 & ~n3709;
  assign n3711 = n3710 ^ x2;
  assign n3724 = n3723 ^ n3711;
  assign n3725 = ~x0 & ~n3724;
  assign n3726 = n3725 ^ n3723;
  assign n3902 = n3901 ^ n3726;
  assign n3705 = n3702 ^ n3537;
  assign n3706 = ~n3703 & ~n3705;
  assign n3707 = n3706 ^ n3537;
  assign n3903 = n3902 ^ n3707;
  assign n4059 = n3824 & n3845;
  assign n4046 = x66 & n3833;
  assign n4047 = x37 ^ x36;
  assign n4048 = n3828 & ~n4047;
  assign n4049 = ~n3496 & n4048;
  assign n4050 = x65 & n4049;
  assign n4051 = ~n4046 & ~n4050;
  assign n4052 = n3496 & ~n3828;
  assign n4053 = x67 & n4052;
  assign n4054 = n4051 & ~n4053;
  assign n4055 = n264 & n3829;
  assign n4056 = n4054 & ~n4055;
  assign n4057 = n4056 ^ x38;
  assign n4044 = x39 ^ x38;
  assign n4045 = x64 & n4044;
  assign n4058 = n4057 ^ n4045;
  assign n4060 = n4059 ^ n4058;
  assign n4036 = n416 & n3330;
  assign n4037 = x68 & n3500;
  assign n4038 = x69 & n3334;
  assign n4039 = ~n4037 & ~n4038;
  assign n4040 = x70 & n3502;
  assign n4041 = n4039 & ~n4040;
  assign n4042 = ~n4036 & n4041;
  assign n4043 = n4042 ^ x35;
  assign n4061 = n4060 ^ n4043;
  assign n4033 = n3846 ^ n3807;
  assign n4034 = n3847 & n4033;
  assign n4035 = n4034 ^ n3807;
  assign n4062 = n4061 ^ n4035;
  assign n4025 = ~n594 & n2836;
  assign n4026 = x72 & n2840;
  assign n4027 = x73 & n2998;
  assign n4028 = ~n4026 & ~n4027;
  assign n4029 = x71 & n2996;
  assign n4030 = n4028 & ~n4029;
  assign n4031 = ~n4025 & n4030;
  assign n4032 = n4031 ^ x32;
  assign n4063 = n4062 ^ n4032;
  assign n4022 = n3848 ^ n3796;
  assign n4023 = ~n3849 & ~n4022;
  assign n4024 = n4023 ^ n3796;
  assign n4064 = n4063 ^ n4024;
  assign n4014 = n799 & n2371;
  assign n4015 = x74 & n2528;
  assign n4016 = x76 & n2531;
  assign n4017 = ~n4015 & ~n4016;
  assign n4018 = x75 & n2377;
  assign n4019 = n4017 & ~n4018;
  assign n4020 = ~n4014 & n4019;
  assign n4021 = n4020 ^ x29;
  assign n4065 = n4064 ^ n4021;
  assign n4011 = n3861 ^ n3850;
  assign n4012 = ~n3862 & n4011;
  assign n4013 = n4012 ^ n3853;
  assign n4066 = n4065 ^ n4013;
  assign n4003 = n1054 & n1969;
  assign n4004 = x77 & n1978;
  assign n4005 = x79 & n2108;
  assign n4006 = ~n4004 & ~n4005;
  assign n4007 = x78 & n1973;
  assign n4008 = n4006 & ~n4007;
  assign n4009 = ~n4003 & n4008;
  assign n4010 = n4009 ^ x26;
  assign n4067 = n4066 ^ n4010;
  assign n4000 = n3874 ^ n3863;
  assign n4001 = ~n3875 & ~n4000;
  assign n4002 = n4001 ^ n3866;
  assign n4068 = n4067 ^ n4002;
  assign n3992 = n1345 & n1624;
  assign n3993 = x80 & n1742;
  assign n3994 = x81 & n1628;
  assign n3995 = ~n3993 & ~n3994;
  assign n3996 = x82 & n1744;
  assign n3997 = n3995 & ~n3996;
  assign n3998 = ~n3992 & n3997;
  assign n3999 = n3998 ^ x23;
  assign n4069 = n4068 ^ n3999;
  assign n3989 = n3887 ^ n3876;
  assign n3990 = ~n3888 & n3989;
  assign n3991 = n3990 ^ n3879;
  assign n4070 = n4069 ^ n3991;
  assign n3981 = n1296 & n1674;
  assign n3982 = x83 & n1403;
  assign n3983 = x84 & n1300;
  assign n3984 = ~n3982 & ~n3983;
  assign n3985 = x85 & n1406;
  assign n3986 = n3984 & ~n3985;
  assign n3987 = ~n3981 & n3986;
  assign n3988 = n3987 ^ x20;
  assign n4071 = n4070 ^ n3988;
  assign n3978 = n3889 ^ n3785;
  assign n3979 = ~n3890 & ~n3978;
  assign n3980 = n3979 ^ n3785;
  assign n4072 = n4071 ^ n3980;
  assign n3970 = n1008 & n2040;
  assign n3971 = x87 & n1012;
  assign n3972 = x86 & n1101;
  assign n3973 = ~n3971 & ~n3972;
  assign n3974 = x88 & n1104;
  assign n3975 = n3973 & ~n3974;
  assign n3976 = ~n3970 & n3975;
  assign n3977 = n3976 ^ x17;
  assign n4073 = n4072 ^ n3977;
  assign n3967 = n3891 ^ n3774;
  assign n3968 = n3892 & n3967;
  assign n3969 = n3968 ^ n3774;
  assign n4074 = n4073 ^ n3969;
  assign n3959 = n752 & n2447;
  assign n3960 = x89 & n825;
  assign n3961 = x91 & n828;
  assign n3962 = ~n3960 & ~n3961;
  assign n3963 = x90 & n757;
  assign n3964 = n3962 & ~n3963;
  assign n3965 = ~n3959 & n3964;
  assign n3966 = n3965 ^ x14;
  assign n4075 = n4074 ^ n3966;
  assign n3956 = n3893 ^ n3763;
  assign n3957 = ~n3894 & ~n3956;
  assign n3958 = n3957 ^ n3763;
  assign n4076 = n4075 ^ n3958;
  assign n3948 = n541 & n2895;
  assign n3949 = x92 & n612;
  assign n3950 = x94 & n615;
  assign n3951 = ~n3949 & ~n3950;
  assign n3952 = x93 & n547;
  assign n3953 = n3951 & ~n3952;
  assign n3954 = ~n3948 & n3953;
  assign n3955 = n3954 ^ x11;
  assign n4077 = n4076 ^ n3955;
  assign n3945 = n3895 ^ n3752;
  assign n3946 = n3896 & n3945;
  assign n3947 = n3946 ^ n3752;
  assign n4078 = n4077 ^ n3947;
  assign n3937 = n372 & n3388;
  assign n3938 = x95 & n433;
  assign n3939 = x97 & n428;
  assign n3940 = ~n3938 & ~n3939;
  assign n3941 = x96 & n376;
  assign n3942 = n3940 & ~n3941;
  assign n3943 = ~n3937 & n3942;
  assign n3944 = n3943 ^ x8;
  assign n4079 = n4078 ^ n3944;
  assign n3934 = n3897 ^ n3741;
  assign n3935 = ~n3898 & ~n3934;
  assign n3936 = n3935 ^ n3741;
  assign n4080 = n4079 ^ n3936;
  assign n3925 = n3374 ^ x100;
  assign n3926 = n210 & n3925;
  assign n3927 = x98 & n219;
  assign n3928 = x99 & n214;
  assign n3929 = ~n3927 & ~n3928;
  assign n3930 = x100 & n259;
  assign n3931 = n3929 & ~n3930;
  assign n3932 = ~n3926 & n3931;
  assign n3933 = n3932 ^ x5;
  assign n4081 = n4080 ^ n3933;
  assign n3922 = n3899 ^ n3729;
  assign n3923 = n3900 & ~n3922;
  assign n3924 = n3923 ^ n3729;
  assign n4082 = n4081 ^ n3924;
  assign n3911 = x101 & n3719;
  assign n3912 = ~x102 & ~n3911;
  assign n3913 = ~x101 & ~n3719;
  assign n3914 = x102 & ~n3913;
  assign n3915 = ~n3912 & ~n3914;
  assign n3916 = n163 & ~n3915;
  assign n3917 = n3916 ^ x1;
  assign n3918 = n3917 ^ x103;
  assign n3907 = ~x101 & n156;
  assign n3908 = x102 ^ x2;
  assign n3909 = x1 & n3908;
  assign n3910 = ~n3907 & ~n3909;
  assign n3919 = n3918 ^ n3910;
  assign n3920 = ~x0 & ~n3919;
  assign n3921 = n3920 ^ n3918;
  assign n4083 = n4082 ^ n3921;
  assign n3904 = n3901 ^ n3707;
  assign n3905 = ~n3902 & n3904;
  assign n3906 = n3905 ^ n3707;
  assign n4084 = n4083 ^ n3906;
  assign n4235 = n467 & n3330;
  assign n4236 = x70 & n3334;
  assign n4237 = x69 & n3500;
  assign n4238 = ~n4236 & ~n4237;
  assign n4239 = x71 & n3502;
  assign n4240 = n4238 & ~n4239;
  assign n4241 = ~n4235 & n4240;
  assign n4242 = n4241 ^ x35;
  assign n4232 = n4060 ^ n4035;
  assign n4233 = ~n4061 & ~n4232;
  assign n4234 = n4233 ^ n4035;
  assign n4243 = n4242 ^ n4234;
  assign n4228 = ~n4045 & ~n4059;
  assign n4229 = ~n4057 & ~n4228;
  assign n4221 = x65 ^ x39;
  assign n4222 = n4044 & ~n4221;
  assign n4223 = n4222 ^ x38;
  assign n4224 = n4223 ^ x40;
  assign n4225 = x64 & n4224;
  assign n4226 = n149 & n4044;
  assign n4227 = ~n4225 & ~n4226;
  assign n4230 = n4229 ^ n4227;
  assign n4213 = n300 & n3829;
  assign n4214 = x67 & n3833;
  assign n4215 = x66 & n4049;
  assign n4216 = ~n4214 & ~n4215;
  assign n4217 = x68 & n4052;
  assign n4218 = n4216 & ~n4217;
  assign n4219 = ~n4213 & n4218;
  assign n4220 = n4219 ^ x38;
  assign n4231 = n4230 ^ n4220;
  assign n4244 = n4243 ^ n4231;
  assign n4205 = ~n656 & n2836;
  assign n4206 = x72 & n2996;
  assign n4207 = x74 & n2998;
  assign n4208 = ~n4206 & ~n4207;
  assign n4209 = x73 & n2840;
  assign n4210 = n4208 & ~n4209;
  assign n4211 = ~n4205 & n4210;
  assign n4212 = n4211 ^ x32;
  assign n4245 = n4244 ^ n4212;
  assign n4202 = n4062 ^ n4024;
  assign n4203 = n4063 & n4202;
  assign n4204 = n4203 ^ n4024;
  assign n4246 = n4245 ^ n4204;
  assign n4194 = n877 & n2371;
  assign n4195 = x76 & n2377;
  assign n4196 = x75 & n2528;
  assign n4197 = ~n4195 & ~n4196;
  assign n4198 = x77 & n2531;
  assign n4199 = n4197 & ~n4198;
  assign n4200 = ~n4194 & n4199;
  assign n4201 = n4200 ^ x29;
  assign n4247 = n4246 ^ n4201;
  assign n4191 = n4064 ^ n4013;
  assign n4192 = ~n4065 & ~n4191;
  assign n4193 = n4192 ^ n4013;
  assign n4248 = n4247 ^ n4193;
  assign n4183 = ~n1141 & n1969;
  assign n4184 = x79 & n1973;
  assign n4185 = x80 & n2108;
  assign n4186 = ~n4184 & ~n4185;
  assign n4187 = x78 & n1978;
  assign n4188 = n4186 & ~n4187;
  assign n4189 = ~n4183 & n4188;
  assign n4190 = n4189 ^ x26;
  assign n4249 = n4248 ^ n4190;
  assign n4180 = n4066 ^ n4002;
  assign n4181 = n4067 & n4180;
  assign n4182 = n4181 ^ n4002;
  assign n4250 = n4249 ^ n4182;
  assign n4172 = n1445 & n1624;
  assign n4173 = x81 & n1742;
  assign n4174 = x82 & n1628;
  assign n4175 = ~n4173 & ~n4174;
  assign n4176 = x83 & n1744;
  assign n4177 = n4175 & ~n4176;
  assign n4178 = ~n4172 & n4177;
  assign n4179 = n4178 ^ x23;
  assign n4251 = n4250 ^ n4179;
  assign n4169 = n4068 ^ n3991;
  assign n4170 = ~n4069 & ~n4169;
  assign n4171 = n4170 ^ n3991;
  assign n4252 = n4251 ^ n4171;
  assign n4161 = n1296 & n1787;
  assign n4162 = x84 & n1403;
  assign n4163 = x86 & n1406;
  assign n4164 = ~n4162 & ~n4163;
  assign n4165 = x85 & n1300;
  assign n4166 = n4164 & ~n4165;
  assign n4167 = ~n4161 & n4166;
  assign n4168 = n4167 ^ x20;
  assign n4253 = n4252 ^ n4168;
  assign n4158 = n4070 ^ n3980;
  assign n4159 = n4071 & n4158;
  assign n4160 = n4159 ^ n3980;
  assign n4254 = n4253 ^ n4160;
  assign n4150 = n1008 & n2164;
  assign n4151 = x88 & n1012;
  assign n4152 = x87 & n1101;
  assign n4153 = ~n4151 & ~n4152;
  assign n4154 = x89 & n1104;
  assign n4155 = n4153 & ~n4154;
  assign n4156 = ~n4150 & n4155;
  assign n4157 = n4156 ^ x17;
  assign n4255 = n4254 ^ n4157;
  assign n4147 = n4072 ^ n3969;
  assign n4148 = ~n4073 & ~n4147;
  assign n4149 = n4148 ^ n3969;
  assign n4256 = n4255 ^ n4149;
  assign n4139 = n752 & n2585;
  assign n4140 = x90 & n825;
  assign n4141 = x91 & n757;
  assign n4142 = ~n4140 & ~n4141;
  assign n4143 = x92 & n828;
  assign n4144 = n4142 & ~n4143;
  assign n4145 = ~n4139 & n4144;
  assign n4146 = n4145 ^ x14;
  assign n4257 = n4256 ^ n4146;
  assign n4136 = n4074 ^ n3958;
  assign n4137 = n4075 & n4136;
  assign n4138 = n4137 ^ n3958;
  assign n4258 = n4257 ^ n4138;
  assign n4128 = n541 & n3054;
  assign n4129 = x93 & n612;
  assign n4130 = x95 & n615;
  assign n4131 = ~n4129 & ~n4130;
  assign n4132 = x94 & n547;
  assign n4133 = n4131 & ~n4132;
  assign n4134 = ~n4128 & n4133;
  assign n4135 = n4134 ^ x11;
  assign n4259 = n4258 ^ n4135;
  assign n4125 = n4076 ^ n3947;
  assign n4126 = ~n4077 & ~n4125;
  assign n4127 = n4126 ^ n3947;
  assign n4260 = n4259 ^ n4127;
  assign n4117 = n372 & n3556;
  assign n4118 = x96 & n433;
  assign n4119 = x98 & n428;
  assign n4120 = ~n4118 & ~n4119;
  assign n4121 = x97 & n376;
  assign n4122 = n4120 & ~n4121;
  assign n4123 = ~n4117 & n4122;
  assign n4124 = n4123 ^ x8;
  assign n4261 = n4260 ^ n4124;
  assign n4114 = n4078 ^ n3936;
  assign n4115 = n4079 & n4114;
  assign n4116 = n4115 ^ n3936;
  assign n4262 = n4261 ^ n4116;
  assign n4105 = n3542 ^ x101;
  assign n4106 = n210 & n4105;
  assign n4107 = x99 & n219;
  assign n4108 = x100 & n214;
  assign n4109 = ~n4107 & ~n4108;
  assign n4110 = x101 & n259;
  assign n4111 = n4109 & ~n4110;
  assign n4112 = ~n4106 & n4111;
  assign n4113 = n4112 ^ x5;
  assign n4263 = n4262 ^ n4113;
  assign n4102 = n4080 ^ n3924;
  assign n4103 = ~n4081 & n4102;
  assign n4104 = n4103 ^ n3924;
  assign n4264 = n4263 ^ n4104;
  assign n4093 = x103 & ~n3912;
  assign n4094 = ~x103 & ~n3914;
  assign n4095 = ~n4093 & ~n4094;
  assign n4096 = n163 & ~n4095;
  assign n4097 = n4096 ^ x1;
  assign n4098 = n4097 ^ x104;
  assign n4089 = x103 ^ x2;
  assign n4088 = x2 & ~x102;
  assign n4090 = n4089 ^ n4088;
  assign n4091 = ~x1 & n4090;
  assign n4092 = n4091 ^ n4089;
  assign n4099 = n4098 ^ n4092;
  assign n4100 = ~x0 & n4099;
  assign n4101 = n4100 ^ n4098;
  assign n4265 = n4264 ^ n4101;
  assign n4085 = n4082 ^ n3906;
  assign n4086 = n4083 & ~n4085;
  assign n4087 = n4086 ^ n3906;
  assign n4266 = n4265 ^ n4087;
  assign n4428 = n358 & n3829;
  assign n4429 = x68 & n3833;
  assign n4430 = x67 & n4049;
  assign n4431 = ~n4429 & ~n4430;
  assign n4432 = x69 & n4052;
  assign n4433 = n4431 & ~n4432;
  assign n4434 = ~n4428 & n4433;
  assign n4435 = n4434 ^ x38;
  assign n4409 = x40 ^ x39;
  assign n4410 = ~n4044 & n4409;
  assign n4414 = x41 ^ x40;
  assign n4415 = n4044 & n4414;
  assign n4416 = n208 & n4415;
  assign n4417 = ~n4410 & ~n4416;
  assign n4418 = x65 & ~n4417;
  assign n4419 = ~n4409 & n4414;
  assign n4420 = ~n4044 & n4419;
  assign n4421 = x64 & n4420;
  assign n4422 = n149 & n4414;
  assign n4423 = x66 & n4044;
  assign n4424 = ~n4422 & n4423;
  assign n4425 = ~n4421 & ~n4424;
  assign n4426 = ~n4418 & n4425;
  assign n4408 = x41 & ~n201;
  assign n4411 = x64 & n4410;
  assign n4412 = n4411 ^ n4044;
  assign n4413 = n4408 & n4412;
  assign n4427 = n4426 ^ n4413;
  assign n4436 = n4435 ^ n4427;
  assign n4405 = n4227 ^ n4220;
  assign n4406 = ~n4230 & ~n4405;
  assign n4407 = n4406 ^ n4229;
  assign n4437 = n4436 ^ n4407;
  assign n4397 = n520 & n3330;
  assign n4398 = x71 & n3334;
  assign n4399 = x72 & n3502;
  assign n4400 = ~n4398 & ~n4399;
  assign n4401 = x70 & n3500;
  assign n4402 = n4400 & ~n4401;
  assign n4403 = ~n4397 & n4402;
  assign n4404 = n4403 ^ x35;
  assign n4438 = n4437 ^ n4404;
  assign n4394 = n4242 ^ n4231;
  assign n4395 = ~n4243 & n4394;
  assign n4396 = n4395 ^ n4234;
  assign n4439 = n4438 ^ n4396;
  assign n4386 = n720 & n2836;
  assign n4387 = x73 & n2996;
  assign n4388 = x74 & n2840;
  assign n4389 = ~n4387 & ~n4388;
  assign n4390 = x75 & n2998;
  assign n4391 = n4389 & ~n4390;
  assign n4392 = ~n4386 & n4391;
  assign n4393 = n4392 ^ x32;
  assign n4440 = n4439 ^ n4393;
  assign n4383 = n4244 ^ n4204;
  assign n4384 = ~n4245 & ~n4383;
  assign n4385 = n4384 ^ n4204;
  assign n4441 = n4440 ^ n4385;
  assign n4375 = n953 & n2371;
  assign n4376 = x76 & n2528;
  assign n4377 = x78 & n2531;
  assign n4378 = ~n4376 & ~n4377;
  assign n4379 = x77 & n2377;
  assign n4380 = n4378 & ~n4379;
  assign n4381 = ~n4375 & n4380;
  assign n4382 = n4381 ^ x29;
  assign n4442 = n4441 ^ n4382;
  assign n4372 = n4246 ^ n4193;
  assign n4373 = n4247 & n4372;
  assign n4374 = n4373 ^ n4193;
  assign n4443 = n4442 ^ n4374;
  assign n4364 = n1230 & n1969;
  assign n4365 = x79 & n1978;
  assign n4366 = x81 & n2108;
  assign n4367 = ~n4365 & ~n4366;
  assign n4368 = x80 & n1973;
  assign n4369 = n4367 & ~n4368;
  assign n4370 = ~n4364 & n4369;
  assign n4371 = n4370 ^ x26;
  assign n4444 = n4443 ^ n4371;
  assign n4361 = n4248 ^ n4182;
  assign n4362 = ~n4249 & ~n4361;
  assign n4363 = n4362 ^ n4182;
  assign n4445 = n4444 ^ n4363;
  assign n4353 = n1547 & n1624;
  assign n4354 = x82 & n1742;
  assign n4355 = x83 & n1628;
  assign n4356 = ~n4354 & ~n4355;
  assign n4357 = x84 & n1744;
  assign n4358 = n4356 & ~n4357;
  assign n4359 = ~n4353 & n4358;
  assign n4360 = n4359 ^ x23;
  assign n4446 = n4445 ^ n4360;
  assign n4350 = n4250 ^ n4171;
  assign n4351 = n4251 & n4350;
  assign n4352 = n4351 ^ n4171;
  assign n4447 = n4446 ^ n4352;
  assign n4342 = n1296 & n1903;
  assign n4343 = x86 & n1300;
  assign n4344 = x85 & n1403;
  assign n4345 = ~n4343 & ~n4344;
  assign n4346 = x87 & n1406;
  assign n4347 = n4345 & ~n4346;
  assign n4348 = ~n4342 & n4347;
  assign n4349 = n4348 ^ x20;
  assign n4448 = n4447 ^ n4349;
  assign n4339 = n4252 ^ n4160;
  assign n4340 = ~n4253 & ~n4339;
  assign n4341 = n4340 ^ n4160;
  assign n4449 = n4448 ^ n4341;
  assign n4331 = n1008 & n2292;
  assign n4332 = x89 & n1012;
  assign n4333 = x88 & n1101;
  assign n4334 = ~n4332 & ~n4333;
  assign n4335 = x90 & n1104;
  assign n4336 = n4334 & ~n4335;
  assign n4337 = ~n4331 & n4336;
  assign n4338 = n4337 ^ x17;
  assign n4450 = n4449 ^ n4338;
  assign n4328 = n4254 ^ n4149;
  assign n4329 = n4255 & n4328;
  assign n4330 = n4329 ^ n4149;
  assign n4451 = n4450 ^ n4330;
  assign n4320 = n752 & n2726;
  assign n4321 = x91 & n825;
  assign n4322 = x93 & n828;
  assign n4323 = ~n4321 & ~n4322;
  assign n4324 = x92 & n757;
  assign n4325 = n4323 & ~n4324;
  assign n4326 = ~n4320 & n4325;
  assign n4327 = n4326 ^ x14;
  assign n4452 = n4451 ^ n4327;
  assign n4317 = n4256 ^ n4138;
  assign n4318 = ~n4257 & ~n4317;
  assign n4319 = n4318 ^ n4138;
  assign n4453 = n4452 ^ n4319;
  assign n4309 = n541 & n3209;
  assign n4310 = x94 & n612;
  assign n4311 = x95 & n547;
  assign n4312 = ~n4310 & ~n4311;
  assign n4313 = x96 & n615;
  assign n4314 = n4312 & ~n4313;
  assign n4315 = ~n4309 & n4314;
  assign n4316 = n4315 ^ x11;
  assign n4454 = n4453 ^ n4316;
  assign n4306 = n4258 ^ n4127;
  assign n4307 = n4259 & n4306;
  assign n4308 = n4307 ^ n4127;
  assign n4455 = n4454 ^ n4308;
  assign n4298 = n372 & n3730;
  assign n4299 = x97 & n433;
  assign n4300 = x98 & n376;
  assign n4301 = ~n4299 & ~n4300;
  assign n4302 = x99 & n428;
  assign n4303 = n4301 & ~n4302;
  assign n4304 = ~n4298 & n4303;
  assign n4305 = n4304 ^ x8;
  assign n4456 = n4455 ^ n4305;
  assign n4295 = n4260 ^ n4116;
  assign n4296 = ~n4261 & ~n4295;
  assign n4297 = n4296 ^ n4116;
  assign n4457 = n4456 ^ n4297;
  assign n4286 = n3720 ^ x102;
  assign n4287 = n210 & n4286;
  assign n4288 = x100 & n219;
  assign n4289 = x102 & n259;
  assign n4290 = ~n4288 & ~n4289;
  assign n4291 = x101 & n214;
  assign n4292 = n4290 & ~n4291;
  assign n4293 = ~n4287 & n4292;
  assign n4294 = n4293 ^ x5;
  assign n4458 = n4457 ^ n4294;
  assign n4283 = n4262 ^ n4104;
  assign n4284 = n4263 & ~n4283;
  assign n4285 = n4284 ^ n4104;
  assign n4459 = n4458 ^ n4285;
  assign n4270 = x104 & ~n4094;
  assign n4271 = ~x104 & ~n4093;
  assign n4272 = ~n4270 & ~n4271;
  assign n4273 = n163 & ~n4272;
  assign n4274 = n4273 ^ x1;
  assign n4275 = n4274 ^ x105;
  assign n4276 = x0 & n4275;
  assign n4277 = x103 & n156;
  assign n4278 = ~x0 & ~n4277;
  assign n4279 = x1 & x104;
  assign n4280 = n4279 ^ x2;
  assign n4281 = n4278 & n4280;
  assign n4282 = ~n4276 & ~n4281;
  assign n4460 = n4459 ^ n4282;
  assign n4267 = n4264 ^ n4087;
  assign n4268 = ~n4265 & n4267;
  assign n4269 = n4268 ^ n4087;
  assign n4461 = n4460 ^ n4269;
  assign n4621 = ~n4413 & n4426;
  assign n4622 = x41 & ~n4621;
  assign n4613 = n264 & n4415;
  assign n4614 = n4044 & ~n4414;
  assign n4615 = x67 & n4614;
  assign n4616 = ~n4613 & ~n4615;
  assign n4617 = x66 & n4410;
  assign n4618 = x65 & n4420;
  assign n4619 = ~n4617 & ~n4618;
  assign n4620 = n4616 & n4619;
  assign n4623 = n4622 ^ n4620;
  assign n4611 = x42 ^ x41;
  assign n4612 = x64 & n4611;
  assign n4624 = n4623 ^ n4612;
  assign n4603 = n416 & n3829;
  assign n4604 = x68 & n4049;
  assign n4605 = x69 & n3833;
  assign n4606 = ~n4604 & ~n4605;
  assign n4607 = x70 & n4052;
  assign n4608 = n4606 & ~n4607;
  assign n4609 = ~n4603 & n4608;
  assign n4610 = n4609 ^ x38;
  assign n4625 = n4624 ^ n4610;
  assign n4600 = n4435 ^ n4407;
  assign n4601 = ~n4436 & ~n4600;
  assign n4602 = n4601 ^ n4407;
  assign n4626 = n4625 ^ n4602;
  assign n4592 = ~n594 & n3330;
  assign n4593 = x72 & n3334;
  assign n4594 = x71 & n3500;
  assign n4595 = ~n4593 & ~n4594;
  assign n4596 = x73 & n3502;
  assign n4597 = n4595 & ~n4596;
  assign n4598 = ~n4592 & n4597;
  assign n4599 = n4598 ^ x35;
  assign n4627 = n4626 ^ n4599;
  assign n4589 = n4437 ^ n4396;
  assign n4590 = n4438 & n4589;
  assign n4591 = n4590 ^ n4396;
  assign n4628 = n4627 ^ n4591;
  assign n4581 = n799 & n2836;
  assign n4582 = x74 & n2996;
  assign n4583 = x75 & n2840;
  assign n4584 = ~n4582 & ~n4583;
  assign n4585 = x76 & n2998;
  assign n4586 = n4584 & ~n4585;
  assign n4587 = ~n4581 & n4586;
  assign n4588 = n4587 ^ x32;
  assign n4629 = n4628 ^ n4588;
  assign n4578 = n4439 ^ n4385;
  assign n4579 = ~n4440 & ~n4578;
  assign n4580 = n4579 ^ n4385;
  assign n4630 = n4629 ^ n4580;
  assign n4570 = n1054 & n2371;
  assign n4571 = x77 & n2528;
  assign n4572 = x79 & n2531;
  assign n4573 = ~n4571 & ~n4572;
  assign n4574 = x78 & n2377;
  assign n4575 = n4573 & ~n4574;
  assign n4576 = ~n4570 & n4575;
  assign n4577 = n4576 ^ x29;
  assign n4631 = n4630 ^ n4577;
  assign n4567 = n4441 ^ n4374;
  assign n4568 = n4442 & n4567;
  assign n4569 = n4568 ^ n4374;
  assign n4632 = n4631 ^ n4569;
  assign n4559 = n1345 & n1969;
  assign n4560 = x81 & n1973;
  assign n4561 = x80 & n1978;
  assign n4562 = ~n4560 & ~n4561;
  assign n4563 = x82 & n2108;
  assign n4564 = n4562 & ~n4563;
  assign n4565 = ~n4559 & n4564;
  assign n4566 = n4565 ^ x26;
  assign n4633 = n4632 ^ n4566;
  assign n4556 = n4443 ^ n4363;
  assign n4557 = ~n4444 & ~n4556;
  assign n4558 = n4557 ^ n4363;
  assign n4634 = n4633 ^ n4558;
  assign n4548 = n1624 & n1674;
  assign n4549 = x83 & n1742;
  assign n4550 = x84 & n1628;
  assign n4551 = ~n4549 & ~n4550;
  assign n4552 = x85 & n1744;
  assign n4553 = n4551 & ~n4552;
  assign n4554 = ~n4548 & n4553;
  assign n4555 = n4554 ^ x23;
  assign n4635 = n4634 ^ n4555;
  assign n4545 = n4445 ^ n4352;
  assign n4546 = n4446 & n4545;
  assign n4547 = n4546 ^ n4352;
  assign n4636 = n4635 ^ n4547;
  assign n4537 = n1296 & n2040;
  assign n4538 = x87 & n1300;
  assign n4539 = x86 & n1403;
  assign n4540 = ~n4538 & ~n4539;
  assign n4541 = x88 & n1406;
  assign n4542 = n4540 & ~n4541;
  assign n4543 = ~n4537 & n4542;
  assign n4544 = n4543 ^ x20;
  assign n4637 = n4636 ^ n4544;
  assign n4534 = n4447 ^ n4341;
  assign n4535 = ~n4448 & ~n4534;
  assign n4536 = n4535 ^ n4341;
  assign n4638 = n4637 ^ n4536;
  assign n4526 = n1008 & n2447;
  assign n4527 = x90 & n1012;
  assign n4528 = x89 & n1101;
  assign n4529 = ~n4527 & ~n4528;
  assign n4530 = x91 & n1104;
  assign n4531 = n4529 & ~n4530;
  assign n4532 = ~n4526 & n4531;
  assign n4533 = n4532 ^ x17;
  assign n4639 = n4638 ^ n4533;
  assign n4523 = n4449 ^ n4330;
  assign n4524 = n4450 & n4523;
  assign n4525 = n4524 ^ n4330;
  assign n4640 = n4639 ^ n4525;
  assign n4515 = n752 & n2895;
  assign n4516 = x92 & n825;
  assign n4517 = x93 & n757;
  assign n4518 = ~n4516 & ~n4517;
  assign n4519 = x94 & n828;
  assign n4520 = n4518 & ~n4519;
  assign n4521 = ~n4515 & n4520;
  assign n4522 = n4521 ^ x14;
  assign n4641 = n4640 ^ n4522;
  assign n4512 = n4451 ^ n4319;
  assign n4513 = ~n4452 & ~n4512;
  assign n4514 = n4513 ^ n4319;
  assign n4642 = n4641 ^ n4514;
  assign n4504 = n541 & n3388;
  assign n4505 = x95 & n612;
  assign n4506 = x96 & n547;
  assign n4507 = ~n4505 & ~n4506;
  assign n4508 = x97 & n615;
  assign n4509 = n4507 & ~n4508;
  assign n4510 = ~n4504 & n4509;
  assign n4511 = n4510 ^ x11;
  assign n4643 = n4642 ^ n4511;
  assign n4501 = n4453 ^ n4308;
  assign n4502 = n4454 & n4501;
  assign n4503 = n4502 ^ n4308;
  assign n4644 = n4643 ^ n4503;
  assign n4493 = n372 & n3925;
  assign n4494 = x98 & n433;
  assign n4495 = x100 & n428;
  assign n4496 = ~n4494 & ~n4495;
  assign n4497 = x99 & n376;
  assign n4498 = n4496 & ~n4497;
  assign n4499 = ~n4493 & n4498;
  assign n4500 = n4499 ^ x8;
  assign n4645 = n4644 ^ n4500;
  assign n4490 = n4455 ^ n4297;
  assign n4491 = ~n4456 & ~n4490;
  assign n4492 = n4491 ^ n4297;
  assign n4646 = n4645 ^ n4492;
  assign n4481 = n3915 ^ x103;
  assign n4482 = n210 & n4481;
  assign n4483 = x101 & n219;
  assign n4484 = x103 & n259;
  assign n4485 = ~n4483 & ~n4484;
  assign n4486 = x102 & n214;
  assign n4487 = n4485 & ~n4486;
  assign n4488 = ~n4482 & n4487;
  assign n4489 = n4488 ^ x5;
  assign n4647 = n4646 ^ n4489;
  assign n4478 = n4457 ^ n4285;
  assign n4479 = n4458 & ~n4478;
  assign n4480 = n4479 ^ n4285;
  assign n4648 = n4647 ^ n4480;
  assign n4469 = x105 & ~n4271;
  assign n4470 = ~x105 & ~n4270;
  assign n4471 = ~n4469 & ~n4470;
  assign n4472 = n163 & ~n4471;
  assign n4473 = n4472 ^ x1;
  assign n4474 = n4473 ^ x106;
  assign n4465 = ~x104 & n156;
  assign n4466 = x105 ^ x2;
  assign n4467 = x1 & n4466;
  assign n4468 = ~n4465 & ~n4467;
  assign n4475 = n4474 ^ n4468;
  assign n4476 = ~x0 & ~n4475;
  assign n4477 = n4476 ^ n4474;
  assign n4649 = n4648 ^ n4477;
  assign n4462 = n4459 ^ n4269;
  assign n4463 = n4460 & n4462;
  assign n4464 = n4463 ^ n4269;
  assign n4650 = n4649 ^ n4464;
  assign n4815 = ~n4612 & ~n4623;
  assign n4816 = n4620 ^ x41;
  assign n4817 = ~n4815 & ~n4816;
  assign n4808 = x65 ^ x42;
  assign n4809 = n4611 & ~n4808;
  assign n4810 = n4809 ^ x41;
  assign n4811 = n4810 ^ x43;
  assign n4812 = x64 & n4811;
  assign n4813 = n149 & n4611;
  assign n4814 = ~n4812 & ~n4813;
  assign n4818 = n4817 ^ n4814;
  assign n4800 = n300 & n4415;
  assign n4801 = x67 & n4410;
  assign n4802 = x66 & n4420;
  assign n4803 = ~n4801 & ~n4802;
  assign n4804 = x68 & n4614;
  assign n4805 = n4803 & ~n4804;
  assign n4806 = ~n4800 & n4805;
  assign n4807 = n4806 ^ x41;
  assign n4819 = n4818 ^ n4807;
  assign n4792 = n467 & n3829;
  assign n4793 = x69 & n4049;
  assign n4794 = x70 & n3833;
  assign n4795 = ~n4793 & ~n4794;
  assign n4796 = x71 & n4052;
  assign n4797 = n4795 & ~n4796;
  assign n4798 = ~n4792 & n4797;
  assign n4799 = n4798 ^ x38;
  assign n4820 = n4819 ^ n4799;
  assign n4789 = n4624 ^ n4602;
  assign n4790 = ~n4625 & ~n4789;
  assign n4791 = n4790 ^ n4602;
  assign n4821 = n4820 ^ n4791;
  assign n4781 = ~n656 & n3330;
  assign n4782 = x73 & n3334;
  assign n4783 = x72 & n3500;
  assign n4784 = ~n4782 & ~n4783;
  assign n4785 = x74 & n3502;
  assign n4786 = n4784 & ~n4785;
  assign n4787 = ~n4781 & n4786;
  assign n4788 = n4787 ^ x35;
  assign n4822 = n4821 ^ n4788;
  assign n4778 = n4626 ^ n4591;
  assign n4779 = n4627 & n4778;
  assign n4780 = n4779 ^ n4591;
  assign n4823 = n4822 ^ n4780;
  assign n4770 = n877 & n2836;
  assign n4771 = x75 & n2996;
  assign n4772 = x76 & n2840;
  assign n4773 = ~n4771 & ~n4772;
  assign n4774 = x77 & n2998;
  assign n4775 = n4773 & ~n4774;
  assign n4776 = ~n4770 & n4775;
  assign n4777 = n4776 ^ x32;
  assign n4824 = n4823 ^ n4777;
  assign n4767 = n4628 ^ n4580;
  assign n4768 = ~n4629 & ~n4767;
  assign n4769 = n4768 ^ n4580;
  assign n4825 = n4824 ^ n4769;
  assign n4759 = ~n1141 & n2371;
  assign n4760 = x78 & n2528;
  assign n4761 = x79 & n2377;
  assign n4762 = ~n4760 & ~n4761;
  assign n4763 = x80 & n2531;
  assign n4764 = n4762 & ~n4763;
  assign n4765 = ~n4759 & n4764;
  assign n4766 = n4765 ^ x29;
  assign n4826 = n4825 ^ n4766;
  assign n4756 = n4630 ^ n4569;
  assign n4757 = n4631 & n4756;
  assign n4758 = n4757 ^ n4569;
  assign n4827 = n4826 ^ n4758;
  assign n4748 = n1445 & n1969;
  assign n4749 = x81 & n1978;
  assign n4750 = x82 & n1973;
  assign n4751 = ~n4749 & ~n4750;
  assign n4752 = x83 & n2108;
  assign n4753 = n4751 & ~n4752;
  assign n4754 = ~n4748 & n4753;
  assign n4755 = n4754 ^ x26;
  assign n4828 = n4827 ^ n4755;
  assign n4745 = n4632 ^ n4558;
  assign n4746 = ~n4633 & ~n4745;
  assign n4747 = n4746 ^ n4558;
  assign n4829 = n4828 ^ n4747;
  assign n4737 = n1624 & n1787;
  assign n4738 = x84 & n1742;
  assign n4739 = x85 & n1628;
  assign n4740 = ~n4738 & ~n4739;
  assign n4741 = x86 & n1744;
  assign n4742 = n4740 & ~n4741;
  assign n4743 = ~n4737 & n4742;
  assign n4744 = n4743 ^ x23;
  assign n4830 = n4829 ^ n4744;
  assign n4734 = n4634 ^ n4547;
  assign n4735 = n4635 & n4734;
  assign n4736 = n4735 ^ n4547;
  assign n4831 = n4830 ^ n4736;
  assign n4726 = n1296 & n2164;
  assign n4727 = x87 & n1403;
  assign n4728 = x88 & n1300;
  assign n4729 = ~n4727 & ~n4728;
  assign n4730 = x89 & n1406;
  assign n4731 = n4729 & ~n4730;
  assign n4732 = ~n4726 & n4731;
  assign n4733 = n4732 ^ x20;
  assign n4832 = n4831 ^ n4733;
  assign n4723 = n4636 ^ n4536;
  assign n4724 = ~n4637 & ~n4723;
  assign n4725 = n4724 ^ n4536;
  assign n4833 = n4832 ^ n4725;
  assign n4715 = n1008 & n2585;
  assign n4716 = x90 & n1101;
  assign n4717 = x91 & n1012;
  assign n4718 = ~n4716 & ~n4717;
  assign n4719 = x92 & n1104;
  assign n4720 = n4718 & ~n4719;
  assign n4721 = ~n4715 & n4720;
  assign n4722 = n4721 ^ x17;
  assign n4834 = n4833 ^ n4722;
  assign n4712 = n4638 ^ n4525;
  assign n4713 = n4639 & n4712;
  assign n4714 = n4713 ^ n4525;
  assign n4835 = n4834 ^ n4714;
  assign n4704 = n752 & n3054;
  assign n4705 = x93 & n825;
  assign n4706 = x94 & n757;
  assign n4707 = ~n4705 & ~n4706;
  assign n4708 = x95 & n828;
  assign n4709 = n4707 & ~n4708;
  assign n4710 = ~n4704 & n4709;
  assign n4711 = n4710 ^ x14;
  assign n4836 = n4835 ^ n4711;
  assign n4701 = n4640 ^ n4514;
  assign n4702 = ~n4641 & ~n4701;
  assign n4703 = n4702 ^ n4514;
  assign n4837 = n4836 ^ n4703;
  assign n4693 = n541 & n3556;
  assign n4694 = x97 & n547;
  assign n4695 = x98 & n615;
  assign n4696 = ~n4694 & ~n4695;
  assign n4697 = x96 & n612;
  assign n4698 = n4696 & ~n4697;
  assign n4699 = ~n4693 & n4698;
  assign n4700 = n4699 ^ x11;
  assign n4838 = n4837 ^ n4700;
  assign n4690 = n4642 ^ n4503;
  assign n4691 = n4643 & n4690;
  assign n4692 = n4691 ^ n4503;
  assign n4839 = n4838 ^ n4692;
  assign n4682 = n372 & n4105;
  assign n4683 = x99 & n433;
  assign n4684 = x100 & n376;
  assign n4685 = ~n4683 & ~n4684;
  assign n4686 = x101 & n428;
  assign n4687 = n4685 & ~n4686;
  assign n4688 = ~n4682 & n4687;
  assign n4689 = n4688 ^ x8;
  assign n4840 = n4839 ^ n4689;
  assign n4679 = n4644 ^ n4492;
  assign n4680 = ~n4645 & ~n4679;
  assign n4681 = n4680 ^ n4492;
  assign n4841 = n4840 ^ n4681;
  assign n4670 = n4095 ^ x104;
  assign n4671 = n210 & n4670;
  assign n4672 = x102 & n219;
  assign n4673 = x103 & n214;
  assign n4674 = ~n4672 & ~n4673;
  assign n4675 = x104 & n259;
  assign n4676 = n4674 & ~n4675;
  assign n4677 = ~n4671 & n4676;
  assign n4678 = n4677 ^ x5;
  assign n4842 = n4841 ^ n4678;
  assign n4667 = n4646 ^ n4480;
  assign n4668 = n4647 & ~n4667;
  assign n4669 = n4668 ^ n4480;
  assign n4843 = n4842 ^ n4669;
  assign n4654 = ~x106 & ~n4469;
  assign n4655 = x106 & ~n4470;
  assign n4656 = ~n4654 & ~n4655;
  assign n4657 = n163 & ~n4656;
  assign n4658 = n4657 ^ x1;
  assign n4659 = n4658 ^ x107;
  assign n4660 = x0 & ~n4659;
  assign n4661 = ~x105 & n156;
  assign n4662 = ~x0 & ~n4661;
  assign n4663 = x106 ^ x2;
  assign n4664 = x1 & n4663;
  assign n4665 = n4662 & ~n4664;
  assign n4666 = ~n4660 & ~n4665;
  assign n4844 = n4843 ^ n4666;
  assign n4651 = n4648 ^ n4464;
  assign n4652 = ~n4649 & n4651;
  assign n4653 = n4652 ^ n4464;
  assign n4845 = n4844 ^ n4653;
  assign n5035 = n720 & n3330;
  assign n5036 = x73 & n3500;
  assign n5037 = x75 & n3502;
  assign n5038 = ~n5036 & ~n5037;
  assign n5039 = x74 & n3334;
  assign n5040 = n5038 & ~n5039;
  assign n5041 = ~n5035 & n5040;
  assign n5042 = n5041 ^ x35;
  assign n5032 = n4821 ^ n4780;
  assign n5033 = ~n4822 & ~n5032;
  assign n5034 = n5033 ^ n4780;
  assign n5043 = n5042 ^ n5034;
  assign n4998 = ~x41 & ~x42;
  assign n5006 = ~x43 & x44;
  assign n5007 = n4998 & n5006;
  assign n5008 = x64 & n5007;
  assign n5009 = x44 ^ x43;
  assign n5010 = n4611 & n5009;
  assign n5011 = n208 & n5010;
  assign n5001 = x41 & x42;
  assign n5012 = n5001 ^ n4998;
  assign n5013 = x43 & n5012;
  assign n5014 = n5013 ^ n5001;
  assign n5015 = ~n5011 & ~n5014;
  assign n5016 = x65 & ~n5015;
  assign n5017 = n149 & n5009;
  assign n5018 = x66 & n4611;
  assign n5019 = ~n5017 & n5018;
  assign n5020 = ~n5016 & ~n5019;
  assign n5021 = n5020 ^ x44;
  assign n4997 = x43 & x64;
  assign n5022 = n4997 & n5001;
  assign n5023 = n5020 & n5022;
  assign n5024 = n5021 & n5023;
  assign n5025 = n5024 ^ n5021;
  assign n5026 = ~n5008 & ~n5025;
  assign n4999 = ~n201 & ~n4998;
  assign n5000 = ~n4997 & ~n4999;
  assign n5002 = ~x43 & x64;
  assign n5003 = n5001 & ~n5002;
  assign n5004 = ~n5000 & ~n5003;
  assign n5005 = x44 & ~n5004;
  assign n5027 = n5026 ^ n5005;
  assign n4989 = n358 & n4415;
  assign n4990 = x67 & n4420;
  assign n4991 = x68 & n4410;
  assign n4992 = ~n4990 & ~n4991;
  assign n4993 = x69 & n4614;
  assign n4994 = n4992 & ~n4993;
  assign n4995 = ~n4989 & n4994;
  assign n4996 = n4995 ^ x41;
  assign n5028 = n5027 ^ n4996;
  assign n4986 = n4814 ^ n4807;
  assign n4987 = ~n4818 & ~n4986;
  assign n4988 = n4987 ^ n4817;
  assign n5029 = n5028 ^ n4988;
  assign n4978 = n520 & n3829;
  assign n4979 = x71 & n3833;
  assign n4980 = x70 & n4049;
  assign n4981 = ~n4979 & ~n4980;
  assign n4982 = x72 & n4052;
  assign n4983 = n4981 & ~n4982;
  assign n4984 = ~n4978 & n4983;
  assign n4985 = n4984 ^ x38;
  assign n5030 = n5029 ^ n4985;
  assign n4975 = n4819 ^ n4791;
  assign n4976 = n4820 & n4975;
  assign n4977 = n4976 ^ n4791;
  assign n5031 = n5030 ^ n4977;
  assign n5044 = n5043 ^ n5031;
  assign n4967 = n953 & n2836;
  assign n4968 = x76 & n2996;
  assign n4969 = x77 & n2840;
  assign n4970 = ~n4968 & ~n4969;
  assign n4971 = x78 & n2998;
  assign n4972 = n4970 & ~n4971;
  assign n4973 = ~n4967 & n4972;
  assign n4974 = n4973 ^ x32;
  assign n5045 = n5044 ^ n4974;
  assign n4964 = n4823 ^ n4769;
  assign n4965 = n4824 & n4964;
  assign n4966 = n4965 ^ n4769;
  assign n5046 = n5045 ^ n4966;
  assign n4956 = n1230 & n2371;
  assign n4957 = x79 & n2528;
  assign n4958 = x80 & n2377;
  assign n4959 = ~n4957 & ~n4958;
  assign n4960 = x81 & n2531;
  assign n4961 = n4959 & ~n4960;
  assign n4962 = ~n4956 & n4961;
  assign n4963 = n4962 ^ x29;
  assign n5047 = n5046 ^ n4963;
  assign n4953 = n4825 ^ n4758;
  assign n4954 = ~n4826 & ~n4953;
  assign n4955 = n4954 ^ n4758;
  assign n5048 = n5047 ^ n4955;
  assign n4945 = n1547 & n1969;
  assign n4946 = x82 & n1978;
  assign n4947 = x84 & n2108;
  assign n4948 = ~n4946 & ~n4947;
  assign n4949 = x83 & n1973;
  assign n4950 = n4948 & ~n4949;
  assign n4951 = ~n4945 & n4950;
  assign n4952 = n4951 ^ x26;
  assign n5049 = n5048 ^ n4952;
  assign n4942 = n4827 ^ n4747;
  assign n4943 = n4828 & n4942;
  assign n4944 = n4943 ^ n4747;
  assign n5050 = n5049 ^ n4944;
  assign n4934 = n1624 & n1903;
  assign n4935 = x85 & n1742;
  assign n4936 = x86 & n1628;
  assign n4937 = ~n4935 & ~n4936;
  assign n4938 = x87 & n1744;
  assign n4939 = n4937 & ~n4938;
  assign n4940 = ~n4934 & n4939;
  assign n4941 = n4940 ^ x23;
  assign n5051 = n5050 ^ n4941;
  assign n4931 = n4829 ^ n4736;
  assign n4932 = ~n4830 & ~n4931;
  assign n4933 = n4932 ^ n4736;
  assign n5052 = n5051 ^ n4933;
  assign n4923 = n1296 & n2292;
  assign n4924 = x89 & n1300;
  assign n4925 = x88 & n1403;
  assign n4926 = ~n4924 & ~n4925;
  assign n4927 = x90 & n1406;
  assign n4928 = n4926 & ~n4927;
  assign n4929 = ~n4923 & n4928;
  assign n4930 = n4929 ^ x20;
  assign n5053 = n5052 ^ n4930;
  assign n4920 = n4831 ^ n4725;
  assign n4921 = n4832 & n4920;
  assign n4922 = n4921 ^ n4725;
  assign n5054 = n5053 ^ n4922;
  assign n4912 = n1008 & n2726;
  assign n4913 = x92 & n1012;
  assign n4914 = x91 & n1101;
  assign n4915 = ~n4913 & ~n4914;
  assign n4916 = x93 & n1104;
  assign n4917 = n4915 & ~n4916;
  assign n4918 = ~n4912 & n4917;
  assign n4919 = n4918 ^ x17;
  assign n5055 = n5054 ^ n4919;
  assign n4909 = n4833 ^ n4714;
  assign n4910 = ~n4834 & ~n4909;
  assign n4911 = n4910 ^ n4714;
  assign n5056 = n5055 ^ n4911;
  assign n4901 = n752 & n3209;
  assign n4902 = x94 & n825;
  assign n4903 = x96 & n828;
  assign n4904 = ~n4902 & ~n4903;
  assign n4905 = x95 & n757;
  assign n4906 = n4904 & ~n4905;
  assign n4907 = ~n4901 & n4906;
  assign n4908 = n4907 ^ x14;
  assign n5057 = n5056 ^ n4908;
  assign n4898 = n4835 ^ n4703;
  assign n4899 = n4836 & n4898;
  assign n4900 = n4899 ^ n4703;
  assign n5058 = n5057 ^ n4900;
  assign n4890 = n541 & n3730;
  assign n4891 = x97 & n612;
  assign n4892 = x99 & n615;
  assign n4893 = ~n4891 & ~n4892;
  assign n4894 = x98 & n547;
  assign n4895 = n4893 & ~n4894;
  assign n4896 = ~n4890 & n4895;
  assign n4897 = n4896 ^ x11;
  assign n5059 = n5058 ^ n4897;
  assign n4887 = n4837 ^ n4692;
  assign n4888 = ~n4838 & ~n4887;
  assign n4889 = n4888 ^ n4692;
  assign n5060 = n5059 ^ n4889;
  assign n4879 = n372 & n4286;
  assign n4880 = x100 & n433;
  assign n4881 = x101 & n376;
  assign n4882 = ~n4880 & ~n4881;
  assign n4883 = x102 & n428;
  assign n4884 = n4882 & ~n4883;
  assign n4885 = ~n4879 & n4884;
  assign n4886 = n4885 ^ x8;
  assign n5061 = n5060 ^ n4886;
  assign n4876 = n4839 ^ n4681;
  assign n4877 = n4840 & n4876;
  assign n4878 = n4877 ^ n4681;
  assign n5062 = n5061 ^ n4878;
  assign n4867 = n4272 ^ x105;
  assign n4868 = n210 & n4867;
  assign n4869 = x103 & n219;
  assign n4870 = x104 & n214;
  assign n4871 = ~n4869 & ~n4870;
  assign n4872 = x105 & n259;
  assign n4873 = n4871 & ~n4872;
  assign n4874 = ~n4868 & n4873;
  assign n4875 = n4874 ^ x5;
  assign n5063 = n5062 ^ n4875;
  assign n4864 = n4841 ^ n4669;
  assign n4865 = ~n4842 & n4864;
  assign n4866 = n4865 ^ n4669;
  assign n5064 = n5063 ^ n4866;
  assign n4853 = x106 & ~x107;
  assign n4854 = ~n4470 & n4853;
  assign n4855 = ~x106 & x107;
  assign n4856 = ~n4469 & n4855;
  assign n4857 = ~n4854 & ~n4856;
  assign n4858 = n163 & n4857;
  assign n4859 = n4858 ^ x1;
  assign n4860 = n4859 ^ x108;
  assign n4849 = ~x106 & n156;
  assign n4850 = x107 ^ x2;
  assign n4851 = x1 & n4850;
  assign n4852 = ~n4849 & ~n4851;
  assign n4861 = n4860 ^ n4852;
  assign n4862 = ~x0 & ~n4861;
  assign n4863 = n4862 ^ n4860;
  assign n5065 = n5064 ^ n4863;
  assign n4846 = n4843 ^ n4653;
  assign n4847 = n4844 & ~n4846;
  assign n4848 = n4847 ^ n4653;
  assign n5066 = n5065 ^ n4848;
  assign n5240 = ~n594 & n3829;
  assign n5241 = x71 & n4049;
  assign n5242 = x73 & n4052;
  assign n5243 = ~n5241 & ~n5242;
  assign n5244 = x72 & n3833;
  assign n5245 = n5243 & ~n5244;
  assign n5246 = ~n5240 & n5245;
  assign n5247 = n5246 ^ x38;
  assign n5237 = n5029 ^ n4977;
  assign n5238 = ~n5030 & ~n5237;
  assign n5239 = n5238 ^ n4977;
  assign n5248 = n5247 ^ n5239;
  assign n5233 = n5005 & n5026;
  assign n5220 = x66 & n5014;
  assign n5221 = x43 ^ x42;
  assign n5222 = n5009 & ~n5221;
  assign n5223 = ~n4611 & n5222;
  assign n5224 = x65 & n5223;
  assign n5225 = ~n5220 & ~n5224;
  assign n5226 = n4611 & ~n5009;
  assign n5227 = x67 & n5226;
  assign n5228 = n5225 & ~n5227;
  assign n5229 = n264 & n5010;
  assign n5230 = n5228 & ~n5229;
  assign n5231 = n5230 ^ x44;
  assign n5218 = x45 ^ x44;
  assign n5219 = x64 & n5218;
  assign n5232 = n5231 ^ n5219;
  assign n5234 = n5233 ^ n5232;
  assign n5210 = n416 & n4415;
  assign n5211 = x69 & n4410;
  assign n5212 = x68 & n4420;
  assign n5213 = ~n5211 & ~n5212;
  assign n5214 = x70 & n4614;
  assign n5215 = n5213 & ~n5214;
  assign n5216 = ~n5210 & n5215;
  assign n5217 = n5216 ^ x41;
  assign n5235 = n5234 ^ n5217;
  assign n5207 = n5027 ^ n4988;
  assign n5208 = n5028 & n5207;
  assign n5209 = n5208 ^ n4988;
  assign n5236 = n5235 ^ n5209;
  assign n5249 = n5248 ^ n5236;
  assign n5199 = n799 & n3330;
  assign n5200 = x74 & n3500;
  assign n5201 = x76 & n3502;
  assign n5202 = ~n5200 & ~n5201;
  assign n5203 = x75 & n3334;
  assign n5204 = n5202 & ~n5203;
  assign n5205 = ~n5199 & n5204;
  assign n5206 = n5205 ^ x35;
  assign n5250 = n5249 ^ n5206;
  assign n5196 = n5042 ^ n5031;
  assign n5197 = ~n5043 & n5196;
  assign n5198 = n5197 ^ n5034;
  assign n5251 = n5250 ^ n5198;
  assign n5188 = n1054 & n2836;
  assign n5189 = x77 & n2996;
  assign n5190 = x78 & n2840;
  assign n5191 = ~n5189 & ~n5190;
  assign n5192 = x79 & n2998;
  assign n5193 = n5191 & ~n5192;
  assign n5194 = ~n5188 & n5193;
  assign n5195 = n5194 ^ x32;
  assign n5252 = n5251 ^ n5195;
  assign n5185 = n5044 ^ n4966;
  assign n5186 = ~n5045 & ~n5185;
  assign n5187 = n5186 ^ n4966;
  assign n5253 = n5252 ^ n5187;
  assign n5177 = n1345 & n2371;
  assign n5178 = x80 & n2528;
  assign n5179 = x81 & n2377;
  assign n5180 = ~n5178 & ~n5179;
  assign n5181 = x82 & n2531;
  assign n5182 = n5180 & ~n5181;
  assign n5183 = ~n5177 & n5182;
  assign n5184 = n5183 ^ x29;
  assign n5254 = n5253 ^ n5184;
  assign n5174 = n5046 ^ n4955;
  assign n5175 = n5047 & n5174;
  assign n5176 = n5175 ^ n4955;
  assign n5255 = n5254 ^ n5176;
  assign n5166 = n1674 & n1969;
  assign n5167 = x83 & n1978;
  assign n5168 = x85 & n2108;
  assign n5169 = ~n5167 & ~n5168;
  assign n5170 = x84 & n1973;
  assign n5171 = n5169 & ~n5170;
  assign n5172 = ~n5166 & n5171;
  assign n5173 = n5172 ^ x26;
  assign n5256 = n5255 ^ n5173;
  assign n5163 = n5048 ^ n4944;
  assign n5164 = ~n5049 & ~n5163;
  assign n5165 = n5164 ^ n4944;
  assign n5257 = n5256 ^ n5165;
  assign n5155 = n1624 & n2040;
  assign n5156 = x86 & n1742;
  assign n5157 = x87 & n1628;
  assign n5158 = ~n5156 & ~n5157;
  assign n5159 = x88 & n1744;
  assign n5160 = n5158 & ~n5159;
  assign n5161 = ~n5155 & n5160;
  assign n5162 = n5161 ^ x23;
  assign n5258 = n5257 ^ n5162;
  assign n5152 = n5050 ^ n4933;
  assign n5153 = n5051 & n5152;
  assign n5154 = n5153 ^ n4933;
  assign n5259 = n5258 ^ n5154;
  assign n5144 = n1296 & n2447;
  assign n5145 = x89 & n1403;
  assign n5146 = x91 & n1406;
  assign n5147 = ~n5145 & ~n5146;
  assign n5148 = x90 & n1300;
  assign n5149 = n5147 & ~n5148;
  assign n5150 = ~n5144 & n5149;
  assign n5151 = n5150 ^ x20;
  assign n5260 = n5259 ^ n5151;
  assign n5141 = n5052 ^ n4922;
  assign n5142 = ~n5053 & ~n5141;
  assign n5143 = n5142 ^ n4922;
  assign n5261 = n5260 ^ n5143;
  assign n5133 = n1008 & n2895;
  assign n5134 = x93 & n1012;
  assign n5135 = x92 & n1101;
  assign n5136 = ~n5134 & ~n5135;
  assign n5137 = x94 & n1104;
  assign n5138 = n5136 & ~n5137;
  assign n5139 = ~n5133 & n5138;
  assign n5140 = n5139 ^ x17;
  assign n5262 = n5261 ^ n5140;
  assign n5130 = n5054 ^ n4911;
  assign n5131 = n5055 & n5130;
  assign n5132 = n5131 ^ n4911;
  assign n5263 = n5262 ^ n5132;
  assign n5122 = n752 & n3388;
  assign n5123 = x95 & n825;
  assign n5124 = x97 & n828;
  assign n5125 = ~n5123 & ~n5124;
  assign n5126 = x96 & n757;
  assign n5127 = n5125 & ~n5126;
  assign n5128 = ~n5122 & n5127;
  assign n5129 = n5128 ^ x14;
  assign n5264 = n5263 ^ n5129;
  assign n5119 = n5056 ^ n4900;
  assign n5120 = ~n5057 & ~n5119;
  assign n5121 = n5120 ^ n4900;
  assign n5265 = n5264 ^ n5121;
  assign n5111 = n541 & n3925;
  assign n5112 = x98 & n612;
  assign n5113 = x100 & n615;
  assign n5114 = ~n5112 & ~n5113;
  assign n5115 = x99 & n547;
  assign n5116 = n5114 & ~n5115;
  assign n5117 = ~n5111 & n5116;
  assign n5118 = n5117 ^ x11;
  assign n5266 = n5265 ^ n5118;
  assign n5108 = n5058 ^ n4889;
  assign n5109 = n5059 & n5108;
  assign n5110 = n5109 ^ n4889;
  assign n5267 = n5266 ^ n5110;
  assign n5100 = n372 & n4481;
  assign n5101 = x101 & n433;
  assign n5102 = x102 & n376;
  assign n5103 = ~n5101 & ~n5102;
  assign n5104 = x103 & n428;
  assign n5105 = n5103 & ~n5104;
  assign n5106 = ~n5100 & n5105;
  assign n5107 = n5106 ^ x8;
  assign n5268 = n5267 ^ n5107;
  assign n5097 = n5060 ^ n4878;
  assign n5098 = ~n5061 & ~n5097;
  assign n5099 = n5098 ^ n4878;
  assign n5269 = n5268 ^ n5099;
  assign n5088 = n4471 ^ x106;
  assign n5089 = n210 & n5088;
  assign n5090 = x104 & n219;
  assign n5091 = x105 & n214;
  assign n5092 = ~n5090 & ~n5091;
  assign n5093 = x106 & n259;
  assign n5094 = n5092 & ~n5093;
  assign n5095 = ~n5089 & n5094;
  assign n5096 = n5095 ^ x5;
  assign n5270 = n5269 ^ n5096;
  assign n5085 = n5062 ^ n4866;
  assign n5086 = n5063 & ~n5085;
  assign n5087 = n5086 ^ n4866;
  assign n5271 = n5270 ^ n5087;
  assign n5070 = ~x107 & x108;
  assign n5071 = ~n4655 & n5070;
  assign n5072 = x107 & ~x108;
  assign n5073 = ~n4654 & n5072;
  assign n5074 = ~n5071 & ~n5073;
  assign n5075 = n163 & n5074;
  assign n5076 = n5075 ^ x1;
  assign n5077 = n5076 ^ x109;
  assign n5078 = x0 & n5077;
  assign n5079 = ~x1 & x107;
  assign n5080 = ~x0 & ~n5079;
  assign n5081 = x1 & x108;
  assign n5082 = n5081 ^ x2;
  assign n5083 = n5080 & n5082;
  assign n5084 = ~n5078 & ~n5083;
  assign n5272 = n5271 ^ n5084;
  assign n5067 = n5064 ^ n4848;
  assign n5068 = ~n5065 & n5067;
  assign n5069 = n5068 ^ n4848;
  assign n5273 = n5272 ^ n5069;
  assign n5453 = n877 & n3330;
  assign n5454 = x75 & n3500;
  assign n5455 = x76 & n3334;
  assign n5456 = ~n5454 & ~n5455;
  assign n5457 = x77 & n3502;
  assign n5458 = n5456 & ~n5457;
  assign n5459 = ~n5453 & n5458;
  assign n5460 = n5459 ^ x35;
  assign n5450 = n5249 ^ n5198;
  assign n5451 = ~n5250 & ~n5450;
  assign n5452 = n5451 ^ n5198;
  assign n5461 = n5460 ^ n5452;
  assign n5438 = n467 & n4415;
  assign n5439 = x70 & n4410;
  assign n5440 = x69 & n4420;
  assign n5441 = ~n5439 & ~n5440;
  assign n5442 = x71 & n4614;
  assign n5443 = n5441 & ~n5442;
  assign n5444 = ~n5438 & n5443;
  assign n5445 = n5444 ^ x41;
  assign n5435 = n5234 ^ n5209;
  assign n5436 = ~n5235 & ~n5435;
  assign n5437 = n5436 ^ n5209;
  assign n5446 = n5445 ^ n5437;
  assign n5432 = ~n5219 & ~n5233;
  assign n5433 = ~n5231 & ~n5432;
  assign n5423 = n300 & n5010;
  assign n5424 = x67 & n5014;
  assign n5425 = x66 & n5223;
  assign n5426 = ~n5424 & ~n5425;
  assign n5427 = x68 & n5226;
  assign n5428 = n5426 & ~n5427;
  assign n5429 = ~n5423 & n5428;
  assign n5430 = n5429 ^ x44;
  assign n5416 = x65 ^ x45;
  assign n5417 = n5218 & ~n5416;
  assign n5418 = n5417 ^ x44;
  assign n5419 = n5418 ^ x46;
  assign n5420 = x64 & n5419;
  assign n5421 = n149 & n5218;
  assign n5422 = ~n5420 & ~n5421;
  assign n5431 = n5430 ^ n5422;
  assign n5434 = n5433 ^ n5431;
  assign n5447 = n5446 ^ n5434;
  assign n5408 = ~n656 & n3829;
  assign n5409 = x73 & n3833;
  assign n5410 = x72 & n4049;
  assign n5411 = ~n5409 & ~n5410;
  assign n5412 = x74 & n4052;
  assign n5413 = n5411 & ~n5412;
  assign n5414 = ~n5408 & n5413;
  assign n5415 = n5414 ^ x38;
  assign n5448 = n5447 ^ n5415;
  assign n5405 = n5247 ^ n5236;
  assign n5406 = ~n5248 & n5405;
  assign n5407 = n5406 ^ n5239;
  assign n5449 = n5448 ^ n5407;
  assign n5462 = n5461 ^ n5449;
  assign n5397 = ~n1141 & n2836;
  assign n5398 = x79 & n2840;
  assign n5399 = x78 & n2996;
  assign n5400 = ~n5398 & ~n5399;
  assign n5401 = x80 & n2998;
  assign n5402 = n5400 & ~n5401;
  assign n5403 = ~n5397 & n5402;
  assign n5404 = n5403 ^ x32;
  assign n5463 = n5462 ^ n5404;
  assign n5394 = n5251 ^ n5187;
  assign n5395 = n5252 & n5394;
  assign n5396 = n5395 ^ n5187;
  assign n5464 = n5463 ^ n5396;
  assign n5386 = n1445 & n2371;
  assign n5387 = x81 & n2528;
  assign n5388 = x82 & n2377;
  assign n5389 = ~n5387 & ~n5388;
  assign n5390 = x83 & n2531;
  assign n5391 = n5389 & ~n5390;
  assign n5392 = ~n5386 & n5391;
  assign n5393 = n5392 ^ x29;
  assign n5465 = n5464 ^ n5393;
  assign n5383 = n5253 ^ n5176;
  assign n5384 = ~n5254 & ~n5383;
  assign n5385 = n5384 ^ n5176;
  assign n5466 = n5465 ^ n5385;
  assign n5375 = n1787 & n1969;
  assign n5376 = x84 & n1978;
  assign n5377 = x85 & n1973;
  assign n5378 = ~n5376 & ~n5377;
  assign n5379 = x86 & n2108;
  assign n5380 = n5378 & ~n5379;
  assign n5381 = ~n5375 & n5380;
  assign n5382 = n5381 ^ x26;
  assign n5467 = n5466 ^ n5382;
  assign n5372 = n5255 ^ n5165;
  assign n5373 = n5256 & n5372;
  assign n5374 = n5373 ^ n5165;
  assign n5468 = n5467 ^ n5374;
  assign n5364 = n1624 & n2164;
  assign n5365 = x88 & n1628;
  assign n5366 = x87 & n1742;
  assign n5367 = ~n5365 & ~n5366;
  assign n5368 = x89 & n1744;
  assign n5369 = n5367 & ~n5368;
  assign n5370 = ~n5364 & n5369;
  assign n5371 = n5370 ^ x23;
  assign n5469 = n5468 ^ n5371;
  assign n5361 = n5257 ^ n5154;
  assign n5362 = ~n5258 & ~n5361;
  assign n5363 = n5362 ^ n5154;
  assign n5470 = n5469 ^ n5363;
  assign n5353 = n1296 & n2585;
  assign n5354 = x91 & n1300;
  assign n5355 = x90 & n1403;
  assign n5356 = ~n5354 & ~n5355;
  assign n5357 = x92 & n1406;
  assign n5358 = n5356 & ~n5357;
  assign n5359 = ~n5353 & n5358;
  assign n5360 = n5359 ^ x20;
  assign n5471 = n5470 ^ n5360;
  assign n5350 = n5259 ^ n5143;
  assign n5351 = n5260 & n5350;
  assign n5352 = n5351 ^ n5143;
  assign n5472 = n5471 ^ n5352;
  assign n5342 = n1008 & n3054;
  assign n5343 = x94 & n1012;
  assign n5344 = x93 & n1101;
  assign n5345 = ~n5343 & ~n5344;
  assign n5346 = x95 & n1104;
  assign n5347 = n5345 & ~n5346;
  assign n5348 = ~n5342 & n5347;
  assign n5349 = n5348 ^ x17;
  assign n5473 = n5472 ^ n5349;
  assign n5339 = n5261 ^ n5132;
  assign n5340 = ~n5262 & ~n5339;
  assign n5341 = n5340 ^ n5132;
  assign n5474 = n5473 ^ n5341;
  assign n5331 = n752 & n3556;
  assign n5332 = x96 & n825;
  assign n5333 = x97 & n757;
  assign n5334 = ~n5332 & ~n5333;
  assign n5335 = x98 & n828;
  assign n5336 = n5334 & ~n5335;
  assign n5337 = ~n5331 & n5336;
  assign n5338 = n5337 ^ x14;
  assign n5475 = n5474 ^ n5338;
  assign n5328 = n5263 ^ n5121;
  assign n5329 = n5264 & n5328;
  assign n5330 = n5329 ^ n5121;
  assign n5476 = n5475 ^ n5330;
  assign n5320 = n541 & n4105;
  assign n5321 = x99 & n612;
  assign n5322 = x101 & n615;
  assign n5323 = ~n5321 & ~n5322;
  assign n5324 = x100 & n547;
  assign n5325 = n5323 & ~n5324;
  assign n5326 = ~n5320 & n5325;
  assign n5327 = n5326 ^ x11;
  assign n5477 = n5476 ^ n5327;
  assign n5317 = n5265 ^ n5110;
  assign n5318 = ~n5266 & ~n5317;
  assign n5319 = n5318 ^ n5110;
  assign n5478 = n5477 ^ n5319;
  assign n5309 = n372 & n4670;
  assign n5310 = x102 & n433;
  assign n5311 = x103 & n376;
  assign n5312 = ~n5310 & ~n5311;
  assign n5313 = x104 & n428;
  assign n5314 = n5312 & ~n5313;
  assign n5315 = ~n5309 & n5314;
  assign n5316 = n5315 ^ x8;
  assign n5479 = n5478 ^ n5316;
  assign n5306 = n5267 ^ n5099;
  assign n5307 = n5268 & n5306;
  assign n5308 = n5307 ^ n5099;
  assign n5480 = n5479 ^ n5308;
  assign n5297 = n4656 ^ x107;
  assign n5298 = n210 & n5297;
  assign n5299 = x105 & n219;
  assign n5300 = x107 & n259;
  assign n5301 = ~n5299 & ~n5300;
  assign n5302 = x106 & n214;
  assign n5303 = n5301 & ~n5302;
  assign n5304 = ~n5298 & n5303;
  assign n5305 = n5304 ^ x5;
  assign n5481 = n5480 ^ n5305;
  assign n5294 = n5269 ^ n5087;
  assign n5295 = ~n5270 & n5294;
  assign n5296 = n5295 ^ n5087;
  assign n5482 = n5481 ^ n5296;
  assign n5277 = x107 & x109;
  assign n5278 = ~n4654 & n5277;
  assign n5279 = ~x108 & ~n5278;
  assign n5280 = ~x107 & ~x109;
  assign n5281 = ~n4655 & n5280;
  assign n5282 = ~n5279 & ~n5281;
  assign n5283 = n5282 ^ x109;
  assign n5284 = n163 & ~n5283;
  assign n5285 = n5284 ^ x1;
  assign n5286 = n5285 ^ x110;
  assign n5287 = x0 & n5286;
  assign n5288 = ~x1 & x108;
  assign n5289 = ~x0 & ~n5288;
  assign n5290 = x1 & x109;
  assign n5291 = n5290 ^ x2;
  assign n5292 = n5289 & n5291;
  assign n5293 = ~n5287 & ~n5292;
  assign n5483 = n5482 ^ n5293;
  assign n5274 = n5271 ^ n5069;
  assign n5275 = ~n5272 & ~n5274;
  assign n5276 = n5275 ^ n5069;
  assign n5484 = n5483 ^ n5276;
  assign n5685 = n5433 ^ n5430;
  assign n5686 = ~n5431 & ~n5685;
  assign n5687 = n5686 ^ n5433;
  assign n5655 = x47 ^ x46;
  assign n5656 = n5218 & n5655;
  assign n5657 = n208 & n5656;
  assign n5659 = x44 & x45;
  assign n5658 = ~x44 & ~x45;
  assign n5660 = n5659 ^ n5658;
  assign n5661 = x46 & n5660;
  assign n5662 = n5661 ^ n5659;
  assign n5663 = ~n5657 & ~n5662;
  assign n5664 = x65 & ~n5663;
  assign n5665 = n149 & n5655;
  assign n5666 = x66 & n5218;
  assign n5667 = ~n5665 & n5666;
  assign n5668 = ~n5664 & ~n5667;
  assign n5677 = ~x46 & x47;
  assign n5678 = n5658 & n5677;
  assign n5679 = x64 & n5678;
  assign n5680 = n5668 & ~n5679;
  assign n5669 = x46 & x64;
  assign n5672 = n5658 & ~n5669;
  assign n5673 = ~n201 & ~n5672;
  assign n5674 = ~x46 & x64;
  assign n5675 = n5659 & ~n5674;
  assign n5676 = n5673 & ~n5675;
  assign n5681 = n5680 ^ n5676;
  assign n5670 = n5659 & n5669;
  assign n5671 = n5668 & ~n5670;
  assign n5682 = n5681 ^ n5671;
  assign n5683 = ~x47 & n5682;
  assign n5684 = n5683 ^ n5681;
  assign n5688 = n5687 ^ n5684;
  assign n5647 = n358 & n5010;
  assign n5648 = x68 & n5014;
  assign n5649 = x67 & n5223;
  assign n5650 = ~n5648 & ~n5649;
  assign n5651 = x69 & n5226;
  assign n5652 = n5650 & ~n5651;
  assign n5653 = ~n5647 & n5652;
  assign n5654 = n5653 ^ x44;
  assign n5689 = n5688 ^ n5654;
  assign n5644 = n5445 ^ n5434;
  assign n5645 = ~n5446 & n5644;
  assign n5646 = n5645 ^ n5437;
  assign n5690 = n5689 ^ n5646;
  assign n5636 = n520 & n4415;
  assign n5637 = x71 & n4410;
  assign n5638 = x70 & n4420;
  assign n5639 = ~n5637 & ~n5638;
  assign n5640 = x72 & n4614;
  assign n5641 = n5639 & ~n5640;
  assign n5642 = ~n5636 & n5641;
  assign n5643 = n5642 ^ x41;
  assign n5691 = n5690 ^ n5643;
  assign n5633 = n5447 ^ n5407;
  assign n5634 = ~n5448 & ~n5633;
  assign n5635 = n5634 ^ n5407;
  assign n5692 = n5691 ^ n5635;
  assign n5625 = n720 & n3829;
  assign n5626 = x74 & n3833;
  assign n5627 = x75 & n4052;
  assign n5628 = ~n5626 & ~n5627;
  assign n5629 = x73 & n4049;
  assign n5630 = n5628 & ~n5629;
  assign n5631 = ~n5625 & n5630;
  assign n5632 = n5631 ^ x38;
  assign n5693 = n5692 ^ n5632;
  assign n5617 = n953 & n3330;
  assign n5618 = x76 & n3500;
  assign n5619 = x78 & n3502;
  assign n5620 = ~n5618 & ~n5619;
  assign n5621 = x77 & n3334;
  assign n5622 = n5620 & ~n5621;
  assign n5623 = ~n5617 & n5622;
  assign n5624 = n5623 ^ x35;
  assign n5694 = n5693 ^ n5624;
  assign n5614 = n5460 ^ n5449;
  assign n5615 = ~n5461 & n5614;
  assign n5616 = n5615 ^ n5452;
  assign n5695 = n5694 ^ n5616;
  assign n5606 = n1230 & n2836;
  assign n5607 = x79 & n2996;
  assign n5608 = x80 & n2840;
  assign n5609 = ~n5607 & ~n5608;
  assign n5610 = x81 & n2998;
  assign n5611 = n5609 & ~n5610;
  assign n5612 = ~n5606 & n5611;
  assign n5613 = n5612 ^ x32;
  assign n5696 = n5695 ^ n5613;
  assign n5603 = n5462 ^ n5396;
  assign n5604 = ~n5463 & ~n5603;
  assign n5605 = n5604 ^ n5396;
  assign n5697 = n5696 ^ n5605;
  assign n5595 = n1547 & n2371;
  assign n5596 = x83 & n2377;
  assign n5597 = x82 & n2528;
  assign n5598 = ~n5596 & ~n5597;
  assign n5599 = x84 & n2531;
  assign n5600 = n5598 & ~n5599;
  assign n5601 = ~n5595 & n5600;
  assign n5602 = n5601 ^ x29;
  assign n5698 = n5697 ^ n5602;
  assign n5592 = n5464 ^ n5385;
  assign n5593 = n5465 & n5592;
  assign n5594 = n5593 ^ n5385;
  assign n5699 = n5698 ^ n5594;
  assign n5584 = n1903 & n1969;
  assign n5585 = x85 & n1978;
  assign n5586 = x86 & n1973;
  assign n5587 = ~n5585 & ~n5586;
  assign n5588 = x87 & n2108;
  assign n5589 = n5587 & ~n5588;
  assign n5590 = ~n5584 & n5589;
  assign n5591 = n5590 ^ x26;
  assign n5700 = n5699 ^ n5591;
  assign n5581 = n5466 ^ n5374;
  assign n5582 = ~n5467 & ~n5581;
  assign n5583 = n5582 ^ n5374;
  assign n5701 = n5700 ^ n5583;
  assign n5573 = n1624 & n2292;
  assign n5574 = x89 & n1628;
  assign n5575 = x88 & n1742;
  assign n5576 = ~n5574 & ~n5575;
  assign n5577 = x90 & n1744;
  assign n5578 = n5576 & ~n5577;
  assign n5579 = ~n5573 & n5578;
  assign n5580 = n5579 ^ x23;
  assign n5702 = n5701 ^ n5580;
  assign n5570 = n5468 ^ n5363;
  assign n5571 = n5469 & n5570;
  assign n5572 = n5571 ^ n5363;
  assign n5703 = n5702 ^ n5572;
  assign n5562 = n1296 & n2726;
  assign n5563 = x92 & n1300;
  assign n5564 = x91 & n1403;
  assign n5565 = ~n5563 & ~n5564;
  assign n5566 = x93 & n1406;
  assign n5567 = n5565 & ~n5566;
  assign n5568 = ~n5562 & n5567;
  assign n5569 = n5568 ^ x20;
  assign n5704 = n5703 ^ n5569;
  assign n5559 = n5470 ^ n5352;
  assign n5560 = ~n5471 & ~n5559;
  assign n5561 = n5560 ^ n5352;
  assign n5705 = n5704 ^ n5561;
  assign n5551 = n1008 & n3209;
  assign n5552 = x94 & n1101;
  assign n5553 = x95 & n1012;
  assign n5554 = ~n5552 & ~n5553;
  assign n5555 = x96 & n1104;
  assign n5556 = n5554 & ~n5555;
  assign n5557 = ~n5551 & n5556;
  assign n5558 = n5557 ^ x17;
  assign n5706 = n5705 ^ n5558;
  assign n5548 = n5472 ^ n5341;
  assign n5549 = n5473 & n5548;
  assign n5550 = n5549 ^ n5341;
  assign n5707 = n5706 ^ n5550;
  assign n5540 = n752 & n3730;
  assign n5541 = x97 & n825;
  assign n5542 = x98 & n757;
  assign n5543 = ~n5541 & ~n5542;
  assign n5544 = x99 & n828;
  assign n5545 = n5543 & ~n5544;
  assign n5546 = ~n5540 & n5545;
  assign n5547 = n5546 ^ x14;
  assign n5708 = n5707 ^ n5547;
  assign n5537 = n5474 ^ n5330;
  assign n5538 = ~n5475 & ~n5537;
  assign n5539 = n5538 ^ n5330;
  assign n5709 = n5708 ^ n5539;
  assign n5529 = n541 & n4286;
  assign n5530 = x100 & n612;
  assign n5531 = x101 & n547;
  assign n5532 = ~n5530 & ~n5531;
  assign n5533 = x102 & n615;
  assign n5534 = n5532 & ~n5533;
  assign n5535 = ~n5529 & n5534;
  assign n5536 = n5535 ^ x11;
  assign n5710 = n5709 ^ n5536;
  assign n5526 = n5476 ^ n5319;
  assign n5527 = n5477 & n5526;
  assign n5528 = n5527 ^ n5319;
  assign n5711 = n5710 ^ n5528;
  assign n5518 = n372 & n4867;
  assign n5519 = x103 & n433;
  assign n5520 = x104 & n376;
  assign n5521 = ~n5519 & ~n5520;
  assign n5522 = x105 & n428;
  assign n5523 = n5521 & ~n5522;
  assign n5524 = ~n5518 & n5523;
  assign n5525 = n5524 ^ x8;
  assign n5712 = n5711 ^ n5525;
  assign n5515 = n5478 ^ n5308;
  assign n5516 = ~n5479 & ~n5515;
  assign n5517 = n5516 ^ n5308;
  assign n5713 = n5712 ^ n5517;
  assign n5506 = n4857 ^ x108;
  assign n5507 = n210 & ~n5506;
  assign n5508 = x106 & n219;
  assign n5509 = x108 & n259;
  assign n5510 = ~n5508 & ~n5509;
  assign n5511 = x107 & n214;
  assign n5512 = n5510 & ~n5511;
  assign n5513 = ~n5507 & n5512;
  assign n5514 = n5513 ^ x5;
  assign n5714 = n5713 ^ n5514;
  assign n5503 = n5480 ^ n5296;
  assign n5504 = n5481 & ~n5503;
  assign n5505 = n5504 ^ n5296;
  assign n5715 = n5714 ^ n5505;
  assign n5492 = x109 & n5282;
  assign n5493 = ~x110 & ~n5492;
  assign n5494 = ~x109 & ~n5282;
  assign n5495 = x110 & ~n5494;
  assign n5496 = ~n5493 & ~n5495;
  assign n5497 = n163 & ~n5496;
  assign n5498 = n5497 ^ x1;
  assign n5499 = n5498 ^ x111;
  assign n5488 = x1 & x110;
  assign n5489 = n5488 ^ x2;
  assign n5490 = ~x1 & x109;
  assign n5491 = n5489 & ~n5490;
  assign n5500 = n5499 ^ n5491;
  assign n5501 = ~x0 & n5500;
  assign n5502 = n5501 ^ n5499;
  assign n5716 = n5715 ^ n5502;
  assign n5485 = n5482 ^ n5276;
  assign n5486 = n5483 & n5485;
  assign n5487 = n5486 ^ n5276;
  assign n5717 = n5716 ^ n5487;
  assign n5902 = ~n5676 & n5680;
  assign n5903 = x47 & n5902;
  assign n5900 = x48 ^ x47;
  assign n5901 = x64 & n5900;
  assign n5904 = n5903 ^ n5901;
  assign n5889 = n162 & n5655;
  assign n5890 = n5889 ^ x67;
  assign n5891 = n5218 & n5890;
  assign n5892 = x66 & n5662;
  assign n5893 = x46 ^ x45;
  assign n5894 = n5655 & ~n5893;
  assign n5895 = ~n5218 & n5894;
  assign n5896 = x65 & n5895;
  assign n5897 = ~n5892 & ~n5896;
  assign n5898 = ~n5891 & n5897;
  assign n5899 = n5898 ^ x47;
  assign n5905 = n5904 ^ n5899;
  assign n5881 = n416 & n5010;
  assign n5882 = x69 & n5014;
  assign n5883 = x68 & n5223;
  assign n5884 = ~n5882 & ~n5883;
  assign n5885 = x70 & n5226;
  assign n5886 = n5884 & ~n5885;
  assign n5887 = ~n5881 & n5886;
  assign n5888 = n5887 ^ x44;
  assign n5906 = n5905 ^ n5888;
  assign n5878 = n5684 ^ n5654;
  assign n5879 = ~n5688 & ~n5878;
  assign n5880 = n5879 ^ n5687;
  assign n5907 = n5906 ^ n5880;
  assign n5875 = n5689 ^ n5643;
  assign n5876 = n5690 & n5875;
  assign n5877 = n5876 ^ n5646;
  assign n5908 = n5907 ^ n5877;
  assign n5867 = ~n594 & n4415;
  assign n5868 = x72 & n4410;
  assign n5869 = x71 & n4420;
  assign n5870 = ~n5868 & ~n5869;
  assign n5871 = x73 & n4614;
  assign n5872 = n5870 & ~n5871;
  assign n5873 = ~n5867 & n5872;
  assign n5874 = n5873 ^ x41;
  assign n5909 = n5908 ^ n5874;
  assign n5859 = n799 & n3829;
  assign n5860 = x74 & n4049;
  assign n5861 = x76 & n4052;
  assign n5862 = ~n5860 & ~n5861;
  assign n5863 = x75 & n3833;
  assign n5864 = n5862 & ~n5863;
  assign n5865 = ~n5859 & n5864;
  assign n5866 = n5865 ^ x38;
  assign n5910 = n5909 ^ n5866;
  assign n5856 = n5691 ^ n5632;
  assign n5857 = ~n5692 & ~n5856;
  assign n5858 = n5857 ^ n5635;
  assign n5911 = n5910 ^ n5858;
  assign n5853 = n5693 ^ n5616;
  assign n5854 = n5694 & n5853;
  assign n5855 = n5854 ^ n5616;
  assign n5912 = n5911 ^ n5855;
  assign n5845 = n1054 & n3330;
  assign n5846 = x77 & n3500;
  assign n5847 = x78 & n3334;
  assign n5848 = ~n5846 & ~n5847;
  assign n5849 = x79 & n3502;
  assign n5850 = n5848 & ~n5849;
  assign n5851 = ~n5845 & n5850;
  assign n5852 = n5851 ^ x35;
  assign n5913 = n5912 ^ n5852;
  assign n5837 = n1345 & n2836;
  assign n5838 = x80 & n2996;
  assign n5839 = x81 & n2840;
  assign n5840 = ~n5838 & ~n5839;
  assign n5841 = x82 & n2998;
  assign n5842 = n5840 & ~n5841;
  assign n5843 = ~n5837 & n5842;
  assign n5844 = n5843 ^ x32;
  assign n5914 = n5913 ^ n5844;
  assign n5834 = n5695 ^ n5605;
  assign n5835 = ~n5696 & ~n5834;
  assign n5836 = n5835 ^ n5605;
  assign n5915 = n5914 ^ n5836;
  assign n5826 = n1674 & n2371;
  assign n5827 = x84 & n2377;
  assign n5828 = x83 & n2528;
  assign n5829 = ~n5827 & ~n5828;
  assign n5830 = x85 & n2531;
  assign n5831 = n5829 & ~n5830;
  assign n5832 = ~n5826 & n5831;
  assign n5833 = n5832 ^ x29;
  assign n5916 = n5915 ^ n5833;
  assign n5823 = n5697 ^ n5594;
  assign n5824 = n5698 & n5823;
  assign n5825 = n5824 ^ n5594;
  assign n5917 = n5916 ^ n5825;
  assign n5815 = n1969 & n2040;
  assign n5816 = x87 & n1973;
  assign n5817 = x86 & n1978;
  assign n5818 = ~n5816 & ~n5817;
  assign n5819 = x88 & n2108;
  assign n5820 = n5818 & ~n5819;
  assign n5821 = ~n5815 & n5820;
  assign n5822 = n5821 ^ x26;
  assign n5918 = n5917 ^ n5822;
  assign n5812 = n5699 ^ n5583;
  assign n5813 = ~n5700 & ~n5812;
  assign n5814 = n5813 ^ n5583;
  assign n5919 = n5918 ^ n5814;
  assign n5804 = n1624 & n2447;
  assign n5805 = x89 & n1742;
  assign n5806 = x90 & n1628;
  assign n5807 = ~n5805 & ~n5806;
  assign n5808 = x91 & n1744;
  assign n5809 = n5807 & ~n5808;
  assign n5810 = ~n5804 & n5809;
  assign n5811 = n5810 ^ x23;
  assign n5920 = n5919 ^ n5811;
  assign n5801 = n5701 ^ n5572;
  assign n5802 = n5702 & n5801;
  assign n5803 = n5802 ^ n5572;
  assign n5921 = n5920 ^ n5803;
  assign n5793 = n1296 & n2895;
  assign n5794 = x93 & n1300;
  assign n5795 = x92 & n1403;
  assign n5796 = ~n5794 & ~n5795;
  assign n5797 = x94 & n1406;
  assign n5798 = n5796 & ~n5797;
  assign n5799 = ~n5793 & n5798;
  assign n5800 = n5799 ^ x20;
  assign n5922 = n5921 ^ n5800;
  assign n5790 = n5703 ^ n5561;
  assign n5791 = ~n5704 & ~n5790;
  assign n5792 = n5791 ^ n5561;
  assign n5923 = n5922 ^ n5792;
  assign n5782 = n1008 & n3388;
  assign n5783 = x96 & n1012;
  assign n5784 = x95 & n1101;
  assign n5785 = ~n5783 & ~n5784;
  assign n5786 = x97 & n1104;
  assign n5787 = n5785 & ~n5786;
  assign n5788 = ~n5782 & n5787;
  assign n5789 = n5788 ^ x17;
  assign n5924 = n5923 ^ n5789;
  assign n5779 = n5705 ^ n5550;
  assign n5780 = n5706 & n5779;
  assign n5781 = n5780 ^ n5550;
  assign n5925 = n5924 ^ n5781;
  assign n5771 = n752 & n3925;
  assign n5772 = x98 & n825;
  assign n5773 = x100 & n828;
  assign n5774 = ~n5772 & ~n5773;
  assign n5775 = x99 & n757;
  assign n5776 = n5774 & ~n5775;
  assign n5777 = ~n5771 & n5776;
  assign n5778 = n5777 ^ x14;
  assign n5926 = n5925 ^ n5778;
  assign n5768 = n5707 ^ n5539;
  assign n5769 = ~n5708 & ~n5768;
  assign n5770 = n5769 ^ n5539;
  assign n5927 = n5926 ^ n5770;
  assign n5760 = n541 & n4481;
  assign n5761 = x101 & n612;
  assign n5762 = x103 & n615;
  assign n5763 = ~n5761 & ~n5762;
  assign n5764 = x102 & n547;
  assign n5765 = n5763 & ~n5764;
  assign n5766 = ~n5760 & n5765;
  assign n5767 = n5766 ^ x11;
  assign n5928 = n5927 ^ n5767;
  assign n5757 = n5709 ^ n5528;
  assign n5758 = n5710 & n5757;
  assign n5759 = n5758 ^ n5528;
  assign n5929 = n5928 ^ n5759;
  assign n5749 = n372 & n5088;
  assign n5750 = x104 & n433;
  assign n5751 = x105 & n376;
  assign n5752 = ~n5750 & ~n5751;
  assign n5753 = x106 & n428;
  assign n5754 = n5752 & ~n5753;
  assign n5755 = ~n5749 & n5754;
  assign n5756 = n5755 ^ x8;
  assign n5930 = n5929 ^ n5756;
  assign n5746 = n5711 ^ n5517;
  assign n5747 = ~n5712 & ~n5746;
  assign n5748 = n5747 ^ n5517;
  assign n5931 = n5930 ^ n5748;
  assign n5737 = n5074 ^ x109;
  assign n5738 = n210 & ~n5737;
  assign n5739 = x107 & n219;
  assign n5740 = x108 & n214;
  assign n5741 = ~n5739 & ~n5740;
  assign n5742 = x109 & n259;
  assign n5743 = n5741 & ~n5742;
  assign n5744 = ~n5738 & n5743;
  assign n5745 = n5744 ^ x5;
  assign n5932 = n5931 ^ n5745;
  assign n5734 = n5713 ^ n5505;
  assign n5735 = n5714 & ~n5734;
  assign n5736 = n5735 ^ n5505;
  assign n5933 = n5932 ^ n5736;
  assign n5725 = ~x111 & ~n5495;
  assign n5726 = x111 & ~n5493;
  assign n5727 = ~n5725 & ~n5726;
  assign n5728 = n163 & ~n5727;
  assign n5729 = n5728 ^ x1;
  assign n5730 = n5729 ^ x112;
  assign n5721 = ~x110 & n156;
  assign n5722 = x111 ^ x2;
  assign n5723 = x1 & n5722;
  assign n5724 = ~n5721 & ~n5723;
  assign n5731 = n5730 ^ n5724;
  assign n5732 = ~x0 & ~n5731;
  assign n5733 = n5732 ^ n5730;
  assign n5934 = n5933 ^ n5733;
  assign n5718 = n5715 ^ n5487;
  assign n5719 = ~n5716 & n5718;
  assign n5720 = n5719 ^ n5487;
  assign n5935 = n5934 ^ n5720;
  assign n6123 = ~n5901 & ~n5903;
  assign n6124 = ~n5899 & ~n6123;
  assign n6116 = x65 ^ x48;
  assign n6117 = n5900 & ~n6116;
  assign n6118 = n6117 ^ x47;
  assign n6119 = n6118 ^ x49;
  assign n6120 = x64 & n6119;
  assign n6121 = n149 & n5900;
  assign n6122 = ~n6120 & ~n6121;
  assign n6125 = n6124 ^ n6122;
  assign n6107 = n300 & n5656;
  assign n6108 = x66 & n5895;
  assign n6109 = x67 & n5662;
  assign n6110 = ~n6108 & ~n6109;
  assign n6111 = n5218 & ~n5655;
  assign n6112 = x68 & n6111;
  assign n6113 = n6110 & ~n6112;
  assign n6114 = ~n6107 & n6113;
  assign n6115 = n6114 ^ x47;
  assign n6126 = n6125 ^ n6115;
  assign n6099 = n467 & n5010;
  assign n6100 = x69 & n5223;
  assign n6101 = x70 & n5014;
  assign n6102 = ~n6100 & ~n6101;
  assign n6103 = x71 & n5226;
  assign n6104 = n6102 & ~n6103;
  assign n6105 = ~n6099 & n6104;
  assign n6106 = n6105 ^ x44;
  assign n6127 = n6126 ^ n6106;
  assign n6096 = n5905 ^ n5880;
  assign n6097 = ~n5906 & ~n6096;
  assign n6098 = n6097 ^ n5880;
  assign n6128 = n6127 ^ n6098;
  assign n6088 = ~n656 & n4415;
  assign n6089 = x73 & n4410;
  assign n6090 = x72 & n4420;
  assign n6091 = ~n6089 & ~n6090;
  assign n6092 = x74 & n4614;
  assign n6093 = n6091 & ~n6092;
  assign n6094 = ~n6088 & n6093;
  assign n6095 = n6094 ^ x41;
  assign n6129 = n6128 ^ n6095;
  assign n6085 = n5907 ^ n5874;
  assign n6086 = n5908 & n6085;
  assign n6087 = n6086 ^ n5877;
  assign n6130 = n6129 ^ n6087;
  assign n6077 = n877 & n3829;
  assign n6078 = x75 & n4049;
  assign n6079 = x76 & n3833;
  assign n6080 = ~n6078 & ~n6079;
  assign n6081 = x77 & n4052;
  assign n6082 = n6080 & ~n6081;
  assign n6083 = ~n6077 & n6082;
  assign n6084 = n6083 ^ x38;
  assign n6131 = n6130 ^ n6084;
  assign n6074 = n5909 ^ n5858;
  assign n6075 = ~n5910 & ~n6074;
  assign n6076 = n6075 ^ n5858;
  assign n6132 = n6131 ^ n6076;
  assign n6066 = ~n1141 & n3330;
  assign n6067 = x78 & n3500;
  assign n6068 = x79 & n3334;
  assign n6069 = ~n6067 & ~n6068;
  assign n6070 = x80 & n3502;
  assign n6071 = n6069 & ~n6070;
  assign n6072 = ~n6066 & n6071;
  assign n6073 = n6072 ^ x35;
  assign n6133 = n6132 ^ n6073;
  assign n6063 = n5911 ^ n5852;
  assign n6064 = n5912 & n6063;
  assign n6065 = n6064 ^ n5855;
  assign n6134 = n6133 ^ n6065;
  assign n6055 = n1445 & n2836;
  assign n6056 = x81 & n2996;
  assign n6057 = x82 & n2840;
  assign n6058 = ~n6056 & ~n6057;
  assign n6059 = x83 & n2998;
  assign n6060 = n6058 & ~n6059;
  assign n6061 = ~n6055 & n6060;
  assign n6062 = n6061 ^ x32;
  assign n6135 = n6134 ^ n6062;
  assign n6052 = n5913 ^ n5836;
  assign n6053 = ~n5914 & ~n6052;
  assign n6054 = n6053 ^ n5836;
  assign n6136 = n6135 ^ n6054;
  assign n6044 = n1787 & n2371;
  assign n6045 = x84 & n2528;
  assign n6046 = x85 & n2377;
  assign n6047 = ~n6045 & ~n6046;
  assign n6048 = x86 & n2531;
  assign n6049 = n6047 & ~n6048;
  assign n6050 = ~n6044 & n6049;
  assign n6051 = n6050 ^ x29;
  assign n6137 = n6136 ^ n6051;
  assign n6041 = n5915 ^ n5825;
  assign n6042 = n5916 & n6041;
  assign n6043 = n6042 ^ n5825;
  assign n6138 = n6137 ^ n6043;
  assign n6033 = n1969 & n2164;
  assign n6034 = x87 & n1978;
  assign n6035 = x88 & n1973;
  assign n6036 = ~n6034 & ~n6035;
  assign n6037 = x89 & n2108;
  assign n6038 = n6036 & ~n6037;
  assign n6039 = ~n6033 & n6038;
  assign n6040 = n6039 ^ x26;
  assign n6139 = n6138 ^ n6040;
  assign n6030 = n5917 ^ n5814;
  assign n6031 = ~n5918 & ~n6030;
  assign n6032 = n6031 ^ n5814;
  assign n6140 = n6139 ^ n6032;
  assign n6022 = n1624 & n2585;
  assign n6023 = x91 & n1628;
  assign n6024 = x90 & n1742;
  assign n6025 = ~n6023 & ~n6024;
  assign n6026 = x92 & n1744;
  assign n6027 = n6025 & ~n6026;
  assign n6028 = ~n6022 & n6027;
  assign n6029 = n6028 ^ x23;
  assign n6141 = n6140 ^ n6029;
  assign n6019 = n5919 ^ n5803;
  assign n6020 = n5920 & n6019;
  assign n6021 = n6020 ^ n5803;
  assign n6142 = n6141 ^ n6021;
  assign n6011 = n1296 & n3054;
  assign n6012 = x93 & n1403;
  assign n6013 = x94 & n1300;
  assign n6014 = ~n6012 & ~n6013;
  assign n6015 = x95 & n1406;
  assign n6016 = n6014 & ~n6015;
  assign n6017 = ~n6011 & n6016;
  assign n6018 = n6017 ^ x20;
  assign n6143 = n6142 ^ n6018;
  assign n6008 = n5921 ^ n5792;
  assign n6009 = ~n5922 & ~n6008;
  assign n6010 = n6009 ^ n5792;
  assign n6144 = n6143 ^ n6010;
  assign n6000 = n1008 & n3556;
  assign n6001 = x97 & n1012;
  assign n6002 = x96 & n1101;
  assign n6003 = ~n6001 & ~n6002;
  assign n6004 = x98 & n1104;
  assign n6005 = n6003 & ~n6004;
  assign n6006 = ~n6000 & n6005;
  assign n6007 = n6006 ^ x17;
  assign n6145 = n6144 ^ n6007;
  assign n5997 = n5923 ^ n5781;
  assign n5998 = n5924 & n5997;
  assign n5999 = n5998 ^ n5781;
  assign n6146 = n6145 ^ n5999;
  assign n5989 = n752 & n4105;
  assign n5990 = x99 & n825;
  assign n5991 = x100 & n757;
  assign n5992 = ~n5990 & ~n5991;
  assign n5993 = x101 & n828;
  assign n5994 = n5992 & ~n5993;
  assign n5995 = ~n5989 & n5994;
  assign n5996 = n5995 ^ x14;
  assign n6147 = n6146 ^ n5996;
  assign n5986 = n5925 ^ n5770;
  assign n5987 = ~n5926 & ~n5986;
  assign n5988 = n5987 ^ n5770;
  assign n6148 = n6147 ^ n5988;
  assign n5978 = n541 & n4670;
  assign n5979 = x102 & n612;
  assign n5980 = x103 & n547;
  assign n5981 = ~n5979 & ~n5980;
  assign n5982 = x104 & n615;
  assign n5983 = n5981 & ~n5982;
  assign n5984 = ~n5978 & n5983;
  assign n5985 = n5984 ^ x11;
  assign n6149 = n6148 ^ n5985;
  assign n5975 = n5927 ^ n5759;
  assign n5976 = n5928 & n5975;
  assign n5977 = n5976 ^ n5759;
  assign n6150 = n6149 ^ n5977;
  assign n5967 = n372 & n5297;
  assign n5968 = x105 & n433;
  assign n5969 = x106 & n376;
  assign n5970 = ~n5968 & ~n5969;
  assign n5971 = x107 & n428;
  assign n5972 = n5970 & ~n5971;
  assign n5973 = ~n5967 & n5972;
  assign n5974 = n5973 ^ x8;
  assign n6151 = n6150 ^ n5974;
  assign n5964 = n5929 ^ n5748;
  assign n5965 = ~n5930 & ~n5964;
  assign n5966 = n5965 ^ n5748;
  assign n6152 = n6151 ^ n5966;
  assign n5954 = x110 ^ x109;
  assign n5955 = n5954 ^ n5282;
  assign n5956 = n210 & n5955;
  assign n5957 = x108 & n219;
  assign n5958 = x109 & n214;
  assign n5959 = ~n5957 & ~n5958;
  assign n5960 = x110 & n259;
  assign n5961 = n5959 & ~n5960;
  assign n5962 = ~n5956 & n5961;
  assign n5963 = n5962 ^ x5;
  assign n6153 = n6152 ^ n5963;
  assign n5951 = n5931 ^ n5736;
  assign n5952 = n5932 & ~n5951;
  assign n5953 = n5952 ^ n5736;
  assign n6154 = n6153 ^ n5953;
  assign n5939 = x112 ^ x111;
  assign n5940 = ~n5727 & n5939;
  assign n5941 = n163 & ~n5940;
  assign n5942 = n5941 ^ x1;
  assign n5943 = n5942 ^ x113;
  assign n5944 = x0 & n5943;
  assign n5945 = x111 & n156;
  assign n5946 = ~x0 & ~n5945;
  assign n5947 = x1 & x112;
  assign n5948 = n5947 ^ x2;
  assign n5949 = n5946 & n5948;
  assign n5950 = ~n5944 & ~n5949;
  assign n6155 = n6154 ^ n5950;
  assign n5936 = n5933 ^ n5720;
  assign n5937 = ~n5934 & n5936;
  assign n5938 = n5937 ^ n5720;
  assign n6156 = n6155 ^ n5938;
  assign n6366 = n720 & n4415;
  assign n6367 = x73 & n4420;
  assign n6368 = x75 & n4614;
  assign n6369 = ~n6367 & ~n6368;
  assign n6370 = x74 & n4410;
  assign n6371 = n6369 & ~n6370;
  assign n6372 = ~n6366 & n6371;
  assign n6373 = n6372 ^ x41;
  assign n6363 = n6128 ^ n6087;
  assign n6364 = ~n6129 & ~n6363;
  assign n6365 = n6364 ^ n6087;
  assign n6374 = n6373 ^ n6365;
  assign n6350 = n358 & n5656;
  assign n6351 = x68 & n5662;
  assign n6352 = x67 & n5895;
  assign n6353 = ~n6351 & ~n6352;
  assign n6354 = x69 & n6111;
  assign n6355 = n6353 & ~n6354;
  assign n6356 = ~n6350 & n6355;
  assign n6357 = n6356 ^ x47;
  assign n6339 = x49 & x64;
  assign n6322 = ~x47 & ~x48;
  assign n6345 = ~n201 & ~n6322;
  assign n6346 = ~n6339 & ~n6345;
  assign n6323 = ~x49 & x64;
  assign n6328 = x47 & x48;
  assign n6347 = ~n6323 & n6328;
  assign n6348 = ~n6346 & ~n6347;
  assign n6349 = x50 & ~n6348;
  assign n6358 = n6357 ^ n6349;
  assign n6324 = n6322 & n6323;
  assign n6325 = x50 ^ x49;
  assign n6326 = n5900 & n6325;
  assign n6327 = n208 & n6326;
  assign n6329 = n6328 ^ n6322;
  assign n6330 = x49 & n6329;
  assign n6331 = n6330 ^ n6328;
  assign n6332 = ~n6327 & ~n6331;
  assign n6333 = x65 & ~n6332;
  assign n6334 = n149 & n6325;
  assign n6335 = x66 & n5900;
  assign n6336 = ~n6334 & n6335;
  assign n6337 = ~n6333 & ~n6336;
  assign n6338 = n6337 ^ x50;
  assign n6340 = n6328 & n6339;
  assign n6341 = n6337 & n6340;
  assign n6342 = n6338 & n6341;
  assign n6343 = n6342 ^ n6338;
  assign n6344 = ~n6324 & ~n6343;
  assign n6359 = n6358 ^ n6344;
  assign n6319 = n6122 ^ n6115;
  assign n6320 = ~n6125 & ~n6319;
  assign n6321 = n6320 ^ n6124;
  assign n6360 = n6359 ^ n6321;
  assign n6316 = n6126 ^ n6098;
  assign n6317 = n6127 & n6316;
  assign n6318 = n6317 ^ n6098;
  assign n6361 = n6360 ^ n6318;
  assign n6308 = n520 & n5010;
  assign n6309 = x71 & n5014;
  assign n6310 = x70 & n5223;
  assign n6311 = ~n6309 & ~n6310;
  assign n6312 = x72 & n5226;
  assign n6313 = n6311 & ~n6312;
  assign n6314 = ~n6308 & n6313;
  assign n6315 = n6314 ^ x44;
  assign n6362 = n6361 ^ n6315;
  assign n6375 = n6374 ^ n6362;
  assign n6300 = n953 & n3829;
  assign n6301 = x76 & n4049;
  assign n6302 = x78 & n4052;
  assign n6303 = ~n6301 & ~n6302;
  assign n6304 = x77 & n3833;
  assign n6305 = n6303 & ~n6304;
  assign n6306 = ~n6300 & n6305;
  assign n6307 = n6306 ^ x38;
  assign n6376 = n6375 ^ n6307;
  assign n6297 = n6130 ^ n6076;
  assign n6298 = n6131 & n6297;
  assign n6299 = n6298 ^ n6076;
  assign n6377 = n6376 ^ n6299;
  assign n6289 = n1230 & n3330;
  assign n6290 = x79 & n3500;
  assign n6291 = x81 & n3502;
  assign n6292 = ~n6290 & ~n6291;
  assign n6293 = x80 & n3334;
  assign n6294 = n6292 & ~n6293;
  assign n6295 = ~n6289 & n6294;
  assign n6296 = n6295 ^ x35;
  assign n6378 = n6377 ^ n6296;
  assign n6286 = n6132 ^ n6065;
  assign n6287 = ~n6133 & ~n6286;
  assign n6288 = n6287 ^ n6065;
  assign n6379 = n6378 ^ n6288;
  assign n6278 = n1547 & n2836;
  assign n6279 = x83 & n2840;
  assign n6280 = x82 & n2996;
  assign n6281 = ~n6279 & ~n6280;
  assign n6282 = x84 & n2998;
  assign n6283 = n6281 & ~n6282;
  assign n6284 = ~n6278 & n6283;
  assign n6285 = n6284 ^ x32;
  assign n6380 = n6379 ^ n6285;
  assign n6275 = n6134 ^ n6054;
  assign n6276 = n6135 & n6275;
  assign n6277 = n6276 ^ n6054;
  assign n6381 = n6380 ^ n6277;
  assign n6267 = n1903 & n2371;
  assign n6268 = x85 & n2528;
  assign n6269 = x86 & n2377;
  assign n6270 = ~n6268 & ~n6269;
  assign n6271 = x87 & n2531;
  assign n6272 = n6270 & ~n6271;
  assign n6273 = ~n6267 & n6272;
  assign n6274 = n6273 ^ x29;
  assign n6382 = n6381 ^ n6274;
  assign n6264 = n6136 ^ n6043;
  assign n6265 = ~n6137 & ~n6264;
  assign n6266 = n6265 ^ n6043;
  assign n6383 = n6382 ^ n6266;
  assign n6256 = n1969 & n2292;
  assign n6257 = x89 & n1973;
  assign n6258 = x88 & n1978;
  assign n6259 = ~n6257 & ~n6258;
  assign n6260 = x90 & n2108;
  assign n6261 = n6259 & ~n6260;
  assign n6262 = ~n6256 & n6261;
  assign n6263 = n6262 ^ x26;
  assign n6384 = n6383 ^ n6263;
  assign n6253 = n6138 ^ n6032;
  assign n6254 = n6139 & n6253;
  assign n6255 = n6254 ^ n6032;
  assign n6385 = n6384 ^ n6255;
  assign n6245 = n1624 & n2726;
  assign n6246 = x92 & n1628;
  assign n6247 = x91 & n1742;
  assign n6248 = ~n6246 & ~n6247;
  assign n6249 = x93 & n1744;
  assign n6250 = n6248 & ~n6249;
  assign n6251 = ~n6245 & n6250;
  assign n6252 = n6251 ^ x23;
  assign n6386 = n6385 ^ n6252;
  assign n6242 = n6140 ^ n6021;
  assign n6243 = ~n6141 & ~n6242;
  assign n6244 = n6243 ^ n6021;
  assign n6387 = n6386 ^ n6244;
  assign n6234 = n1296 & n3209;
  assign n6235 = x94 & n1403;
  assign n6236 = x95 & n1300;
  assign n6237 = ~n6235 & ~n6236;
  assign n6238 = x96 & n1406;
  assign n6239 = n6237 & ~n6238;
  assign n6240 = ~n6234 & n6239;
  assign n6241 = n6240 ^ x20;
  assign n6388 = n6387 ^ n6241;
  assign n6231 = n6142 ^ n6010;
  assign n6232 = n6143 & n6231;
  assign n6233 = n6232 ^ n6010;
  assign n6389 = n6388 ^ n6233;
  assign n6223 = n1008 & n3730;
  assign n6224 = x98 & n1012;
  assign n6225 = x97 & n1101;
  assign n6226 = ~n6224 & ~n6225;
  assign n6227 = x99 & n1104;
  assign n6228 = n6226 & ~n6227;
  assign n6229 = ~n6223 & n6228;
  assign n6230 = n6229 ^ x17;
  assign n6390 = n6389 ^ n6230;
  assign n6220 = n6144 ^ n5999;
  assign n6221 = ~n6145 & ~n6220;
  assign n6222 = n6221 ^ n5999;
  assign n6391 = n6390 ^ n6222;
  assign n6212 = n752 & n4286;
  assign n6213 = x100 & n825;
  assign n6214 = x101 & n757;
  assign n6215 = ~n6213 & ~n6214;
  assign n6216 = x102 & n828;
  assign n6217 = n6215 & ~n6216;
  assign n6218 = ~n6212 & n6217;
  assign n6219 = n6218 ^ x14;
  assign n6392 = n6391 ^ n6219;
  assign n6209 = n6146 ^ n5988;
  assign n6210 = n6147 & n6209;
  assign n6211 = n6210 ^ n5988;
  assign n6393 = n6392 ^ n6211;
  assign n6201 = n541 & n4867;
  assign n6202 = x104 & n547;
  assign n6203 = x103 & n612;
  assign n6204 = ~n6202 & ~n6203;
  assign n6205 = x105 & n615;
  assign n6206 = n6204 & ~n6205;
  assign n6207 = ~n6201 & n6206;
  assign n6208 = n6207 ^ x11;
  assign n6394 = n6393 ^ n6208;
  assign n6198 = n6148 ^ n5977;
  assign n6199 = ~n6149 & ~n6198;
  assign n6200 = n6199 ^ n5977;
  assign n6395 = n6394 ^ n6200;
  assign n6190 = n372 & ~n5506;
  assign n6191 = x106 & n433;
  assign n6192 = x108 & n428;
  assign n6193 = ~n6191 & ~n6192;
  assign n6194 = x107 & n376;
  assign n6195 = n6193 & ~n6194;
  assign n6196 = ~n6190 & n6195;
  assign n6197 = n6196 ^ x8;
  assign n6396 = n6395 ^ n6197;
  assign n6187 = n6150 ^ n5966;
  assign n6188 = n6151 & n6187;
  assign n6189 = n6188 ^ n5966;
  assign n6397 = n6396 ^ n6189;
  assign n6178 = n5496 ^ x111;
  assign n6179 = n210 & n6178;
  assign n6180 = x109 & n219;
  assign n6181 = x110 & n214;
  assign n6182 = ~n6180 & ~n6181;
  assign n6183 = x111 & n259;
  assign n6184 = n6182 & ~n6183;
  assign n6185 = ~n6179 & n6184;
  assign n6186 = n6185 ^ x5;
  assign n6398 = n6397 ^ n6186;
  assign n6175 = n6152 ^ n5953;
  assign n6176 = ~n6153 & n6175;
  assign n6177 = n6176 ^ n5953;
  assign n6399 = n6398 ^ n6177;
  assign n6164 = ~x112 & ~n5726;
  assign n6165 = x113 & ~n6164;
  assign n6166 = x112 & ~n5725;
  assign n6167 = ~x113 & ~n6166;
  assign n6168 = ~n6165 & ~n6167;
  assign n6169 = n163 & ~n6168;
  assign n6170 = n6169 ^ x1;
  assign n6171 = n6170 ^ x114;
  assign n6160 = x113 ^ x2;
  assign n6161 = x1 & n6160;
  assign n6162 = ~x112 & n156;
  assign n6163 = ~n6161 & ~n6162;
  assign n6172 = n6171 ^ n6163;
  assign n6173 = ~x0 & ~n6172;
  assign n6174 = n6173 ^ n6171;
  assign n6400 = n6399 ^ n6174;
  assign n6157 = n6154 ^ n5938;
  assign n6158 = ~n6155 & ~n6157;
  assign n6159 = n6158 ^ n5938;
  assign n6401 = n6400 ^ n6159;
  assign n6601 = n1054 & n3829;
  assign n6602 = x77 & n4049;
  assign n6603 = x78 & n3833;
  assign n6604 = ~n6602 & ~n6603;
  assign n6605 = x79 & n4052;
  assign n6606 = n6604 & ~n6605;
  assign n6607 = ~n6601 & n6606;
  assign n6608 = n6607 ^ x38;
  assign n6598 = n6375 ^ n6299;
  assign n6599 = ~n6376 & ~n6598;
  assign n6600 = n6599 ^ n6299;
  assign n6609 = n6608 ^ n6600;
  assign n6589 = ~n6344 & ~n6349;
  assign n6590 = n6360 & ~n6589;
  assign n6585 = n6321 & ~n6357;
  assign n6587 = n6344 & n6349;
  assign n6591 = ~n6585 & ~n6587;
  assign n6592 = n6590 & n6591;
  assign n6576 = n416 & n5656;
  assign n6577 = x69 & n5662;
  assign n6578 = x68 & n5895;
  assign n6579 = ~n6577 & ~n6578;
  assign n6580 = x70 & n6111;
  assign n6581 = n6579 & ~n6580;
  assign n6582 = ~n6576 & n6581;
  assign n6583 = n6582 ^ x47;
  assign n6563 = x49 ^ x48;
  assign n6564 = n6325 & ~n6563;
  assign n6565 = ~n5900 & n6564;
  assign n6566 = x65 & n6565;
  assign n6567 = x66 & n6331;
  assign n6568 = ~n6566 & ~n6567;
  assign n6569 = n5900 & ~n6325;
  assign n6570 = x67 & n6569;
  assign n6571 = n6568 & ~n6570;
  assign n6572 = n264 & n6326;
  assign n6573 = n6571 & ~n6572;
  assign n6574 = n6573 ^ x50;
  assign n6561 = x51 ^ x50;
  assign n6562 = x64 & n6561;
  assign n6575 = n6574 ^ n6562;
  assign n6584 = n6583 ^ n6575;
  assign n6586 = n6585 ^ n6584;
  assign n6588 = n6587 ^ n6586;
  assign n6593 = n6592 ^ n6588;
  assign n6553 = ~n594 & n5010;
  assign n6554 = x72 & n5014;
  assign n6555 = x71 & n5223;
  assign n6556 = ~n6554 & ~n6555;
  assign n6557 = x73 & n5226;
  assign n6558 = n6556 & ~n6557;
  assign n6559 = ~n6553 & n6558;
  assign n6560 = n6559 ^ x44;
  assign n6594 = n6593 ^ n6560;
  assign n6550 = n6360 ^ n6315;
  assign n6551 = ~n6361 & ~n6550;
  assign n6552 = n6551 ^ n6318;
  assign n6595 = n6594 ^ n6552;
  assign n6542 = n799 & n4415;
  assign n6543 = x74 & n4420;
  assign n6544 = x75 & n4410;
  assign n6545 = ~n6543 & ~n6544;
  assign n6546 = x76 & n4614;
  assign n6547 = n6545 & ~n6546;
  assign n6548 = ~n6542 & n6547;
  assign n6549 = n6548 ^ x41;
  assign n6596 = n6595 ^ n6549;
  assign n6539 = n6373 ^ n6362;
  assign n6540 = ~n6374 & n6539;
  assign n6541 = n6540 ^ n6365;
  assign n6597 = n6596 ^ n6541;
  assign n6610 = n6609 ^ n6597;
  assign n6531 = n1345 & n3330;
  assign n6532 = x80 & n3500;
  assign n6533 = x82 & n3502;
  assign n6534 = ~n6532 & ~n6533;
  assign n6535 = x81 & n3334;
  assign n6536 = n6534 & ~n6535;
  assign n6537 = ~n6531 & n6536;
  assign n6538 = n6537 ^ x35;
  assign n6611 = n6610 ^ n6538;
  assign n6528 = n6377 ^ n6288;
  assign n6529 = n6378 & n6528;
  assign n6530 = n6529 ^ n6288;
  assign n6612 = n6611 ^ n6530;
  assign n6520 = n1674 & n2836;
  assign n6521 = x83 & n2996;
  assign n6522 = x84 & n2840;
  assign n6523 = ~n6521 & ~n6522;
  assign n6524 = x85 & n2998;
  assign n6525 = n6523 & ~n6524;
  assign n6526 = ~n6520 & n6525;
  assign n6527 = n6526 ^ x32;
  assign n6613 = n6612 ^ n6527;
  assign n6517 = n6285 ^ n6277;
  assign n6518 = n6380 & n6517;
  assign n6519 = n6518 ^ n6379;
  assign n6614 = n6613 ^ n6519;
  assign n6509 = n2040 & n2371;
  assign n6510 = x86 & n2528;
  assign n6511 = x87 & n2377;
  assign n6512 = ~n6510 & ~n6511;
  assign n6513 = x88 & n2531;
  assign n6514 = n6512 & ~n6513;
  assign n6515 = ~n6509 & n6514;
  assign n6516 = n6515 ^ x29;
  assign n6615 = n6614 ^ n6516;
  assign n6506 = n6381 ^ n6266;
  assign n6507 = n6382 & n6506;
  assign n6508 = n6507 ^ n6266;
  assign n6616 = n6615 ^ n6508;
  assign n6498 = n1969 & n2447;
  assign n6499 = x89 & n1978;
  assign n6500 = x91 & n2108;
  assign n6501 = ~n6499 & ~n6500;
  assign n6502 = x90 & n1973;
  assign n6503 = n6501 & ~n6502;
  assign n6504 = ~n6498 & n6503;
  assign n6505 = n6504 ^ x26;
  assign n6617 = n6616 ^ n6505;
  assign n6495 = n6383 ^ n6255;
  assign n6496 = ~n6384 & ~n6495;
  assign n6497 = n6496 ^ n6255;
  assign n6618 = n6617 ^ n6497;
  assign n6487 = n1624 & n2895;
  assign n6488 = x93 & n1628;
  assign n6489 = x92 & n1742;
  assign n6490 = ~n6488 & ~n6489;
  assign n6491 = x94 & n1744;
  assign n6492 = n6490 & ~n6491;
  assign n6493 = ~n6487 & n6492;
  assign n6494 = n6493 ^ x23;
  assign n6619 = n6618 ^ n6494;
  assign n6484 = n6385 ^ n6244;
  assign n6485 = n6386 & n6484;
  assign n6486 = n6485 ^ n6244;
  assign n6620 = n6619 ^ n6486;
  assign n6476 = n1296 & n3388;
  assign n6477 = x96 & n1300;
  assign n6478 = x95 & n1403;
  assign n6479 = ~n6477 & ~n6478;
  assign n6480 = x97 & n1406;
  assign n6481 = n6479 & ~n6480;
  assign n6482 = ~n6476 & n6481;
  assign n6483 = n6482 ^ x20;
  assign n6621 = n6620 ^ n6483;
  assign n6473 = n6387 ^ n6233;
  assign n6474 = ~n6388 & ~n6473;
  assign n6475 = n6474 ^ n6233;
  assign n6622 = n6621 ^ n6475;
  assign n6465 = n1008 & n3925;
  assign n6466 = x98 & n1101;
  assign n6467 = x99 & n1012;
  assign n6468 = ~n6466 & ~n6467;
  assign n6469 = x100 & n1104;
  assign n6470 = n6468 & ~n6469;
  assign n6471 = ~n6465 & n6470;
  assign n6472 = n6471 ^ x17;
  assign n6623 = n6622 ^ n6472;
  assign n6462 = n6389 ^ n6222;
  assign n6463 = n6390 & n6462;
  assign n6464 = n6463 ^ n6222;
  assign n6624 = n6623 ^ n6464;
  assign n6454 = n752 & n4481;
  assign n6455 = x101 & n825;
  assign n6456 = x102 & n757;
  assign n6457 = ~n6455 & ~n6456;
  assign n6458 = x103 & n828;
  assign n6459 = n6457 & ~n6458;
  assign n6460 = ~n6454 & n6459;
  assign n6461 = n6460 ^ x14;
  assign n6625 = n6624 ^ n6461;
  assign n6451 = n6391 ^ n6211;
  assign n6452 = ~n6392 & ~n6451;
  assign n6453 = n6452 ^ n6211;
  assign n6626 = n6625 ^ n6453;
  assign n6443 = n541 & n5088;
  assign n6444 = x104 & n612;
  assign n6445 = x105 & n547;
  assign n6446 = ~n6444 & ~n6445;
  assign n6447 = x106 & n615;
  assign n6448 = n6446 & ~n6447;
  assign n6449 = ~n6443 & n6448;
  assign n6450 = n6449 ^ x11;
  assign n6627 = n6626 ^ n6450;
  assign n6440 = n6393 ^ n6200;
  assign n6441 = n6394 & n6440;
  assign n6442 = n6441 ^ n6200;
  assign n6628 = n6627 ^ n6442;
  assign n6432 = n372 & ~n5737;
  assign n6433 = x107 & n433;
  assign n6434 = x108 & n376;
  assign n6435 = ~n6433 & ~n6434;
  assign n6436 = x109 & n428;
  assign n6437 = n6435 & ~n6436;
  assign n6438 = ~n6432 & n6437;
  assign n6439 = n6438 ^ x8;
  assign n6629 = n6628 ^ n6439;
  assign n6429 = n6395 ^ n6189;
  assign n6430 = ~n6396 & ~n6429;
  assign n6431 = n6430 ^ n6189;
  assign n6630 = n6629 ^ n6431;
  assign n6420 = n5727 ^ x112;
  assign n6421 = n210 & n6420;
  assign n6422 = x110 & n219;
  assign n6423 = x111 & n214;
  assign n6424 = ~n6422 & ~n6423;
  assign n6425 = x112 & n259;
  assign n6426 = n6424 & ~n6425;
  assign n6427 = ~n6421 & n6426;
  assign n6428 = n6427 ^ x5;
  assign n6631 = n6630 ^ n6428;
  assign n6417 = n6397 ^ n6177;
  assign n6418 = n6398 & ~n6417;
  assign n6419 = n6418 ^ n6177;
  assign n6632 = n6631 ^ n6419;
  assign n6409 = x114 ^ x113;
  assign n6410 = ~n6168 & n6409;
  assign n6411 = n163 & ~n6410;
  assign n6412 = n6411 ^ x1;
  assign n6413 = n6412 ^ x115;
  assign n6405 = ~x113 & n156;
  assign n6406 = x114 ^ x2;
  assign n6407 = x1 & n6406;
  assign n6408 = ~n6405 & ~n6407;
  assign n6414 = n6413 ^ n6408;
  assign n6415 = ~x0 & ~n6414;
  assign n6416 = n6415 ^ n6413;
  assign n6633 = n6632 ^ n6416;
  assign n6402 = n6399 ^ n6159;
  assign n6403 = ~n6400 & n6402;
  assign n6404 = n6403 ^ n6159;
  assign n6634 = n6633 ^ n6404;
  assign n6837 = n877 & n4415;
  assign n6838 = x75 & n4420;
  assign n6839 = x76 & n4410;
  assign n6840 = ~n6838 & ~n6839;
  assign n6841 = x77 & n4614;
  assign n6842 = n6840 & ~n6841;
  assign n6843 = ~n6837 & n6842;
  assign n6844 = n6843 ^ x41;
  assign n6834 = n6595 ^ n6541;
  assign n6835 = ~n6596 & ~n6834;
  assign n6836 = n6835 ^ n6541;
  assign n6845 = n6844 ^ n6836;
  assign n6824 = ~n6590 & n6591;
  assign n6825 = n6584 & n6824;
  assign n6812 = ~n6575 & ~n6587;
  assign n6826 = ~n6575 & ~n6585;
  assign n6827 = ~n6583 & ~n6826;
  assign n6828 = ~n6812 & ~n6827;
  assign n6829 = ~n6825 & ~n6828;
  assign n6816 = n467 & n5656;
  assign n6817 = x70 & n5662;
  assign n6818 = x69 & n5895;
  assign n6819 = ~n6817 & ~n6818;
  assign n6820 = x71 & n6111;
  assign n6821 = n6819 & ~n6820;
  assign n6822 = ~n6816 & n6821;
  assign n6823 = n6822 ^ x47;
  assign n6830 = n6829 ^ n6823;
  assign n6813 = ~n6574 & ~n6812;
  assign n6805 = x65 ^ x51;
  assign n6806 = n6561 & ~n6805;
  assign n6807 = n6806 ^ x50;
  assign n6808 = n6807 ^ x52;
  assign n6809 = x64 & n6808;
  assign n6810 = n149 & n6561;
  assign n6811 = ~n6809 & ~n6810;
  assign n6814 = n6813 ^ n6811;
  assign n6797 = n300 & n6326;
  assign n6798 = x67 & n6331;
  assign n6799 = x66 & n6565;
  assign n6800 = ~n6798 & ~n6799;
  assign n6801 = x68 & n6569;
  assign n6802 = n6800 & ~n6801;
  assign n6803 = ~n6797 & n6802;
  assign n6804 = n6803 ^ x50;
  assign n6815 = n6814 ^ n6804;
  assign n6831 = n6830 ^ n6815;
  assign n6789 = ~n656 & n5010;
  assign n6790 = x73 & n5014;
  assign n6791 = x72 & n5223;
  assign n6792 = ~n6790 & ~n6791;
  assign n6793 = x74 & n5226;
  assign n6794 = n6792 & ~n6793;
  assign n6795 = ~n6789 & n6794;
  assign n6796 = n6795 ^ x44;
  assign n6832 = n6831 ^ n6796;
  assign n6786 = n6593 ^ n6552;
  assign n6787 = n6594 & n6786;
  assign n6788 = n6787 ^ n6552;
  assign n6833 = n6832 ^ n6788;
  assign n6846 = n6845 ^ n6833;
  assign n6778 = ~n1141 & n3829;
  assign n6779 = x78 & n4049;
  assign n6780 = x80 & n4052;
  assign n6781 = ~n6779 & ~n6780;
  assign n6782 = x79 & n3833;
  assign n6783 = n6781 & ~n6782;
  assign n6784 = ~n6778 & n6783;
  assign n6785 = n6784 ^ x38;
  assign n6847 = n6846 ^ n6785;
  assign n6775 = n6608 ^ n6597;
  assign n6776 = ~n6609 & n6775;
  assign n6777 = n6776 ^ n6600;
  assign n6848 = n6847 ^ n6777;
  assign n6767 = n1445 & n3330;
  assign n6768 = x81 & n3500;
  assign n6769 = x82 & n3334;
  assign n6770 = ~n6768 & ~n6769;
  assign n6771 = x83 & n3502;
  assign n6772 = n6770 & ~n6771;
  assign n6773 = ~n6767 & n6772;
  assign n6774 = n6773 ^ x35;
  assign n6849 = n6848 ^ n6774;
  assign n6764 = n6610 ^ n6530;
  assign n6765 = ~n6611 & ~n6764;
  assign n6766 = n6765 ^ n6530;
  assign n6850 = n6849 ^ n6766;
  assign n6756 = n1787 & n2836;
  assign n6757 = x85 & n2840;
  assign n6758 = x84 & n2996;
  assign n6759 = ~n6757 & ~n6758;
  assign n6760 = x86 & n2998;
  assign n6761 = n6759 & ~n6760;
  assign n6762 = ~n6756 & n6761;
  assign n6763 = n6762 ^ x32;
  assign n6851 = n6850 ^ n6763;
  assign n6753 = n6527 ^ n6519;
  assign n6754 = ~n6613 & ~n6753;
  assign n6755 = n6754 ^ n6612;
  assign n6852 = n6851 ^ n6755;
  assign n6745 = n2164 & n2371;
  assign n6746 = x88 & n2377;
  assign n6747 = x87 & n2528;
  assign n6748 = ~n6746 & ~n6747;
  assign n6749 = x89 & n2531;
  assign n6750 = n6748 & ~n6749;
  assign n6751 = ~n6745 & n6750;
  assign n6752 = n6751 ^ x29;
  assign n6853 = n6852 ^ n6752;
  assign n6742 = n6614 ^ n6508;
  assign n6743 = n6615 & n6742;
  assign n6744 = n6743 ^ n6508;
  assign n6854 = n6853 ^ n6744;
  assign n6734 = n1969 & n2585;
  assign n6735 = x90 & n1978;
  assign n6736 = x92 & n2108;
  assign n6737 = ~n6735 & ~n6736;
  assign n6738 = x91 & n1973;
  assign n6739 = n6737 & ~n6738;
  assign n6740 = ~n6734 & n6739;
  assign n6741 = n6740 ^ x26;
  assign n6855 = n6854 ^ n6741;
  assign n6731 = n6616 ^ n6497;
  assign n6732 = ~n6617 & ~n6731;
  assign n6733 = n6732 ^ n6497;
  assign n6856 = n6855 ^ n6733;
  assign n6723 = n1624 & n3054;
  assign n6724 = x94 & n1628;
  assign n6725 = x93 & n1742;
  assign n6726 = ~n6724 & ~n6725;
  assign n6727 = x95 & n1744;
  assign n6728 = n6726 & ~n6727;
  assign n6729 = ~n6723 & n6728;
  assign n6730 = n6729 ^ x23;
  assign n6857 = n6856 ^ n6730;
  assign n6720 = n6618 ^ n6486;
  assign n6721 = n6619 & n6720;
  assign n6722 = n6721 ^ n6486;
  assign n6858 = n6857 ^ n6722;
  assign n6712 = n1296 & n3556;
  assign n6713 = x96 & n1403;
  assign n6714 = x98 & n1406;
  assign n6715 = ~n6713 & ~n6714;
  assign n6716 = x97 & n1300;
  assign n6717 = n6715 & ~n6716;
  assign n6718 = ~n6712 & n6717;
  assign n6719 = n6718 ^ x20;
  assign n6859 = n6858 ^ n6719;
  assign n6709 = n6620 ^ n6475;
  assign n6710 = ~n6621 & ~n6709;
  assign n6711 = n6710 ^ n6475;
  assign n6860 = n6859 ^ n6711;
  assign n6701 = n1008 & n4105;
  assign n6702 = x100 & n1012;
  assign n6703 = x99 & n1101;
  assign n6704 = ~n6702 & ~n6703;
  assign n6705 = x101 & n1104;
  assign n6706 = n6704 & ~n6705;
  assign n6707 = ~n6701 & n6706;
  assign n6708 = n6707 ^ x17;
  assign n6861 = n6860 ^ n6708;
  assign n6698 = n6622 ^ n6464;
  assign n6699 = n6623 & n6698;
  assign n6700 = n6699 ^ n6464;
  assign n6862 = n6861 ^ n6700;
  assign n6690 = n752 & n4670;
  assign n6691 = x103 & n757;
  assign n6692 = x102 & n825;
  assign n6693 = ~n6691 & ~n6692;
  assign n6694 = x104 & n828;
  assign n6695 = n6693 & ~n6694;
  assign n6696 = ~n6690 & n6695;
  assign n6697 = n6696 ^ x14;
  assign n6863 = n6862 ^ n6697;
  assign n6687 = n6624 ^ n6453;
  assign n6688 = ~n6625 & ~n6687;
  assign n6689 = n6688 ^ n6453;
  assign n6864 = n6863 ^ n6689;
  assign n6679 = n541 & n5297;
  assign n6680 = x105 & n612;
  assign n6681 = x106 & n547;
  assign n6682 = ~n6680 & ~n6681;
  assign n6683 = x107 & n615;
  assign n6684 = n6682 & ~n6683;
  assign n6685 = ~n6679 & n6684;
  assign n6686 = n6685 ^ x11;
  assign n6865 = n6864 ^ n6686;
  assign n6676 = n6626 ^ n6442;
  assign n6677 = n6627 & n6676;
  assign n6678 = n6677 ^ n6442;
  assign n6866 = n6865 ^ n6678;
  assign n6668 = n372 & n5955;
  assign n6669 = x108 & n433;
  assign n6670 = x109 & n376;
  assign n6671 = ~n6669 & ~n6670;
  assign n6672 = x110 & n428;
  assign n6673 = n6671 & ~n6672;
  assign n6674 = ~n6668 & n6673;
  assign n6675 = n6674 ^ x8;
  assign n6867 = n6866 ^ n6675;
  assign n6665 = n6628 ^ n6431;
  assign n6666 = ~n6629 & ~n6665;
  assign n6667 = n6666 ^ n6431;
  assign n6868 = n6867 ^ n6667;
  assign n6656 = n5940 ^ x113;
  assign n6657 = n210 & n6656;
  assign n6658 = x111 & n219;
  assign n6659 = x112 & n214;
  assign n6660 = ~n6658 & ~n6659;
  assign n6661 = x113 & n259;
  assign n6662 = n6660 & ~n6661;
  assign n6663 = ~n6657 & n6662;
  assign n6664 = n6663 ^ x5;
  assign n6869 = n6868 ^ n6664;
  assign n6653 = n6630 ^ n6419;
  assign n6654 = n6631 & ~n6653;
  assign n6655 = n6654 ^ n6419;
  assign n6870 = n6869 ^ n6655;
  assign n6638 = ~x114 & ~n6165;
  assign n6639 = x115 & ~n6638;
  assign n6640 = x114 & ~n6167;
  assign n6641 = ~x115 & ~n6640;
  assign n6642 = ~n6639 & ~n6641;
  assign n6643 = n163 & ~n6642;
  assign n6644 = n6643 ^ x1;
  assign n6645 = n6644 ^ x116;
  assign n6646 = x0 & n6645;
  assign n6647 = ~x1 & x114;
  assign n6648 = ~x0 & ~n6647;
  assign n6649 = x1 & x115;
  assign n6650 = n6649 ^ x2;
  assign n6651 = n6648 & n6650;
  assign n6652 = ~n6646 & ~n6651;
  assign n6871 = n6870 ^ n6652;
  assign n6635 = n6632 ^ n6404;
  assign n6636 = ~n6633 & n6635;
  assign n6637 = n6636 ^ n6404;
  assign n6872 = n6871 ^ n6637;
  assign n7075 = x53 ^ x52;
  assign n7076 = n6561 & n7075;
  assign n7077 = n208 & n7076;
  assign n7070 = x50 & x51;
  assign n7066 = ~x50 & ~x51;
  assign n7078 = n7070 ^ n7066;
  assign n7079 = x52 & n7078;
  assign n7080 = n7079 ^ n7070;
  assign n7081 = ~n7077 & ~n7080;
  assign n7082 = x65 & ~n7081;
  assign n7083 = n149 & n7075;
  assign n7084 = x66 & n6561;
  assign n7085 = ~n7083 & n7084;
  assign n7086 = ~n7082 & ~n7085;
  assign n7087 = ~x53 & ~n7086;
  assign n7088 = x52 & ~x53;
  assign n7089 = n7070 & n7088;
  assign n7090 = x64 & n7089;
  assign n7091 = ~n7087 & ~n7090;
  assign n7071 = ~x52 & x64;
  assign n7092 = n7066 & n7071;
  assign n7093 = x53 & ~n7092;
  assign n7094 = n7086 & n7093;
  assign n7095 = n7091 & ~n7094;
  assign n7067 = x52 & x64;
  assign n7068 = n7066 & ~n7067;
  assign n7069 = ~n201 & ~n7068;
  assign n7072 = n7070 & ~n7071;
  assign n7073 = n7069 & ~n7072;
  assign n7074 = x53 & ~n7073;
  assign n7096 = n7095 ^ n7074;
  assign n7058 = n358 & n6326;
  assign n7059 = x68 & n6331;
  assign n7060 = x67 & n6565;
  assign n7061 = ~n7059 & ~n7060;
  assign n7062 = x69 & n6569;
  assign n7063 = n7061 & ~n7062;
  assign n7064 = ~n7058 & n7063;
  assign n7065 = n7064 ^ x50;
  assign n7097 = n7096 ^ n7065;
  assign n7055 = n6811 ^ n6804;
  assign n7056 = ~n6814 & ~n7055;
  assign n7057 = n7056 ^ n6813;
  assign n7098 = n7097 ^ n7057;
  assign n7047 = n520 & n5656;
  assign n7048 = x71 & n5662;
  assign n7049 = x70 & n5895;
  assign n7050 = ~n7048 & ~n7049;
  assign n7051 = x72 & n6111;
  assign n7052 = n7050 & ~n7051;
  assign n7053 = ~n7047 & n7052;
  assign n7054 = n7053 ^ x47;
  assign n7099 = n7098 ^ n7054;
  assign n7044 = n6823 ^ n6815;
  assign n7045 = ~n6830 & n7044;
  assign n7046 = n7045 ^ n6829;
  assign n7100 = n7099 ^ n7046;
  assign n7036 = n720 & n5010;
  assign n7037 = x74 & n5014;
  assign n7038 = x75 & n5226;
  assign n7039 = ~n7037 & ~n7038;
  assign n7040 = x73 & n5223;
  assign n7041 = n7039 & ~n7040;
  assign n7042 = ~n7036 & n7041;
  assign n7043 = n7042 ^ x44;
  assign n7101 = n7100 ^ n7043;
  assign n7033 = n6831 ^ n6788;
  assign n7034 = ~n6832 & ~n7033;
  assign n7035 = n7034 ^ n6788;
  assign n7102 = n7101 ^ n7035;
  assign n7025 = n953 & n4415;
  assign n7026 = x76 & n4420;
  assign n7027 = x78 & n4614;
  assign n7028 = ~n7026 & ~n7027;
  assign n7029 = x77 & n4410;
  assign n7030 = n7028 & ~n7029;
  assign n7031 = ~n7025 & n7030;
  assign n7032 = n7031 ^ x41;
  assign n7103 = n7102 ^ n7032;
  assign n7022 = n6844 ^ n6833;
  assign n7023 = ~n6845 & n7022;
  assign n7024 = n7023 ^ n6836;
  assign n7104 = n7103 ^ n7024;
  assign n7019 = n6846 ^ n6777;
  assign n7020 = ~n6847 & ~n7019;
  assign n7021 = n7020 ^ n6777;
  assign n7105 = n7104 ^ n7021;
  assign n7011 = n1230 & n3829;
  assign n7012 = x80 & n3833;
  assign n7013 = x81 & n4052;
  assign n7014 = ~n7012 & ~n7013;
  assign n7015 = x79 & n4049;
  assign n7016 = n7014 & ~n7015;
  assign n7017 = ~n7011 & n7016;
  assign n7018 = n7017 ^ x38;
  assign n7106 = n7105 ^ n7018;
  assign n7003 = n1547 & n3330;
  assign n7004 = x82 & n3500;
  assign n7005 = x83 & n3334;
  assign n7006 = ~n7004 & ~n7005;
  assign n7007 = x84 & n3502;
  assign n7008 = n7006 & ~n7007;
  assign n7009 = ~n7003 & n7008;
  assign n7010 = n7009 ^ x35;
  assign n7107 = n7106 ^ n7010;
  assign n7000 = n6848 ^ n6766;
  assign n7001 = n6849 & n7000;
  assign n7002 = n7001 ^ n6766;
  assign n7108 = n7107 ^ n7002;
  assign n6992 = n1903 & n2836;
  assign n6993 = x86 & n2840;
  assign n6994 = x85 & n2996;
  assign n6995 = ~n6993 & ~n6994;
  assign n6996 = x87 & n2998;
  assign n6997 = n6995 & ~n6996;
  assign n6998 = ~n6992 & n6997;
  assign n6999 = n6998 ^ x32;
  assign n7109 = n7108 ^ n6999;
  assign n6989 = n6763 ^ n6755;
  assign n6990 = n6851 & n6989;
  assign n6991 = n6990 ^ n6850;
  assign n7110 = n7109 ^ n6991;
  assign n6981 = n2292 & n2371;
  assign n6982 = x88 & n2528;
  assign n6983 = x90 & n2531;
  assign n6984 = ~n6982 & ~n6983;
  assign n6985 = x89 & n2377;
  assign n6986 = n6984 & ~n6985;
  assign n6987 = ~n6981 & n6986;
  assign n6988 = n6987 ^ x29;
  assign n7111 = n7110 ^ n6988;
  assign n6978 = n6852 ^ n6744;
  assign n6979 = n6853 & n6978;
  assign n6980 = n6979 ^ n6744;
  assign n7112 = n7111 ^ n6980;
  assign n6970 = n1969 & n2726;
  assign n6971 = x91 & n1978;
  assign n6972 = x93 & n2108;
  assign n6973 = ~n6971 & ~n6972;
  assign n6974 = x92 & n1973;
  assign n6975 = n6973 & ~n6974;
  assign n6976 = ~n6970 & n6975;
  assign n6977 = n6976 ^ x26;
  assign n7113 = n7112 ^ n6977;
  assign n6967 = n6854 ^ n6733;
  assign n6968 = ~n6855 & ~n6967;
  assign n6969 = n6968 ^ n6733;
  assign n7114 = n7113 ^ n6969;
  assign n6959 = n1624 & n3209;
  assign n6960 = x94 & n1742;
  assign n6961 = x95 & n1628;
  assign n6962 = ~n6960 & ~n6961;
  assign n6963 = x96 & n1744;
  assign n6964 = n6962 & ~n6963;
  assign n6965 = ~n6959 & n6964;
  assign n6966 = n6965 ^ x23;
  assign n7115 = n7114 ^ n6966;
  assign n6956 = n6856 ^ n6722;
  assign n6957 = n6857 & n6956;
  assign n6958 = n6957 ^ n6722;
  assign n7116 = n7115 ^ n6958;
  assign n6948 = n1296 & n3730;
  assign n6949 = x98 & n1300;
  assign n6950 = x97 & n1403;
  assign n6951 = ~n6949 & ~n6950;
  assign n6952 = x99 & n1406;
  assign n6953 = n6951 & ~n6952;
  assign n6954 = ~n6948 & n6953;
  assign n6955 = n6954 ^ x20;
  assign n7117 = n7116 ^ n6955;
  assign n6945 = n6858 ^ n6711;
  assign n6946 = ~n6859 & ~n6945;
  assign n6947 = n6946 ^ n6711;
  assign n7118 = n7117 ^ n6947;
  assign n6937 = n1008 & n4286;
  assign n6938 = x101 & n1012;
  assign n6939 = x100 & n1101;
  assign n6940 = ~n6938 & ~n6939;
  assign n6941 = x102 & n1104;
  assign n6942 = n6940 & ~n6941;
  assign n6943 = ~n6937 & n6942;
  assign n6944 = n6943 ^ x17;
  assign n7119 = n7118 ^ n6944;
  assign n6934 = n6860 ^ n6700;
  assign n6935 = n6861 & n6934;
  assign n6936 = n6935 ^ n6700;
  assign n7120 = n7119 ^ n6936;
  assign n6926 = n752 & n4867;
  assign n6927 = x103 & n825;
  assign n6928 = x105 & n828;
  assign n6929 = ~n6927 & ~n6928;
  assign n6930 = x104 & n757;
  assign n6931 = n6929 & ~n6930;
  assign n6932 = ~n6926 & n6931;
  assign n6933 = n6932 ^ x14;
  assign n7121 = n7120 ^ n6933;
  assign n6923 = n6862 ^ n6689;
  assign n6924 = ~n6863 & ~n6923;
  assign n6925 = n6924 ^ n6689;
  assign n7122 = n7121 ^ n6925;
  assign n6915 = n541 & ~n5506;
  assign n6916 = x106 & n612;
  assign n6917 = x107 & n547;
  assign n6918 = ~n6916 & ~n6917;
  assign n6919 = x108 & n615;
  assign n6920 = n6918 & ~n6919;
  assign n6921 = ~n6915 & n6920;
  assign n6922 = n6921 ^ x11;
  assign n7123 = n7122 ^ n6922;
  assign n6912 = n6864 ^ n6678;
  assign n6913 = n6865 & n6912;
  assign n6914 = n6913 ^ n6678;
  assign n7124 = n7123 ^ n6914;
  assign n6904 = n372 & n6178;
  assign n6905 = x109 & n433;
  assign n6906 = x111 & n428;
  assign n6907 = ~n6905 & ~n6906;
  assign n6908 = x110 & n376;
  assign n6909 = n6907 & ~n6908;
  assign n6910 = ~n6904 & n6909;
  assign n6911 = n6910 ^ x8;
  assign n7125 = n7124 ^ n6911;
  assign n6901 = n6866 ^ n6667;
  assign n6902 = ~n6867 & ~n6901;
  assign n6903 = n6902 ^ n6667;
  assign n7126 = n7125 ^ n6903;
  assign n6892 = n6168 ^ x114;
  assign n6893 = n210 & n6892;
  assign n6894 = x112 & n219;
  assign n6895 = x114 & n259;
  assign n6896 = ~n6894 & ~n6895;
  assign n6897 = x113 & n214;
  assign n6898 = n6896 & ~n6897;
  assign n6899 = ~n6893 & n6898;
  assign n6900 = n6899 ^ x5;
  assign n7127 = n7126 ^ n6900;
  assign n6889 = n6868 ^ n6655;
  assign n6890 = n6869 & ~n6889;
  assign n6891 = n6890 ^ n6655;
  assign n7128 = n7127 ^ n6891;
  assign n6876 = ~x116 & ~n6639;
  assign n6877 = x116 & ~n6641;
  assign n6878 = ~n6876 & ~n6877;
  assign n6879 = n163 & ~n6878;
  assign n6880 = n6879 ^ x1;
  assign n6881 = n6880 ^ x117;
  assign n6882 = x0 & n6881;
  assign n6883 = ~x1 & x115;
  assign n6884 = ~x0 & ~n6883;
  assign n6885 = x1 & x116;
  assign n6886 = n6885 ^ x2;
  assign n6887 = n6884 & n6886;
  assign n6888 = ~n6882 & ~n6887;
  assign n7129 = n7128 ^ n6888;
  assign n6873 = n6870 ^ n6637;
  assign n6874 = n6871 & n6873;
  assign n6875 = n6874 ^ n6637;
  assign n7130 = n7129 ^ n6875;
  assign n7339 = n1054 & n4415;
  assign n7340 = x77 & n4420;
  assign n7341 = x79 & n4614;
  assign n7342 = ~n7340 & ~n7341;
  assign n7343 = x78 & n4410;
  assign n7344 = n7342 & ~n7343;
  assign n7345 = ~n7339 & n7344;
  assign n7346 = n7345 ^ x41;
  assign n7336 = n7102 ^ n7024;
  assign n7337 = n7103 & n7336;
  assign n7338 = n7337 ^ n7024;
  assign n7347 = n7346 ^ n7338;
  assign n7328 = n7074 & ~n7095;
  assign n7315 = x52 ^ x51;
  assign n7316 = n7075 & ~n7315;
  assign n7317 = ~n6561 & n7316;
  assign n7318 = x65 & n7317;
  assign n7319 = n6561 & ~n7075;
  assign n7320 = x67 & n7319;
  assign n7321 = ~n7318 & ~n7320;
  assign n7322 = x66 & n7080;
  assign n7323 = n7321 & ~n7322;
  assign n7324 = n264 & n7076;
  assign n7325 = n7323 & ~n7324;
  assign n7326 = n7325 ^ x53;
  assign n7313 = x54 ^ x53;
  assign n7314 = x64 & n7313;
  assign n7327 = n7326 ^ n7314;
  assign n7329 = n7328 ^ n7327;
  assign n7305 = n416 & n6326;
  assign n7306 = x68 & n6565;
  assign n7307 = x69 & n6331;
  assign n7308 = ~n7306 & ~n7307;
  assign n7309 = x70 & n6569;
  assign n7310 = n7308 & ~n7309;
  assign n7311 = ~n7305 & n7310;
  assign n7312 = n7311 ^ x50;
  assign n7330 = n7329 ^ n7312;
  assign n7302 = n7096 ^ n7057;
  assign n7303 = ~n7097 & ~n7302;
  assign n7304 = n7303 ^ n7057;
  assign n7331 = n7330 ^ n7304;
  assign n7294 = ~n594 & n5656;
  assign n7295 = x72 & n5662;
  assign n7296 = x71 & n5895;
  assign n7297 = ~n7295 & ~n7296;
  assign n7298 = x73 & n6111;
  assign n7299 = n7297 & ~n7298;
  assign n7300 = ~n7294 & n7299;
  assign n7301 = n7300 ^ x47;
  assign n7332 = n7331 ^ n7301;
  assign n7291 = n7098 ^ n7046;
  assign n7292 = n7099 & n7291;
  assign n7293 = n7292 ^ n7046;
  assign n7333 = n7332 ^ n7293;
  assign n7283 = n799 & n5010;
  assign n7284 = x74 & n5223;
  assign n7285 = x75 & n5014;
  assign n7286 = ~n7284 & ~n7285;
  assign n7287 = x76 & n5226;
  assign n7288 = n7286 & ~n7287;
  assign n7289 = ~n7283 & n7288;
  assign n7290 = n7289 ^ x44;
  assign n7334 = n7333 ^ n7290;
  assign n7280 = n7100 ^ n7035;
  assign n7281 = ~n7101 & ~n7280;
  assign n7282 = n7281 ^ n7035;
  assign n7335 = n7334 ^ n7282;
  assign n7348 = n7347 ^ n7335;
  assign n7272 = n1345 & n3829;
  assign n7273 = x80 & n4049;
  assign n7274 = x82 & n4052;
  assign n7275 = ~n7273 & ~n7274;
  assign n7276 = x81 & n3833;
  assign n7277 = n7275 & ~n7276;
  assign n7278 = ~n7272 & n7277;
  assign n7279 = n7278 ^ x38;
  assign n7349 = n7348 ^ n7279;
  assign n7269 = n7104 ^ n7018;
  assign n7270 = ~n7105 & ~n7269;
  assign n7271 = n7270 ^ n7021;
  assign n7350 = n7349 ^ n7271;
  assign n7261 = n1674 & n3330;
  assign n7262 = x83 & n3500;
  assign n7263 = x85 & n3502;
  assign n7264 = ~n7262 & ~n7263;
  assign n7265 = x84 & n3334;
  assign n7266 = n7264 & ~n7265;
  assign n7267 = ~n7261 & n7266;
  assign n7268 = n7267 ^ x35;
  assign n7351 = n7350 ^ n7268;
  assign n7258 = n7106 ^ n7002;
  assign n7259 = n7107 & n7258;
  assign n7260 = n7259 ^ n7002;
  assign n7352 = n7351 ^ n7260;
  assign n7250 = n2040 & n2836;
  assign n7251 = x87 & n2840;
  assign n7252 = x86 & n2996;
  assign n7253 = ~n7251 & ~n7252;
  assign n7254 = x88 & n2998;
  assign n7255 = n7253 & ~n7254;
  assign n7256 = ~n7250 & n7255;
  assign n7257 = n7256 ^ x32;
  assign n7353 = n7352 ^ n7257;
  assign n7247 = n7108 ^ n6991;
  assign n7248 = ~n7109 & n7247;
  assign n7249 = n7248 ^ n6991;
  assign n7354 = n7353 ^ n7249;
  assign n7239 = n2371 & n2447;
  assign n7240 = x89 & n2528;
  assign n7241 = x90 & n2377;
  assign n7242 = ~n7240 & ~n7241;
  assign n7243 = x91 & n2531;
  assign n7244 = n7242 & ~n7243;
  assign n7245 = ~n7239 & n7244;
  assign n7246 = n7245 ^ x29;
  assign n7355 = n7354 ^ n7246;
  assign n7236 = n7110 ^ n6980;
  assign n7237 = ~n7111 & ~n7236;
  assign n7238 = n7237 ^ n6980;
  assign n7356 = n7355 ^ n7238;
  assign n7228 = n1969 & n2895;
  assign n7229 = x93 & n1973;
  assign n7230 = x92 & n1978;
  assign n7231 = ~n7229 & ~n7230;
  assign n7232 = x94 & n2108;
  assign n7233 = n7231 & ~n7232;
  assign n7234 = ~n7228 & n7233;
  assign n7235 = n7234 ^ x26;
  assign n7357 = n7356 ^ n7235;
  assign n7225 = n7112 ^ n6969;
  assign n7226 = n7113 & n7225;
  assign n7227 = n7226 ^ n6969;
  assign n7358 = n7357 ^ n7227;
  assign n7217 = n1624 & n3388;
  assign n7218 = x96 & n1628;
  assign n7219 = x95 & n1742;
  assign n7220 = ~n7218 & ~n7219;
  assign n7221 = x97 & n1744;
  assign n7222 = n7220 & ~n7221;
  assign n7223 = ~n7217 & n7222;
  assign n7224 = n7223 ^ x23;
  assign n7359 = n7358 ^ n7224;
  assign n7214 = n7114 ^ n6958;
  assign n7215 = ~n7115 & ~n7214;
  assign n7216 = n7215 ^ n6958;
  assign n7360 = n7359 ^ n7216;
  assign n7206 = n1296 & n3925;
  assign n7207 = x98 & n1403;
  assign n7208 = x99 & n1300;
  assign n7209 = ~n7207 & ~n7208;
  assign n7210 = x100 & n1406;
  assign n7211 = n7209 & ~n7210;
  assign n7212 = ~n7206 & n7211;
  assign n7213 = n7212 ^ x20;
  assign n7361 = n7360 ^ n7213;
  assign n7203 = n7116 ^ n6947;
  assign n7204 = n7117 & n7203;
  assign n7205 = n7204 ^ n6947;
  assign n7362 = n7361 ^ n7205;
  assign n7195 = n1008 & n4481;
  assign n7196 = x102 & n1012;
  assign n7197 = x101 & n1101;
  assign n7198 = ~n7196 & ~n7197;
  assign n7199 = x103 & n1104;
  assign n7200 = n7198 & ~n7199;
  assign n7201 = ~n7195 & n7200;
  assign n7202 = n7201 ^ x17;
  assign n7363 = n7362 ^ n7202;
  assign n7192 = n7118 ^ n6936;
  assign n7193 = ~n7119 & ~n7192;
  assign n7194 = n7193 ^ n6936;
  assign n7364 = n7363 ^ n7194;
  assign n7184 = n752 & n5088;
  assign n7185 = x104 & n825;
  assign n7186 = x106 & n828;
  assign n7187 = ~n7185 & ~n7186;
  assign n7188 = x105 & n757;
  assign n7189 = n7187 & ~n7188;
  assign n7190 = ~n7184 & n7189;
  assign n7191 = n7190 ^ x14;
  assign n7365 = n7364 ^ n7191;
  assign n7176 = n541 & ~n5737;
  assign n7177 = x107 & n612;
  assign n7178 = x108 & n547;
  assign n7179 = ~n7177 & ~n7178;
  assign n7180 = x109 & n615;
  assign n7181 = n7179 & ~n7180;
  assign n7182 = ~n7176 & n7181;
  assign n7183 = n7182 ^ x11;
  assign n7366 = n7365 ^ n7183;
  assign n7173 = n7120 ^ n6925;
  assign n7174 = n7121 & n7173;
  assign n7175 = n7174 ^ n6925;
  assign n7367 = n7366 ^ n7175;
  assign n7170 = n7122 ^ n6914;
  assign n7171 = ~n7123 & ~n7170;
  assign n7172 = n7171 ^ n6914;
  assign n7368 = n7367 ^ n7172;
  assign n7162 = n372 & n6420;
  assign n7163 = x110 & n433;
  assign n7164 = x112 & n428;
  assign n7165 = ~n7163 & ~n7164;
  assign n7166 = x111 & n376;
  assign n7167 = n7165 & ~n7166;
  assign n7168 = ~n7162 & n7167;
  assign n7169 = n7168 ^ x8;
  assign n7369 = n7368 ^ n7169;
  assign n7159 = n7124 ^ n6903;
  assign n7160 = n7125 & n7159;
  assign n7161 = n7160 ^ n6903;
  assign n7370 = n7369 ^ n7161;
  assign n7150 = n6410 ^ x115;
  assign n7151 = n210 & n7150;
  assign n7152 = x113 & n219;
  assign n7153 = x115 & n259;
  assign n7154 = ~n7152 & ~n7153;
  assign n7155 = x114 & n214;
  assign n7156 = n7154 & ~n7155;
  assign n7157 = ~n7151 & n7156;
  assign n7158 = n7157 ^ x5;
  assign n7371 = n7370 ^ n7158;
  assign n7147 = n7126 ^ n6891;
  assign n7148 = ~n7127 & n7147;
  assign n7149 = n7148 ^ n6891;
  assign n7372 = n7371 ^ n7149;
  assign n7134 = x117 & ~n6876;
  assign n7135 = ~x117 & ~n6877;
  assign n7136 = ~n7134 & ~n7135;
  assign n7137 = n163 & ~n7136;
  assign n7138 = n7137 ^ x1;
  assign n7139 = n7138 ^ x118;
  assign n7140 = x0 & ~n7139;
  assign n7141 = x117 ^ x2;
  assign n7142 = x1 & n7141;
  assign n7143 = ~x0 & ~n7142;
  assign n7144 = ~x116 & n156;
  assign n7145 = n7143 & ~n7144;
  assign n7146 = ~n7140 & ~n7145;
  assign n7373 = n7372 ^ n7146;
  assign n7131 = n7128 ^ n6875;
  assign n7132 = ~n7129 & ~n7131;
  assign n7133 = n7132 ^ n6875;
  assign n7374 = n7373 ^ n7133;
  assign n7584 = n877 & n5010;
  assign n7585 = x75 & n5223;
  assign n7586 = x77 & n5226;
  assign n7587 = ~n7585 & ~n7586;
  assign n7588 = x76 & n5014;
  assign n7589 = n7587 & ~n7588;
  assign n7590 = ~n7584 & n7589;
  assign n7591 = n7590 ^ x44;
  assign n7581 = n7333 ^ n7282;
  assign n7582 = ~n7334 & ~n7581;
  assign n7583 = n7582 ^ n7282;
  assign n7592 = n7591 ^ n7583;
  assign n7574 = ~n7314 & ~n7328;
  assign n7575 = ~n7326 & ~n7574;
  assign n7565 = n300 & n7076;
  assign n7566 = x67 & n7080;
  assign n7567 = x66 & n7317;
  assign n7568 = ~n7566 & ~n7567;
  assign n7569 = x68 & n7319;
  assign n7570 = n7568 & ~n7569;
  assign n7571 = ~n7565 & n7570;
  assign n7572 = n7571 ^ x53;
  assign n7558 = x65 ^ x54;
  assign n7559 = n7313 & ~n7558;
  assign n7560 = n7559 ^ x53;
  assign n7561 = n7560 ^ x55;
  assign n7562 = x64 & n7561;
  assign n7563 = n149 & n7313;
  assign n7564 = ~n7562 & ~n7563;
  assign n7573 = n7572 ^ n7564;
  assign n7576 = n7575 ^ n7573;
  assign n7550 = n467 & n6326;
  assign n7551 = x70 & n6331;
  assign n7552 = x69 & n6565;
  assign n7553 = ~n7551 & ~n7552;
  assign n7554 = x71 & n6569;
  assign n7555 = n7553 & ~n7554;
  assign n7556 = ~n7550 & n7555;
  assign n7557 = n7556 ^ x50;
  assign n7577 = n7576 ^ n7557;
  assign n7547 = n7329 ^ n7304;
  assign n7548 = ~n7330 & ~n7547;
  assign n7549 = n7548 ^ n7304;
  assign n7578 = n7577 ^ n7549;
  assign n7539 = ~n656 & n5656;
  assign n7540 = x73 & n5662;
  assign n7541 = x72 & n5895;
  assign n7542 = ~n7540 & ~n7541;
  assign n7543 = x74 & n6111;
  assign n7544 = n7542 & ~n7543;
  assign n7545 = ~n7539 & n7544;
  assign n7546 = n7545 ^ x47;
  assign n7579 = n7578 ^ n7546;
  assign n7536 = n7331 ^ n7293;
  assign n7537 = n7332 & n7536;
  assign n7538 = n7537 ^ n7293;
  assign n7580 = n7579 ^ n7538;
  assign n7593 = n7592 ^ n7580;
  assign n7528 = ~n1141 & n4415;
  assign n7529 = x78 & n4420;
  assign n7530 = x79 & n4410;
  assign n7531 = ~n7529 & ~n7530;
  assign n7532 = x80 & n4614;
  assign n7533 = n7531 & ~n7532;
  assign n7534 = ~n7528 & n7533;
  assign n7535 = n7534 ^ x41;
  assign n7594 = n7593 ^ n7535;
  assign n7525 = n7346 ^ n7335;
  assign n7526 = ~n7347 & n7525;
  assign n7527 = n7526 ^ n7338;
  assign n7595 = n7594 ^ n7527;
  assign n7517 = n1445 & n3829;
  assign n7518 = x81 & n4049;
  assign n7519 = x82 & n3833;
  assign n7520 = ~n7518 & ~n7519;
  assign n7521 = x83 & n4052;
  assign n7522 = n7520 & ~n7521;
  assign n7523 = ~n7517 & n7522;
  assign n7524 = n7523 ^ x38;
  assign n7596 = n7595 ^ n7524;
  assign n7514 = n7348 ^ n7271;
  assign n7515 = ~n7349 & ~n7514;
  assign n7516 = n7515 ^ n7271;
  assign n7597 = n7596 ^ n7516;
  assign n7506 = n1787 & n3330;
  assign n7507 = x84 & n3500;
  assign n7508 = x86 & n3502;
  assign n7509 = ~n7507 & ~n7508;
  assign n7510 = x85 & n3334;
  assign n7511 = n7509 & ~n7510;
  assign n7512 = ~n7506 & n7511;
  assign n7513 = n7512 ^ x35;
  assign n7598 = n7597 ^ n7513;
  assign n7503 = n7350 ^ n7260;
  assign n7504 = n7351 & n7503;
  assign n7505 = n7504 ^ n7260;
  assign n7599 = n7598 ^ n7505;
  assign n7495 = n2164 & n2836;
  assign n7496 = x87 & n2996;
  assign n7497 = x88 & n2840;
  assign n7498 = ~n7496 & ~n7497;
  assign n7499 = x89 & n2998;
  assign n7500 = n7498 & ~n7499;
  assign n7501 = ~n7495 & n7500;
  assign n7502 = n7501 ^ x32;
  assign n7600 = n7599 ^ n7502;
  assign n7492 = n7352 ^ n7249;
  assign n7493 = ~n7353 & n7492;
  assign n7494 = n7493 ^ n7249;
  assign n7601 = n7600 ^ n7494;
  assign n7484 = n2371 & n2585;
  assign n7485 = x90 & n2528;
  assign n7486 = x91 & n2377;
  assign n7487 = ~n7485 & ~n7486;
  assign n7488 = x92 & n2531;
  assign n7489 = n7487 & ~n7488;
  assign n7490 = ~n7484 & n7489;
  assign n7491 = n7490 ^ x29;
  assign n7602 = n7601 ^ n7491;
  assign n7481 = n7354 ^ n7238;
  assign n7482 = ~n7355 & ~n7481;
  assign n7483 = n7482 ^ n7238;
  assign n7603 = n7602 ^ n7483;
  assign n7473 = n1969 & n3054;
  assign n7474 = x93 & n1978;
  assign n7475 = x95 & n2108;
  assign n7476 = ~n7474 & ~n7475;
  assign n7477 = x94 & n1973;
  assign n7478 = n7476 & ~n7477;
  assign n7479 = ~n7473 & n7478;
  assign n7480 = n7479 ^ x26;
  assign n7604 = n7603 ^ n7480;
  assign n7470 = n7356 ^ n7227;
  assign n7471 = n7357 & n7470;
  assign n7472 = n7471 ^ n7227;
  assign n7605 = n7604 ^ n7472;
  assign n7462 = n1624 & n3556;
  assign n7463 = x96 & n1742;
  assign n7464 = x97 & n1628;
  assign n7465 = ~n7463 & ~n7464;
  assign n7466 = x98 & n1744;
  assign n7467 = n7465 & ~n7466;
  assign n7468 = ~n7462 & n7467;
  assign n7469 = n7468 ^ x23;
  assign n7606 = n7605 ^ n7469;
  assign n7459 = n7358 ^ n7216;
  assign n7460 = ~n7359 & ~n7459;
  assign n7461 = n7460 ^ n7216;
  assign n7607 = n7606 ^ n7461;
  assign n7451 = n1296 & n4105;
  assign n7452 = x100 & n1300;
  assign n7453 = x99 & n1403;
  assign n7454 = ~n7452 & ~n7453;
  assign n7455 = x101 & n1406;
  assign n7456 = n7454 & ~n7455;
  assign n7457 = ~n7451 & n7456;
  assign n7458 = n7457 ^ x20;
  assign n7608 = n7607 ^ n7458;
  assign n7448 = n7360 ^ n7205;
  assign n7449 = n7361 & n7448;
  assign n7450 = n7449 ^ n7205;
  assign n7609 = n7608 ^ n7450;
  assign n7440 = n1008 & n4670;
  assign n7441 = x103 & n1012;
  assign n7442 = x102 & n1101;
  assign n7443 = ~n7441 & ~n7442;
  assign n7444 = x104 & n1104;
  assign n7445 = n7443 & ~n7444;
  assign n7446 = ~n7440 & n7445;
  assign n7447 = n7446 ^ x17;
  assign n7610 = n7609 ^ n7447;
  assign n7437 = n7362 ^ n7194;
  assign n7438 = ~n7363 & ~n7437;
  assign n7439 = n7438 ^ n7194;
  assign n7611 = n7610 ^ n7439;
  assign n7429 = n752 & n5297;
  assign n7430 = x105 & n825;
  assign n7431 = x106 & n757;
  assign n7432 = ~n7430 & ~n7431;
  assign n7433 = x107 & n828;
  assign n7434 = n7432 & ~n7433;
  assign n7435 = ~n7429 & n7434;
  assign n7436 = n7435 ^ x14;
  assign n7612 = n7611 ^ n7436;
  assign n7426 = n7364 ^ n7175;
  assign n7427 = n7365 & n7426;
  assign n7428 = n7427 ^ n7175;
  assign n7613 = n7612 ^ n7428;
  assign n7418 = n541 & n5955;
  assign n7419 = x109 & n547;
  assign n7420 = x110 & n615;
  assign n7421 = ~n7419 & ~n7420;
  assign n7422 = x108 & n612;
  assign n7423 = n7421 & ~n7422;
  assign n7424 = ~n7418 & n7423;
  assign n7425 = n7424 ^ x11;
  assign n7614 = n7613 ^ n7425;
  assign n7413 = n7365 ^ n7175;
  assign n7414 = n7413 ^ n7183;
  assign n7415 = n7183 ^ n7172;
  assign n7416 = ~n7414 & ~n7415;
  assign n7417 = n7416 ^ n7172;
  assign n7615 = n7614 ^ n7417;
  assign n7405 = n372 & n6656;
  assign n7406 = x111 & n433;
  assign n7407 = x113 & n428;
  assign n7408 = ~n7406 & ~n7407;
  assign n7409 = x112 & n376;
  assign n7410 = n7408 & ~n7409;
  assign n7411 = ~n7405 & n7410;
  assign n7412 = n7411 ^ x8;
  assign n7616 = n7615 ^ n7412;
  assign n7402 = n7368 ^ n7161;
  assign n7403 = n7369 & n7402;
  assign n7404 = n7403 ^ n7161;
  assign n7617 = n7616 ^ n7404;
  assign n7393 = n6642 ^ x116;
  assign n7394 = n210 & n7393;
  assign n7395 = x114 & n219;
  assign n7396 = x115 & n214;
  assign n7397 = ~n7395 & ~n7396;
  assign n7398 = x116 & n259;
  assign n7399 = n7397 & ~n7398;
  assign n7400 = ~n7394 & n7399;
  assign n7401 = n7400 ^ x5;
  assign n7618 = n7617 ^ n7401;
  assign n7390 = n7370 ^ n7149;
  assign n7391 = ~n7371 & n7390;
  assign n7392 = n7391 ^ n7149;
  assign n7619 = n7618 ^ n7392;
  assign n7378 = x118 ^ x117;
  assign n7379 = ~n7136 & n7378;
  assign n7380 = n163 & ~n7379;
  assign n7381 = n7380 ^ x1;
  assign n7382 = n7381 ^ x119;
  assign n7383 = x0 & ~n7382;
  assign n7384 = ~x117 & n156;
  assign n7385 = ~x0 & ~n7384;
  assign n7386 = x118 ^ x2;
  assign n7387 = x1 & n7386;
  assign n7388 = n7385 & ~n7387;
  assign n7389 = ~n7383 & ~n7388;
  assign n7620 = n7619 ^ n7389;
  assign n7375 = n7372 ^ n7133;
  assign n7376 = n7373 & ~n7375;
  assign n7377 = n7376 ^ n7133;
  assign n7621 = n7620 ^ n7377;
  assign n7847 = n358 & n7076;
  assign n7848 = x67 & n7317;
  assign n7849 = x69 & n7319;
  assign n7850 = ~n7848 & ~n7849;
  assign n7851 = x68 & n7080;
  assign n7852 = n7850 & ~n7851;
  assign n7853 = ~n7847 & n7852;
  assign n7854 = n7853 ^ x53;
  assign n7829 = x56 ^ x55;
  assign n7830 = n7313 & n7829;
  assign n7831 = n208 & n7830;
  assign n7824 = x53 & x54;
  assign n7820 = ~x53 & ~x54;
  assign n7832 = n7824 ^ n7820;
  assign n7833 = x55 & n7832;
  assign n7834 = n7833 ^ n7824;
  assign n7835 = ~n7831 & ~n7834;
  assign n7836 = x65 & ~n7835;
  assign n7837 = x55 ^ x54;
  assign n7838 = n7829 & ~n7837;
  assign n7839 = ~n7313 & n7838;
  assign n7840 = x64 & n7839;
  assign n7841 = n149 & n7829;
  assign n7842 = x66 & n7313;
  assign n7843 = ~n7841 & n7842;
  assign n7844 = ~n7840 & ~n7843;
  assign n7845 = ~n7836 & n7844;
  assign n7821 = x55 & x64;
  assign n7822 = n7820 & ~n7821;
  assign n7823 = ~n201 & ~n7822;
  assign n7825 = ~x55 & x64;
  assign n7826 = n7824 & ~n7825;
  assign n7827 = n7823 & ~n7826;
  assign n7828 = x56 & n7827;
  assign n7846 = n7845 ^ n7828;
  assign n7855 = n7854 ^ n7846;
  assign n7817 = n7575 ^ n7572;
  assign n7818 = ~n7573 & ~n7817;
  assign n7819 = n7818 ^ n7575;
  assign n7856 = n7855 ^ n7819;
  assign n7809 = n520 & n6326;
  assign n7810 = x71 & n6331;
  assign n7811 = x70 & n6565;
  assign n7812 = ~n7810 & ~n7811;
  assign n7813 = x72 & n6569;
  assign n7814 = n7812 & ~n7813;
  assign n7815 = ~n7809 & n7814;
  assign n7816 = n7815 ^ x50;
  assign n7857 = n7856 ^ n7816;
  assign n7806 = n7576 ^ n7549;
  assign n7807 = n7577 & n7806;
  assign n7808 = n7807 ^ n7549;
  assign n7858 = n7857 ^ n7808;
  assign n7798 = n720 & n5656;
  assign n7799 = x74 & n5662;
  assign n7800 = x73 & n5895;
  assign n7801 = ~n7799 & ~n7800;
  assign n7802 = x75 & n6111;
  assign n7803 = n7801 & ~n7802;
  assign n7804 = ~n7798 & n7803;
  assign n7805 = n7804 ^ x47;
  assign n7859 = n7858 ^ n7805;
  assign n7795 = n7578 ^ n7538;
  assign n7796 = ~n7579 & ~n7795;
  assign n7797 = n7796 ^ n7538;
  assign n7860 = n7859 ^ n7797;
  assign n7787 = n953 & n5010;
  assign n7788 = x76 & n5223;
  assign n7789 = x77 & n5014;
  assign n7790 = ~n7788 & ~n7789;
  assign n7791 = x78 & n5226;
  assign n7792 = n7790 & ~n7791;
  assign n7793 = ~n7787 & n7792;
  assign n7794 = n7793 ^ x44;
  assign n7861 = n7860 ^ n7794;
  assign n7779 = n1230 & n4415;
  assign n7780 = x79 & n4420;
  assign n7781 = x80 & n4410;
  assign n7782 = ~n7780 & ~n7781;
  assign n7783 = x81 & n4614;
  assign n7784 = n7782 & ~n7783;
  assign n7785 = ~n7779 & n7784;
  assign n7786 = n7785 ^ x41;
  assign n7862 = n7861 ^ n7786;
  assign n7776 = n7591 ^ n7580;
  assign n7777 = ~n7592 & n7776;
  assign n7778 = n7777 ^ n7583;
  assign n7863 = n7862 ^ n7778;
  assign n7773 = n7593 ^ n7527;
  assign n7774 = ~n7594 & ~n7773;
  assign n7775 = n7774 ^ n7527;
  assign n7864 = n7863 ^ n7775;
  assign n7765 = n1547 & n3829;
  assign n7766 = x82 & n4049;
  assign n7767 = x83 & n3833;
  assign n7768 = ~n7766 & ~n7767;
  assign n7769 = x84 & n4052;
  assign n7770 = n7768 & ~n7769;
  assign n7771 = ~n7765 & n7770;
  assign n7772 = n7771 ^ x38;
  assign n7865 = n7864 ^ n7772;
  assign n7762 = n7595 ^ n7516;
  assign n7763 = n7596 & n7762;
  assign n7764 = n7763 ^ n7516;
  assign n7866 = n7865 ^ n7764;
  assign n7754 = n1903 & n3330;
  assign n7755 = x85 & n3500;
  assign n7756 = x86 & n3334;
  assign n7757 = ~n7755 & ~n7756;
  assign n7758 = x87 & n3502;
  assign n7759 = n7757 & ~n7758;
  assign n7760 = ~n7754 & n7759;
  assign n7761 = n7760 ^ x35;
  assign n7867 = n7866 ^ n7761;
  assign n7751 = n7597 ^ n7505;
  assign n7752 = ~n7598 & ~n7751;
  assign n7753 = n7752 ^ n7505;
  assign n7868 = n7867 ^ n7753;
  assign n7743 = n2292 & n2836;
  assign n7744 = x89 & n2840;
  assign n7745 = x88 & n2996;
  assign n7746 = ~n7744 & ~n7745;
  assign n7747 = x90 & n2998;
  assign n7748 = n7746 & ~n7747;
  assign n7749 = ~n7743 & n7748;
  assign n7750 = n7749 ^ x32;
  assign n7869 = n7868 ^ n7750;
  assign n7740 = n7599 ^ n7494;
  assign n7741 = n7600 & ~n7740;
  assign n7742 = n7741 ^ n7494;
  assign n7870 = n7869 ^ n7742;
  assign n7732 = n2371 & n2726;
  assign n7733 = x91 & n2528;
  assign n7734 = x92 & n2377;
  assign n7735 = ~n7733 & ~n7734;
  assign n7736 = x93 & n2531;
  assign n7737 = n7735 & ~n7736;
  assign n7738 = ~n7732 & n7737;
  assign n7739 = n7738 ^ x29;
  assign n7871 = n7870 ^ n7739;
  assign n7729 = n7601 ^ n7483;
  assign n7730 = n7602 & n7729;
  assign n7731 = n7730 ^ n7483;
  assign n7872 = n7871 ^ n7731;
  assign n7721 = n1969 & n3209;
  assign n7722 = x94 & n1978;
  assign n7723 = x95 & n1973;
  assign n7724 = ~n7722 & ~n7723;
  assign n7725 = x96 & n2108;
  assign n7726 = n7724 & ~n7725;
  assign n7727 = ~n7721 & n7726;
  assign n7728 = n7727 ^ x26;
  assign n7873 = n7872 ^ n7728;
  assign n7718 = n7603 ^ n7472;
  assign n7719 = ~n7604 & ~n7718;
  assign n7720 = n7719 ^ n7472;
  assign n7874 = n7873 ^ n7720;
  assign n7710 = n1624 & n3730;
  assign n7711 = x97 & n1742;
  assign n7712 = x98 & n1628;
  assign n7713 = ~n7711 & ~n7712;
  assign n7714 = x99 & n1744;
  assign n7715 = n7713 & ~n7714;
  assign n7716 = ~n7710 & n7715;
  assign n7717 = n7716 ^ x23;
  assign n7875 = n7874 ^ n7717;
  assign n7707 = n7605 ^ n7461;
  assign n7708 = n7606 & n7707;
  assign n7709 = n7708 ^ n7461;
  assign n7876 = n7875 ^ n7709;
  assign n7699 = n1296 & n4286;
  assign n7700 = x100 & n1403;
  assign n7701 = x101 & n1300;
  assign n7702 = ~n7700 & ~n7701;
  assign n7703 = x102 & n1406;
  assign n7704 = n7702 & ~n7703;
  assign n7705 = ~n7699 & n7704;
  assign n7706 = n7705 ^ x20;
  assign n7877 = n7876 ^ n7706;
  assign n7696 = n7607 ^ n7450;
  assign n7697 = ~n7608 & ~n7696;
  assign n7698 = n7697 ^ n7450;
  assign n7878 = n7877 ^ n7698;
  assign n7688 = n1008 & n4867;
  assign n7689 = x103 & n1101;
  assign n7690 = x104 & n1012;
  assign n7691 = ~n7689 & ~n7690;
  assign n7692 = x105 & n1104;
  assign n7693 = n7691 & ~n7692;
  assign n7694 = ~n7688 & n7693;
  assign n7695 = n7694 ^ x17;
  assign n7879 = n7878 ^ n7695;
  assign n7685 = n7609 ^ n7439;
  assign n7686 = n7610 & n7685;
  assign n7687 = n7686 ^ n7439;
  assign n7880 = n7879 ^ n7687;
  assign n7677 = n752 & ~n5506;
  assign n7678 = x106 & n825;
  assign n7679 = x107 & n757;
  assign n7680 = ~n7678 & ~n7679;
  assign n7681 = x108 & n828;
  assign n7682 = n7680 & ~n7681;
  assign n7683 = ~n7677 & n7682;
  assign n7684 = n7683 ^ x14;
  assign n7881 = n7880 ^ n7684;
  assign n7674 = n7611 ^ n7428;
  assign n7675 = ~n7612 & ~n7674;
  assign n7676 = n7675 ^ n7428;
  assign n7882 = n7881 ^ n7676;
  assign n7666 = n541 & n6178;
  assign n7667 = x109 & n612;
  assign n7668 = x111 & n615;
  assign n7669 = ~n7667 & ~n7668;
  assign n7670 = x110 & n547;
  assign n7671 = n7669 & ~n7670;
  assign n7672 = ~n7666 & n7671;
  assign n7673 = n7672 ^ x11;
  assign n7883 = n7882 ^ n7673;
  assign n7663 = n7613 ^ n7417;
  assign n7664 = n7614 & n7663;
  assign n7665 = n7664 ^ n7417;
  assign n7884 = n7883 ^ n7665;
  assign n7655 = n372 & n6892;
  assign n7656 = x112 & n433;
  assign n7657 = x113 & n376;
  assign n7658 = ~n7656 & ~n7657;
  assign n7659 = x114 & n428;
  assign n7660 = n7658 & ~n7659;
  assign n7661 = ~n7655 & n7660;
  assign n7662 = n7661 ^ x8;
  assign n7885 = n7884 ^ n7662;
  assign n7652 = n7615 ^ n7404;
  assign n7653 = ~n7616 & ~n7652;
  assign n7654 = n7653 ^ n7404;
  assign n7886 = n7885 ^ n7654;
  assign n7643 = n6878 ^ x117;
  assign n7644 = n210 & n7643;
  assign n7645 = x115 & n219;
  assign n7646 = x116 & n214;
  assign n7647 = ~n7645 & ~n7646;
  assign n7648 = x117 & n259;
  assign n7649 = n7647 & ~n7648;
  assign n7650 = ~n7644 & n7649;
  assign n7651 = n7650 ^ x5;
  assign n7887 = n7886 ^ n7651;
  assign n7640 = n7617 ^ n7392;
  assign n7641 = n7618 & ~n7640;
  assign n7642 = n7641 ^ n7392;
  assign n7888 = n7887 ^ n7642;
  assign n7625 = ~x118 & x119;
  assign n7626 = ~n7134 & n7625;
  assign n7627 = x118 & ~x119;
  assign n7628 = ~n7135 & n7627;
  assign n7629 = ~n7626 & ~n7628;
  assign n7630 = n163 & n7629;
  assign n7631 = n7630 ^ x1;
  assign n7632 = n7631 ^ x120;
  assign n7633 = x0 & ~n7632;
  assign n7634 = x119 ^ x2;
  assign n7635 = x1 & n7634;
  assign n7636 = ~x0 & ~n7635;
  assign n7637 = ~x118 & n156;
  assign n7638 = n7636 & ~n7637;
  assign n7639 = ~n7633 & ~n7638;
  assign n7889 = n7888 ^ n7639;
  assign n7622 = n7619 ^ n7377;
  assign n7623 = ~n7620 & n7622;
  assign n7624 = n7623 ^ n7377;
  assign n7890 = n7889 ^ n7624;
  assign n8125 = n1054 & n5010;
  assign n8126 = x77 & n5223;
  assign n8127 = x79 & n5226;
  assign n8128 = ~n8126 & ~n8127;
  assign n8129 = x78 & n5014;
  assign n8130 = n8128 & ~n8129;
  assign n8131 = ~n8125 & n8130;
  assign n8132 = n8131 ^ x44;
  assign n8122 = n7860 ^ n7778;
  assign n8123 = n7861 & n8122;
  assign n8124 = n8123 ^ n7778;
  assign n8133 = n8132 ^ n8124;
  assign n8110 = ~n594 & n6326;
  assign n8111 = x72 & n6331;
  assign n8112 = x71 & n6565;
  assign n8113 = ~n8111 & ~n8112;
  assign n8114 = x73 & n6569;
  assign n8115 = n8113 & ~n8114;
  assign n8116 = ~n8110 & n8115;
  assign n8117 = n8116 ^ x50;
  assign n8107 = n7856 ^ n7808;
  assign n8108 = n7857 & n8107;
  assign n8109 = n8108 ^ n7808;
  assign n8118 = n8117 ^ n8109;
  assign n8097 = n416 & n7076;
  assign n8098 = x68 & n7317;
  assign n8099 = x69 & n7080;
  assign n8100 = ~n8098 & ~n8099;
  assign n8101 = x70 & n7319;
  assign n8102 = n8100 & ~n8101;
  assign n8103 = ~n8097 & n8102;
  assign n8104 = n8103 ^ x53;
  assign n8094 = n7854 ^ n7819;
  assign n8095 = ~n7855 & ~n8094;
  assign n8096 = n8095 ^ n7819;
  assign n8105 = n8104 ^ n8096;
  assign n8071 = n7845 ^ x57;
  assign n8072 = x56 & ~n7827;
  assign n8073 = x64 & n8072;
  assign n8074 = n8071 & n8073;
  assign n8075 = x57 ^ x56;
  assign n8076 = ~n8072 & ~n8075;
  assign n8077 = ~n8074 & ~n8076;
  assign n8078 = n162 & n7829;
  assign n8079 = n8078 ^ x67;
  assign n8080 = n7313 & n8079;
  assign n8081 = x65 & n7839;
  assign n8082 = x66 & n7834;
  assign n8083 = ~n8081 & ~n8082;
  assign n8084 = ~n8080 & n8083;
  assign n8085 = n8084 ^ x56;
  assign n8086 = n7845 & n8072;
  assign n8087 = ~x64 & ~n8086;
  assign n8088 = ~n8085 & ~n8087;
  assign n8089 = n8077 & n8088;
  assign n8090 = x64 & n8075;
  assign n8091 = ~n8086 & ~n8090;
  assign n8092 = n8085 & n8091;
  assign n8093 = ~n8089 & ~n8092;
  assign n8106 = n8105 ^ n8093;
  assign n8119 = n8118 ^ n8106;
  assign n8063 = n799 & n5656;
  assign n8064 = x74 & n5895;
  assign n8065 = x76 & n6111;
  assign n8066 = ~n8064 & ~n8065;
  assign n8067 = x75 & n5662;
  assign n8068 = n8066 & ~n8067;
  assign n8069 = ~n8063 & n8068;
  assign n8070 = n8069 ^ x47;
  assign n8120 = n8119 ^ n8070;
  assign n8060 = n7858 ^ n7797;
  assign n8061 = ~n7859 & ~n8060;
  assign n8062 = n8061 ^ n7797;
  assign n8121 = n8120 ^ n8062;
  assign n8134 = n8133 ^ n8121;
  assign n8052 = n1345 & n4415;
  assign n8053 = x80 & n4420;
  assign n8054 = x81 & n4410;
  assign n8055 = ~n8053 & ~n8054;
  assign n8056 = x82 & n4614;
  assign n8057 = n8055 & ~n8056;
  assign n8058 = ~n8052 & n8057;
  assign n8059 = n8058 ^ x41;
  assign n8135 = n8134 ^ n8059;
  assign n8049 = n7786 ^ n7775;
  assign n8050 = ~n7863 & ~n8049;
  assign n8051 = n8050 ^ n7775;
  assign n8136 = n8135 ^ n8051;
  assign n8041 = n1674 & n3829;
  assign n8042 = x83 & n4049;
  assign n8043 = x85 & n4052;
  assign n8044 = ~n8042 & ~n8043;
  assign n8045 = x84 & n3833;
  assign n8046 = n8044 & ~n8045;
  assign n8047 = ~n8041 & n8046;
  assign n8048 = n8047 ^ x38;
  assign n8137 = n8136 ^ n8048;
  assign n8038 = n7864 ^ n7764;
  assign n8039 = n7865 & n8038;
  assign n8040 = n8039 ^ n7764;
  assign n8138 = n8137 ^ n8040;
  assign n8030 = n2040 & n3330;
  assign n8031 = x86 & n3500;
  assign n8032 = x87 & n3334;
  assign n8033 = ~n8031 & ~n8032;
  assign n8034 = x88 & n3502;
  assign n8035 = n8033 & ~n8034;
  assign n8036 = ~n8030 & n8035;
  assign n8037 = n8036 ^ x35;
  assign n8139 = n8138 ^ n8037;
  assign n8027 = n7866 ^ n7753;
  assign n8028 = ~n7867 & ~n8027;
  assign n8029 = n8028 ^ n7753;
  assign n8140 = n8139 ^ n8029;
  assign n8019 = n2447 & n2836;
  assign n8020 = x89 & n2996;
  assign n8021 = x90 & n2840;
  assign n8022 = ~n8020 & ~n8021;
  assign n8023 = x91 & n2998;
  assign n8024 = n8022 & ~n8023;
  assign n8025 = ~n8019 & n8024;
  assign n8026 = n8025 ^ x32;
  assign n8141 = n8140 ^ n8026;
  assign n8016 = n7868 ^ n7742;
  assign n8017 = n7869 & ~n8016;
  assign n8018 = n8017 ^ n7742;
  assign n8142 = n8141 ^ n8018;
  assign n8008 = n2371 & n2895;
  assign n8009 = x92 & n2528;
  assign n8010 = x93 & n2377;
  assign n8011 = ~n8009 & ~n8010;
  assign n8012 = x94 & n2531;
  assign n8013 = n8011 & ~n8012;
  assign n8014 = ~n8008 & n8013;
  assign n8015 = n8014 ^ x29;
  assign n8143 = n8142 ^ n8015;
  assign n8005 = n7870 ^ n7731;
  assign n8006 = n7871 & n8005;
  assign n8007 = n8006 ^ n7731;
  assign n8144 = n8143 ^ n8007;
  assign n7997 = n1969 & n3388;
  assign n7998 = x95 & n1978;
  assign n7999 = x97 & n2108;
  assign n8000 = ~n7998 & ~n7999;
  assign n8001 = x96 & n1973;
  assign n8002 = n8000 & ~n8001;
  assign n8003 = ~n7997 & n8002;
  assign n8004 = n8003 ^ x26;
  assign n8145 = n8144 ^ n8004;
  assign n7994 = n7872 ^ n7720;
  assign n7995 = ~n7873 & ~n7994;
  assign n7996 = n7995 ^ n7720;
  assign n8146 = n8145 ^ n7996;
  assign n7986 = n1624 & n3925;
  assign n7987 = x98 & n1742;
  assign n7988 = x99 & n1628;
  assign n7989 = ~n7987 & ~n7988;
  assign n7990 = x100 & n1744;
  assign n7991 = n7989 & ~n7990;
  assign n7992 = ~n7986 & n7991;
  assign n7993 = n7992 ^ x23;
  assign n8147 = n8146 ^ n7993;
  assign n7983 = n7874 ^ n7709;
  assign n7984 = n7875 & n7983;
  assign n7985 = n7984 ^ n7709;
  assign n8148 = n8147 ^ n7985;
  assign n7975 = n1296 & n4481;
  assign n7976 = x101 & n1403;
  assign n7977 = x103 & n1406;
  assign n7978 = ~n7976 & ~n7977;
  assign n7979 = x102 & n1300;
  assign n7980 = n7978 & ~n7979;
  assign n7981 = ~n7975 & n7980;
  assign n7982 = n7981 ^ x20;
  assign n8149 = n8148 ^ n7982;
  assign n7972 = n7876 ^ n7698;
  assign n7973 = ~n7877 & ~n7972;
  assign n7974 = n7973 ^ n7698;
  assign n8150 = n8149 ^ n7974;
  assign n7964 = n1008 & n5088;
  assign n7965 = x104 & n1101;
  assign n7966 = x105 & n1012;
  assign n7967 = ~n7965 & ~n7966;
  assign n7968 = x106 & n1104;
  assign n7969 = n7967 & ~n7968;
  assign n7970 = ~n7964 & n7969;
  assign n7971 = n7970 ^ x17;
  assign n8151 = n8150 ^ n7971;
  assign n7961 = n7878 ^ n7687;
  assign n7962 = n7879 & n7961;
  assign n7963 = n7962 ^ n7687;
  assign n8152 = n8151 ^ n7963;
  assign n7953 = n752 & ~n5737;
  assign n7954 = x107 & n825;
  assign n7955 = x108 & n757;
  assign n7956 = ~n7954 & ~n7955;
  assign n7957 = x109 & n828;
  assign n7958 = n7956 & ~n7957;
  assign n7959 = ~n7953 & n7958;
  assign n7960 = n7959 ^ x14;
  assign n8153 = n8152 ^ n7960;
  assign n7950 = n7880 ^ n7676;
  assign n7951 = ~n7881 & ~n7950;
  assign n7952 = n7951 ^ n7676;
  assign n8154 = n8153 ^ n7952;
  assign n7942 = n541 & n6420;
  assign n7943 = x110 & n612;
  assign n7944 = x112 & n615;
  assign n7945 = ~n7943 & ~n7944;
  assign n7946 = x111 & n547;
  assign n7947 = n7945 & ~n7946;
  assign n7948 = ~n7942 & n7947;
  assign n7949 = n7948 ^ x11;
  assign n8155 = n8154 ^ n7949;
  assign n7939 = n7882 ^ n7665;
  assign n7940 = n7883 & n7939;
  assign n7941 = n7940 ^ n7665;
  assign n8156 = n8155 ^ n7941;
  assign n7931 = n372 & n7150;
  assign n7932 = x113 & n433;
  assign n7933 = x114 & n376;
  assign n7934 = ~n7932 & ~n7933;
  assign n7935 = x115 & n428;
  assign n7936 = n7934 & ~n7935;
  assign n7937 = ~n7931 & n7936;
  assign n7938 = n7937 ^ x8;
  assign n8157 = n8156 ^ n7938;
  assign n7928 = n7884 ^ n7654;
  assign n7929 = ~n7885 & ~n7928;
  assign n7930 = n7929 ^ n7654;
  assign n8158 = n8157 ^ n7930;
  assign n7894 = ~n6876 & ~n7135;
  assign n7919 = n7894 ^ n7378;
  assign n7920 = n210 & n7919;
  assign n7921 = x116 & n219;
  assign n7922 = x118 & n259;
  assign n7923 = ~n7921 & ~n7922;
  assign n7924 = x117 & n214;
  assign n7925 = n7923 & ~n7924;
  assign n7926 = ~n7920 & n7925;
  assign n7927 = n7926 ^ x5;
  assign n8159 = n8158 ^ n7927;
  assign n7916 = n7886 ^ n7642;
  assign n7917 = n7887 & ~n7916;
  assign n7918 = n7917 ^ n7642;
  assign n8160 = n8159 ^ n7918;
  assign n7895 = ~x118 & ~x120;
  assign n7896 = ~x117 & ~x119;
  assign n7897 = ~n7895 & ~n7896;
  assign n7898 = ~n7894 & ~n7897;
  assign n7899 = ~x117 & n7895;
  assign n7900 = ~x119 & x120;
  assign n7901 = x118 & n7900;
  assign n7902 = n7901 ^ x119;
  assign n7903 = ~n7899 & n7902;
  assign n7904 = ~n7898 & n7903;
  assign n7905 = n7904 ^ x120;
  assign n7906 = n163 & ~n7905;
  assign n7907 = n7906 ^ x1;
  assign n7908 = n7907 ^ x121;
  assign n7909 = x0 & ~n7908;
  assign n7910 = ~x119 & n156;
  assign n7911 = ~x0 & ~n7910;
  assign n7912 = x120 ^ x2;
  assign n7913 = x1 & n7912;
  assign n7914 = n7911 & ~n7913;
  assign n7915 = ~n7909 & ~n7914;
  assign n8161 = n8160 ^ n7915;
  assign n7891 = n7888 ^ n7624;
  assign n7892 = ~n7889 & n7891;
  assign n7893 = n7892 ^ n7624;
  assign n8162 = n8161 ^ n7893;
  assign n8386 = ~n8085 & ~n8091;
  assign n8379 = x65 ^ x57;
  assign n8380 = n8075 & ~n8379;
  assign n8381 = n8380 ^ x56;
  assign n8382 = n8381 ^ x58;
  assign n8383 = x64 & n8382;
  assign n8384 = n149 & n8075;
  assign n8385 = ~n8383 & ~n8384;
  assign n8387 = n8386 ^ n8385;
  assign n8370 = n300 & n7830;
  assign n8371 = x67 & n7834;
  assign n8372 = x66 & n7839;
  assign n8373 = ~n8371 & ~n8372;
  assign n8374 = n7313 & ~n7829;
  assign n8375 = x68 & n8374;
  assign n8376 = n8373 & ~n8375;
  assign n8377 = ~n8370 & n8376;
  assign n8378 = n8377 ^ x56;
  assign n8388 = n8387 ^ n8378;
  assign n8362 = n467 & n7076;
  assign n8363 = x70 & n7080;
  assign n8364 = x69 & n7317;
  assign n8365 = ~n8363 & ~n8364;
  assign n8366 = x71 & n7319;
  assign n8367 = n8365 & ~n8366;
  assign n8368 = ~n8362 & n8367;
  assign n8369 = n8368 ^ x53;
  assign n8389 = n8388 ^ n8369;
  assign n8359 = n8104 ^ n8093;
  assign n8360 = ~n8105 & n8359;
  assign n8361 = n8360 ^ n8096;
  assign n8390 = n8389 ^ n8361;
  assign n8351 = ~n656 & n6326;
  assign n8352 = x73 & n6331;
  assign n8353 = x72 & n6565;
  assign n8354 = ~n8352 & ~n8353;
  assign n8355 = x74 & n6569;
  assign n8356 = n8354 & ~n8355;
  assign n8357 = ~n8351 & n8356;
  assign n8358 = n8357 ^ x50;
  assign n8391 = n8390 ^ n8358;
  assign n8348 = n8117 ^ n8106;
  assign n8349 = ~n8118 & ~n8348;
  assign n8350 = n8349 ^ n8109;
  assign n8392 = n8391 ^ n8350;
  assign n8340 = n877 & n5656;
  assign n8341 = x75 & n5895;
  assign n8342 = x76 & n5662;
  assign n8343 = ~n8341 & ~n8342;
  assign n8344 = x77 & n6111;
  assign n8345 = n8343 & ~n8344;
  assign n8346 = ~n8340 & n8345;
  assign n8347 = n8346 ^ x47;
  assign n8393 = n8392 ^ n8347;
  assign n8337 = n8119 ^ n8062;
  assign n8338 = n8120 & n8337;
  assign n8339 = n8338 ^ n8062;
  assign n8394 = n8393 ^ n8339;
  assign n8329 = ~n1141 & n5010;
  assign n8330 = x79 & n5014;
  assign n8331 = x80 & n5226;
  assign n8332 = ~n8330 & ~n8331;
  assign n8333 = x78 & n5223;
  assign n8334 = n8332 & ~n8333;
  assign n8335 = ~n8329 & n8334;
  assign n8336 = n8335 ^ x44;
  assign n8395 = n8394 ^ n8336;
  assign n8326 = n8132 ^ n8121;
  assign n8327 = ~n8133 & ~n8326;
  assign n8328 = n8327 ^ n8124;
  assign n8396 = n8395 ^ n8328;
  assign n8318 = n1445 & n4415;
  assign n8319 = x81 & n4420;
  assign n8320 = x82 & n4410;
  assign n8321 = ~n8319 & ~n8320;
  assign n8322 = x83 & n4614;
  assign n8323 = n8321 & ~n8322;
  assign n8324 = ~n8318 & n8323;
  assign n8325 = n8324 ^ x41;
  assign n8397 = n8396 ^ n8325;
  assign n8315 = n8134 ^ n8051;
  assign n8316 = n8135 & n8315;
  assign n8317 = n8316 ^ n8051;
  assign n8398 = n8397 ^ n8317;
  assign n8307 = n1787 & n3829;
  assign n8308 = x84 & n4049;
  assign n8309 = x86 & n4052;
  assign n8310 = ~n8308 & ~n8309;
  assign n8311 = x85 & n3833;
  assign n8312 = n8310 & ~n8311;
  assign n8313 = ~n8307 & n8312;
  assign n8314 = n8313 ^ x38;
  assign n8399 = n8398 ^ n8314;
  assign n8304 = n8136 ^ n8040;
  assign n8305 = ~n8137 & ~n8304;
  assign n8306 = n8305 ^ n8040;
  assign n8400 = n8399 ^ n8306;
  assign n8296 = n2164 & n3330;
  assign n8297 = x87 & n3500;
  assign n8298 = x89 & n3502;
  assign n8299 = ~n8297 & ~n8298;
  assign n8300 = x88 & n3334;
  assign n8301 = n8299 & ~n8300;
  assign n8302 = ~n8296 & n8301;
  assign n8303 = n8302 ^ x35;
  assign n8401 = n8400 ^ n8303;
  assign n8293 = n8138 ^ n8029;
  assign n8294 = n8139 & n8293;
  assign n8295 = n8294 ^ n8029;
  assign n8402 = n8401 ^ n8295;
  assign n8285 = n2585 & n2836;
  assign n8286 = x91 & n2840;
  assign n8287 = x90 & n2996;
  assign n8288 = ~n8286 & ~n8287;
  assign n8289 = x92 & n2998;
  assign n8290 = n8288 & ~n8289;
  assign n8291 = ~n8285 & n8290;
  assign n8292 = n8291 ^ x32;
  assign n8403 = n8402 ^ n8292;
  assign n8282 = n8140 ^ n8018;
  assign n8283 = ~n8141 & n8282;
  assign n8284 = n8283 ^ n8018;
  assign n8404 = n8403 ^ n8284;
  assign n8274 = n2371 & n3054;
  assign n8275 = x93 & n2528;
  assign n8276 = x94 & n2377;
  assign n8277 = ~n8275 & ~n8276;
  assign n8278 = x95 & n2531;
  assign n8279 = n8277 & ~n8278;
  assign n8280 = ~n8274 & n8279;
  assign n8281 = n8280 ^ x29;
  assign n8405 = n8404 ^ n8281;
  assign n8271 = n8142 ^ n8007;
  assign n8272 = ~n8143 & ~n8271;
  assign n8273 = n8272 ^ n8007;
  assign n8406 = n8405 ^ n8273;
  assign n8263 = n1969 & n3556;
  assign n8264 = x96 & n1978;
  assign n8265 = x97 & n1973;
  assign n8266 = ~n8264 & ~n8265;
  assign n8267 = x98 & n2108;
  assign n8268 = n8266 & ~n8267;
  assign n8269 = ~n8263 & n8268;
  assign n8270 = n8269 ^ x26;
  assign n8407 = n8406 ^ n8270;
  assign n8260 = n8144 ^ n7996;
  assign n8261 = n8145 & n8260;
  assign n8262 = n8261 ^ n7996;
  assign n8408 = n8407 ^ n8262;
  assign n8252 = n1624 & n4105;
  assign n8253 = x100 & n1628;
  assign n8254 = x99 & n1742;
  assign n8255 = ~n8253 & ~n8254;
  assign n8256 = x101 & n1744;
  assign n8257 = n8255 & ~n8256;
  assign n8258 = ~n8252 & n8257;
  assign n8259 = n8258 ^ x23;
  assign n8409 = n8408 ^ n8259;
  assign n8249 = n8146 ^ n7985;
  assign n8250 = ~n8147 & ~n8249;
  assign n8251 = n8250 ^ n7985;
  assign n8410 = n8409 ^ n8251;
  assign n8241 = n1296 & n4670;
  assign n8242 = x102 & n1403;
  assign n8243 = x103 & n1300;
  assign n8244 = ~n8242 & ~n8243;
  assign n8245 = x104 & n1406;
  assign n8246 = n8244 & ~n8245;
  assign n8247 = ~n8241 & n8246;
  assign n8248 = n8247 ^ x20;
  assign n8411 = n8410 ^ n8248;
  assign n8238 = n8148 ^ n7974;
  assign n8239 = n8149 & n8238;
  assign n8240 = n8239 ^ n7974;
  assign n8412 = n8411 ^ n8240;
  assign n8230 = n1008 & n5297;
  assign n8231 = x105 & n1101;
  assign n8232 = x106 & n1012;
  assign n8233 = ~n8231 & ~n8232;
  assign n8234 = x107 & n1104;
  assign n8235 = n8233 & ~n8234;
  assign n8236 = ~n8230 & n8235;
  assign n8237 = n8236 ^ x17;
  assign n8413 = n8412 ^ n8237;
  assign n8227 = n8150 ^ n7963;
  assign n8228 = ~n8151 & ~n8227;
  assign n8229 = n8228 ^ n7963;
  assign n8414 = n8413 ^ n8229;
  assign n8219 = n752 & n5955;
  assign n8220 = x108 & n825;
  assign n8221 = x109 & n757;
  assign n8222 = ~n8220 & ~n8221;
  assign n8223 = x110 & n828;
  assign n8224 = n8222 & ~n8223;
  assign n8225 = ~n8219 & n8224;
  assign n8226 = n8225 ^ x14;
  assign n8415 = n8414 ^ n8226;
  assign n8216 = n8152 ^ n7952;
  assign n8217 = n8153 & n8216;
  assign n8218 = n8217 ^ n7952;
  assign n8416 = n8415 ^ n8218;
  assign n8208 = n541 & n6656;
  assign n8209 = x111 & n612;
  assign n8210 = x112 & n547;
  assign n8211 = ~n8209 & ~n8210;
  assign n8212 = x113 & n615;
  assign n8213 = n8211 & ~n8212;
  assign n8214 = ~n8208 & n8213;
  assign n8215 = n8214 ^ x11;
  assign n8417 = n8416 ^ n8215;
  assign n8205 = n8154 ^ n7941;
  assign n8206 = ~n8155 & ~n8205;
  assign n8207 = n8206 ^ n7941;
  assign n8418 = n8417 ^ n8207;
  assign n8197 = n372 & n7393;
  assign n8198 = x114 & n433;
  assign n8199 = x115 & n376;
  assign n8200 = ~n8198 & ~n8199;
  assign n8201 = x116 & n428;
  assign n8202 = n8200 & ~n8201;
  assign n8203 = ~n8197 & n8202;
  assign n8204 = n8203 ^ x8;
  assign n8419 = n8418 ^ n8204;
  assign n8194 = n8156 ^ n7930;
  assign n8195 = n8157 & n8194;
  assign n8196 = n8195 ^ n7930;
  assign n8420 = n8419 ^ n8196;
  assign n8178 = x120 & n7904;
  assign n8179 = ~x121 & ~n8178;
  assign n8180 = ~x120 & ~n7904;
  assign n8181 = x121 & ~n8180;
  assign n8182 = ~n8179 & ~n8181;
  assign n8183 = n163 & ~n8182;
  assign n8184 = n8183 ^ x1;
  assign n8185 = n8184 ^ x122;
  assign n8186 = x0 & ~n8185;
  assign n8187 = x121 ^ x2;
  assign n8188 = x1 & n8187;
  assign n8189 = ~x0 & ~n8188;
  assign n8190 = ~x120 & n156;
  assign n8191 = n8189 & ~n8190;
  assign n8192 = ~n8186 & ~n8191;
  assign n8169 = n7379 ^ x119;
  assign n8170 = n210 & n8169;
  assign n8171 = x117 & n219;
  assign n8172 = x119 & n259;
  assign n8173 = ~n8171 & ~n8172;
  assign n8174 = x118 & n214;
  assign n8175 = n8173 & ~n8174;
  assign n8176 = ~n8170 & n8175;
  assign n8177 = n8176 ^ x5;
  assign n8193 = n8192 ^ n8177;
  assign n8421 = n8420 ^ n8193;
  assign n8166 = n8158 ^ n7918;
  assign n8167 = ~n8159 & n8166;
  assign n8168 = n8167 ^ n7918;
  assign n8422 = n8421 ^ n8168;
  assign n8163 = n8160 ^ n7893;
  assign n8164 = n8161 & ~n8163;
  assign n8165 = n8164 ^ n7893;
  assign n8423 = n8422 ^ n8165;
  assign n8696 = n8420 ^ n8192;
  assign n8697 = n8193 & ~n8696;
  assign n8698 = n8697 ^ n8420;
  assign n8699 = n8168 & n8698;
  assign n8700 = n8177 & ~n8192;
  assign n8701 = n8420 & n8700;
  assign n8702 = ~n8699 & ~n8701;
  assign n8703 = ~n8165 & ~n8702;
  assign n8704 = ~n8177 & n8192;
  assign n8705 = ~n8420 & n8704;
  assign n8706 = ~n8168 & n8705;
  assign n8707 = n8168 & n8701;
  assign n8708 = ~n8706 & ~n8707;
  assign n8709 = ~n8703 & n8708;
  assign n8710 = n8168 & ~n8705;
  assign n8711 = ~n8698 & ~n8710;
  assign n8712 = n8165 & n8711;
  assign n8713 = n8709 & ~n8712;
  assign n8659 = n953 & n5656;
  assign n8660 = x77 & n5662;
  assign n8661 = x76 & n5895;
  assign n8662 = ~n8660 & ~n8661;
  assign n8663 = x78 & n6111;
  assign n8664 = n8662 & ~n8663;
  assign n8665 = ~n8659 & n8664;
  assign n8666 = n8665 ^ x47;
  assign n8656 = n8392 ^ n8339;
  assign n8657 = n8393 & n8656;
  assign n8658 = n8657 ^ n8339;
  assign n8667 = n8666 ^ n8658;
  assign n8646 = n720 & n6326;
  assign n8647 = x73 & n6565;
  assign n8648 = x75 & n6569;
  assign n8649 = ~n8647 & ~n8648;
  assign n8650 = x74 & n6331;
  assign n8651 = n8649 & ~n8650;
  assign n8652 = ~n8646 & n8651;
  assign n8653 = n8652 ^ x50;
  assign n8643 = n8390 ^ n8350;
  assign n8644 = ~n8391 & ~n8643;
  assign n8645 = n8644 ^ n8350;
  assign n8654 = n8653 ^ n8645;
  assign n8621 = x59 ^ x58;
  assign n8622 = n8075 & n8621;
  assign n8623 = n208 & n8622;
  assign n8616 = x56 & x57;
  assign n8612 = ~x56 & ~x57;
  assign n8624 = n8616 ^ n8612;
  assign n8625 = x58 & n8624;
  assign n8626 = n8625 ^ n8616;
  assign n8627 = ~n8623 & ~n8626;
  assign n8628 = x65 & ~n8627;
  assign n8629 = x58 ^ x57;
  assign n8630 = n8621 & ~n8629;
  assign n8631 = ~n8075 & n8630;
  assign n8632 = x64 & n8631;
  assign n8633 = n149 & n8621;
  assign n8634 = x66 & n8075;
  assign n8635 = ~n8633 & n8634;
  assign n8636 = ~n8632 & ~n8635;
  assign n8637 = ~n8628 & n8636;
  assign n8613 = x58 & x64;
  assign n8614 = n8612 & ~n8613;
  assign n8615 = ~n201 & ~n8614;
  assign n8617 = ~x58 & x64;
  assign n8618 = n8616 & ~n8617;
  assign n8619 = n8615 & ~n8618;
  assign n8620 = x59 & n8619;
  assign n8638 = n8637 ^ n8620;
  assign n8609 = n8385 ^ n8378;
  assign n8610 = ~n8387 & ~n8609;
  assign n8611 = n8610 ^ n8386;
  assign n8639 = n8638 ^ n8611;
  assign n8601 = n358 & n7830;
  assign n8602 = x68 & n7834;
  assign n8603 = x67 & n7839;
  assign n8604 = ~n8602 & ~n8603;
  assign n8605 = x69 & n8374;
  assign n8606 = n8604 & ~n8605;
  assign n8607 = ~n8601 & n8606;
  assign n8608 = n8607 ^ x56;
  assign n8640 = n8639 ^ n8608;
  assign n8593 = n520 & n7076;
  assign n8594 = x70 & n7317;
  assign n8595 = x72 & n7319;
  assign n8596 = ~n8594 & ~n8595;
  assign n8597 = x71 & n7080;
  assign n8598 = n8596 & ~n8597;
  assign n8599 = ~n8593 & n8598;
  assign n8600 = n8599 ^ x53;
  assign n8641 = n8640 ^ n8600;
  assign n8590 = n8388 ^ n8361;
  assign n8591 = n8389 & n8590;
  assign n8592 = n8591 ^ n8361;
  assign n8642 = n8641 ^ n8592;
  assign n8655 = n8654 ^ n8642;
  assign n8668 = n8667 ^ n8655;
  assign n8582 = n1230 & n5010;
  assign n8583 = x79 & n5223;
  assign n8584 = x80 & n5014;
  assign n8585 = ~n8583 & ~n8584;
  assign n8586 = x81 & n5226;
  assign n8587 = n8585 & ~n8586;
  assign n8588 = ~n8582 & n8587;
  assign n8589 = n8588 ^ x44;
  assign n8669 = n8668 ^ n8589;
  assign n8579 = n8394 ^ n8328;
  assign n8580 = ~n8395 & ~n8579;
  assign n8581 = n8580 ^ n8328;
  assign n8670 = n8669 ^ n8581;
  assign n8571 = n1547 & n4415;
  assign n8572 = x82 & n4420;
  assign n8573 = x83 & n4410;
  assign n8574 = ~n8572 & ~n8573;
  assign n8575 = x84 & n4614;
  assign n8576 = n8574 & ~n8575;
  assign n8577 = ~n8571 & n8576;
  assign n8578 = n8577 ^ x41;
  assign n8671 = n8670 ^ n8578;
  assign n8568 = n8396 ^ n8317;
  assign n8569 = n8397 & n8568;
  assign n8570 = n8569 ^ n8317;
  assign n8672 = n8671 ^ n8570;
  assign n8560 = n1903 & n3829;
  assign n8561 = x85 & n4049;
  assign n8562 = x86 & n3833;
  assign n8563 = ~n8561 & ~n8562;
  assign n8564 = x87 & n4052;
  assign n8565 = n8563 & ~n8564;
  assign n8566 = ~n8560 & n8565;
  assign n8567 = n8566 ^ x38;
  assign n8673 = n8672 ^ n8567;
  assign n8557 = n8398 ^ n8306;
  assign n8558 = ~n8399 & ~n8557;
  assign n8559 = n8558 ^ n8306;
  assign n8674 = n8673 ^ n8559;
  assign n8549 = n2292 & n3330;
  assign n8550 = x88 & n3500;
  assign n8551 = x90 & n3502;
  assign n8552 = ~n8550 & ~n8551;
  assign n8553 = x89 & n3334;
  assign n8554 = n8552 & ~n8553;
  assign n8555 = ~n8549 & n8554;
  assign n8556 = n8555 ^ x35;
  assign n8675 = n8674 ^ n8556;
  assign n8546 = n8400 ^ n8295;
  assign n8547 = n8401 & n8546;
  assign n8548 = n8547 ^ n8295;
  assign n8676 = n8675 ^ n8548;
  assign n8538 = n2726 & n2836;
  assign n8539 = x92 & n2840;
  assign n8540 = x91 & n2996;
  assign n8541 = ~n8539 & ~n8540;
  assign n8542 = x93 & n2998;
  assign n8543 = n8541 & ~n8542;
  assign n8544 = ~n8538 & n8543;
  assign n8545 = n8544 ^ x32;
  assign n8677 = n8676 ^ n8545;
  assign n8535 = n8402 ^ n8284;
  assign n8536 = ~n8403 & n8535;
  assign n8537 = n8536 ^ n8284;
  assign n8678 = n8677 ^ n8537;
  assign n8527 = n2371 & n3209;
  assign n8528 = x94 & n2528;
  assign n8529 = x95 & n2377;
  assign n8530 = ~n8528 & ~n8529;
  assign n8531 = x96 & n2531;
  assign n8532 = n8530 & ~n8531;
  assign n8533 = ~n8527 & n8532;
  assign n8534 = n8533 ^ x29;
  assign n8679 = n8678 ^ n8534;
  assign n8524 = n8281 ^ n8273;
  assign n8525 = n8405 & n8524;
  assign n8526 = n8525 ^ n8404;
  assign n8680 = n8679 ^ n8526;
  assign n8516 = n1969 & n3730;
  assign n8517 = x97 & n1978;
  assign n8518 = x99 & n2108;
  assign n8519 = ~n8517 & ~n8518;
  assign n8520 = x98 & n1973;
  assign n8521 = n8519 & ~n8520;
  assign n8522 = ~n8516 & n8521;
  assign n8523 = n8522 ^ x26;
  assign n8681 = n8680 ^ n8523;
  assign n8513 = n8406 ^ n8262;
  assign n8514 = n8407 & n8513;
  assign n8515 = n8514 ^ n8262;
  assign n8682 = n8681 ^ n8515;
  assign n8505 = n1624 & n4286;
  assign n8506 = x100 & n1742;
  assign n8507 = x101 & n1628;
  assign n8508 = ~n8506 & ~n8507;
  assign n8509 = x102 & n1744;
  assign n8510 = n8508 & ~n8509;
  assign n8511 = ~n8505 & n8510;
  assign n8512 = n8511 ^ x23;
  assign n8683 = n8682 ^ n8512;
  assign n8502 = n8408 ^ n8251;
  assign n8503 = ~n8409 & ~n8502;
  assign n8504 = n8503 ^ n8251;
  assign n8684 = n8683 ^ n8504;
  assign n8494 = n1296 & n4867;
  assign n8495 = x104 & n1300;
  assign n8496 = x103 & n1403;
  assign n8497 = ~n8495 & ~n8496;
  assign n8498 = x105 & n1406;
  assign n8499 = n8497 & ~n8498;
  assign n8500 = ~n8494 & n8499;
  assign n8501 = n8500 ^ x20;
  assign n8685 = n8684 ^ n8501;
  assign n8491 = n8410 ^ n8240;
  assign n8492 = n8411 & n8491;
  assign n8493 = n8492 ^ n8240;
  assign n8686 = n8685 ^ n8493;
  assign n8483 = n1008 & ~n5506;
  assign n8484 = x106 & n1101;
  assign n8485 = x107 & n1012;
  assign n8486 = ~n8484 & ~n8485;
  assign n8487 = x108 & n1104;
  assign n8488 = n8486 & ~n8487;
  assign n8489 = ~n8483 & n8488;
  assign n8490 = n8489 ^ x17;
  assign n8687 = n8686 ^ n8490;
  assign n8480 = n8412 ^ n8229;
  assign n8481 = ~n8413 & ~n8480;
  assign n8482 = n8481 ^ n8229;
  assign n8688 = n8687 ^ n8482;
  assign n8472 = n752 & n6178;
  assign n8473 = x109 & n825;
  assign n8474 = x111 & n828;
  assign n8475 = ~n8473 & ~n8474;
  assign n8476 = x110 & n757;
  assign n8477 = n8475 & ~n8476;
  assign n8478 = ~n8472 & n8477;
  assign n8479 = n8478 ^ x14;
  assign n8689 = n8688 ^ n8479;
  assign n8469 = n8414 ^ n8218;
  assign n8470 = n8415 & n8469;
  assign n8471 = n8470 ^ n8218;
  assign n8690 = n8689 ^ n8471;
  assign n8461 = n541 & n6892;
  assign n8462 = x112 & n612;
  assign n8463 = x114 & n615;
  assign n8464 = ~n8462 & ~n8463;
  assign n8465 = x113 & n547;
  assign n8466 = n8464 & ~n8465;
  assign n8467 = ~n8461 & n8466;
  assign n8468 = n8467 ^ x11;
  assign n8691 = n8690 ^ n8468;
  assign n8458 = n8416 ^ n8207;
  assign n8459 = ~n8417 & ~n8458;
  assign n8460 = n8459 ^ n8207;
  assign n8692 = n8691 ^ n8460;
  assign n8450 = n372 & n7643;
  assign n8451 = x115 & n433;
  assign n8452 = x116 & n376;
  assign n8453 = ~n8451 & ~n8452;
  assign n8454 = x117 & n428;
  assign n8455 = n8453 & ~n8454;
  assign n8456 = ~n8450 & n8455;
  assign n8457 = n8456 ^ x8;
  assign n8693 = n8692 ^ n8457;
  assign n8447 = n8418 ^ n8196;
  assign n8448 = n8419 & n8447;
  assign n8449 = n8448 ^ n8196;
  assign n8694 = n8693 ^ n8449;
  assign n8433 = ~x122 & ~n8181;
  assign n8434 = x122 & ~n8179;
  assign n8435 = ~n8433 & ~n8434;
  assign n8436 = n163 & ~n8435;
  assign n8437 = n8436 ^ x1;
  assign n8438 = n8437 ^ x123;
  assign n8439 = x0 & ~n8438;
  assign n8440 = ~x121 & n156;
  assign n8441 = ~x0 & ~n8440;
  assign n8442 = x122 ^ x2;
  assign n8443 = x1 & n8442;
  assign n8444 = n8441 & ~n8443;
  assign n8445 = ~n8439 & ~n8444;
  assign n8424 = n7629 ^ x120;
  assign n8425 = n210 & ~n8424;
  assign n8426 = x118 & n219;
  assign n8427 = x119 & n214;
  assign n8428 = ~n8426 & ~n8427;
  assign n8429 = x120 & n259;
  assign n8430 = n8428 & ~n8429;
  assign n8431 = ~n8425 & n8430;
  assign n8432 = n8431 ^ x5;
  assign n8446 = n8445 ^ n8432;
  assign n8695 = n8694 ^ n8446;
  assign n8714 = n8713 ^ n8695;
  assign n8983 = ~n8695 & ~n8707;
  assign n8984 = ~n8711 & ~n8983;
  assign n8985 = n8165 & ~n8984;
  assign n8986 = ~n8695 & n8702;
  assign n8987 = ~n8706 & ~n8986;
  assign n8988 = ~n8985 & n8987;
  assign n8939 = n416 & n7830;
  assign n8940 = x69 & n7834;
  assign n8941 = x68 & n7839;
  assign n8942 = ~n8940 & ~n8941;
  assign n8943 = x70 & n8374;
  assign n8944 = n8942 & ~n8943;
  assign n8945 = ~n8939 & n8944;
  assign n8946 = n8945 ^ x56;
  assign n8927 = x59 & ~n8619;
  assign n8928 = n8637 & n8927;
  assign n8929 = x60 ^ x59;
  assign n8930 = x64 & n8929;
  assign n8931 = ~n8928 & ~n8930;
  assign n8919 = n162 & n8621;
  assign n8920 = n8919 ^ x67;
  assign n8921 = n8075 & n8920;
  assign n8922 = x66 & n8626;
  assign n8923 = x65 & n8631;
  assign n8924 = ~n8922 & ~n8923;
  assign n8925 = ~n8921 & n8924;
  assign n8926 = n8925 ^ x59;
  assign n8932 = n8931 ^ n8926;
  assign n8933 = n8637 ^ x60;
  assign n8934 = x64 & n8927;
  assign n8935 = n8933 & n8934;
  assign n8936 = ~n8926 & n8935;
  assign n8937 = ~n8932 & n8936;
  assign n8938 = n8937 ^ n8932;
  assign n8947 = n8946 ^ n8938;
  assign n8916 = n8638 ^ n8608;
  assign n8917 = ~n8639 & ~n8916;
  assign n8918 = n8917 ^ n8611;
  assign n8948 = n8947 ^ n8918;
  assign n8908 = ~n594 & n7076;
  assign n8909 = x72 & n7080;
  assign n8910 = x71 & n7317;
  assign n8911 = ~n8909 & ~n8910;
  assign n8912 = x73 & n7319;
  assign n8913 = n8911 & ~n8912;
  assign n8914 = ~n8908 & n8913;
  assign n8915 = n8914 ^ x53;
  assign n8949 = n8948 ^ n8915;
  assign n8905 = n8640 ^ n8592;
  assign n8906 = n8641 & n8905;
  assign n8907 = n8906 ^ n8592;
  assign n8950 = n8949 ^ n8907;
  assign n8897 = n799 & n6326;
  assign n8898 = x74 & n6565;
  assign n8899 = x76 & n6569;
  assign n8900 = ~n8898 & ~n8899;
  assign n8901 = x75 & n6331;
  assign n8902 = n8900 & ~n8901;
  assign n8903 = ~n8897 & n8902;
  assign n8904 = n8903 ^ x50;
  assign n8951 = n8950 ^ n8904;
  assign n8894 = n8653 ^ n8642;
  assign n8895 = ~n8654 & ~n8894;
  assign n8896 = n8895 ^ n8645;
  assign n8952 = n8951 ^ n8896;
  assign n8886 = n1054 & n5656;
  assign n8887 = x77 & n5895;
  assign n8888 = x78 & n5662;
  assign n8889 = ~n8887 & ~n8888;
  assign n8890 = x79 & n6111;
  assign n8891 = n8889 & ~n8890;
  assign n8892 = ~n8886 & n8891;
  assign n8893 = n8892 ^ x47;
  assign n8953 = n8952 ^ n8893;
  assign n8883 = n8666 ^ n8655;
  assign n8884 = ~n8667 & n8883;
  assign n8885 = n8884 ^ n8658;
  assign n8954 = n8953 ^ n8885;
  assign n8875 = n1345 & n5010;
  assign n8876 = x80 & n5223;
  assign n8877 = x81 & n5014;
  assign n8878 = ~n8876 & ~n8877;
  assign n8879 = x82 & n5226;
  assign n8880 = n8878 & ~n8879;
  assign n8881 = ~n8875 & n8880;
  assign n8882 = n8881 ^ x44;
  assign n8955 = n8954 ^ n8882;
  assign n8872 = n8668 ^ n8581;
  assign n8873 = ~n8669 & ~n8872;
  assign n8874 = n8873 ^ n8581;
  assign n8956 = n8955 ^ n8874;
  assign n8864 = n1674 & n4415;
  assign n8865 = x83 & n4420;
  assign n8866 = x85 & n4614;
  assign n8867 = ~n8865 & ~n8866;
  assign n8868 = x84 & n4410;
  assign n8869 = n8867 & ~n8868;
  assign n8870 = ~n8864 & n8869;
  assign n8871 = n8870 ^ x41;
  assign n8957 = n8956 ^ n8871;
  assign n8861 = n8670 ^ n8570;
  assign n8862 = n8671 & n8861;
  assign n8863 = n8862 ^ n8570;
  assign n8958 = n8957 ^ n8863;
  assign n8853 = n2040 & n3829;
  assign n8854 = x86 & n4049;
  assign n8855 = x88 & n4052;
  assign n8856 = ~n8854 & ~n8855;
  assign n8857 = x87 & n3833;
  assign n8858 = n8856 & ~n8857;
  assign n8859 = ~n8853 & n8858;
  assign n8860 = n8859 ^ x38;
  assign n8959 = n8958 ^ n8860;
  assign n8850 = n8672 ^ n8559;
  assign n8851 = ~n8673 & ~n8850;
  assign n8852 = n8851 ^ n8559;
  assign n8960 = n8959 ^ n8852;
  assign n8842 = n2447 & n3330;
  assign n8843 = x89 & n3500;
  assign n8844 = x90 & n3334;
  assign n8845 = ~n8843 & ~n8844;
  assign n8846 = x91 & n3502;
  assign n8847 = n8845 & ~n8846;
  assign n8848 = ~n8842 & n8847;
  assign n8849 = n8848 ^ x35;
  assign n8961 = n8960 ^ n8849;
  assign n8839 = n8674 ^ n8548;
  assign n8840 = n8675 & n8839;
  assign n8841 = n8840 ^ n8548;
  assign n8962 = n8961 ^ n8841;
  assign n8831 = n2836 & n2895;
  assign n8832 = x92 & n2996;
  assign n8833 = x93 & n2840;
  assign n8834 = ~n8832 & ~n8833;
  assign n8835 = x94 & n2998;
  assign n8836 = n8834 & ~n8835;
  assign n8837 = ~n8831 & n8836;
  assign n8838 = n8837 ^ x32;
  assign n8963 = n8962 ^ n8838;
  assign n8828 = n8676 ^ n8537;
  assign n8829 = ~n8677 & n8828;
  assign n8830 = n8829 ^ n8537;
  assign n8964 = n8963 ^ n8830;
  assign n8820 = n2371 & n3388;
  assign n8821 = x95 & n2528;
  assign n8822 = x96 & n2377;
  assign n8823 = ~n8821 & ~n8822;
  assign n8824 = x97 & n2531;
  assign n8825 = n8823 & ~n8824;
  assign n8826 = ~n8820 & n8825;
  assign n8827 = n8826 ^ x29;
  assign n8965 = n8964 ^ n8827;
  assign n8817 = n8534 ^ n8526;
  assign n8818 = n8679 & ~n8817;
  assign n8819 = n8818 ^ n8678;
  assign n8966 = n8965 ^ n8819;
  assign n8809 = n1969 & n3925;
  assign n8810 = x98 & n1978;
  assign n8811 = x99 & n1973;
  assign n8812 = ~n8810 & ~n8811;
  assign n8813 = x100 & n2108;
  assign n8814 = n8812 & ~n8813;
  assign n8815 = ~n8809 & n8814;
  assign n8816 = n8815 ^ x26;
  assign n8967 = n8966 ^ n8816;
  assign n8806 = n8680 ^ n8515;
  assign n8807 = ~n8681 & ~n8806;
  assign n8808 = n8807 ^ n8515;
  assign n8968 = n8967 ^ n8808;
  assign n8798 = n1624 & n4481;
  assign n8799 = x101 & n1742;
  assign n8800 = x102 & n1628;
  assign n8801 = ~n8799 & ~n8800;
  assign n8802 = x103 & n1744;
  assign n8803 = n8801 & ~n8802;
  assign n8804 = ~n8798 & n8803;
  assign n8805 = n8804 ^ x23;
  assign n8969 = n8968 ^ n8805;
  assign n8795 = n8682 ^ n8504;
  assign n8796 = n8683 & n8795;
  assign n8797 = n8796 ^ n8504;
  assign n8970 = n8969 ^ n8797;
  assign n8787 = n1296 & n5088;
  assign n8788 = x104 & n1403;
  assign n8789 = x105 & n1300;
  assign n8790 = ~n8788 & ~n8789;
  assign n8791 = x106 & n1406;
  assign n8792 = n8790 & ~n8791;
  assign n8793 = ~n8787 & n8792;
  assign n8794 = n8793 ^ x20;
  assign n8971 = n8970 ^ n8794;
  assign n8784 = n8684 ^ n8493;
  assign n8785 = ~n8685 & ~n8784;
  assign n8786 = n8785 ^ n8493;
  assign n8972 = n8971 ^ n8786;
  assign n8776 = n1008 & ~n5737;
  assign n8777 = x107 & n1101;
  assign n8778 = x108 & n1012;
  assign n8779 = ~n8777 & ~n8778;
  assign n8780 = x109 & n1104;
  assign n8781 = n8779 & ~n8780;
  assign n8782 = ~n8776 & n8781;
  assign n8783 = n8782 ^ x17;
  assign n8973 = n8972 ^ n8783;
  assign n8773 = n8686 ^ n8482;
  assign n8774 = n8687 & n8773;
  assign n8775 = n8774 ^ n8482;
  assign n8974 = n8973 ^ n8775;
  assign n8765 = n752 & n6420;
  assign n8766 = x110 & n825;
  assign n8767 = x111 & n757;
  assign n8768 = ~n8766 & ~n8767;
  assign n8769 = x112 & n828;
  assign n8770 = n8768 & ~n8769;
  assign n8771 = ~n8765 & n8770;
  assign n8772 = n8771 ^ x14;
  assign n8975 = n8974 ^ n8772;
  assign n8762 = n8688 ^ n8471;
  assign n8763 = ~n8689 & ~n8762;
  assign n8764 = n8763 ^ n8471;
  assign n8976 = n8975 ^ n8764;
  assign n8754 = n541 & n7150;
  assign n8755 = x113 & n612;
  assign n8756 = x114 & n547;
  assign n8757 = ~n8755 & ~n8756;
  assign n8758 = x115 & n615;
  assign n8759 = n8757 & ~n8758;
  assign n8760 = ~n8754 & n8759;
  assign n8761 = n8760 ^ x11;
  assign n8977 = n8976 ^ n8761;
  assign n8751 = n8690 ^ n8460;
  assign n8752 = n8691 & n8751;
  assign n8753 = n8752 ^ n8460;
  assign n8978 = n8977 ^ n8753;
  assign n8743 = n372 & n7919;
  assign n8744 = x116 & n433;
  assign n8745 = x117 & n376;
  assign n8746 = ~n8744 & ~n8745;
  assign n8747 = x118 & n428;
  assign n8748 = n8746 & ~n8747;
  assign n8749 = ~n8743 & n8748;
  assign n8750 = n8749 ^ x8;
  assign n8979 = n8978 ^ n8750;
  assign n8740 = n8692 ^ n8449;
  assign n8741 = ~n8693 & ~n8740;
  assign n8742 = n8741 ^ n8449;
  assign n8980 = n8979 ^ n8742;
  assign n8737 = n8694 ^ n8445;
  assign n8738 = n8446 & n8737;
  assign n8739 = n8738 ^ n8694;
  assign n8981 = n8980 ^ n8739;
  assign n8724 = x123 ^ x122;
  assign n8725 = ~n8435 & n8724;
  assign n8726 = n163 & ~n8725;
  assign n8727 = n8726 ^ x1;
  assign n8728 = n8727 ^ x124;
  assign n8729 = x0 & n8728;
  assign n8730 = x122 & n156;
  assign n8731 = ~x0 & ~n8730;
  assign n8732 = x1 & x123;
  assign n8733 = n8732 ^ x2;
  assign n8734 = n8731 & n8733;
  assign n8735 = ~n8729 & ~n8734;
  assign n8715 = n7905 ^ x121;
  assign n8716 = n210 & n8715;
  assign n8717 = x119 & n219;
  assign n8718 = x121 & n259;
  assign n8719 = ~n8717 & ~n8718;
  assign n8720 = x120 & n214;
  assign n8721 = n8719 & ~n8720;
  assign n8722 = ~n8716 & n8721;
  assign n8723 = n8722 ^ x5;
  assign n8736 = n8735 ^ n8723;
  assign n8982 = n8981 ^ n8736;
  assign n8989 = n8988 ^ n8982;
  assign n9256 = n8739 & ~n8980;
  assign n9257 = ~n8723 & ~n8735;
  assign n9258 = n9256 & n9257;
  assign n9259 = ~n8739 & n8980;
  assign n9260 = n8723 & n8735;
  assign n9261 = n9259 & n9260;
  assign n9262 = ~n9258 & ~n9261;
  assign n9263 = n8739 ^ n8723;
  assign n9264 = ~n8981 & n9263;
  assign n9265 = n9264 ^ n8980;
  assign n9269 = n8723 & n9259;
  assign n9270 = ~n8735 & ~n9269;
  assign n9271 = n9265 & ~n9270;
  assign n9266 = ~n8723 & n9256;
  assign n9267 = n8735 & ~n9266;
  assign n9268 = ~n9265 & ~n9267;
  assign n9272 = n9271 ^ n9268;
  assign n9273 = ~n8988 & n9272;
  assign n9274 = n9273 ^ n9271;
  assign n9275 = n9262 & ~n9274;
  assign n9218 = n877 & n6326;
  assign n9219 = x75 & n6565;
  assign n9220 = x76 & n6331;
  assign n9221 = ~n9219 & ~n9220;
  assign n9222 = x77 & n6569;
  assign n9223 = n9221 & ~n9222;
  assign n9224 = ~n9218 & n9223;
  assign n9225 = n9224 ^ x50;
  assign n9215 = n8950 ^ n8896;
  assign n9216 = n8951 & n9215;
  assign n9217 = n9216 ^ n8896;
  assign n9226 = n9225 ^ n9217;
  assign n9203 = n467 & n7830;
  assign n9204 = x70 & n7834;
  assign n9205 = x69 & n7839;
  assign n9206 = ~n9204 & ~n9205;
  assign n9207 = x71 & n8374;
  assign n9208 = n9206 & ~n9207;
  assign n9209 = ~n9203 & n9208;
  assign n9210 = n9209 ^ x56;
  assign n9200 = ~n8926 & ~n8931;
  assign n9193 = x65 ^ x60;
  assign n9194 = n8929 & ~n9193;
  assign n9195 = n9194 ^ x59;
  assign n9196 = n9195 ^ x61;
  assign n9197 = x64 & n9196;
  assign n9198 = n149 & n8929;
  assign n9199 = ~n9197 & ~n9198;
  assign n9201 = n9200 ^ n9199;
  assign n9184 = n300 & n8622;
  assign n9185 = x66 & n8631;
  assign n9186 = n8075 & ~n8621;
  assign n9187 = x68 & n9186;
  assign n9188 = ~n9185 & ~n9187;
  assign n9189 = x67 & n8626;
  assign n9190 = n9188 & ~n9189;
  assign n9191 = ~n9184 & n9190;
  assign n9192 = n9191 ^ x59;
  assign n9202 = n9201 ^ n9192;
  assign n9211 = n9210 ^ n9202;
  assign n9181 = n8938 ^ n8918;
  assign n9182 = n8947 & n9181;
  assign n9183 = n9182 ^ n8918;
  assign n9212 = n9211 ^ n9183;
  assign n9173 = ~n656 & n7076;
  assign n9174 = x72 & n7317;
  assign n9175 = x73 & n7080;
  assign n9176 = ~n9174 & ~n9175;
  assign n9177 = x74 & n7319;
  assign n9178 = n9176 & ~n9177;
  assign n9179 = ~n9173 & n9178;
  assign n9180 = n9179 ^ x53;
  assign n9213 = n9212 ^ n9180;
  assign n9170 = n8948 ^ n8907;
  assign n9171 = ~n8949 & ~n9170;
  assign n9172 = n9171 ^ n8907;
  assign n9214 = n9213 ^ n9172;
  assign n9227 = n9226 ^ n9214;
  assign n9162 = ~n1141 & n5656;
  assign n9163 = x78 & n5895;
  assign n9164 = x79 & n5662;
  assign n9165 = ~n9163 & ~n9164;
  assign n9166 = x80 & n6111;
  assign n9167 = n9165 & ~n9166;
  assign n9168 = ~n9162 & n9167;
  assign n9169 = n9168 ^ x47;
  assign n9228 = n9227 ^ n9169;
  assign n9159 = n8952 ^ n8885;
  assign n9160 = ~n8953 & ~n9159;
  assign n9161 = n9160 ^ n8885;
  assign n9229 = n9228 ^ n9161;
  assign n9151 = n1445 & n5010;
  assign n9152 = x81 & n5223;
  assign n9153 = x82 & n5014;
  assign n9154 = ~n9152 & ~n9153;
  assign n9155 = x83 & n5226;
  assign n9156 = n9154 & ~n9155;
  assign n9157 = ~n9151 & n9156;
  assign n9158 = n9157 ^ x44;
  assign n9230 = n9229 ^ n9158;
  assign n9148 = n8954 ^ n8874;
  assign n9149 = n8955 & n9148;
  assign n9150 = n9149 ^ n8874;
  assign n9231 = n9230 ^ n9150;
  assign n9140 = n1787 & n4415;
  assign n9141 = x84 & n4420;
  assign n9142 = x86 & n4614;
  assign n9143 = ~n9141 & ~n9142;
  assign n9144 = x85 & n4410;
  assign n9145 = n9143 & ~n9144;
  assign n9146 = ~n9140 & n9145;
  assign n9147 = n9146 ^ x41;
  assign n9232 = n9231 ^ n9147;
  assign n9137 = n8956 ^ n8863;
  assign n9138 = ~n8957 & ~n9137;
  assign n9139 = n9138 ^ n8863;
  assign n9233 = n9232 ^ n9139;
  assign n9129 = n2164 & n3829;
  assign n9130 = x87 & n4049;
  assign n9131 = x89 & n4052;
  assign n9132 = ~n9130 & ~n9131;
  assign n9133 = x88 & n3833;
  assign n9134 = n9132 & ~n9133;
  assign n9135 = ~n9129 & n9134;
  assign n9136 = n9135 ^ x38;
  assign n9234 = n9233 ^ n9136;
  assign n9126 = n8958 ^ n8852;
  assign n9127 = n8959 & n9126;
  assign n9128 = n9127 ^ n8852;
  assign n9235 = n9234 ^ n9128;
  assign n9118 = n2585 & n3330;
  assign n9119 = x90 & n3500;
  assign n9120 = x91 & n3334;
  assign n9121 = ~n9119 & ~n9120;
  assign n9122 = x92 & n3502;
  assign n9123 = n9121 & ~n9122;
  assign n9124 = ~n9118 & n9123;
  assign n9125 = n9124 ^ x35;
  assign n9236 = n9235 ^ n9125;
  assign n9115 = n8960 ^ n8841;
  assign n9116 = ~n8961 & ~n9115;
  assign n9117 = n9116 ^ n8841;
  assign n9237 = n9236 ^ n9117;
  assign n9107 = n2836 & n3054;
  assign n9108 = x93 & n2996;
  assign n9109 = x94 & n2840;
  assign n9110 = ~n9108 & ~n9109;
  assign n9111 = x95 & n2998;
  assign n9112 = n9110 & ~n9111;
  assign n9113 = ~n9107 & n9112;
  assign n9114 = n9113 ^ x32;
  assign n9238 = n9237 ^ n9114;
  assign n9104 = n8962 ^ n8830;
  assign n9105 = n8963 & ~n9104;
  assign n9106 = n9105 ^ n8830;
  assign n9239 = n9238 ^ n9106;
  assign n9096 = n2371 & n3556;
  assign n9097 = x96 & n2528;
  assign n9098 = x97 & n2377;
  assign n9099 = ~n9097 & ~n9098;
  assign n9100 = x98 & n2531;
  assign n9101 = n9099 & ~n9100;
  assign n9102 = ~n9096 & n9101;
  assign n9103 = n9102 ^ x29;
  assign n9240 = n9239 ^ n9103;
  assign n9093 = n8827 ^ n8819;
  assign n9094 = ~n8965 & ~n9093;
  assign n9095 = n9094 ^ n8964;
  assign n9241 = n9240 ^ n9095;
  assign n9085 = n1969 & n4105;
  assign n9086 = x99 & n1978;
  assign n9087 = x100 & n1973;
  assign n9088 = ~n9086 & ~n9087;
  assign n9089 = x101 & n2108;
  assign n9090 = n9088 & ~n9089;
  assign n9091 = ~n9085 & n9090;
  assign n9092 = n9091 ^ x26;
  assign n9242 = n9241 ^ n9092;
  assign n9082 = n8966 ^ n8808;
  assign n9083 = n8967 & n9082;
  assign n9084 = n9083 ^ n8808;
  assign n9243 = n9242 ^ n9084;
  assign n9074 = n1624 & n4670;
  assign n9075 = x102 & n1742;
  assign n9076 = x103 & n1628;
  assign n9077 = ~n9075 & ~n9076;
  assign n9078 = x104 & n1744;
  assign n9079 = n9077 & ~n9078;
  assign n9080 = ~n9074 & n9079;
  assign n9081 = n9080 ^ x23;
  assign n9244 = n9243 ^ n9081;
  assign n9071 = n8968 ^ n8797;
  assign n9072 = ~n8969 & ~n9071;
  assign n9073 = n9072 ^ n8797;
  assign n9245 = n9244 ^ n9073;
  assign n9063 = n1296 & n5297;
  assign n9064 = x105 & n1403;
  assign n9065 = x106 & n1300;
  assign n9066 = ~n9064 & ~n9065;
  assign n9067 = x107 & n1406;
  assign n9068 = n9066 & ~n9067;
  assign n9069 = ~n9063 & n9068;
  assign n9070 = n9069 ^ x20;
  assign n9246 = n9245 ^ n9070;
  assign n9060 = n8970 ^ n8786;
  assign n9061 = n8971 & n9060;
  assign n9062 = n9061 ^ n8786;
  assign n9247 = n9246 ^ n9062;
  assign n9052 = n1008 & n5955;
  assign n9053 = x108 & n1101;
  assign n9054 = x109 & n1012;
  assign n9055 = ~n9053 & ~n9054;
  assign n9056 = x110 & n1104;
  assign n9057 = n9055 & ~n9056;
  assign n9058 = ~n9052 & n9057;
  assign n9059 = n9058 ^ x17;
  assign n9248 = n9247 ^ n9059;
  assign n9049 = n8972 ^ n8775;
  assign n9050 = ~n8973 & ~n9049;
  assign n9051 = n9050 ^ n8775;
  assign n9249 = n9248 ^ n9051;
  assign n9041 = n752 & n6656;
  assign n9042 = x111 & n825;
  assign n9043 = x112 & n757;
  assign n9044 = ~n9042 & ~n9043;
  assign n9045 = x113 & n828;
  assign n9046 = n9044 & ~n9045;
  assign n9047 = ~n9041 & n9046;
  assign n9048 = n9047 ^ x14;
  assign n9250 = n9249 ^ n9048;
  assign n9038 = n8974 ^ n8764;
  assign n9039 = n8975 & n9038;
  assign n9040 = n9039 ^ n8764;
  assign n9251 = n9250 ^ n9040;
  assign n9030 = n541 & n7393;
  assign n9031 = x114 & n612;
  assign n9032 = x116 & n615;
  assign n9033 = ~n9031 & ~n9032;
  assign n9034 = x115 & n547;
  assign n9035 = n9033 & ~n9034;
  assign n9036 = ~n9030 & n9035;
  assign n9037 = n9036 ^ x11;
  assign n9252 = n9251 ^ n9037;
  assign n9027 = n8976 ^ n8753;
  assign n9028 = ~n8977 & ~n9027;
  assign n9029 = n9028 ^ n8753;
  assign n9253 = n9252 ^ n9029;
  assign n9011 = x124 & n8434;
  assign n9012 = ~x123 & ~n9011;
  assign n9013 = ~x124 & n8433;
  assign n9014 = ~n9012 & ~n9013;
  assign n9015 = n9014 ^ x124;
  assign n9016 = n163 & ~n9015;
  assign n9017 = n9016 ^ x1;
  assign n9018 = n9017 ^ x125;
  assign n9019 = x0 & ~n9018;
  assign n9020 = ~x123 & n156;
  assign n9021 = ~x0 & ~n9020;
  assign n9022 = x124 ^ x2;
  assign n9023 = x1 & n9022;
  assign n9024 = n9021 & ~n9023;
  assign n9025 = ~n9019 & ~n9024;
  assign n9001 = n8182 ^ x122;
  assign n9002 = n210 & n9001;
  assign n9003 = x120 & n219;
  assign n9004 = x121 & n214;
  assign n9005 = ~n9003 & ~n9004;
  assign n9006 = x122 & n259;
  assign n9007 = n9005 & ~n9006;
  assign n9008 = ~n9002 & n9007;
  assign n9009 = n9008 ^ x5;
  assign n8993 = n372 & n8169;
  assign n8994 = x117 & n433;
  assign n8995 = x119 & n428;
  assign n8996 = ~n8994 & ~n8995;
  assign n8997 = x118 & n376;
  assign n8998 = n8996 & ~n8997;
  assign n8999 = ~n8993 & n8998;
  assign n9000 = n8999 ^ x8;
  assign n9010 = n9009 ^ n9000;
  assign n9026 = n9025 ^ n9010;
  assign n9254 = n9253 ^ n9026;
  assign n8990 = n8978 ^ n8742;
  assign n8991 = n8979 & n8990;
  assign n8992 = n8991 ^ n8742;
  assign n9255 = n9254 ^ n8992;
  assign n9276 = n9275 ^ n9255;
  assign n9571 = n9255 & ~n9256;
  assign n9572 = n9257 & ~n9571;
  assign n9573 = n8988 & ~n9572;
  assign n9574 = ~n9255 & ~n9261;
  assign n9575 = ~n9268 & ~n9574;
  assign n9576 = ~n9573 & ~n9575;
  assign n9577 = ~n9255 & ~n9259;
  assign n9578 = ~n9256 & n9260;
  assign n9579 = n9577 & ~n9578;
  assign n9580 = ~n9576 & ~n9579;
  assign n9530 = n720 & n7076;
  assign n9531 = x74 & n7080;
  assign n9532 = x73 & n7317;
  assign n9533 = ~n9531 & ~n9532;
  assign n9534 = x75 & n7319;
  assign n9535 = n9533 & ~n9534;
  assign n9536 = ~n9530 & n9535;
  assign n9537 = n9536 ^ x53;
  assign n9527 = n9212 ^ n9172;
  assign n9528 = ~n9213 & ~n9527;
  assign n9529 = n9528 ^ n9172;
  assign n9538 = n9537 ^ n9529;
  assign n9516 = n358 & n8622;
  assign n9517 = x67 & n8631;
  assign n9518 = x69 & n9186;
  assign n9519 = ~n9517 & ~n9518;
  assign n9520 = x68 & n8626;
  assign n9521 = n9519 & ~n9520;
  assign n9522 = ~n9516 & n9521;
  assign n9498 = x62 ^ x61;
  assign n9499 = n8929 & n9498;
  assign n9500 = n208 & n9499;
  assign n9493 = x59 & x60;
  assign n9489 = ~x59 & ~x60;
  assign n9501 = n9493 ^ n9489;
  assign n9502 = x61 & n9501;
  assign n9503 = n9502 ^ n9493;
  assign n9504 = ~n9500 & ~n9503;
  assign n9505 = x65 & ~n9504;
  assign n9506 = x61 ^ x60;
  assign n9507 = n9498 & ~n9506;
  assign n9508 = ~n8929 & n9507;
  assign n9509 = x64 & n9508;
  assign n9510 = n149 & n9498;
  assign n9511 = x66 & n8929;
  assign n9512 = ~n9510 & n9511;
  assign n9513 = ~n9509 & ~n9512;
  assign n9514 = ~n9505 & n9513;
  assign n9490 = x61 & x64;
  assign n9491 = n9489 & ~n9490;
  assign n9492 = ~n201 & ~n9491;
  assign n9494 = ~x61 & x64;
  assign n9495 = n9493 & ~n9494;
  assign n9496 = n9492 & ~n9495;
  assign n9497 = x62 & n9496;
  assign n9515 = n9514 ^ n9497;
  assign n9523 = n9522 ^ n9515;
  assign n9485 = n9199 ^ x59;
  assign n9486 = n9485 ^ n9191;
  assign n9487 = n9201 & n9486;
  assign n9488 = n9487 ^ n9191;
  assign n9524 = n9523 ^ n9488;
  assign n9477 = n520 & n7830;
  assign n9478 = x71 & n7834;
  assign n9479 = x70 & n7839;
  assign n9480 = ~n9478 & ~n9479;
  assign n9481 = x72 & n8374;
  assign n9482 = n9480 & ~n9481;
  assign n9483 = ~n9477 & n9482;
  assign n9484 = n9483 ^ x56;
  assign n9525 = n9524 ^ n9484;
  assign n9474 = n9210 ^ n9183;
  assign n9475 = n9211 & ~n9474;
  assign n9476 = n9475 ^ n9183;
  assign n9526 = n9525 ^ n9476;
  assign n9539 = n9538 ^ n9526;
  assign n9465 = n1230 & n5656;
  assign n9466 = x79 & n5895;
  assign n9467 = x81 & n6111;
  assign n9468 = ~n9466 & ~n9467;
  assign n9469 = x80 & n5662;
  assign n9470 = n9468 & ~n9469;
  assign n9471 = ~n9465 & n9470;
  assign n9472 = n9471 ^ x47;
  assign n9457 = n953 & n6326;
  assign n9458 = x77 & n6331;
  assign n9459 = x76 & n6565;
  assign n9460 = ~n9458 & ~n9459;
  assign n9461 = x78 & n6569;
  assign n9462 = n9460 & ~n9461;
  assign n9463 = ~n9457 & n9462;
  assign n9464 = n9463 ^ x50;
  assign n9473 = n9472 ^ n9464;
  assign n9540 = n9539 ^ n9473;
  assign n9454 = n9225 ^ n9214;
  assign n9455 = ~n9226 & n9454;
  assign n9456 = n9455 ^ n9217;
  assign n9541 = n9540 ^ n9456;
  assign n9451 = n9227 ^ n9161;
  assign n9452 = ~n9228 & ~n9451;
  assign n9453 = n9452 ^ n9161;
  assign n9542 = n9541 ^ n9453;
  assign n9443 = n1547 & n5010;
  assign n9444 = x82 & n5223;
  assign n9445 = x84 & n5226;
  assign n9446 = ~n9444 & ~n9445;
  assign n9447 = x83 & n5014;
  assign n9448 = n9446 & ~n9447;
  assign n9449 = ~n9443 & n9448;
  assign n9450 = n9449 ^ x44;
  assign n9543 = n9542 ^ n9450;
  assign n9440 = n9229 ^ n9150;
  assign n9441 = n9230 & n9440;
  assign n9442 = n9441 ^ n9150;
  assign n9544 = n9543 ^ n9442;
  assign n9432 = n1903 & n4415;
  assign n9433 = x85 & n4420;
  assign n9434 = x86 & n4410;
  assign n9435 = ~n9433 & ~n9434;
  assign n9436 = x87 & n4614;
  assign n9437 = n9435 & ~n9436;
  assign n9438 = ~n9432 & n9437;
  assign n9439 = n9438 ^ x41;
  assign n9545 = n9544 ^ n9439;
  assign n9429 = n9231 ^ n9139;
  assign n9430 = ~n9232 & ~n9429;
  assign n9431 = n9430 ^ n9139;
  assign n9546 = n9545 ^ n9431;
  assign n9421 = n2292 & n3829;
  assign n9422 = x88 & n4049;
  assign n9423 = x90 & n4052;
  assign n9424 = ~n9422 & ~n9423;
  assign n9425 = x89 & n3833;
  assign n9426 = n9424 & ~n9425;
  assign n9427 = ~n9421 & n9426;
  assign n9428 = n9427 ^ x38;
  assign n9547 = n9546 ^ n9428;
  assign n9418 = n9233 ^ n9128;
  assign n9419 = n9234 & n9418;
  assign n9420 = n9419 ^ n9128;
  assign n9548 = n9547 ^ n9420;
  assign n9410 = n2726 & n3330;
  assign n9411 = x91 & n3500;
  assign n9412 = x93 & n3502;
  assign n9413 = ~n9411 & ~n9412;
  assign n9414 = x92 & n3334;
  assign n9415 = n9413 & ~n9414;
  assign n9416 = ~n9410 & n9415;
  assign n9417 = n9416 ^ x35;
  assign n9549 = n9548 ^ n9417;
  assign n9407 = n9235 ^ n9117;
  assign n9408 = ~n9236 & ~n9407;
  assign n9409 = n9408 ^ n9117;
  assign n9550 = n9549 ^ n9409;
  assign n9399 = n2836 & n3209;
  assign n9400 = x94 & n2996;
  assign n9401 = x95 & n2840;
  assign n9402 = ~n9400 & ~n9401;
  assign n9403 = x96 & n2998;
  assign n9404 = n9402 & ~n9403;
  assign n9405 = ~n9399 & n9404;
  assign n9406 = n9405 ^ x32;
  assign n9551 = n9550 ^ n9406;
  assign n9396 = n9237 ^ n9106;
  assign n9397 = n9238 & ~n9396;
  assign n9398 = n9397 ^ n9106;
  assign n9552 = n9551 ^ n9398;
  assign n9388 = n2371 & n3730;
  assign n9389 = x97 & n2528;
  assign n9390 = x98 & n2377;
  assign n9391 = ~n9389 & ~n9390;
  assign n9392 = x99 & n2531;
  assign n9393 = n9391 & ~n9392;
  assign n9394 = ~n9388 & n9393;
  assign n9395 = n9394 ^ x29;
  assign n9553 = n9552 ^ n9395;
  assign n9385 = n9103 ^ n9095;
  assign n9386 = ~n9240 & n9385;
  assign n9387 = n9386 ^ n9239;
  assign n9554 = n9553 ^ n9387;
  assign n9377 = n1969 & n4286;
  assign n9378 = x100 & n1978;
  assign n9379 = x102 & n2108;
  assign n9380 = ~n9378 & ~n9379;
  assign n9381 = x101 & n1973;
  assign n9382 = n9380 & ~n9381;
  assign n9383 = ~n9377 & n9382;
  assign n9384 = n9383 ^ x26;
  assign n9555 = n9554 ^ n9384;
  assign n9374 = n9241 ^ n9084;
  assign n9375 = ~n9242 & ~n9374;
  assign n9376 = n9375 ^ n9084;
  assign n9556 = n9555 ^ n9376;
  assign n9366 = n1624 & n4867;
  assign n9367 = x103 & n1742;
  assign n9368 = x104 & n1628;
  assign n9369 = ~n9367 & ~n9368;
  assign n9370 = x105 & n1744;
  assign n9371 = n9369 & ~n9370;
  assign n9372 = ~n9366 & n9371;
  assign n9373 = n9372 ^ x23;
  assign n9557 = n9556 ^ n9373;
  assign n9363 = n9243 ^ n9073;
  assign n9364 = n9244 & n9363;
  assign n9365 = n9364 ^ n9073;
  assign n9558 = n9557 ^ n9365;
  assign n9355 = n1296 & ~n5506;
  assign n9356 = x106 & n1403;
  assign n9357 = x107 & n1300;
  assign n9358 = ~n9356 & ~n9357;
  assign n9359 = x108 & n1406;
  assign n9360 = n9358 & ~n9359;
  assign n9361 = ~n9355 & n9360;
  assign n9362 = n9361 ^ x20;
  assign n9559 = n9558 ^ n9362;
  assign n9352 = n9245 ^ n9062;
  assign n9353 = ~n9246 & ~n9352;
  assign n9354 = n9353 ^ n9062;
  assign n9560 = n9559 ^ n9354;
  assign n9344 = n1008 & n6178;
  assign n9345 = x109 & n1101;
  assign n9346 = x110 & n1012;
  assign n9347 = ~n9345 & ~n9346;
  assign n9348 = x111 & n1104;
  assign n9349 = n9347 & ~n9348;
  assign n9350 = ~n9344 & n9349;
  assign n9351 = n9350 ^ x17;
  assign n9561 = n9560 ^ n9351;
  assign n9341 = n9247 ^ n9051;
  assign n9342 = n9248 & n9341;
  assign n9343 = n9342 ^ n9051;
  assign n9562 = n9561 ^ n9343;
  assign n9333 = n752 & n6892;
  assign n9334 = x112 & n825;
  assign n9335 = x114 & n828;
  assign n9336 = ~n9334 & ~n9335;
  assign n9337 = x113 & n757;
  assign n9338 = n9336 & ~n9337;
  assign n9339 = ~n9333 & n9338;
  assign n9340 = n9339 ^ x14;
  assign n9563 = n9562 ^ n9340;
  assign n9330 = n9249 ^ n9040;
  assign n9331 = ~n9250 & ~n9330;
  assign n9332 = n9331 ^ n9040;
  assign n9564 = n9563 ^ n9332;
  assign n9322 = n541 & n7643;
  assign n9323 = x115 & n612;
  assign n9324 = x117 & n615;
  assign n9325 = ~n9323 & ~n9324;
  assign n9326 = x116 & n547;
  assign n9327 = n9325 & ~n9326;
  assign n9328 = ~n9322 & n9327;
  assign n9329 = n9328 ^ x11;
  assign n9565 = n9564 ^ n9329;
  assign n9319 = n9251 ^ n9029;
  assign n9320 = n9252 & n9319;
  assign n9321 = n9320 ^ n9029;
  assign n9566 = n9565 ^ n9321;
  assign n9309 = n8435 ^ x123;
  assign n9310 = n210 & n9309;
  assign n9311 = x121 & n219;
  assign n9312 = x123 & n259;
  assign n9313 = ~n9311 & ~n9312;
  assign n9314 = x122 & n214;
  assign n9315 = n9313 & ~n9314;
  assign n9316 = ~n9310 & n9315;
  assign n9317 = n9316 ^ x5;
  assign n9301 = n372 & ~n8424;
  assign n9302 = x118 & n433;
  assign n9303 = x119 & n376;
  assign n9304 = ~n9302 & ~n9303;
  assign n9305 = x120 & n428;
  assign n9306 = n9304 & ~n9305;
  assign n9307 = ~n9301 & n9306;
  assign n9308 = n9307 ^ x8;
  assign n9318 = n9317 ^ n9308;
  assign n9567 = n9566 ^ n9318;
  assign n9286 = ~x124 & x125;
  assign n9287 = ~n9014 & n9286;
  assign n9288 = x124 & ~x125;
  assign n9289 = ~n9012 & n9288;
  assign n9290 = ~n9287 & ~n9289;
  assign n9291 = n163 & n9290;
  assign n9292 = n9291 ^ x1;
  assign n9293 = n9292 ^ x126;
  assign n9294 = x0 & n9293;
  assign n9295 = ~x1 & x124;
  assign n9296 = ~x0 & ~n9295;
  assign n9297 = x1 & x125;
  assign n9298 = n9297 ^ x2;
  assign n9299 = n9296 & n9298;
  assign n9300 = ~n9294 & ~n9299;
  assign n9568 = n9567 ^ n9300;
  assign n9278 = n9253 ^ n9000;
  assign n9283 = n9253 ^ n8992;
  assign n9284 = ~n9278 & ~n9283;
  assign n9285 = n9284 ^ n8992;
  assign n9569 = n9568 ^ n9285;
  assign n9277 = n9025 ^ n9009;
  assign n9279 = n9278 ^ n8992;
  assign n9280 = n9279 ^ n9009;
  assign n9281 = ~n9277 & n9280;
  assign n9282 = n9281 ^ n9025;
  assign n9570 = n9569 ^ n9282;
  assign n9581 = n9580 ^ n9570;
  assign n9831 = ~n594 & n7830;
  assign n9832 = x72 & n7834;
  assign n9833 = x71 & n7839;
  assign n9834 = ~n9832 & ~n9833;
  assign n9835 = x73 & n8374;
  assign n9836 = n9834 & ~n9835;
  assign n9837 = ~n9831 & n9836;
  assign n9838 = n9837 ^ x56;
  assign n9828 = n9524 ^ n9476;
  assign n9829 = ~n9525 & ~n9828;
  assign n9830 = n9829 ^ n9476;
  assign n9839 = n9838 ^ n9830;
  assign n9816 = n9199 & ~n9200;
  assign n9817 = n9523 ^ n9191;
  assign n9818 = ~n9192 & n9817;
  assign n9819 = ~n9816 & n9818;
  assign n9820 = ~n9199 & n9200;
  assign n9821 = n9820 ^ n9515;
  assign n9822 = n9522 ^ x59;
  assign n9823 = n9822 ^ n9515;
  assign n9824 = ~n9821 & ~n9823;
  assign n9825 = n9824 ^ n9820;
  assign n9826 = ~n9819 & ~n9825;
  assign n9800 = n162 & n9498;
  assign n9801 = n9800 ^ x67;
  assign n9802 = n8929 & n9801;
  assign n9803 = x65 & n9508;
  assign n9804 = x66 & n9503;
  assign n9805 = ~n9803 & ~n9804;
  assign n9806 = ~n9802 & n9805;
  assign n9807 = n9806 ^ x62;
  assign n9798 = x63 ^ x62;
  assign n9799 = x64 & n9798;
  assign n9808 = n9807 ^ n9799;
  assign n9809 = x62 & ~n9496;
  assign n9810 = n9514 & n9809;
  assign n9811 = n9808 & ~n9810;
  assign n9812 = n9806 & n9810;
  assign n9813 = ~n9799 & n9812;
  assign n9814 = ~n9811 & ~n9813;
  assign n9790 = n416 & n8622;
  assign n9791 = x68 & n8631;
  assign n9792 = x70 & n9186;
  assign n9793 = ~n9791 & ~n9792;
  assign n9794 = x69 & n8626;
  assign n9795 = n9793 & ~n9794;
  assign n9796 = ~n9790 & n9795;
  assign n9797 = n9796 ^ x59;
  assign n9815 = n9814 ^ n9797;
  assign n9827 = n9826 ^ n9815;
  assign n9840 = n9839 ^ n9827;
  assign n9782 = n799 & n7076;
  assign n9783 = x74 & n7317;
  assign n9784 = x75 & n7080;
  assign n9785 = ~n9783 & ~n9784;
  assign n9786 = x76 & n7319;
  assign n9787 = n9785 & ~n9786;
  assign n9788 = ~n9782 & n9787;
  assign n9789 = n9788 ^ x53;
  assign n9841 = n9840 ^ n9789;
  assign n9779 = n9537 ^ n9526;
  assign n9780 = ~n9538 & n9779;
  assign n9781 = n9780 ^ n9529;
  assign n9842 = n9841 ^ n9781;
  assign n9775 = n9539 ^ n9456;
  assign n9776 = n9539 ^ n9464;
  assign n9777 = ~n9775 & ~n9776;
  assign n9778 = n9777 ^ n9456;
  assign n9843 = n9842 ^ n9778;
  assign n9767 = n1054 & n6326;
  assign n9768 = x77 & n6565;
  assign n9769 = x79 & n6569;
  assign n9770 = ~n9768 & ~n9769;
  assign n9771 = x78 & n6331;
  assign n9772 = n9770 & ~n9771;
  assign n9773 = ~n9767 & n9772;
  assign n9774 = n9773 ^ x50;
  assign n9844 = n9843 ^ n9774;
  assign n9759 = n1345 & n5656;
  assign n9760 = x80 & n5895;
  assign n9761 = x82 & n6111;
  assign n9762 = ~n9760 & ~n9761;
  assign n9763 = x81 & n5662;
  assign n9764 = n9762 & ~n9763;
  assign n9765 = ~n9759 & n9764;
  assign n9766 = n9765 ^ x47;
  assign n9845 = n9844 ^ n9766;
  assign n9756 = n9472 ^ n9453;
  assign n9757 = n9541 & ~n9756;
  assign n9758 = n9757 ^ n9453;
  assign n9846 = n9845 ^ n9758;
  assign n9748 = n1674 & n5010;
  assign n9749 = x83 & n5223;
  assign n9750 = x84 & n5014;
  assign n9751 = ~n9749 & ~n9750;
  assign n9752 = x85 & n5226;
  assign n9753 = n9751 & ~n9752;
  assign n9754 = ~n9748 & n9753;
  assign n9755 = n9754 ^ x44;
  assign n9847 = n9846 ^ n9755;
  assign n9745 = n9542 ^ n9442;
  assign n9746 = ~n9543 & ~n9745;
  assign n9747 = n9746 ^ n9442;
  assign n9848 = n9847 ^ n9747;
  assign n9737 = n2040 & n4415;
  assign n9738 = x86 & n4420;
  assign n9739 = x88 & n4614;
  assign n9740 = ~n9738 & ~n9739;
  assign n9741 = x87 & n4410;
  assign n9742 = n9740 & ~n9741;
  assign n9743 = ~n9737 & n9742;
  assign n9744 = n9743 ^ x41;
  assign n9849 = n9848 ^ n9744;
  assign n9734 = n9544 ^ n9431;
  assign n9735 = n9545 & n9734;
  assign n9736 = n9735 ^ n9431;
  assign n9850 = n9849 ^ n9736;
  assign n9726 = n2447 & n3829;
  assign n9727 = x89 & n4049;
  assign n9728 = x91 & n4052;
  assign n9729 = ~n9727 & ~n9728;
  assign n9730 = x90 & n3833;
  assign n9731 = n9729 & ~n9730;
  assign n9732 = ~n9726 & n9731;
  assign n9733 = n9732 ^ x38;
  assign n9851 = n9850 ^ n9733;
  assign n9723 = n9546 ^ n9420;
  assign n9724 = ~n9547 & ~n9723;
  assign n9725 = n9724 ^ n9420;
  assign n9852 = n9851 ^ n9725;
  assign n9715 = n2895 & n3330;
  assign n9716 = x92 & n3500;
  assign n9717 = x94 & n3502;
  assign n9718 = ~n9716 & ~n9717;
  assign n9719 = x93 & n3334;
  assign n9720 = n9718 & ~n9719;
  assign n9721 = ~n9715 & n9720;
  assign n9722 = n9721 ^ x35;
  assign n9853 = n9852 ^ n9722;
  assign n9712 = n9548 ^ n9409;
  assign n9713 = n9549 & n9712;
  assign n9714 = n9713 ^ n9409;
  assign n9854 = n9853 ^ n9714;
  assign n9704 = n2836 & n3388;
  assign n9705 = x95 & n2996;
  assign n9706 = x96 & n2840;
  assign n9707 = ~n9705 & ~n9706;
  assign n9708 = x97 & n2998;
  assign n9709 = n9707 & ~n9708;
  assign n9710 = ~n9704 & n9709;
  assign n9711 = n9710 ^ x32;
  assign n9855 = n9854 ^ n9711;
  assign n9701 = n9550 ^ n9398;
  assign n9702 = ~n9551 & n9701;
  assign n9703 = n9702 ^ n9398;
  assign n9856 = n9855 ^ n9703;
  assign n9693 = n2371 & n3925;
  assign n9694 = x98 & n2528;
  assign n9695 = x99 & n2377;
  assign n9696 = ~n9694 & ~n9695;
  assign n9697 = x100 & n2531;
  assign n9698 = n9696 & ~n9697;
  assign n9699 = ~n9693 & n9698;
  assign n9700 = n9699 ^ x29;
  assign n9857 = n9856 ^ n9700;
  assign n9690 = n9395 ^ n9387;
  assign n9691 = n9553 & n9690;
  assign n9692 = n9691 ^ n9552;
  assign n9858 = n9857 ^ n9692;
  assign n9682 = n1969 & n4481;
  assign n9683 = x101 & n1978;
  assign n9684 = x102 & n1973;
  assign n9685 = ~n9683 & ~n9684;
  assign n9686 = x103 & n2108;
  assign n9687 = n9685 & ~n9686;
  assign n9688 = ~n9682 & n9687;
  assign n9689 = n9688 ^ x26;
  assign n9859 = n9858 ^ n9689;
  assign n9679 = n9554 ^ n9376;
  assign n9680 = n9555 & n9679;
  assign n9681 = n9680 ^ n9376;
  assign n9860 = n9859 ^ n9681;
  assign n9671 = n1624 & n5088;
  assign n9672 = x105 & n1628;
  assign n9673 = x104 & n1742;
  assign n9674 = ~n9672 & ~n9673;
  assign n9675 = x106 & n1744;
  assign n9676 = n9674 & ~n9675;
  assign n9677 = ~n9671 & n9676;
  assign n9678 = n9677 ^ x23;
  assign n9861 = n9860 ^ n9678;
  assign n9668 = n9556 ^ n9365;
  assign n9669 = ~n9557 & ~n9668;
  assign n9670 = n9669 ^ n9365;
  assign n9862 = n9861 ^ n9670;
  assign n9660 = n1296 & ~n5737;
  assign n9661 = x107 & n1403;
  assign n9662 = x108 & n1300;
  assign n9663 = ~n9661 & ~n9662;
  assign n9664 = x109 & n1406;
  assign n9665 = n9663 & ~n9664;
  assign n9666 = ~n9660 & n9665;
  assign n9667 = n9666 ^ x20;
  assign n9863 = n9862 ^ n9667;
  assign n9657 = n9558 ^ n9354;
  assign n9658 = n9559 & n9657;
  assign n9659 = n9658 ^ n9354;
  assign n9864 = n9863 ^ n9659;
  assign n9649 = n1008 & n6420;
  assign n9650 = x110 & n1101;
  assign n9651 = x111 & n1012;
  assign n9652 = ~n9650 & ~n9651;
  assign n9653 = x112 & n1104;
  assign n9654 = n9652 & ~n9653;
  assign n9655 = ~n9649 & n9654;
  assign n9656 = n9655 ^ x17;
  assign n9865 = n9864 ^ n9656;
  assign n9646 = n9560 ^ n9343;
  assign n9647 = ~n9561 & ~n9646;
  assign n9648 = n9647 ^ n9343;
  assign n9866 = n9865 ^ n9648;
  assign n9638 = n752 & n7150;
  assign n9639 = x113 & n825;
  assign n9640 = x115 & n828;
  assign n9641 = ~n9639 & ~n9640;
  assign n9642 = x114 & n757;
  assign n9643 = n9641 & ~n9642;
  assign n9644 = ~n9638 & n9643;
  assign n9645 = n9644 ^ x14;
  assign n9867 = n9866 ^ n9645;
  assign n9635 = n9562 ^ n9332;
  assign n9636 = n9563 & n9635;
  assign n9637 = n9636 ^ n9332;
  assign n9868 = n9867 ^ n9637;
  assign n9627 = n541 & n7919;
  assign n9628 = x116 & n612;
  assign n9629 = x118 & n615;
  assign n9630 = ~n9628 & ~n9629;
  assign n9631 = x117 & n547;
  assign n9632 = n9630 & ~n9631;
  assign n9633 = ~n9627 & n9632;
  assign n9634 = n9633 ^ x11;
  assign n9869 = n9868 ^ n9634;
  assign n9624 = n9564 ^ n9321;
  assign n9625 = ~n9565 & ~n9624;
  assign n9626 = n9625 ^ n9321;
  assign n9870 = n9869 ^ n9626;
  assign n9614 = n8725 ^ x124;
  assign n9615 = n210 & n9614;
  assign n9616 = x122 & n219;
  assign n9617 = x123 & n214;
  assign n9618 = ~n9616 & ~n9617;
  assign n9619 = x124 & n259;
  assign n9620 = n9618 & ~n9619;
  assign n9621 = ~n9615 & n9620;
  assign n9622 = n9621 ^ x5;
  assign n9606 = n372 & n8715;
  assign n9607 = x119 & n433;
  assign n9608 = x121 & n428;
  assign n9609 = ~n9607 & ~n9608;
  assign n9610 = x120 & n376;
  assign n9611 = n9609 & ~n9610;
  assign n9612 = ~n9606 & n9611;
  assign n9613 = n9612 ^ x8;
  assign n9623 = n9622 ^ n9613;
  assign n9871 = n9870 ^ n9623;
  assign n9595 = x125 & ~x126;
  assign n9596 = ~n9287 & n9595;
  assign n9597 = ~x125 & x126;
  assign n9598 = ~n9289 & n9597;
  assign n9599 = ~n9596 & ~n9598;
  assign n9600 = n163 & n9599;
  assign n9601 = n9600 ^ x1;
  assign n9602 = n9601 ^ x127;
  assign n9591 = ~x125 & n156;
  assign n9592 = x126 ^ x2;
  assign n9593 = x1 & n9592;
  assign n9594 = ~n9591 & ~n9593;
  assign n9603 = n9602 ^ n9594;
  assign n9604 = ~x0 & ~n9603;
  assign n9605 = n9604 ^ n9602;
  assign n9872 = n9871 ^ n9605;
  assign n9588 = n9566 ^ n9317;
  assign n9589 = ~n9318 & ~n9588;
  assign n9590 = n9589 ^ n9566;
  assign n9873 = n9872 ^ n9590;
  assign n9585 = n9567 ^ n9285;
  assign n9586 = n9568 & n9585;
  assign n9587 = n9586 ^ n9285;
  assign n9874 = n9873 ^ n9587;
  assign n9582 = n9580 ^ n9569;
  assign n9583 = n9570 & n9582;
  assign n9584 = n9583 ^ n9580;
  assign n9875 = n9874 ^ n9584;
  assign n10122 = n877 & n7076;
  assign n10123 = x76 & n7080;
  assign n10124 = x75 & n7317;
  assign n10125 = ~n10123 & ~n10124;
  assign n10126 = x77 & n7319;
  assign n10127 = n10125 & ~n10126;
  assign n10128 = ~n10122 & n10127;
  assign n10129 = n10128 ^ x53;
  assign n10119 = n9840 ^ n9781;
  assign n10120 = ~n9841 & ~n10119;
  assign n10121 = n10120 ^ n9781;
  assign n10130 = n10129 ^ n10121;
  assign n10112 = n9799 & ~n9807;
  assign n10113 = ~n9812 & ~n10112;
  assign n10102 = n300 & n9499;
  assign n10103 = x67 & n9503;
  assign n10104 = x66 & n9508;
  assign n10105 = ~n10103 & ~n10104;
  assign n10106 = n8929 & ~n9498;
  assign n10107 = x68 & n10106;
  assign n10108 = n10105 & ~n10107;
  assign n10109 = ~n10102 & n10108;
  assign n10110 = n10109 ^ x62;
  assign n10098 = x65 & n9798;
  assign n10099 = x62 & x63;
  assign n10100 = x64 & n10099;
  assign n10101 = ~n10098 & ~n10100;
  assign n10111 = n10110 ^ n10101;
  assign n10114 = n10113 ^ n10111;
  assign n10090 = n467 & n8622;
  assign n10091 = x69 & n8631;
  assign n10092 = x71 & n9186;
  assign n10093 = ~n10091 & ~n10092;
  assign n10094 = x70 & n8626;
  assign n10095 = n10093 & ~n10094;
  assign n10096 = ~n10090 & n10095;
  assign n10097 = n10096 ^ x59;
  assign n10115 = n10114 ^ n10097;
  assign n10087 = n9826 ^ n9814;
  assign n10088 = n9815 & ~n10087;
  assign n10089 = n10088 ^ n9826;
  assign n10116 = n10115 ^ n10089;
  assign n10079 = ~n656 & n7830;
  assign n10080 = x73 & n7834;
  assign n10081 = x72 & n7839;
  assign n10082 = ~n10080 & ~n10081;
  assign n10083 = x74 & n8374;
  assign n10084 = n10082 & ~n10083;
  assign n10085 = ~n10079 & n10084;
  assign n10086 = n10085 ^ x56;
  assign n10117 = n10116 ^ n10086;
  assign n10076 = n9838 ^ n9827;
  assign n10077 = ~n9839 & n10076;
  assign n10078 = n10077 ^ n9830;
  assign n10118 = n10117 ^ n10078;
  assign n10131 = n10130 ^ n10118;
  assign n10068 = ~n1141 & n6326;
  assign n10069 = x78 & n6565;
  assign n10070 = x79 & n6331;
  assign n10071 = ~n10069 & ~n10070;
  assign n10072 = x80 & n6569;
  assign n10073 = n10071 & ~n10072;
  assign n10074 = ~n10068 & n10073;
  assign n10075 = n10074 ^ x50;
  assign n10132 = n10131 ^ n10075;
  assign n10065 = n9842 ^ n9774;
  assign n10066 = n9843 & n10065;
  assign n10067 = n10066 ^ n9778;
  assign n10133 = n10132 ^ n10067;
  assign n10057 = n1445 & n5656;
  assign n10058 = x81 & n5895;
  assign n10059 = x82 & n5662;
  assign n10060 = ~n10058 & ~n10059;
  assign n10061 = x83 & n6111;
  assign n10062 = n10060 & ~n10061;
  assign n10063 = ~n10057 & n10062;
  assign n10064 = n10063 ^ x47;
  assign n10134 = n10133 ^ n10064;
  assign n10054 = n9844 ^ n9758;
  assign n10055 = ~n9845 & ~n10054;
  assign n10056 = n10055 ^ n9758;
  assign n10135 = n10134 ^ n10056;
  assign n10046 = n1787 & n5010;
  assign n10047 = x85 & n5014;
  assign n10048 = x86 & n5226;
  assign n10049 = ~n10047 & ~n10048;
  assign n10050 = x84 & n5223;
  assign n10051 = n10049 & ~n10050;
  assign n10052 = ~n10046 & n10051;
  assign n10053 = n10052 ^ x44;
  assign n10136 = n10135 ^ n10053;
  assign n10043 = n9846 ^ n9747;
  assign n10044 = n9847 & n10043;
  assign n10045 = n10044 ^ n9747;
  assign n10137 = n10136 ^ n10045;
  assign n10035 = n2164 & n4415;
  assign n10036 = x87 & n4420;
  assign n10037 = x88 & n4410;
  assign n10038 = ~n10036 & ~n10037;
  assign n10039 = x89 & n4614;
  assign n10040 = n10038 & ~n10039;
  assign n10041 = ~n10035 & n10040;
  assign n10042 = n10041 ^ x41;
  assign n10138 = n10137 ^ n10042;
  assign n10032 = n9848 ^ n9736;
  assign n10033 = ~n9849 & ~n10032;
  assign n10034 = n10033 ^ n9736;
  assign n10139 = n10138 ^ n10034;
  assign n10024 = n2585 & n3829;
  assign n10025 = x90 & n4049;
  assign n10026 = x91 & n3833;
  assign n10027 = ~n10025 & ~n10026;
  assign n10028 = x92 & n4052;
  assign n10029 = n10027 & ~n10028;
  assign n10030 = ~n10024 & n10029;
  assign n10031 = n10030 ^ x38;
  assign n10140 = n10139 ^ n10031;
  assign n10021 = n9850 ^ n9725;
  assign n10022 = n9851 & n10021;
  assign n10023 = n10022 ^ n9725;
  assign n10141 = n10140 ^ n10023;
  assign n10013 = n3054 & n3330;
  assign n10014 = x93 & n3500;
  assign n10015 = x94 & n3334;
  assign n10016 = ~n10014 & ~n10015;
  assign n10017 = x95 & n3502;
  assign n10018 = n10016 & ~n10017;
  assign n10019 = ~n10013 & n10018;
  assign n10020 = n10019 ^ x35;
  assign n10142 = n10141 ^ n10020;
  assign n10010 = n9852 ^ n9714;
  assign n10011 = ~n9853 & ~n10010;
  assign n10012 = n10011 ^ n9714;
  assign n10143 = n10142 ^ n10012;
  assign n10002 = n2836 & n3556;
  assign n10003 = x96 & n2996;
  assign n10004 = x97 & n2840;
  assign n10005 = ~n10003 & ~n10004;
  assign n10006 = x98 & n2998;
  assign n10007 = n10005 & ~n10006;
  assign n10008 = ~n10002 & n10007;
  assign n10009 = n10008 ^ x32;
  assign n10144 = n10143 ^ n10009;
  assign n9999 = n9854 ^ n9703;
  assign n10000 = n9855 & ~n9999;
  assign n10001 = n10000 ^ n9703;
  assign n10145 = n10144 ^ n10001;
  assign n9991 = n2371 & n4105;
  assign n9992 = x100 & n2377;
  assign n9993 = x99 & n2528;
  assign n9994 = ~n9992 & ~n9993;
  assign n9995 = x101 & n2531;
  assign n9996 = n9994 & ~n9995;
  assign n9997 = ~n9991 & n9996;
  assign n9998 = n9997 ^ x29;
  assign n10146 = n10145 ^ n9998;
  assign n9988 = n9856 ^ n9692;
  assign n9989 = n9857 & ~n9988;
  assign n9990 = n9989 ^ n9692;
  assign n10147 = n10146 ^ n9990;
  assign n9980 = n1969 & n4670;
  assign n9981 = x102 & n1978;
  assign n9982 = x103 & n1973;
  assign n9983 = ~n9981 & ~n9982;
  assign n9984 = x104 & n2108;
  assign n9985 = n9983 & ~n9984;
  assign n9986 = ~n9980 & n9985;
  assign n9987 = n9986 ^ x26;
  assign n10148 = n10147 ^ n9987;
  assign n9977 = n9858 ^ n9681;
  assign n9978 = n9859 & n9977;
  assign n9979 = n9978 ^ n9681;
  assign n10149 = n10148 ^ n9979;
  assign n9969 = n1624 & n5297;
  assign n9970 = x106 & n1628;
  assign n9971 = x105 & n1742;
  assign n9972 = ~n9970 & ~n9971;
  assign n9973 = x107 & n1744;
  assign n9974 = n9972 & ~n9973;
  assign n9975 = ~n9969 & n9974;
  assign n9976 = n9975 ^ x23;
  assign n10150 = n10149 ^ n9976;
  assign n9966 = n9860 ^ n9670;
  assign n9967 = ~n9861 & ~n9966;
  assign n9968 = n9967 ^ n9670;
  assign n10151 = n10150 ^ n9968;
  assign n9958 = n1296 & n5955;
  assign n9959 = x109 & n1300;
  assign n9960 = x108 & n1403;
  assign n9961 = ~n9959 & ~n9960;
  assign n9962 = x110 & n1406;
  assign n9963 = n9961 & ~n9962;
  assign n9964 = ~n9958 & n9963;
  assign n9965 = n9964 ^ x20;
  assign n10152 = n10151 ^ n9965;
  assign n9955 = n9862 ^ n9659;
  assign n9956 = n9863 & n9955;
  assign n9957 = n9956 ^ n9659;
  assign n10153 = n10152 ^ n9957;
  assign n9947 = n1008 & n6656;
  assign n9948 = x111 & n1101;
  assign n9949 = x112 & n1012;
  assign n9950 = ~n9948 & ~n9949;
  assign n9951 = x113 & n1104;
  assign n9952 = n9950 & ~n9951;
  assign n9953 = ~n9947 & n9952;
  assign n9954 = n9953 ^ x17;
  assign n10154 = n10153 ^ n9954;
  assign n9944 = n9864 ^ n9648;
  assign n9945 = ~n9865 & ~n9944;
  assign n9946 = n9945 ^ n9648;
  assign n10155 = n10154 ^ n9946;
  assign n9936 = n752 & n7393;
  assign n9937 = x115 & n757;
  assign n9938 = x114 & n825;
  assign n9939 = ~n9937 & ~n9938;
  assign n9940 = x116 & n828;
  assign n9941 = n9939 & ~n9940;
  assign n9942 = ~n9936 & n9941;
  assign n9943 = n9942 ^ x14;
  assign n10156 = n10155 ^ n9943;
  assign n9933 = n9866 ^ n9637;
  assign n9934 = n9867 & n9933;
  assign n9935 = n9934 ^ n9637;
  assign n10157 = n10156 ^ n9935;
  assign n9925 = n541 & n8169;
  assign n9926 = x117 & n612;
  assign n9927 = x118 & n547;
  assign n9928 = ~n9926 & ~n9927;
  assign n9929 = x119 & n615;
  assign n9930 = n9928 & ~n9929;
  assign n9931 = ~n9925 & n9930;
  assign n9932 = n9931 ^ x11;
  assign n10158 = n10157 ^ n9932;
  assign n9922 = n9868 ^ n9626;
  assign n9923 = ~n9869 & ~n9922;
  assign n9924 = n9923 ^ n9626;
  assign n10159 = n10158 ^ n9924;
  assign n9911 = x125 ^ x124;
  assign n9912 = n9911 ^ n9014;
  assign n9913 = n210 & n9912;
  assign n9914 = x123 & n219;
  assign n9915 = x125 & n259;
  assign n9916 = ~n9914 & ~n9915;
  assign n9917 = x124 & n214;
  assign n9918 = n9916 & ~n9917;
  assign n9919 = ~n9913 & n9918;
  assign n9920 = n9919 ^ x5;
  assign n9903 = n372 & n9001;
  assign n9904 = x120 & n433;
  assign n9905 = x121 & n376;
  assign n9906 = ~n9904 & ~n9905;
  assign n9907 = x122 & n428;
  assign n9908 = n9906 & ~n9907;
  assign n9909 = ~n9903 & n9908;
  assign n9910 = n9909 ^ x8;
  assign n9921 = n9920 ^ n9910;
  assign n10160 = n10159 ^ n9921;
  assign n9885 = ~x126 & x127;
  assign n9886 = ~n9596 & n9885;
  assign n9887 = x126 & ~x127;
  assign n9888 = ~n9598 & n9887;
  assign n9889 = ~n9886 & ~n9888;
  assign n9890 = n163 & n9889;
  assign n9891 = n9890 ^ x1;
  assign n9892 = x0 & n9891;
  assign n9893 = ~x126 & n156;
  assign n9894 = x1 & ~x2;
  assign n9895 = x127 & n9894;
  assign n9896 = ~n9893 & ~n9895;
  assign n9897 = ~x0 & ~n9896;
  assign n9898 = ~x1 & x126;
  assign n9899 = x2 & ~x127;
  assign n9900 = ~n9898 & n9899;
  assign n9901 = ~n9897 & ~n9900;
  assign n9902 = ~n9892 & n9901;
  assign n10161 = n10160 ^ n9902;
  assign n9882 = n9870 ^ n9622;
  assign n9883 = ~n9623 & ~n9882;
  assign n9884 = n9883 ^ n9870;
  assign n10162 = n10161 ^ n9884;
  assign n9879 = n9605 ^ n9590;
  assign n9880 = n9872 & ~n9879;
  assign n9881 = n9880 ^ n9871;
  assign n10163 = n10162 ^ n9881;
  assign n9876 = n9587 ^ n9584;
  assign n9877 = ~n9874 & ~n9876;
  assign n9878 = n9877 ^ n9584;
  assign n10164 = n10163 ^ n9878;
  assign n10430 = x127 & ~n9886;
  assign n10431 = x0 & n10430;
  assign n10432 = ~x2 & ~n10431;
  assign n10433 = x0 & n9886;
  assign n10434 = ~x1 & x127;
  assign n10435 = ~n10433 & n10434;
  assign n10436 = ~n10432 & ~n10435;
  assign n10427 = n10159 ^ n9920;
  assign n10428 = ~n9921 & n10427;
  assign n10429 = n10428 ^ n10159;
  assign n10437 = n10436 ^ n10429;
  assign n10388 = n953 & n7076;
  assign n10389 = x77 & n7080;
  assign n10390 = x76 & n7317;
  assign n10391 = ~n10389 & ~n10390;
  assign n10392 = x78 & n7319;
  assign n10393 = n10391 & ~n10392;
  assign n10394 = ~n10388 & n10393;
  assign n10395 = n10394 ^ x53;
  assign n10385 = n10129 ^ n10118;
  assign n10386 = ~n10130 & n10385;
  assign n10387 = n10386 ^ n10121;
  assign n10396 = n10395 ^ n10387;
  assign n10375 = n720 & n7830;
  assign n10376 = x74 & n7834;
  assign n10377 = x73 & n7839;
  assign n10378 = ~n10376 & ~n10377;
  assign n10379 = x75 & n8374;
  assign n10380 = n10378 & ~n10379;
  assign n10381 = ~n10375 & n10380;
  assign n10382 = n10381 ^ x56;
  assign n10372 = n10116 ^ n10078;
  assign n10373 = ~n10117 & ~n10372;
  assign n10374 = n10373 ^ n10078;
  assign n10383 = n10382 ^ n10374;
  assign n10365 = x66 & n9798;
  assign n10366 = x65 & n10099;
  assign n10367 = ~n10365 & ~n10366;
  assign n10362 = n10113 ^ n10110;
  assign n10363 = ~n10111 & n10362;
  assign n10364 = n10363 ^ n10113;
  assign n10368 = n10367 ^ n10364;
  assign n10354 = n358 & n9499;
  assign n10355 = x68 & n9503;
  assign n10356 = x67 & n9508;
  assign n10357 = ~n10355 & ~n10356;
  assign n10358 = x69 & n10106;
  assign n10359 = n10357 & ~n10358;
  assign n10360 = ~n10354 & n10359;
  assign n10361 = n10360 ^ x62;
  assign n10369 = n10368 ^ n10361;
  assign n10346 = n520 & n8622;
  assign n10347 = x70 & n8631;
  assign n10348 = x71 & n8626;
  assign n10349 = ~n10347 & ~n10348;
  assign n10350 = x72 & n9186;
  assign n10351 = n10349 & ~n10350;
  assign n10352 = ~n10346 & n10351;
  assign n10353 = n10352 ^ x59;
  assign n10370 = n10369 ^ n10353;
  assign n10343 = n10114 ^ n10089;
  assign n10344 = ~n10115 & n10343;
  assign n10345 = n10344 ^ n10089;
  assign n10371 = n10370 ^ n10345;
  assign n10384 = n10383 ^ n10371;
  assign n10397 = n10396 ^ n10384;
  assign n10335 = n1230 & n6326;
  assign n10336 = x79 & n6565;
  assign n10337 = x80 & n6331;
  assign n10338 = ~n10336 & ~n10337;
  assign n10339 = x81 & n6569;
  assign n10340 = n10338 & ~n10339;
  assign n10341 = ~n10335 & n10340;
  assign n10342 = n10341 ^ x50;
  assign n10398 = n10397 ^ n10342;
  assign n10332 = n10131 ^ n10067;
  assign n10333 = ~n10132 & ~n10332;
  assign n10334 = n10333 ^ n10067;
  assign n10399 = n10398 ^ n10334;
  assign n10324 = n1547 & n5656;
  assign n10325 = x82 & n5895;
  assign n10326 = x84 & n6111;
  assign n10327 = ~n10325 & ~n10326;
  assign n10328 = x83 & n5662;
  assign n10329 = n10327 & ~n10328;
  assign n10330 = ~n10324 & n10329;
  assign n10331 = n10330 ^ x47;
  assign n10400 = n10399 ^ n10331;
  assign n10321 = n10133 ^ n10056;
  assign n10322 = n10134 & n10321;
  assign n10323 = n10322 ^ n10056;
  assign n10401 = n10400 ^ n10323;
  assign n10313 = n1903 & n5010;
  assign n10314 = x85 & n5223;
  assign n10315 = x86 & n5014;
  assign n10316 = ~n10314 & ~n10315;
  assign n10317 = x87 & n5226;
  assign n10318 = n10316 & ~n10317;
  assign n10319 = ~n10313 & n10318;
  assign n10320 = n10319 ^ x44;
  assign n10402 = n10401 ^ n10320;
  assign n10310 = n10135 ^ n10045;
  assign n10311 = ~n10136 & ~n10310;
  assign n10312 = n10311 ^ n10045;
  assign n10403 = n10402 ^ n10312;
  assign n10302 = n2292 & n4415;
  assign n10303 = x88 & n4420;
  assign n10304 = x90 & n4614;
  assign n10305 = ~n10303 & ~n10304;
  assign n10306 = x89 & n4410;
  assign n10307 = n10305 & ~n10306;
  assign n10308 = ~n10302 & n10307;
  assign n10309 = n10308 ^ x41;
  assign n10404 = n10403 ^ n10309;
  assign n10299 = n10137 ^ n10034;
  assign n10300 = n10138 & n10299;
  assign n10301 = n10300 ^ n10034;
  assign n10405 = n10404 ^ n10301;
  assign n10291 = n2726 & n3829;
  assign n10292 = x91 & n4049;
  assign n10293 = x93 & n4052;
  assign n10294 = ~n10292 & ~n10293;
  assign n10295 = x92 & n3833;
  assign n10296 = n10294 & ~n10295;
  assign n10297 = ~n10291 & n10296;
  assign n10298 = n10297 ^ x38;
  assign n10406 = n10405 ^ n10298;
  assign n10288 = n10139 ^ n10023;
  assign n10289 = ~n10140 & ~n10288;
  assign n10290 = n10289 ^ n10023;
  assign n10407 = n10406 ^ n10290;
  assign n10280 = n3209 & n3330;
  assign n10281 = x94 & n3500;
  assign n10282 = x96 & n3502;
  assign n10283 = ~n10281 & ~n10282;
  assign n10284 = x95 & n3334;
  assign n10285 = n10283 & ~n10284;
  assign n10286 = ~n10280 & n10285;
  assign n10287 = n10286 ^ x35;
  assign n10408 = n10407 ^ n10287;
  assign n10277 = n10141 ^ n10012;
  assign n10278 = n10142 & n10277;
  assign n10279 = n10278 ^ n10012;
  assign n10409 = n10408 ^ n10279;
  assign n10269 = n2836 & n3730;
  assign n10270 = x97 & n2996;
  assign n10271 = x98 & n2840;
  assign n10272 = ~n10270 & ~n10271;
  assign n10273 = x99 & n2998;
  assign n10274 = n10272 & ~n10273;
  assign n10275 = ~n10269 & n10274;
  assign n10276 = n10275 ^ x32;
  assign n10410 = n10409 ^ n10276;
  assign n10266 = n10143 ^ n10001;
  assign n10267 = ~n10144 & n10266;
  assign n10268 = n10267 ^ n10001;
  assign n10411 = n10410 ^ n10268;
  assign n10258 = n2371 & n4286;
  assign n10259 = x101 & n2377;
  assign n10260 = x100 & n2528;
  assign n10261 = ~n10259 & ~n10260;
  assign n10262 = x102 & n2531;
  assign n10263 = n10261 & ~n10262;
  assign n10264 = ~n10258 & n10263;
  assign n10265 = n10264 ^ x29;
  assign n10412 = n10411 ^ n10265;
  assign n10255 = n10145 ^ n9990;
  assign n10256 = ~n10146 & n10255;
  assign n10257 = n10256 ^ n9990;
  assign n10413 = n10412 ^ n10257;
  assign n10247 = n1969 & n4867;
  assign n10248 = x103 & n1978;
  assign n10249 = x105 & n2108;
  assign n10250 = ~n10248 & ~n10249;
  assign n10251 = x104 & n1973;
  assign n10252 = n10250 & ~n10251;
  assign n10253 = ~n10247 & n10252;
  assign n10254 = n10253 ^ x26;
  assign n10414 = n10413 ^ n10254;
  assign n10244 = n10147 ^ n9979;
  assign n10245 = ~n10148 & ~n10244;
  assign n10246 = n10245 ^ n9979;
  assign n10415 = n10414 ^ n10246;
  assign n10236 = n1624 & ~n5506;
  assign n10237 = x106 & n1742;
  assign n10238 = x108 & n1744;
  assign n10239 = ~n10237 & ~n10238;
  assign n10240 = x107 & n1628;
  assign n10241 = n10239 & ~n10240;
  assign n10242 = ~n10236 & n10241;
  assign n10243 = n10242 ^ x23;
  assign n10416 = n10415 ^ n10243;
  assign n10233 = n10149 ^ n9968;
  assign n10234 = n10150 & n10233;
  assign n10235 = n10234 ^ n9968;
  assign n10417 = n10416 ^ n10235;
  assign n10225 = n1296 & n6178;
  assign n10226 = x109 & n1403;
  assign n10227 = x110 & n1300;
  assign n10228 = ~n10226 & ~n10227;
  assign n10229 = x111 & n1406;
  assign n10230 = n10228 & ~n10229;
  assign n10231 = ~n10225 & n10230;
  assign n10232 = n10231 ^ x20;
  assign n10418 = n10417 ^ n10232;
  assign n10222 = n10151 ^ n9957;
  assign n10223 = ~n10152 & ~n10222;
  assign n10224 = n10223 ^ n9957;
  assign n10419 = n10418 ^ n10224;
  assign n10214 = n1008 & n6892;
  assign n10215 = x113 & n1012;
  assign n10216 = x112 & n1101;
  assign n10217 = ~n10215 & ~n10216;
  assign n10218 = x114 & n1104;
  assign n10219 = n10217 & ~n10218;
  assign n10220 = ~n10214 & n10219;
  assign n10221 = n10220 ^ x17;
  assign n10420 = n10419 ^ n10221;
  assign n10211 = n10153 ^ n9946;
  assign n10212 = n10154 & n10211;
  assign n10213 = n10212 ^ n9946;
  assign n10421 = n10420 ^ n10213;
  assign n10203 = n752 & n7643;
  assign n10204 = x115 & n825;
  assign n10205 = x116 & n757;
  assign n10206 = ~n10204 & ~n10205;
  assign n10207 = x117 & n828;
  assign n10208 = n10206 & ~n10207;
  assign n10209 = ~n10203 & n10208;
  assign n10210 = n10209 ^ x14;
  assign n10422 = n10421 ^ n10210;
  assign n10200 = n10155 ^ n9935;
  assign n10201 = ~n10156 & ~n10200;
  assign n10202 = n10201 ^ n9935;
  assign n10423 = n10422 ^ n10202;
  assign n10191 = n372 & n9309;
  assign n10192 = x121 & n433;
  assign n10193 = x123 & n428;
  assign n10194 = ~n10192 & ~n10193;
  assign n10195 = x122 & n376;
  assign n10196 = n10194 & ~n10195;
  assign n10197 = ~n10191 & n10196;
  assign n10198 = n10197 ^ x8;
  assign n10183 = n541 & ~n8424;
  assign n10184 = x119 & n547;
  assign n10185 = x118 & n612;
  assign n10186 = ~n10184 & ~n10185;
  assign n10187 = x120 & n615;
  assign n10188 = n10186 & ~n10187;
  assign n10189 = ~n10183 & n10188;
  assign n10190 = n10189 ^ x11;
  assign n10199 = n10198 ^ n10190;
  assign n10424 = n10423 ^ n10199;
  assign n10174 = n9290 ^ x126;
  assign n10175 = n210 & ~n10174;
  assign n10176 = x124 & n219;
  assign n10177 = x125 & n214;
  assign n10178 = ~n10176 & ~n10177;
  assign n10179 = x126 & n259;
  assign n10180 = n10178 & ~n10179;
  assign n10181 = ~n10175 & n10180;
  assign n10182 = n10181 ^ x5;
  assign n10425 = n10424 ^ n10182;
  assign n10171 = n10157 ^ n9924;
  assign n10172 = n10158 & n10171;
  assign n10173 = n10172 ^ n9924;
  assign n10426 = n10425 ^ n10173;
  assign n10438 = n10437 ^ n10426;
  assign n10168 = n9902 ^ n9884;
  assign n10169 = n10161 & n10168;
  assign n10170 = n10169 ^ n10160;
  assign n10439 = n10438 ^ n10170;
  assign n10165 = n10162 ^ n9878;
  assign n10166 = ~n10163 & ~n10165;
  assign n10167 = n10166 ^ n9878;
  assign n10440 = n10439 ^ n10167;
  assign n10665 = ~n594 & n8622;
  assign n10666 = x72 & n8626;
  assign n10667 = x71 & n8631;
  assign n10668 = ~n10666 & ~n10667;
  assign n10669 = x73 & n9186;
  assign n10670 = n10668 & ~n10669;
  assign n10671 = ~n10665 & n10670;
  assign n10672 = n10671 ^ x59;
  assign n10657 = n416 & n9499;
  assign n10658 = x68 & n9508;
  assign n10659 = x70 & n10106;
  assign n10660 = ~n10658 & ~n10659;
  assign n10661 = x69 & n9503;
  assign n10662 = n10660 & ~n10661;
  assign n10663 = ~n10657 & n10662;
  assign n10652 = x63 & x67;
  assign n10649 = x67 ^ x66;
  assign n10650 = ~x63 & n10649;
  assign n10651 = n10650 ^ x66;
  assign n10653 = n10652 ^ n10651;
  assign n10654 = ~x62 & ~n10653;
  assign n10655 = n10654 ^ n10651;
  assign n10656 = n10655 ^ x2;
  assign n10664 = n10663 ^ n10656;
  assign n10673 = n10672 ^ n10664;
  assign n10646 = n10367 ^ n10361;
  assign n10647 = n10368 & ~n10646;
  assign n10648 = n10647 ^ n10364;
  assign n10674 = n10673 ^ n10648;
  assign n10638 = n799 & n7830;
  assign n10639 = x74 & n7839;
  assign n10640 = x75 & n7834;
  assign n10641 = ~n10639 & ~n10640;
  assign n10642 = x76 & n8374;
  assign n10643 = n10641 & ~n10642;
  assign n10644 = ~n10638 & n10643;
  assign n10645 = n10644 ^ x56;
  assign n10675 = n10674 ^ n10645;
  assign n10635 = n10369 ^ n10345;
  assign n10636 = ~n10370 & n10635;
  assign n10637 = n10636 ^ n10345;
  assign n10676 = n10675 ^ n10637;
  assign n10627 = n1054 & n7076;
  assign n10628 = x78 & n7080;
  assign n10629 = x77 & n7317;
  assign n10630 = ~n10628 & ~n10629;
  assign n10631 = x79 & n7319;
  assign n10632 = n10630 & ~n10631;
  assign n10633 = ~n10627 & n10632;
  assign n10634 = n10633 ^ x53;
  assign n10677 = n10676 ^ n10634;
  assign n10624 = n10382 ^ n10371;
  assign n10625 = ~n10383 & ~n10624;
  assign n10626 = n10625 ^ n10374;
  assign n10678 = n10677 ^ n10626;
  assign n10616 = n1345 & n6326;
  assign n10617 = x80 & n6565;
  assign n10618 = x81 & n6331;
  assign n10619 = ~n10617 & ~n10618;
  assign n10620 = x82 & n6569;
  assign n10621 = n10619 & ~n10620;
  assign n10622 = ~n10616 & n10621;
  assign n10623 = n10622 ^ x50;
  assign n10679 = n10678 ^ n10623;
  assign n10613 = n10395 ^ n10384;
  assign n10614 = ~n10396 & n10613;
  assign n10615 = n10614 ^ n10387;
  assign n10680 = n10679 ^ n10615;
  assign n10605 = n1674 & n5656;
  assign n10606 = x83 & n5895;
  assign n10607 = x85 & n6111;
  assign n10608 = ~n10606 & ~n10607;
  assign n10609 = x84 & n5662;
  assign n10610 = n10608 & ~n10609;
  assign n10611 = ~n10605 & n10610;
  assign n10612 = n10611 ^ x47;
  assign n10681 = n10680 ^ n10612;
  assign n10602 = n10397 ^ n10334;
  assign n10603 = ~n10398 & ~n10602;
  assign n10604 = n10603 ^ n10334;
  assign n10682 = n10681 ^ n10604;
  assign n10594 = n2040 & n5010;
  assign n10595 = x86 & n5223;
  assign n10596 = x88 & n5226;
  assign n10597 = ~n10595 & ~n10596;
  assign n10598 = x87 & n5014;
  assign n10599 = n10597 & ~n10598;
  assign n10600 = ~n10594 & n10599;
  assign n10601 = n10600 ^ x44;
  assign n10683 = n10682 ^ n10601;
  assign n10591 = n10399 ^ n10323;
  assign n10592 = n10400 & n10591;
  assign n10593 = n10592 ^ n10323;
  assign n10684 = n10683 ^ n10593;
  assign n10583 = n2447 & n4415;
  assign n10584 = x89 & n4420;
  assign n10585 = x90 & n4410;
  assign n10586 = ~n10584 & ~n10585;
  assign n10587 = x91 & n4614;
  assign n10588 = n10586 & ~n10587;
  assign n10589 = ~n10583 & n10588;
  assign n10590 = n10589 ^ x41;
  assign n10685 = n10684 ^ n10590;
  assign n10580 = n10401 ^ n10312;
  assign n10581 = ~n10402 & ~n10580;
  assign n10582 = n10581 ^ n10312;
  assign n10686 = n10685 ^ n10582;
  assign n10572 = n2895 & n3829;
  assign n10573 = x93 & n3833;
  assign n10574 = x92 & n4049;
  assign n10575 = ~n10573 & ~n10574;
  assign n10576 = x94 & n4052;
  assign n10577 = n10575 & ~n10576;
  assign n10578 = ~n10572 & n10577;
  assign n10579 = n10578 ^ x38;
  assign n10687 = n10686 ^ n10579;
  assign n10569 = n10403 ^ n10301;
  assign n10570 = n10404 & n10569;
  assign n10571 = n10570 ^ n10301;
  assign n10688 = n10687 ^ n10571;
  assign n10561 = n3330 & n3388;
  assign n10562 = x95 & n3500;
  assign n10563 = x96 & n3334;
  assign n10564 = ~n10562 & ~n10563;
  assign n10565 = x97 & n3502;
  assign n10566 = n10564 & ~n10565;
  assign n10567 = ~n10561 & n10566;
  assign n10568 = n10567 ^ x35;
  assign n10689 = n10688 ^ n10568;
  assign n10558 = n10405 ^ n10290;
  assign n10559 = ~n10406 & ~n10558;
  assign n10560 = n10559 ^ n10290;
  assign n10690 = n10689 ^ n10560;
  assign n10550 = n2836 & n3925;
  assign n10551 = x99 & n2840;
  assign n10552 = x98 & n2996;
  assign n10553 = ~n10551 & ~n10552;
  assign n10554 = x100 & n2998;
  assign n10555 = n10553 & ~n10554;
  assign n10556 = ~n10550 & n10555;
  assign n10557 = n10556 ^ x32;
  assign n10691 = n10690 ^ n10557;
  assign n10547 = n10407 ^ n10279;
  assign n10548 = n10408 & n10547;
  assign n10549 = n10548 ^ n10279;
  assign n10692 = n10691 ^ n10549;
  assign n10539 = n2371 & n4481;
  assign n10540 = x101 & n2528;
  assign n10541 = x103 & n2531;
  assign n10542 = ~n10540 & ~n10541;
  assign n10543 = x102 & n2377;
  assign n10544 = n10542 & ~n10543;
  assign n10545 = ~n10539 & n10544;
  assign n10546 = n10545 ^ x29;
  assign n10693 = n10692 ^ n10546;
  assign n10536 = n10409 ^ n10268;
  assign n10537 = ~n10410 & n10536;
  assign n10538 = n10537 ^ n10268;
  assign n10694 = n10693 ^ n10538;
  assign n10528 = n1969 & n5088;
  assign n10529 = x104 & n1978;
  assign n10530 = x106 & n2108;
  assign n10531 = ~n10529 & ~n10530;
  assign n10532 = x105 & n1973;
  assign n10533 = n10531 & ~n10532;
  assign n10534 = ~n10528 & n10533;
  assign n10535 = n10534 ^ x26;
  assign n10695 = n10694 ^ n10535;
  assign n10525 = n10411 ^ n10257;
  assign n10526 = ~n10412 & n10525;
  assign n10527 = n10526 ^ n10257;
  assign n10696 = n10695 ^ n10527;
  assign n10517 = n1624 & ~n5737;
  assign n10518 = x107 & n1742;
  assign n10519 = x108 & n1628;
  assign n10520 = ~n10518 & ~n10519;
  assign n10521 = x109 & n1744;
  assign n10522 = n10520 & ~n10521;
  assign n10523 = ~n10517 & n10522;
  assign n10524 = n10523 ^ x23;
  assign n10697 = n10696 ^ n10524;
  assign n10514 = n10413 ^ n10246;
  assign n10515 = ~n10414 & ~n10514;
  assign n10516 = n10515 ^ n10246;
  assign n10698 = n10697 ^ n10516;
  assign n10506 = n1296 & n6420;
  assign n10507 = x110 & n1403;
  assign n10508 = x111 & n1300;
  assign n10509 = ~n10507 & ~n10508;
  assign n10510 = x112 & n1406;
  assign n10511 = n10509 & ~n10510;
  assign n10512 = ~n10506 & n10511;
  assign n10513 = n10512 ^ x20;
  assign n10699 = n10698 ^ n10513;
  assign n10503 = n10415 ^ n10235;
  assign n10504 = n10416 & n10503;
  assign n10505 = n10504 ^ n10235;
  assign n10700 = n10699 ^ n10505;
  assign n10495 = n1008 & n7150;
  assign n10496 = x114 & n1012;
  assign n10497 = x113 & n1101;
  assign n10498 = ~n10496 & ~n10497;
  assign n10499 = x115 & n1104;
  assign n10500 = n10498 & ~n10499;
  assign n10501 = ~n10495 & n10500;
  assign n10502 = n10501 ^ x17;
  assign n10701 = n10700 ^ n10502;
  assign n10492 = n10417 ^ n10224;
  assign n10493 = ~n10418 & ~n10492;
  assign n10494 = n10493 ^ n10224;
  assign n10702 = n10701 ^ n10494;
  assign n10484 = n752 & n7919;
  assign n10485 = x116 & n825;
  assign n10486 = x117 & n757;
  assign n10487 = ~n10485 & ~n10486;
  assign n10488 = x118 & n828;
  assign n10489 = n10487 & ~n10488;
  assign n10490 = ~n10484 & n10489;
  assign n10491 = n10490 ^ x14;
  assign n10703 = n10702 ^ n10491;
  assign n10481 = n10419 ^ n10213;
  assign n10482 = n10420 & n10481;
  assign n10483 = n10482 ^ n10213;
  assign n10704 = n10703 ^ n10483;
  assign n10473 = n541 & n8715;
  assign n10474 = x119 & n612;
  assign n10475 = x121 & n615;
  assign n10476 = ~n10474 & ~n10475;
  assign n10477 = x120 & n547;
  assign n10478 = n10476 & ~n10477;
  assign n10479 = ~n10473 & n10478;
  assign n10480 = n10479 ^ x11;
  assign n10705 = n10704 ^ n10480;
  assign n10470 = n10421 ^ n10202;
  assign n10471 = ~n10422 & ~n10470;
  assign n10472 = n10471 ^ n10202;
  assign n10706 = n10705 ^ n10472;
  assign n10467 = n10423 ^ n10198;
  assign n10468 = ~n10199 & ~n10467;
  assign n10469 = n10468 ^ n10423;
  assign n10707 = n10706 ^ n10469;
  assign n10459 = n372 & n9614;
  assign n10460 = x122 & n433;
  assign n10461 = x124 & n428;
  assign n10462 = ~n10460 & ~n10461;
  assign n10463 = x123 & n376;
  assign n10464 = n10462 & ~n10463;
  assign n10465 = ~n10459 & n10464;
  assign n10466 = n10465 ^ x8;
  assign n10708 = n10707 ^ n10466;
  assign n10456 = n10424 ^ n10173;
  assign n10457 = n10425 & n10456;
  assign n10458 = n10457 ^ n10173;
  assign n10709 = n10708 ^ n10458;
  assign n10447 = n9599 ^ x127;
  assign n10448 = n210 & ~n10447;
  assign n10449 = x125 & n219;
  assign n10450 = x127 & n259;
  assign n10451 = ~n10449 & ~n10450;
  assign n10452 = x126 & n214;
  assign n10453 = n10451 & ~n10452;
  assign n10454 = ~n10448 & n10453;
  assign n10455 = n10454 ^ x5;
  assign n10710 = n10709 ^ n10455;
  assign n10444 = n10436 ^ n10426;
  assign n10445 = ~n10437 & n10444;
  assign n10446 = n10445 ^ n10429;
  assign n10711 = n10710 ^ n10446;
  assign n10441 = n10438 ^ n10167;
  assign n10442 = n10439 & ~n10441;
  assign n10443 = n10442 ^ n10167;
  assign n10712 = n10711 ^ n10443;
  assign n10948 = n1445 & n6326;
  assign n10949 = x81 & n6565;
  assign n10950 = x83 & n6569;
  assign n10951 = ~n10949 & ~n10950;
  assign n10952 = x82 & n6331;
  assign n10953 = n10951 & ~n10952;
  assign n10954 = ~n10948 & n10953;
  assign n10955 = n10954 ^ x50;
  assign n10945 = n10676 ^ n10626;
  assign n10946 = n10677 & n10945;
  assign n10947 = n10946 ^ n10626;
  assign n10956 = n10955 ^ n10947;
  assign n10935 = ~n1141 & n7076;
  assign n10936 = x79 & n7080;
  assign n10937 = x80 & n7319;
  assign n10938 = ~n10936 & ~n10937;
  assign n10939 = x78 & n7317;
  assign n10940 = n10938 & ~n10939;
  assign n10941 = ~n10935 & n10940;
  assign n10942 = n10941 ^ x53;
  assign n10925 = n877 & n7830;
  assign n10926 = x75 & n7839;
  assign n10927 = x77 & n8374;
  assign n10928 = ~n10926 & ~n10927;
  assign n10929 = x76 & n7834;
  assign n10930 = n10928 & ~n10929;
  assign n10931 = ~n10925 & n10930;
  assign n10932 = n10931 ^ x56;
  assign n10912 = ~x2 & ~n10663;
  assign n10913 = n10651 & ~n10912;
  assign n10914 = x2 & n10663;
  assign n10915 = x62 & ~n10914;
  assign n10916 = ~n10913 & n10915;
  assign n10917 = ~x2 & ~n10652;
  assign n10918 = ~n10663 & ~n10917;
  assign n10919 = x2 & n10652;
  assign n10920 = ~x62 & ~n10919;
  assign n10921 = ~n10918 & n10920;
  assign n10922 = ~n10916 & ~n10921;
  assign n10904 = n467 & n9499;
  assign n10905 = x69 & n9508;
  assign n10906 = x71 & n10106;
  assign n10907 = ~n10905 & ~n10906;
  assign n10908 = x70 & n9503;
  assign n10909 = n10907 & ~n10908;
  assign n10910 = ~n10904 & n10909;
  assign n10899 = x63 & x68;
  assign n10896 = x68 ^ x67;
  assign n10897 = ~x63 & n10896;
  assign n10898 = n10897 ^ x67;
  assign n10900 = n10899 ^ n10898;
  assign n10901 = ~x62 & ~n10900;
  assign n10902 = n10901 ^ n10898;
  assign n10903 = n10902 ^ x2;
  assign n10911 = n10910 ^ n10903;
  assign n10923 = n10922 ^ n10911;
  assign n10888 = ~n656 & n8622;
  assign n10889 = x73 & n8626;
  assign n10890 = x72 & n8631;
  assign n10891 = ~n10889 & ~n10890;
  assign n10892 = x74 & n9186;
  assign n10893 = n10891 & ~n10892;
  assign n10894 = ~n10888 & n10893;
  assign n10895 = n10894 ^ x59;
  assign n10924 = n10923 ^ n10895;
  assign n10933 = n10932 ^ n10924;
  assign n10885 = n10672 ^ n10648;
  assign n10886 = n10673 & n10885;
  assign n10887 = n10886 ^ n10648;
  assign n10934 = n10933 ^ n10887;
  assign n10943 = n10942 ^ n10934;
  assign n10882 = n10674 ^ n10637;
  assign n10883 = n10675 & ~n10882;
  assign n10884 = n10883 ^ n10637;
  assign n10944 = n10943 ^ n10884;
  assign n10957 = n10956 ^ n10944;
  assign n10874 = n1787 & n5656;
  assign n10875 = x84 & n5895;
  assign n10876 = x86 & n6111;
  assign n10877 = ~n10875 & ~n10876;
  assign n10878 = x85 & n5662;
  assign n10879 = n10877 & ~n10878;
  assign n10880 = ~n10874 & n10879;
  assign n10881 = n10880 ^ x47;
  assign n10958 = n10957 ^ n10881;
  assign n10871 = n10678 ^ n10615;
  assign n10872 = ~n10679 & ~n10871;
  assign n10873 = n10872 ^ n10615;
  assign n10959 = n10958 ^ n10873;
  assign n10863 = n2164 & n5010;
  assign n10864 = x87 & n5223;
  assign n10865 = x88 & n5014;
  assign n10866 = ~n10864 & ~n10865;
  assign n10867 = x89 & n5226;
  assign n10868 = n10866 & ~n10867;
  assign n10869 = ~n10863 & n10868;
  assign n10870 = n10869 ^ x44;
  assign n10960 = n10959 ^ n10870;
  assign n10860 = n10680 ^ n10604;
  assign n10861 = n10681 & n10860;
  assign n10862 = n10861 ^ n10604;
  assign n10961 = n10960 ^ n10862;
  assign n10852 = n2585 & n4415;
  assign n10853 = x90 & n4420;
  assign n10854 = x91 & n4410;
  assign n10855 = ~n10853 & ~n10854;
  assign n10856 = x92 & n4614;
  assign n10857 = n10855 & ~n10856;
  assign n10858 = ~n10852 & n10857;
  assign n10859 = n10858 ^ x41;
  assign n10962 = n10961 ^ n10859;
  assign n10849 = n10682 ^ n10593;
  assign n10850 = ~n10683 & ~n10849;
  assign n10851 = n10850 ^ n10593;
  assign n10963 = n10962 ^ n10851;
  assign n10841 = n3054 & n3829;
  assign n10842 = x93 & n4049;
  assign n10843 = x95 & n4052;
  assign n10844 = ~n10842 & ~n10843;
  assign n10845 = x94 & n3833;
  assign n10846 = n10844 & ~n10845;
  assign n10847 = ~n10841 & n10846;
  assign n10848 = n10847 ^ x38;
  assign n10964 = n10963 ^ n10848;
  assign n10838 = n10684 ^ n10582;
  assign n10839 = n10685 & n10838;
  assign n10840 = n10839 ^ n10582;
  assign n10965 = n10964 ^ n10840;
  assign n10830 = n3330 & n3556;
  assign n10831 = x96 & n3500;
  assign n10832 = x97 & n3334;
  assign n10833 = ~n10831 & ~n10832;
  assign n10834 = x98 & n3502;
  assign n10835 = n10833 & ~n10834;
  assign n10836 = ~n10830 & n10835;
  assign n10837 = n10836 ^ x35;
  assign n10966 = n10965 ^ n10837;
  assign n10827 = n10686 ^ n10571;
  assign n10828 = ~n10687 & ~n10827;
  assign n10829 = n10828 ^ n10571;
  assign n10967 = n10966 ^ n10829;
  assign n10819 = n2836 & n4105;
  assign n10820 = x100 & n2840;
  assign n10821 = x99 & n2996;
  assign n10822 = ~n10820 & ~n10821;
  assign n10823 = x101 & n2998;
  assign n10824 = n10822 & ~n10823;
  assign n10825 = ~n10819 & n10824;
  assign n10826 = n10825 ^ x32;
  assign n10968 = n10967 ^ n10826;
  assign n10816 = n10688 ^ n10560;
  assign n10817 = n10689 & n10816;
  assign n10818 = n10817 ^ n10560;
  assign n10969 = n10968 ^ n10818;
  assign n10808 = n2371 & n4670;
  assign n10809 = x103 & n2377;
  assign n10810 = x102 & n2528;
  assign n10811 = ~n10809 & ~n10810;
  assign n10812 = x104 & n2531;
  assign n10813 = n10811 & ~n10812;
  assign n10814 = ~n10808 & n10813;
  assign n10815 = n10814 ^ x29;
  assign n10970 = n10969 ^ n10815;
  assign n10805 = n10690 ^ n10549;
  assign n10806 = ~n10691 & ~n10805;
  assign n10807 = n10806 ^ n10549;
  assign n10971 = n10970 ^ n10807;
  assign n10797 = n1969 & n5297;
  assign n10798 = x105 & n1978;
  assign n10799 = x106 & n1973;
  assign n10800 = ~n10798 & ~n10799;
  assign n10801 = x107 & n2108;
  assign n10802 = n10800 & ~n10801;
  assign n10803 = ~n10797 & n10802;
  assign n10804 = n10803 ^ x26;
  assign n10972 = n10971 ^ n10804;
  assign n10794 = n10692 ^ n10538;
  assign n10795 = n10693 & ~n10794;
  assign n10796 = n10795 ^ n10538;
  assign n10973 = n10972 ^ n10796;
  assign n10786 = n1624 & n5955;
  assign n10787 = x108 & n1742;
  assign n10788 = x109 & n1628;
  assign n10789 = ~n10787 & ~n10788;
  assign n10790 = x110 & n1744;
  assign n10791 = n10789 & ~n10790;
  assign n10792 = ~n10786 & n10791;
  assign n10793 = n10792 ^ x23;
  assign n10974 = n10973 ^ n10793;
  assign n10783 = n10694 ^ n10527;
  assign n10784 = n10695 & ~n10783;
  assign n10785 = n10784 ^ n10527;
  assign n10975 = n10974 ^ n10785;
  assign n10775 = n1296 & n6656;
  assign n10776 = x112 & n1300;
  assign n10777 = x111 & n1403;
  assign n10778 = ~n10776 & ~n10777;
  assign n10779 = x113 & n1406;
  assign n10780 = n10778 & ~n10779;
  assign n10781 = ~n10775 & n10780;
  assign n10782 = n10781 ^ x20;
  assign n10976 = n10975 ^ n10782;
  assign n10772 = n10696 ^ n10516;
  assign n10773 = n10697 & n10772;
  assign n10774 = n10773 ^ n10516;
  assign n10977 = n10976 ^ n10774;
  assign n10764 = n1008 & n7393;
  assign n10765 = x114 & n1101;
  assign n10766 = x115 & n1012;
  assign n10767 = ~n10765 & ~n10766;
  assign n10768 = x116 & n1104;
  assign n10769 = n10767 & ~n10768;
  assign n10770 = ~n10764 & n10769;
  assign n10771 = n10770 ^ x17;
  assign n10978 = n10977 ^ n10771;
  assign n10761 = n10698 ^ n10505;
  assign n10762 = ~n10699 & ~n10761;
  assign n10763 = n10762 ^ n10505;
  assign n10979 = n10978 ^ n10763;
  assign n10753 = n752 & n8169;
  assign n10754 = x117 & n825;
  assign n10755 = x119 & n828;
  assign n10756 = ~n10754 & ~n10755;
  assign n10757 = x118 & n757;
  assign n10758 = n10756 & ~n10757;
  assign n10759 = ~n10753 & n10758;
  assign n10760 = n10759 ^ x14;
  assign n10980 = n10979 ^ n10760;
  assign n10750 = n10700 ^ n10494;
  assign n10751 = n10701 & n10750;
  assign n10752 = n10751 ^ n10494;
  assign n10981 = n10980 ^ n10752;
  assign n10742 = n541 & n9001;
  assign n10743 = x120 & n612;
  assign n10744 = x121 & n547;
  assign n10745 = ~n10743 & ~n10744;
  assign n10746 = x122 & n615;
  assign n10747 = n10745 & ~n10746;
  assign n10748 = ~n10742 & n10747;
  assign n10749 = n10748 ^ x11;
  assign n10982 = n10981 ^ n10749;
  assign n10739 = n10702 ^ n10483;
  assign n10740 = ~n10703 & ~n10739;
  assign n10741 = n10740 ^ n10483;
  assign n10983 = n10982 ^ n10741;
  assign n10731 = n372 & n9912;
  assign n10732 = x123 & n433;
  assign n10733 = x124 & n376;
  assign n10734 = ~n10732 & ~n10733;
  assign n10735 = x125 & n428;
  assign n10736 = n10734 & ~n10735;
  assign n10737 = ~n10731 & n10736;
  assign n10738 = n10737 ^ x8;
  assign n10984 = n10983 ^ n10738;
  assign n10728 = n10704 ^ n10472;
  assign n10729 = n10705 & n10728;
  assign n10730 = n10729 ^ n10472;
  assign n10985 = n10984 ^ n10730;
  assign n10722 = n210 & ~n9889;
  assign n10723 = x127 & n214;
  assign n10724 = x126 & n219;
  assign n10725 = ~n10723 & ~n10724;
  assign n10726 = ~n10722 & n10725;
  assign n10727 = n10726 ^ x5;
  assign n10986 = n10985 ^ n10727;
  assign n10719 = n10706 ^ n10466;
  assign n10720 = ~n10707 & ~n10719;
  assign n10721 = n10720 ^ n10469;
  assign n10987 = n10986 ^ n10721;
  assign n10716 = n10708 ^ n10455;
  assign n10717 = n10709 & n10716;
  assign n10718 = n10717 ^ n10458;
  assign n10988 = n10987 ^ n10718;
  assign n10713 = n10710 ^ n10443;
  assign n10714 = ~n10711 & n10713;
  assign n10715 = n10714 ^ n10443;
  assign n10989 = n10988 ^ n10715;
  assign n11229 = n1547 & n6326;
  assign n11230 = x82 & n6565;
  assign n11231 = x83 & n6331;
  assign n11232 = ~n11230 & ~n11231;
  assign n11233 = x84 & n6569;
  assign n11234 = n11232 & ~n11233;
  assign n11235 = ~n11229 & n11234;
  assign n11236 = n11235 ^ x50;
  assign n11219 = n1230 & n7076;
  assign n11220 = x80 & n7080;
  assign n11221 = x79 & n7317;
  assign n11222 = ~n11220 & ~n11221;
  assign n11223 = x81 & n7319;
  assign n11224 = n11222 & ~n11223;
  assign n11225 = ~n11219 & n11224;
  assign n11226 = n11225 ^ x53;
  assign n11209 = n953 & n7830;
  assign n11210 = x76 & n7839;
  assign n11211 = x78 & n8374;
  assign n11212 = ~n11210 & ~n11211;
  assign n11213 = x77 & n7834;
  assign n11214 = n11212 & ~n11213;
  assign n11215 = ~n11209 & n11214;
  assign n11216 = n11215 ^ x56;
  assign n11206 = n10911 ^ n10895;
  assign n11207 = n10923 & n11206;
  assign n11208 = n11207 ^ n10922;
  assign n11217 = n11216 ^ n11208;
  assign n11196 = n720 & n8622;
  assign n11197 = x73 & n8631;
  assign n11198 = x74 & n8626;
  assign n11199 = ~n11197 & ~n11198;
  assign n11200 = x75 & n9186;
  assign n11201 = n11199 & ~n11200;
  assign n11202 = ~n11196 & n11201;
  assign n11203 = n11202 ^ x59;
  assign n11184 = ~x2 & ~n10910;
  assign n11185 = n10898 & ~n11184;
  assign n11186 = x2 & n10910;
  assign n11187 = x62 & ~n11186;
  assign n11188 = ~n11185 & n11187;
  assign n11189 = ~x2 & ~n10899;
  assign n11190 = ~n10910 & ~n11189;
  assign n11191 = ~x62 & n10899;
  assign n11192 = x2 & n11191;
  assign n11193 = n11192 ^ x62;
  assign n11194 = ~n11190 & ~n11193;
  assign n11195 = ~n11188 & ~n11194;
  assign n11204 = n11203 ^ n11195;
  assign n11176 = n520 & n9499;
  assign n11177 = x70 & n9508;
  assign n11178 = x72 & n10106;
  assign n11179 = ~n11177 & ~n11178;
  assign n11180 = x71 & n9503;
  assign n11181 = n11179 & ~n11180;
  assign n11182 = ~n11176 & n11181;
  assign n11171 = x63 & x69;
  assign n11168 = x69 ^ x68;
  assign n11169 = ~x63 & n11168;
  assign n11170 = n11169 ^ x68;
  assign n11172 = n11171 ^ n11170;
  assign n11173 = ~x62 & ~n11172;
  assign n11174 = n11173 ^ n11170;
  assign n11175 = n11174 ^ x2;
  assign n11183 = n11182 ^ n11175;
  assign n11205 = n11204 ^ n11183;
  assign n11218 = n11217 ^ n11205;
  assign n11227 = n11226 ^ n11218;
  assign n11165 = n10924 ^ n10887;
  assign n11166 = n10933 & ~n11165;
  assign n11167 = n11166 ^ n10932;
  assign n11228 = n11227 ^ n11167;
  assign n11237 = n11236 ^ n11228;
  assign n11162 = n10942 ^ n10884;
  assign n11163 = ~n10943 & n11162;
  assign n11164 = n11163 ^ n10884;
  assign n11238 = n11237 ^ n11164;
  assign n11159 = n10955 ^ n10944;
  assign n11160 = ~n10956 & ~n11159;
  assign n11161 = n11160 ^ n10947;
  assign n11239 = n11238 ^ n11161;
  assign n11151 = n1903 & n5656;
  assign n11152 = x85 & n5895;
  assign n11153 = x87 & n6111;
  assign n11154 = ~n11152 & ~n11153;
  assign n11155 = x86 & n5662;
  assign n11156 = n11154 & ~n11155;
  assign n11157 = ~n11151 & n11156;
  assign n11158 = n11157 ^ x47;
  assign n11240 = n11239 ^ n11158;
  assign n11143 = n2292 & n5010;
  assign n11144 = x88 & n5223;
  assign n11145 = x89 & n5014;
  assign n11146 = ~n11144 & ~n11145;
  assign n11147 = x90 & n5226;
  assign n11148 = n11146 & ~n11147;
  assign n11149 = ~n11143 & n11148;
  assign n11150 = n11149 ^ x44;
  assign n11241 = n11240 ^ n11150;
  assign n11140 = n10957 ^ n10873;
  assign n11141 = n10958 & n11140;
  assign n11142 = n11141 ^ n10873;
  assign n11242 = n11241 ^ n11142;
  assign n11132 = n2726 & n4415;
  assign n11133 = x91 & n4420;
  assign n11134 = x93 & n4614;
  assign n11135 = ~n11133 & ~n11134;
  assign n11136 = x92 & n4410;
  assign n11137 = n11135 & ~n11136;
  assign n11138 = ~n11132 & n11137;
  assign n11139 = n11138 ^ x41;
  assign n11243 = n11242 ^ n11139;
  assign n11129 = n10959 ^ n10862;
  assign n11130 = ~n10960 & ~n11129;
  assign n11131 = n11130 ^ n10862;
  assign n11244 = n11243 ^ n11131;
  assign n11121 = n3209 & n3829;
  assign n11122 = x94 & n4049;
  assign n11123 = x95 & n3833;
  assign n11124 = ~n11122 & ~n11123;
  assign n11125 = x96 & n4052;
  assign n11126 = n11124 & ~n11125;
  assign n11127 = ~n11121 & n11126;
  assign n11128 = n11127 ^ x38;
  assign n11245 = n11244 ^ n11128;
  assign n11118 = n10961 ^ n10851;
  assign n11119 = n10962 & n11118;
  assign n11120 = n11119 ^ n10851;
  assign n11246 = n11245 ^ n11120;
  assign n11110 = n3330 & n3730;
  assign n11111 = x97 & n3500;
  assign n11112 = x98 & n3334;
  assign n11113 = ~n11111 & ~n11112;
  assign n11114 = x99 & n3502;
  assign n11115 = n11113 & ~n11114;
  assign n11116 = ~n11110 & n11115;
  assign n11117 = n11116 ^ x35;
  assign n11247 = n11246 ^ n11117;
  assign n11107 = n10963 ^ n10840;
  assign n11108 = ~n10964 & ~n11107;
  assign n11109 = n11108 ^ n10840;
  assign n11248 = n11247 ^ n11109;
  assign n11099 = n2836 & n4286;
  assign n11100 = x100 & n2996;
  assign n11101 = x102 & n2998;
  assign n11102 = ~n11100 & ~n11101;
  assign n11103 = x101 & n2840;
  assign n11104 = n11102 & ~n11103;
  assign n11105 = ~n11099 & n11104;
  assign n11106 = n11105 ^ x32;
  assign n11249 = n11248 ^ n11106;
  assign n11096 = n10965 ^ n10829;
  assign n11097 = n10966 & n11096;
  assign n11098 = n11097 ^ n10829;
  assign n11250 = n11249 ^ n11098;
  assign n11088 = n2371 & n4867;
  assign n11089 = x103 & n2528;
  assign n11090 = x104 & n2377;
  assign n11091 = ~n11089 & ~n11090;
  assign n11092 = x105 & n2531;
  assign n11093 = n11091 & ~n11092;
  assign n11094 = ~n11088 & n11093;
  assign n11095 = n11094 ^ x29;
  assign n11251 = n11250 ^ n11095;
  assign n11085 = n10967 ^ n10818;
  assign n11086 = ~n10968 & ~n11085;
  assign n11087 = n11086 ^ n10818;
  assign n11252 = n11251 ^ n11087;
  assign n11077 = n1969 & ~n5506;
  assign n11078 = x106 & n1978;
  assign n11079 = x107 & n1973;
  assign n11080 = ~n11078 & ~n11079;
  assign n11081 = x108 & n2108;
  assign n11082 = n11080 & ~n11081;
  assign n11083 = ~n11077 & n11082;
  assign n11084 = n11083 ^ x26;
  assign n11253 = n11252 ^ n11084;
  assign n11074 = n10969 ^ n10807;
  assign n11075 = n10970 & n11074;
  assign n11076 = n11075 ^ n10807;
  assign n11254 = n11253 ^ n11076;
  assign n11066 = n1624 & n6178;
  assign n11067 = x109 & n1742;
  assign n11068 = x110 & n1628;
  assign n11069 = ~n11067 & ~n11068;
  assign n11070 = x111 & n1744;
  assign n11071 = n11069 & ~n11070;
  assign n11072 = ~n11066 & n11071;
  assign n11073 = n11072 ^ x23;
  assign n11255 = n11254 ^ n11073;
  assign n11063 = n10971 ^ n10796;
  assign n11064 = ~n10972 & n11063;
  assign n11065 = n11064 ^ n10796;
  assign n11256 = n11255 ^ n11065;
  assign n11055 = n1296 & n6892;
  assign n11056 = x112 & n1403;
  assign n11057 = x113 & n1300;
  assign n11058 = ~n11056 & ~n11057;
  assign n11059 = x114 & n1406;
  assign n11060 = n11058 & ~n11059;
  assign n11061 = ~n11055 & n11060;
  assign n11062 = n11061 ^ x20;
  assign n11257 = n11256 ^ n11062;
  assign n11052 = n10973 ^ n10785;
  assign n11053 = ~n10974 & n11052;
  assign n11054 = n11053 ^ n10785;
  assign n11258 = n11257 ^ n11054;
  assign n11044 = n1008 & n7643;
  assign n11045 = x115 & n1101;
  assign n11046 = x116 & n1012;
  assign n11047 = ~n11045 & ~n11046;
  assign n11048 = x117 & n1104;
  assign n11049 = n11047 & ~n11048;
  assign n11050 = ~n11044 & n11049;
  assign n11051 = n11050 ^ x17;
  assign n11259 = n11258 ^ n11051;
  assign n11041 = n10975 ^ n10774;
  assign n11042 = ~n10976 & ~n11041;
  assign n11043 = n11042 ^ n10774;
  assign n11260 = n11259 ^ n11043;
  assign n11033 = n752 & ~n8424;
  assign n11034 = x118 & n825;
  assign n11035 = x120 & n828;
  assign n11036 = ~n11034 & ~n11035;
  assign n11037 = x119 & n757;
  assign n11038 = n11036 & ~n11037;
  assign n11039 = ~n11033 & n11038;
  assign n11040 = n11039 ^ x14;
  assign n11261 = n11260 ^ n11040;
  assign n11030 = n10977 ^ n10763;
  assign n11031 = n10978 & n11030;
  assign n11032 = n11031 ^ n10763;
  assign n11262 = n11261 ^ n11032;
  assign n11022 = n541 & n9309;
  assign n11023 = x121 & n612;
  assign n11024 = x122 & n547;
  assign n11025 = ~n11023 & ~n11024;
  assign n11026 = x123 & n615;
  assign n11027 = n11025 & ~n11026;
  assign n11028 = ~n11022 & n11027;
  assign n11029 = n11028 ^ x11;
  assign n11263 = n11262 ^ n11029;
  assign n11019 = n10979 ^ n10752;
  assign n11020 = ~n10980 & ~n11019;
  assign n11021 = n11020 ^ n10752;
  assign n11264 = n11263 ^ n11021;
  assign n11011 = n372 & ~n10174;
  assign n11012 = x124 & n433;
  assign n11013 = x125 & n376;
  assign n11014 = ~n11012 & ~n11013;
  assign n11015 = x126 & n428;
  assign n11016 = n11014 & ~n11015;
  assign n11017 = ~n11011 & n11016;
  assign n11018 = n11017 ^ x8;
  assign n11265 = n11264 ^ n11018;
  assign n11008 = n10981 ^ n10741;
  assign n11009 = n10982 & n11008;
  assign n11010 = n11009 ^ n10741;
  assign n11266 = n11265 ^ n11010;
  assign n10999 = n172 & n10430;
  assign n11000 = x127 & n198;
  assign n11001 = x5 & ~n11000;
  assign n11002 = ~n10999 & n11001;
  assign n11003 = ~x4 & ~n11002;
  assign n11004 = x127 & n203;
  assign n11005 = ~x5 & ~n11004;
  assign n11006 = ~n10999 & n11005;
  assign n11007 = ~n11003 & ~n11006;
  assign n11267 = n11266 ^ n11007;
  assign n10996 = n10983 ^ n10730;
  assign n10997 = ~n10984 & ~n10996;
  assign n10998 = n10997 ^ n10730;
  assign n11268 = n11267 ^ n10998;
  assign n10993 = n10985 ^ n10721;
  assign n10994 = n10986 & n10993;
  assign n10995 = n10994 ^ n10721;
  assign n11269 = n11268 ^ n10995;
  assign n10990 = n10718 ^ n10715;
  assign n10991 = n10988 & ~n10990;
  assign n10992 = n10991 ^ n10715;
  assign n11270 = n11269 ^ n10992;
  assign n11531 = n10995 & n11266;
  assign n11532 = ~n10998 & ~n11007;
  assign n11538 = ~n11531 & n11532;
  assign n11534 = ~n10995 & ~n11266;
  assign n11535 = n10998 & n11007;
  assign n11539 = n11534 & ~n11535;
  assign n11540 = ~n11538 & ~n11539;
  assign n11533 = n11531 & ~n11532;
  assign n11536 = ~n11534 & n11535;
  assign n11537 = ~n11533 & ~n11536;
  assign n11541 = n11540 ^ n11537;
  assign n11542 = ~n10992 & n11541;
  assign n11543 = n11542 ^ n11540;
  assign n11544 = n10998 ^ n10995;
  assign n11545 = n11266 ^ n10998;
  assign n11546 = ~n11267 & ~n11545;
  assign n11547 = ~n11544 & n11546;
  assign n11548 = n11543 & ~n11547;
  assign n11489 = n1054 & n7830;
  assign n11490 = x77 & n7839;
  assign n11491 = x78 & n7834;
  assign n11492 = ~n11490 & ~n11491;
  assign n11493 = x79 & n8374;
  assign n11494 = n11492 & ~n11493;
  assign n11495 = ~n11489 & n11494;
  assign n11496 = n11495 ^ x56;
  assign n11486 = n11208 ^ n11205;
  assign n11487 = ~n11217 & n11486;
  assign n11488 = n11487 ^ n11216;
  assign n11497 = n11496 ^ n11488;
  assign n11471 = x2 & n11182;
  assign n11472 = ~n11170 & ~n11471;
  assign n11473 = ~x2 & ~n11182;
  assign n11474 = x62 & ~n11473;
  assign n11475 = ~n11472 & n11474;
  assign n11476 = x2 & n11171;
  assign n11477 = n11182 & ~n11476;
  assign n11478 = ~x2 & ~n11171;
  assign n11479 = ~x62 & ~n11478;
  assign n11480 = ~n11477 & n11479;
  assign n11481 = ~n11475 & ~n11480;
  assign n11467 = x70 & n9798;
  assign n11468 = x69 & n10099;
  assign n11469 = ~n11467 & ~n11468;
  assign n11466 = x5 ^ x2;
  assign n11470 = n11469 ^ n11466;
  assign n11482 = n11481 ^ n11470;
  assign n11458 = ~n594 & n9499;
  assign n11459 = x71 & n9508;
  assign n11460 = x73 & n10106;
  assign n11461 = ~n11459 & ~n11460;
  assign n11462 = x72 & n9503;
  assign n11463 = n11461 & ~n11462;
  assign n11464 = ~n11458 & n11463;
  assign n11465 = n11464 ^ x62;
  assign n11483 = n11482 ^ n11465;
  assign n11450 = n799 & n8622;
  assign n11451 = x74 & n8631;
  assign n11452 = x75 & n8626;
  assign n11453 = ~n11451 & ~n11452;
  assign n11454 = x76 & n9186;
  assign n11455 = n11453 & ~n11454;
  assign n11456 = ~n11450 & n11455;
  assign n11457 = n11456 ^ x59;
  assign n11484 = n11483 ^ n11457;
  assign n11447 = n11195 ^ n11183;
  assign n11448 = ~n11204 & ~n11447;
  assign n11449 = n11448 ^ n11203;
  assign n11485 = n11484 ^ n11449;
  assign n11498 = n11497 ^ n11485;
  assign n11439 = n1345 & n7076;
  assign n11440 = x80 & n7317;
  assign n11441 = x81 & n7080;
  assign n11442 = ~n11440 & ~n11441;
  assign n11443 = x82 & n7319;
  assign n11444 = n11442 & ~n11443;
  assign n11445 = ~n11439 & n11444;
  assign n11446 = n11445 ^ x53;
  assign n11499 = n11498 ^ n11446;
  assign n11436 = n11218 ^ n11167;
  assign n11437 = ~n11227 & n11436;
  assign n11438 = n11437 ^ n11226;
  assign n11500 = n11499 ^ n11438;
  assign n11428 = n1674 & n6326;
  assign n11429 = x83 & n6565;
  assign n11430 = x85 & n6569;
  assign n11431 = ~n11429 & ~n11430;
  assign n11432 = x84 & n6331;
  assign n11433 = n11431 & ~n11432;
  assign n11434 = ~n11428 & n11433;
  assign n11435 = n11434 ^ x50;
  assign n11501 = n11500 ^ n11435;
  assign n11425 = n11236 ^ n11164;
  assign n11426 = n11237 & n11425;
  assign n11427 = n11426 ^ n11164;
  assign n11502 = n11501 ^ n11427;
  assign n11422 = n11238 ^ n11158;
  assign n11423 = n11239 & n11422;
  assign n11424 = n11423 ^ n11161;
  assign n11503 = n11502 ^ n11424;
  assign n11414 = n2040 & n5656;
  assign n11415 = x86 & n5895;
  assign n11416 = x88 & n6111;
  assign n11417 = ~n11415 & ~n11416;
  assign n11418 = x87 & n5662;
  assign n11419 = n11417 & ~n11418;
  assign n11420 = ~n11414 & n11419;
  assign n11421 = n11420 ^ x47;
  assign n11504 = n11503 ^ n11421;
  assign n11406 = n2447 & n5010;
  assign n11407 = x89 & n5223;
  assign n11408 = x91 & n5226;
  assign n11409 = ~n11407 & ~n11408;
  assign n11410 = x90 & n5014;
  assign n11411 = n11409 & ~n11410;
  assign n11412 = ~n11406 & n11411;
  assign n11413 = n11412 ^ x44;
  assign n11505 = n11504 ^ n11413;
  assign n11403 = n11240 ^ n11142;
  assign n11404 = ~n11241 & ~n11403;
  assign n11405 = n11404 ^ n11142;
  assign n11506 = n11505 ^ n11405;
  assign n11395 = n2895 & n4415;
  assign n11396 = x92 & n4420;
  assign n11397 = x93 & n4410;
  assign n11398 = ~n11396 & ~n11397;
  assign n11399 = x94 & n4614;
  assign n11400 = n11398 & ~n11399;
  assign n11401 = ~n11395 & n11400;
  assign n11402 = n11401 ^ x41;
  assign n11507 = n11506 ^ n11402;
  assign n11392 = n11242 ^ n11131;
  assign n11393 = n11243 & n11392;
  assign n11394 = n11393 ^ n11131;
  assign n11508 = n11507 ^ n11394;
  assign n11384 = n3388 & n3829;
  assign n11385 = x95 & n4049;
  assign n11386 = x97 & n4052;
  assign n11387 = ~n11385 & ~n11386;
  assign n11388 = x96 & n3833;
  assign n11389 = n11387 & ~n11388;
  assign n11390 = ~n11384 & n11389;
  assign n11391 = n11390 ^ x38;
  assign n11509 = n11508 ^ n11391;
  assign n11381 = n11244 ^ n11120;
  assign n11382 = ~n11245 & ~n11381;
  assign n11383 = n11382 ^ n11120;
  assign n11510 = n11509 ^ n11383;
  assign n11373 = n3330 & n3925;
  assign n11374 = x98 & n3500;
  assign n11375 = x99 & n3334;
  assign n11376 = ~n11374 & ~n11375;
  assign n11377 = x100 & n3502;
  assign n11378 = n11376 & ~n11377;
  assign n11379 = ~n11373 & n11378;
  assign n11380 = n11379 ^ x35;
  assign n11511 = n11510 ^ n11380;
  assign n11370 = n11246 ^ n11109;
  assign n11371 = n11247 & n11370;
  assign n11372 = n11371 ^ n11109;
  assign n11512 = n11511 ^ n11372;
  assign n11362 = n2836 & n4481;
  assign n11363 = x101 & n2996;
  assign n11364 = x102 & n2840;
  assign n11365 = ~n11363 & ~n11364;
  assign n11366 = x103 & n2998;
  assign n11367 = n11365 & ~n11366;
  assign n11368 = ~n11362 & n11367;
  assign n11369 = n11368 ^ x32;
  assign n11513 = n11512 ^ n11369;
  assign n11359 = n11248 ^ n11098;
  assign n11360 = ~n11249 & ~n11359;
  assign n11361 = n11360 ^ n11098;
  assign n11514 = n11513 ^ n11361;
  assign n11351 = n2371 & n5088;
  assign n11352 = x104 & n2528;
  assign n11353 = x105 & n2377;
  assign n11354 = ~n11352 & ~n11353;
  assign n11355 = x106 & n2531;
  assign n11356 = n11354 & ~n11355;
  assign n11357 = ~n11351 & n11356;
  assign n11358 = n11357 ^ x29;
  assign n11515 = n11514 ^ n11358;
  assign n11348 = n11250 ^ n11087;
  assign n11349 = n11251 & n11348;
  assign n11350 = n11349 ^ n11087;
  assign n11516 = n11515 ^ n11350;
  assign n11340 = n1969 & ~n5737;
  assign n11341 = x107 & n1978;
  assign n11342 = x108 & n1973;
  assign n11343 = ~n11341 & ~n11342;
  assign n11344 = x109 & n2108;
  assign n11345 = n11343 & ~n11344;
  assign n11346 = ~n11340 & n11345;
  assign n11347 = n11346 ^ x26;
  assign n11517 = n11516 ^ n11347;
  assign n11337 = n11252 ^ n11076;
  assign n11338 = ~n11253 & ~n11337;
  assign n11339 = n11338 ^ n11076;
  assign n11518 = n11517 ^ n11339;
  assign n11329 = n1624 & n6420;
  assign n11330 = x111 & n1628;
  assign n11331 = x110 & n1742;
  assign n11332 = ~n11330 & ~n11331;
  assign n11333 = x112 & n1744;
  assign n11334 = n11332 & ~n11333;
  assign n11335 = ~n11329 & n11334;
  assign n11336 = n11335 ^ x23;
  assign n11519 = n11518 ^ n11336;
  assign n11326 = n11254 ^ n11065;
  assign n11327 = n11255 & ~n11326;
  assign n11328 = n11327 ^ n11065;
  assign n11520 = n11519 ^ n11328;
  assign n11318 = n1296 & n7150;
  assign n11319 = x113 & n1403;
  assign n11320 = x114 & n1300;
  assign n11321 = ~n11319 & ~n11320;
  assign n11322 = x115 & n1406;
  assign n11323 = n11321 & ~n11322;
  assign n11324 = ~n11318 & n11323;
  assign n11325 = n11324 ^ x20;
  assign n11521 = n11520 ^ n11325;
  assign n11315 = n11256 ^ n11054;
  assign n11316 = n11257 & ~n11315;
  assign n11317 = n11316 ^ n11054;
  assign n11522 = n11521 ^ n11317;
  assign n11307 = n1008 & n7919;
  assign n11308 = x116 & n1101;
  assign n11309 = x117 & n1012;
  assign n11310 = ~n11308 & ~n11309;
  assign n11311 = x118 & n1104;
  assign n11312 = n11310 & ~n11311;
  assign n11313 = ~n11307 & n11312;
  assign n11314 = n11313 ^ x17;
  assign n11523 = n11522 ^ n11314;
  assign n11304 = n11258 ^ n11043;
  assign n11305 = n11259 & n11304;
  assign n11306 = n11305 ^ n11043;
  assign n11524 = n11523 ^ n11306;
  assign n11296 = n752 & n8715;
  assign n11297 = x120 & n757;
  assign n11298 = x119 & n825;
  assign n11299 = ~n11297 & ~n11298;
  assign n11300 = x121 & n828;
  assign n11301 = n11299 & ~n11300;
  assign n11302 = ~n11296 & n11301;
  assign n11303 = n11302 ^ x14;
  assign n11525 = n11524 ^ n11303;
  assign n11293 = n11260 ^ n11032;
  assign n11294 = ~n11261 & ~n11293;
  assign n11295 = n11294 ^ n11032;
  assign n11526 = n11525 ^ n11295;
  assign n11285 = n541 & n9614;
  assign n11286 = x122 & n612;
  assign n11287 = x123 & n547;
  assign n11288 = ~n11286 & ~n11287;
  assign n11289 = x124 & n615;
  assign n11290 = n11288 & ~n11289;
  assign n11291 = ~n11285 & n11290;
  assign n11292 = n11291 ^ x11;
  assign n11527 = n11526 ^ n11292;
  assign n11282 = n11262 ^ n11021;
  assign n11283 = n11263 & n11282;
  assign n11284 = n11283 ^ n11021;
  assign n11528 = n11527 ^ n11284;
  assign n11274 = n372 & ~n10447;
  assign n11275 = x125 & n433;
  assign n11276 = x126 & n376;
  assign n11277 = ~n11275 & ~n11276;
  assign n11278 = x127 & n428;
  assign n11279 = n11277 & ~n11278;
  assign n11280 = ~n11274 & n11279;
  assign n11281 = n11280 ^ x8;
  assign n11529 = n11528 ^ n11281;
  assign n11271 = n11264 ^ n11010;
  assign n11272 = ~n11265 & ~n11271;
  assign n11273 = n11272 ^ n11010;
  assign n11530 = n11529 ^ n11273;
  assign n11549 = n11548 ^ n11530;
  assign n11802 = ~n11530 & ~n11534;
  assign n11803 = n10992 & ~n11802;
  assign n11804 = n11530 & ~n11531;
  assign n11805 = ~n11532 & ~n11804;
  assign n11806 = ~n11803 & n11805;
  assign n11807 = ~n11530 & n11535;
  assign n11808 = ~n11806 & ~n11807;
  assign n11809 = n10992 & ~n11531;
  assign n11810 = ~n11536 & ~n11802;
  assign n11811 = ~n11809 & ~n11810;
  assign n11812 = n11808 & ~n11811;
  assign n11767 = n2585 & n5010;
  assign n11768 = x90 & n5223;
  assign n11769 = x92 & n5226;
  assign n11770 = ~n11768 & ~n11769;
  assign n11771 = x91 & n5014;
  assign n11772 = n11770 & ~n11771;
  assign n11773 = ~n11767 & n11772;
  assign n11774 = n11773 ^ x44;
  assign n11757 = n2164 & n5656;
  assign n11758 = x87 & n5895;
  assign n11759 = x88 & n5662;
  assign n11760 = ~n11758 & ~n11759;
  assign n11761 = x89 & n6111;
  assign n11762 = n11760 & ~n11761;
  assign n11763 = ~n11757 & n11762;
  assign n11764 = n11763 ^ x47;
  assign n11747 = n1787 & n6326;
  assign n11748 = x84 & n6565;
  assign n11749 = x86 & n6569;
  assign n11750 = ~n11748 & ~n11749;
  assign n11751 = x85 & n6331;
  assign n11752 = n11750 & ~n11751;
  assign n11753 = ~n11747 & n11752;
  assign n11754 = n11753 ^ x50;
  assign n11737 = n1445 & n7076;
  assign n11738 = x81 & n7317;
  assign n11739 = x82 & n7080;
  assign n11740 = ~n11738 & ~n11739;
  assign n11741 = x83 & n7319;
  assign n11742 = n11740 & ~n11741;
  assign n11743 = ~n11737 & n11742;
  assign n11744 = n11743 ^ x53;
  assign n11725 = n877 & n8622;
  assign n11726 = x75 & n8631;
  assign n11727 = x77 & n9186;
  assign n11728 = ~n11726 & ~n11727;
  assign n11729 = x76 & n8626;
  assign n11730 = n11728 & ~n11729;
  assign n11731 = ~n11725 & n11730;
  assign n11732 = n11731 ^ x59;
  assign n11716 = ~n656 & n9499;
  assign n11717 = x73 & n9503;
  assign n11718 = x72 & n9508;
  assign n11719 = ~n11717 & ~n11718;
  assign n11720 = x74 & n10106;
  assign n11721 = n11719 & ~n11720;
  assign n11722 = ~n11716 & n11721;
  assign n11723 = n11722 ^ x62;
  assign n11712 = x71 & n9798;
  assign n11713 = x70 & n10099;
  assign n11714 = ~n11712 & ~n11713;
  assign n11709 = n11469 ^ x5;
  assign n11710 = n11466 & ~n11709;
  assign n11711 = n11710 ^ x2;
  assign n11715 = n11714 ^ n11711;
  assign n11724 = n11723 ^ n11715;
  assign n11733 = n11732 ^ n11724;
  assign n11706 = n11470 ^ n11465;
  assign n11707 = n11482 & ~n11706;
  assign n11708 = n11707 ^ n11481;
  assign n11734 = n11733 ^ n11708;
  assign n11698 = ~n1141 & n7830;
  assign n11699 = x78 & n7839;
  assign n11700 = x79 & n7834;
  assign n11701 = ~n11699 & ~n11700;
  assign n11702 = x80 & n8374;
  assign n11703 = n11701 & ~n11702;
  assign n11704 = ~n11698 & n11703;
  assign n11705 = n11704 ^ x56;
  assign n11735 = n11734 ^ n11705;
  assign n11695 = n11483 ^ n11449;
  assign n11696 = ~n11484 & n11695;
  assign n11697 = n11696 ^ n11449;
  assign n11736 = n11735 ^ n11697;
  assign n11745 = n11744 ^ n11736;
  assign n11692 = n11496 ^ n11485;
  assign n11693 = n11497 & ~n11692;
  assign n11694 = n11693 ^ n11488;
  assign n11746 = n11745 ^ n11694;
  assign n11755 = n11754 ^ n11746;
  assign n11689 = n11446 ^ n11438;
  assign n11690 = n11499 & ~n11689;
  assign n11691 = n11690 ^ n11498;
  assign n11756 = n11755 ^ n11691;
  assign n11765 = n11764 ^ n11756;
  assign n11686 = n11500 ^ n11427;
  assign n11687 = ~n11501 & n11686;
  assign n11688 = n11687 ^ n11427;
  assign n11766 = n11765 ^ n11688;
  assign n11775 = n11774 ^ n11766;
  assign n11683 = n11502 ^ n11421;
  assign n11684 = ~n11503 & ~n11683;
  assign n11685 = n11684 ^ n11424;
  assign n11776 = n11775 ^ n11685;
  assign n11675 = n3054 & n4415;
  assign n11676 = x93 & n4420;
  assign n11677 = x95 & n4614;
  assign n11678 = ~n11676 & ~n11677;
  assign n11679 = x94 & n4410;
  assign n11680 = n11678 & ~n11679;
  assign n11681 = ~n11675 & n11680;
  assign n11682 = n11681 ^ x41;
  assign n11777 = n11776 ^ n11682;
  assign n11672 = n11504 ^ n11405;
  assign n11673 = n11505 & n11672;
  assign n11674 = n11673 ^ n11405;
  assign n11778 = n11777 ^ n11674;
  assign n11664 = n3556 & n3829;
  assign n11665 = x96 & n4049;
  assign n11666 = x98 & n4052;
  assign n11667 = ~n11665 & ~n11666;
  assign n11668 = x97 & n3833;
  assign n11669 = n11667 & ~n11668;
  assign n11670 = ~n11664 & n11669;
  assign n11671 = n11670 ^ x38;
  assign n11779 = n11778 ^ n11671;
  assign n11661 = n11506 ^ n11394;
  assign n11662 = ~n11507 & ~n11661;
  assign n11663 = n11662 ^ n11394;
  assign n11780 = n11779 ^ n11663;
  assign n11653 = n3330 & n4105;
  assign n11654 = x99 & n3500;
  assign n11655 = x100 & n3334;
  assign n11656 = ~n11654 & ~n11655;
  assign n11657 = x101 & n3502;
  assign n11658 = n11656 & ~n11657;
  assign n11659 = ~n11653 & n11658;
  assign n11660 = n11659 ^ x35;
  assign n11781 = n11780 ^ n11660;
  assign n11650 = n11508 ^ n11383;
  assign n11651 = n11509 & n11650;
  assign n11652 = n11651 ^ n11383;
  assign n11782 = n11781 ^ n11652;
  assign n11642 = n2836 & n4670;
  assign n11643 = x103 & n2840;
  assign n11644 = x102 & n2996;
  assign n11645 = ~n11643 & ~n11644;
  assign n11646 = x104 & n2998;
  assign n11647 = n11645 & ~n11646;
  assign n11648 = ~n11642 & n11647;
  assign n11649 = n11648 ^ x32;
  assign n11783 = n11782 ^ n11649;
  assign n11639 = n11510 ^ n11372;
  assign n11640 = ~n11511 & ~n11639;
  assign n11641 = n11640 ^ n11372;
  assign n11784 = n11783 ^ n11641;
  assign n11631 = n2371 & n5297;
  assign n11632 = x105 & n2528;
  assign n11633 = x106 & n2377;
  assign n11634 = ~n11632 & ~n11633;
  assign n11635 = x107 & n2531;
  assign n11636 = n11634 & ~n11635;
  assign n11637 = ~n11631 & n11636;
  assign n11638 = n11637 ^ x29;
  assign n11785 = n11784 ^ n11638;
  assign n11628 = n11512 ^ n11361;
  assign n11629 = n11513 & n11628;
  assign n11630 = n11629 ^ n11361;
  assign n11786 = n11785 ^ n11630;
  assign n11620 = n1969 & n5955;
  assign n11621 = x108 & n1978;
  assign n11622 = x109 & n1973;
  assign n11623 = ~n11621 & ~n11622;
  assign n11624 = x110 & n2108;
  assign n11625 = n11623 & ~n11624;
  assign n11626 = ~n11620 & n11625;
  assign n11627 = n11626 ^ x26;
  assign n11787 = n11786 ^ n11627;
  assign n11617 = n11514 ^ n11350;
  assign n11618 = ~n11515 & ~n11617;
  assign n11619 = n11618 ^ n11350;
  assign n11788 = n11787 ^ n11619;
  assign n11609 = n1624 & n6656;
  assign n11610 = x112 & n1628;
  assign n11611 = x111 & n1742;
  assign n11612 = ~n11610 & ~n11611;
  assign n11613 = x113 & n1744;
  assign n11614 = n11612 & ~n11613;
  assign n11615 = ~n11609 & n11614;
  assign n11616 = n11615 ^ x23;
  assign n11789 = n11788 ^ n11616;
  assign n11606 = n11516 ^ n11339;
  assign n11607 = n11517 & n11606;
  assign n11608 = n11607 ^ n11339;
  assign n11790 = n11789 ^ n11608;
  assign n11598 = n1296 & n7393;
  assign n11599 = x114 & n1403;
  assign n11600 = x115 & n1300;
  assign n11601 = ~n11599 & ~n11600;
  assign n11602 = x116 & n1406;
  assign n11603 = n11601 & ~n11602;
  assign n11604 = ~n11598 & n11603;
  assign n11605 = n11604 ^ x20;
  assign n11791 = n11790 ^ n11605;
  assign n11595 = n11518 ^ n11328;
  assign n11596 = ~n11519 & n11595;
  assign n11597 = n11596 ^ n11328;
  assign n11792 = n11791 ^ n11597;
  assign n11587 = n1008 & n8169;
  assign n11588 = x117 & n1101;
  assign n11589 = x118 & n1012;
  assign n11590 = ~n11588 & ~n11589;
  assign n11591 = x119 & n1104;
  assign n11592 = n11590 & ~n11591;
  assign n11593 = ~n11587 & n11592;
  assign n11594 = n11593 ^ x17;
  assign n11793 = n11792 ^ n11594;
  assign n11584 = n11520 ^ n11317;
  assign n11585 = ~n11521 & n11584;
  assign n11586 = n11585 ^ n11317;
  assign n11794 = n11793 ^ n11586;
  assign n11576 = n752 & n9001;
  assign n11577 = x120 & n825;
  assign n11578 = x121 & n757;
  assign n11579 = ~n11577 & ~n11578;
  assign n11580 = x122 & n828;
  assign n11581 = n11579 & ~n11580;
  assign n11582 = ~n11576 & n11581;
  assign n11583 = n11582 ^ x14;
  assign n11795 = n11794 ^ n11583;
  assign n11573 = n11522 ^ n11306;
  assign n11574 = ~n11523 & ~n11573;
  assign n11575 = n11574 ^ n11306;
  assign n11796 = n11795 ^ n11575;
  assign n11565 = n541 & n9912;
  assign n11566 = x123 & n612;
  assign n11567 = x124 & n547;
  assign n11568 = ~n11566 & ~n11567;
  assign n11569 = x125 & n615;
  assign n11570 = n11568 & ~n11569;
  assign n11571 = ~n11565 & n11570;
  assign n11572 = n11571 ^ x11;
  assign n11797 = n11796 ^ n11572;
  assign n11562 = n11524 ^ n11295;
  assign n11563 = n11525 & n11562;
  assign n11564 = n11563 ^ n11295;
  assign n11798 = n11797 ^ n11564;
  assign n11556 = n372 & ~n9889;
  assign n11557 = x126 & n433;
  assign n11558 = x127 & n376;
  assign n11559 = ~n11557 & ~n11558;
  assign n11560 = ~n11556 & n11559;
  assign n11561 = n11560 ^ x8;
  assign n11799 = n11798 ^ n11561;
  assign n11553 = n11526 ^ n11284;
  assign n11554 = ~n11527 & ~n11553;
  assign n11555 = n11554 ^ n11284;
  assign n11800 = n11799 ^ n11555;
  assign n11550 = n11528 ^ n11273;
  assign n11551 = n11529 & n11550;
  assign n11552 = n11551 ^ n11273;
  assign n11801 = n11800 ^ n11552;
  assign n11813 = n11812 ^ n11801;
  assign n12037 = n3209 & n4415;
  assign n12038 = x94 & n4420;
  assign n12039 = x95 & n4410;
  assign n12040 = ~n12038 & ~n12039;
  assign n12041 = x96 & n4614;
  assign n12042 = n12040 & ~n12041;
  assign n12043 = ~n12037 & n12042;
  assign n12044 = n12043 ^ x41;
  assign n12027 = n2726 & n5010;
  assign n12028 = x91 & n5223;
  assign n12029 = x92 & n5014;
  assign n12030 = ~n12028 & ~n12029;
  assign n12031 = x93 & n5226;
  assign n12032 = n12030 & ~n12031;
  assign n12033 = ~n12027 & n12032;
  assign n12034 = n12033 ^ x44;
  assign n12017 = n2292 & n5656;
  assign n12018 = x88 & n5895;
  assign n12019 = x90 & n6111;
  assign n12020 = ~n12018 & ~n12019;
  assign n12021 = x89 & n5662;
  assign n12022 = n12020 & ~n12021;
  assign n12023 = ~n12017 & n12022;
  assign n12024 = n12023 ^ x47;
  assign n12014 = n11754 ^ n11691;
  assign n12015 = n11755 & n12014;
  assign n12016 = n12015 ^ n11691;
  assign n12025 = n12024 ^ n12016;
  assign n12004 = n1903 & n6326;
  assign n12005 = x85 & n6565;
  assign n12006 = x87 & n6569;
  assign n12007 = ~n12005 & ~n12006;
  assign n12008 = x86 & n6331;
  assign n12009 = n12007 & ~n12008;
  assign n12010 = ~n12004 & n12009;
  assign n12011 = n12010 ^ x50;
  assign n11994 = n1547 & n7076;
  assign n11995 = x82 & n7317;
  assign n11996 = x83 & n7080;
  assign n11997 = ~n11995 & ~n11996;
  assign n11998 = x84 & n7319;
  assign n11999 = n11997 & ~n11998;
  assign n12000 = ~n11994 & n11999;
  assign n12001 = n12000 ^ x53;
  assign n11982 = n953 & n8622;
  assign n11983 = x76 & n8631;
  assign n11984 = x77 & n8626;
  assign n11985 = ~n11983 & ~n11984;
  assign n11986 = x78 & n9186;
  assign n11987 = n11985 & ~n11986;
  assign n11988 = ~n11982 & n11987;
  assign n11989 = n11988 ^ x59;
  assign n11974 = n720 & n9499;
  assign n11975 = x73 & n9508;
  assign n11976 = x74 & n9503;
  assign n11977 = ~n11975 & ~n11976;
  assign n11978 = x75 & n10106;
  assign n11979 = n11977 & ~n11978;
  assign n11980 = ~n11974 & n11979;
  assign n11981 = n11980 ^ x62;
  assign n11990 = n11989 ^ n11981;
  assign n11969 = n344 & n10099;
  assign n11970 = x72 ^ x71;
  assign n11971 = n9798 & n11970;
  assign n11972 = ~n11969 & ~n11971;
  assign n11966 = n11723 ^ n11711;
  assign n11967 = n11715 & n11966;
  assign n11968 = n11967 ^ n11723;
  assign n11973 = n11972 ^ n11968;
  assign n11991 = n11990 ^ n11973;
  assign n11958 = n1230 & n7830;
  assign n11959 = x79 & n7839;
  assign n11960 = x81 & n8374;
  assign n11961 = ~n11959 & ~n11960;
  assign n11962 = x80 & n7834;
  assign n11963 = n11961 & ~n11962;
  assign n11964 = ~n11958 & n11963;
  assign n11965 = n11964 ^ x56;
  assign n11992 = n11991 ^ n11965;
  assign n11955 = n11732 ^ n11708;
  assign n11956 = n11733 & n11955;
  assign n11957 = n11956 ^ n11708;
  assign n11993 = n11992 ^ n11957;
  assign n12002 = n12001 ^ n11993;
  assign n11952 = n11734 ^ n11697;
  assign n11953 = n11735 & ~n11952;
  assign n11954 = n11953 ^ n11697;
  assign n12003 = n12002 ^ n11954;
  assign n12012 = n12011 ^ n12003;
  assign n11949 = n11744 ^ n11694;
  assign n11950 = n11745 & n11949;
  assign n11951 = n11950 ^ n11694;
  assign n12013 = n12012 ^ n11951;
  assign n12026 = n12025 ^ n12013;
  assign n12035 = n12034 ^ n12026;
  assign n11946 = n11756 ^ n11688;
  assign n11947 = ~n11765 & n11946;
  assign n11948 = n11947 ^ n11764;
  assign n12036 = n12035 ^ n11948;
  assign n12045 = n12044 ^ n12036;
  assign n11943 = n11774 ^ n11685;
  assign n11944 = n11775 & ~n11943;
  assign n11945 = n11944 ^ n11685;
  assign n12046 = n12045 ^ n11945;
  assign n11935 = n3730 & n3829;
  assign n11936 = x97 & n4049;
  assign n11937 = x99 & n4052;
  assign n11938 = ~n11936 & ~n11937;
  assign n11939 = x98 & n3833;
  assign n11940 = n11938 & ~n11939;
  assign n11941 = ~n11935 & n11940;
  assign n11942 = n11941 ^ x38;
  assign n12047 = n12046 ^ n11942;
  assign n11932 = n11776 ^ n11674;
  assign n11933 = ~n11777 & ~n11932;
  assign n11934 = n11933 ^ n11674;
  assign n12048 = n12047 ^ n11934;
  assign n11924 = n3330 & n4286;
  assign n11925 = x100 & n3500;
  assign n11926 = x102 & n3502;
  assign n11927 = ~n11925 & ~n11926;
  assign n11928 = x101 & n3334;
  assign n11929 = n11927 & ~n11928;
  assign n11930 = ~n11924 & n11929;
  assign n11931 = n11930 ^ x35;
  assign n12049 = n12048 ^ n11931;
  assign n11921 = n11778 ^ n11663;
  assign n11922 = n11779 & n11921;
  assign n11923 = n11922 ^ n11663;
  assign n12050 = n12049 ^ n11923;
  assign n11913 = n2836 & n4867;
  assign n11914 = x103 & n2996;
  assign n11915 = x104 & n2840;
  assign n11916 = ~n11914 & ~n11915;
  assign n11917 = x105 & n2998;
  assign n11918 = n11916 & ~n11917;
  assign n11919 = ~n11913 & n11918;
  assign n11920 = n11919 ^ x32;
  assign n12051 = n12050 ^ n11920;
  assign n11910 = n11780 ^ n11652;
  assign n11911 = ~n11781 & ~n11910;
  assign n11912 = n11911 ^ n11652;
  assign n12052 = n12051 ^ n11912;
  assign n11902 = n2371 & ~n5506;
  assign n11903 = x107 & n2377;
  assign n11904 = x106 & n2528;
  assign n11905 = ~n11903 & ~n11904;
  assign n11906 = x108 & n2531;
  assign n11907 = n11905 & ~n11906;
  assign n11908 = ~n11902 & n11907;
  assign n11909 = n11908 ^ x29;
  assign n12053 = n12052 ^ n11909;
  assign n11899 = n11782 ^ n11641;
  assign n11900 = n11783 & n11899;
  assign n11901 = n11900 ^ n11641;
  assign n12054 = n12053 ^ n11901;
  assign n11891 = n1969 & n6178;
  assign n11892 = x109 & n1978;
  assign n11893 = x111 & n2108;
  assign n11894 = ~n11892 & ~n11893;
  assign n11895 = x110 & n1973;
  assign n11896 = n11894 & ~n11895;
  assign n11897 = ~n11891 & n11896;
  assign n11898 = n11897 ^ x26;
  assign n12055 = n12054 ^ n11898;
  assign n11888 = n11784 ^ n11630;
  assign n11889 = ~n11785 & ~n11888;
  assign n11890 = n11889 ^ n11630;
  assign n12056 = n12055 ^ n11890;
  assign n11880 = n1624 & n6892;
  assign n11881 = x113 & n1628;
  assign n11882 = x112 & n1742;
  assign n11883 = ~n11881 & ~n11882;
  assign n11884 = x114 & n1744;
  assign n11885 = n11883 & ~n11884;
  assign n11886 = ~n11880 & n11885;
  assign n11887 = n11886 ^ x23;
  assign n12057 = n12056 ^ n11887;
  assign n11877 = n11786 ^ n11619;
  assign n11878 = n11787 & n11877;
  assign n11879 = n11878 ^ n11619;
  assign n12058 = n12057 ^ n11879;
  assign n11869 = n1296 & n7643;
  assign n11870 = x116 & n1300;
  assign n11871 = x115 & n1403;
  assign n11872 = ~n11870 & ~n11871;
  assign n11873 = x117 & n1406;
  assign n11874 = n11872 & ~n11873;
  assign n11875 = ~n11869 & n11874;
  assign n11876 = n11875 ^ x20;
  assign n12059 = n12058 ^ n11876;
  assign n11866 = n11788 ^ n11608;
  assign n11867 = ~n11789 & ~n11866;
  assign n11868 = n11867 ^ n11608;
  assign n12060 = n12059 ^ n11868;
  assign n11858 = n1008 & ~n8424;
  assign n11859 = x119 & n1012;
  assign n11860 = x118 & n1101;
  assign n11861 = ~n11859 & ~n11860;
  assign n11862 = x120 & n1104;
  assign n11863 = n11861 & ~n11862;
  assign n11864 = ~n11858 & n11863;
  assign n11865 = n11864 ^ x17;
  assign n12061 = n12060 ^ n11865;
  assign n11855 = n11790 ^ n11597;
  assign n11856 = n11791 & ~n11855;
  assign n11857 = n11856 ^ n11597;
  assign n12062 = n12061 ^ n11857;
  assign n11847 = n752 & n9309;
  assign n11848 = x121 & n825;
  assign n11849 = x123 & n828;
  assign n11850 = ~n11848 & ~n11849;
  assign n11851 = x122 & n757;
  assign n11852 = n11850 & ~n11851;
  assign n11853 = ~n11847 & n11852;
  assign n11854 = n11853 ^ x14;
  assign n12063 = n12062 ^ n11854;
  assign n11844 = n11792 ^ n11586;
  assign n11845 = n11793 & ~n11844;
  assign n11846 = n11845 ^ n11586;
  assign n12064 = n12063 ^ n11846;
  assign n11836 = n541 & ~n10174;
  assign n11837 = x124 & n612;
  assign n11838 = x126 & n615;
  assign n11839 = ~n11837 & ~n11838;
  assign n11840 = x125 & n547;
  assign n11841 = n11839 & ~n11840;
  assign n11842 = ~n11836 & n11841;
  assign n11843 = n11842 ^ x11;
  assign n12065 = n12064 ^ n11843;
  assign n11833 = n11583 ^ n11575;
  assign n11834 = ~n11795 & n11833;
  assign n11835 = n11834 ^ n11794;
  assign n12066 = n12065 ^ n11835;
  assign n11823 = x8 & n9886;
  assign n11824 = ~n314 & ~n11823;
  assign n11825 = ~x7 & n10430;
  assign n11826 = n11825 ^ n9886;
  assign n11827 = n11824 & n11826;
  assign n11828 = n310 ^ x7;
  assign n11829 = n371 & n11828;
  assign n11830 = x127 & n11829;
  assign n11831 = n11830 ^ x8;
  assign n11832 = ~n11827 & n11831;
  assign n12067 = n12066 ^ n11832;
  assign n11820 = n11796 ^ n11564;
  assign n11821 = ~n11797 & ~n11820;
  assign n11822 = n11821 ^ n11564;
  assign n12068 = n12067 ^ n11822;
  assign n11817 = n11798 ^ n11555;
  assign n11818 = n11799 & n11817;
  assign n11819 = n11818 ^ n11555;
  assign n12069 = n12068 ^ n11819;
  assign n11814 = n11812 ^ n11552;
  assign n11815 = n11801 & ~n11814;
  assign n11816 = n11815 ^ n11812;
  assign n12070 = n12069 ^ n11816;
  assign n12316 = n12066 ^ n11822;
  assign n12317 = ~n12067 & n12316;
  assign n12318 = n12317 ^ n11822;
  assign n12319 = n11819 & n12318;
  assign n12320 = n11832 & n12066;
  assign n12321 = n11822 & n12320;
  assign n12322 = ~n12319 & ~n12321;
  assign n12323 = ~n11816 & ~n12322;
  assign n12324 = ~n11832 & ~n12066;
  assign n12325 = ~n11822 & n12324;
  assign n12326 = n12325 ^ n12321;
  assign n12327 = ~n11819 & n12326;
  assign n12328 = n12327 ^ n12321;
  assign n12329 = ~n12323 & ~n12328;
  assign n12330 = n11819 & ~n12325;
  assign n12331 = ~n12318 & ~n12330;
  assign n12332 = n11816 & n12331;
  assign n12333 = n12329 & ~n12332;
  assign n12286 = n3388 & n4415;
  assign n12287 = x95 & n4420;
  assign n12288 = x96 & n4410;
  assign n12289 = ~n12287 & ~n12288;
  assign n12290 = x97 & n4614;
  assign n12291 = n12289 & ~n12290;
  assign n12292 = ~n12286 & n12291;
  assign n12293 = n12292 ^ x41;
  assign n12274 = n2447 & n5656;
  assign n12275 = x89 & n5895;
  assign n12276 = x90 & n5662;
  assign n12277 = ~n12275 & ~n12276;
  assign n12278 = x91 & n6111;
  assign n12279 = n12277 & ~n12278;
  assign n12280 = ~n12274 & n12279;
  assign n12281 = n12280 ^ x47;
  assign n12264 = n2040 & n6326;
  assign n12265 = x86 & n6565;
  assign n12266 = x88 & n6569;
  assign n12267 = ~n12265 & ~n12266;
  assign n12268 = x87 & n6331;
  assign n12269 = n12267 & ~n12268;
  assign n12270 = ~n12264 & n12269;
  assign n12271 = n12270 ^ x50;
  assign n12250 = n1054 & n8622;
  assign n12251 = x77 & n8631;
  assign n12252 = x78 & n8626;
  assign n12253 = ~n12251 & ~n12252;
  assign n12254 = x79 & n9186;
  assign n12255 = n12253 & ~n12254;
  assign n12256 = ~n12250 & n12255;
  assign n12257 = n12256 ^ x59;
  assign n12247 = n11981 ^ n11973;
  assign n12248 = n11990 & ~n12247;
  assign n12249 = n12248 ^ n11989;
  assign n12258 = n12257 ^ n12249;
  assign n12237 = ~x71 & n11713;
  assign n12238 = n402 & n9798;
  assign n12239 = ~n12237 & ~n12238;
  assign n12240 = n11968 & n12239;
  assign n12241 = x71 & n10099;
  assign n12242 = ~x70 & n12241;
  assign n12243 = n404 & n9798;
  assign n12244 = ~n12242 & ~n12243;
  assign n12245 = ~n12240 & n12244;
  assign n12228 = n799 & n9499;
  assign n12229 = x74 & n9508;
  assign n12230 = x76 & n10106;
  assign n12231 = ~n12229 & ~n12230;
  assign n12232 = x75 & n9503;
  assign n12233 = n12231 & ~n12232;
  assign n12234 = ~n12228 & n12233;
  assign n12235 = n12234 ^ x62;
  assign n12223 = n10099 & n11970;
  assign n12224 = x73 ^ x72;
  assign n12225 = n9798 & n12224;
  assign n12226 = ~n12223 & ~n12225;
  assign n12227 = n12226 ^ x8;
  assign n12236 = n12235 ^ n12227;
  assign n12246 = n12245 ^ n12236;
  assign n12259 = n12258 ^ n12246;
  assign n12215 = n1345 & n7830;
  assign n12216 = x80 & n7839;
  assign n12217 = x82 & n8374;
  assign n12218 = ~n12216 & ~n12217;
  assign n12219 = x81 & n7834;
  assign n12220 = n12218 & ~n12219;
  assign n12221 = ~n12215 & n12220;
  assign n12222 = n12221 ^ x56;
  assign n12260 = n12259 ^ n12222;
  assign n12212 = n11965 ^ n11957;
  assign n12213 = n11992 & ~n12212;
  assign n12214 = n12213 ^ n11991;
  assign n12261 = n12260 ^ n12214;
  assign n12204 = n1674 & n7076;
  assign n12205 = x83 & n7317;
  assign n12206 = x84 & n7080;
  assign n12207 = ~n12205 & ~n12206;
  assign n12208 = x85 & n7319;
  assign n12209 = n12207 & ~n12208;
  assign n12210 = ~n12204 & n12209;
  assign n12211 = n12210 ^ x53;
  assign n12262 = n12261 ^ n12211;
  assign n12201 = n11993 ^ n11954;
  assign n12202 = n12002 & ~n12201;
  assign n12203 = n12202 ^ n12001;
  assign n12263 = n12262 ^ n12203;
  assign n12272 = n12271 ^ n12263;
  assign n12198 = n12003 ^ n11951;
  assign n12199 = n12012 & ~n12198;
  assign n12200 = n12199 ^ n12011;
  assign n12273 = n12272 ^ n12200;
  assign n12282 = n12281 ^ n12273;
  assign n12195 = n12016 ^ n12013;
  assign n12196 = n12025 & ~n12195;
  assign n12197 = n12196 ^ n12024;
  assign n12283 = n12282 ^ n12197;
  assign n12192 = n12026 ^ n11948;
  assign n12193 = n12035 & ~n12192;
  assign n12194 = n12193 ^ n12034;
  assign n12284 = n12283 ^ n12194;
  assign n12184 = n2895 & n5010;
  assign n12185 = x92 & n5223;
  assign n12186 = x94 & n5226;
  assign n12187 = ~n12185 & ~n12186;
  assign n12188 = x93 & n5014;
  assign n12189 = n12187 & ~n12188;
  assign n12190 = ~n12184 & n12189;
  assign n12191 = n12190 ^ x44;
  assign n12285 = n12284 ^ n12191;
  assign n12294 = n12293 ^ n12285;
  assign n12181 = n12044 ^ n11945;
  assign n12182 = ~n12045 & ~n12181;
  assign n12183 = n12182 ^ n11945;
  assign n12295 = n12294 ^ n12183;
  assign n12173 = n3829 & n3925;
  assign n12174 = x98 & n4049;
  assign n12175 = x99 & n3833;
  assign n12176 = ~n12174 & ~n12175;
  assign n12177 = x100 & n4052;
  assign n12178 = n12176 & ~n12177;
  assign n12179 = ~n12173 & n12178;
  assign n12180 = n12179 ^ x38;
  assign n12296 = n12295 ^ n12180;
  assign n12170 = n12046 ^ n11934;
  assign n12171 = n12047 & n12170;
  assign n12172 = n12171 ^ n11934;
  assign n12297 = n12296 ^ n12172;
  assign n12162 = n3330 & n4481;
  assign n12163 = x101 & n3500;
  assign n12164 = x103 & n3502;
  assign n12165 = ~n12163 & ~n12164;
  assign n12166 = x102 & n3334;
  assign n12167 = n12165 & ~n12166;
  assign n12168 = ~n12162 & n12167;
  assign n12169 = n12168 ^ x35;
  assign n12298 = n12297 ^ n12169;
  assign n12159 = n12048 ^ n11923;
  assign n12160 = ~n12049 & ~n12159;
  assign n12161 = n12160 ^ n11923;
  assign n12299 = n12298 ^ n12161;
  assign n12151 = n2836 & n5088;
  assign n12152 = x104 & n2996;
  assign n12153 = x105 & n2840;
  assign n12154 = ~n12152 & ~n12153;
  assign n12155 = x106 & n2998;
  assign n12156 = n12154 & ~n12155;
  assign n12157 = ~n12151 & n12156;
  assign n12158 = n12157 ^ x32;
  assign n12300 = n12299 ^ n12158;
  assign n12148 = n12050 ^ n11912;
  assign n12149 = n12051 & n12148;
  assign n12150 = n12149 ^ n11912;
  assign n12301 = n12300 ^ n12150;
  assign n12140 = n2371 & ~n5737;
  assign n12141 = x107 & n2528;
  assign n12142 = x109 & n2531;
  assign n12143 = ~n12141 & ~n12142;
  assign n12144 = x108 & n2377;
  assign n12145 = n12143 & ~n12144;
  assign n12146 = ~n12140 & n12145;
  assign n12147 = n12146 ^ x29;
  assign n12302 = n12301 ^ n12147;
  assign n12137 = n12052 ^ n11901;
  assign n12138 = ~n12053 & ~n12137;
  assign n12139 = n12138 ^ n11901;
  assign n12303 = n12302 ^ n12139;
  assign n12129 = n1969 & n6420;
  assign n12130 = x110 & n1978;
  assign n12131 = x112 & n2108;
  assign n12132 = ~n12130 & ~n12131;
  assign n12133 = x111 & n1973;
  assign n12134 = n12132 & ~n12133;
  assign n12135 = ~n12129 & n12134;
  assign n12136 = n12135 ^ x26;
  assign n12304 = n12303 ^ n12136;
  assign n12126 = n12054 ^ n11890;
  assign n12127 = n12055 & n12126;
  assign n12128 = n12127 ^ n11890;
  assign n12305 = n12304 ^ n12128;
  assign n12118 = n1624 & n7150;
  assign n12119 = x113 & n1742;
  assign n12120 = x114 & n1628;
  assign n12121 = ~n12119 & ~n12120;
  assign n12122 = x115 & n1744;
  assign n12123 = n12121 & ~n12122;
  assign n12124 = ~n12118 & n12123;
  assign n12125 = n12124 ^ x23;
  assign n12306 = n12305 ^ n12125;
  assign n12115 = n12056 ^ n11879;
  assign n12116 = ~n12057 & ~n12115;
  assign n12117 = n12116 ^ n11879;
  assign n12307 = n12306 ^ n12117;
  assign n12107 = n1296 & n7919;
  assign n12108 = x117 & n1300;
  assign n12109 = x116 & n1403;
  assign n12110 = ~n12108 & ~n12109;
  assign n12111 = x118 & n1406;
  assign n12112 = n12110 & ~n12111;
  assign n12113 = ~n12107 & n12112;
  assign n12114 = n12113 ^ x20;
  assign n12308 = n12307 ^ n12114;
  assign n12104 = n12058 ^ n11868;
  assign n12105 = n12059 & n12104;
  assign n12106 = n12105 ^ n11868;
  assign n12309 = n12308 ^ n12106;
  assign n12096 = n1008 & n8715;
  assign n12097 = x120 & n1012;
  assign n12098 = x119 & n1101;
  assign n12099 = ~n12097 & ~n12098;
  assign n12100 = x121 & n1104;
  assign n12101 = n12099 & ~n12100;
  assign n12102 = ~n12096 & n12101;
  assign n12103 = n12102 ^ x17;
  assign n12310 = n12309 ^ n12103;
  assign n12093 = n12060 ^ n11857;
  assign n12094 = ~n12061 & n12093;
  assign n12095 = n12094 ^ n11857;
  assign n12311 = n12310 ^ n12095;
  assign n12085 = n752 & n9614;
  assign n12086 = x122 & n825;
  assign n12087 = x124 & n828;
  assign n12088 = ~n12086 & ~n12087;
  assign n12089 = x123 & n757;
  assign n12090 = n12088 & ~n12089;
  assign n12091 = ~n12085 & n12090;
  assign n12092 = n12091 ^ x14;
  assign n12312 = n12311 ^ n12092;
  assign n12082 = n12062 ^ n11846;
  assign n12083 = ~n12063 & n12082;
  assign n12084 = n12083 ^ n11846;
  assign n12313 = n12312 ^ n12084;
  assign n12074 = n541 & ~n10447;
  assign n12075 = x125 & n612;
  assign n12076 = x126 & n547;
  assign n12077 = ~n12075 & ~n12076;
  assign n12078 = x127 & n615;
  assign n12079 = n12077 & ~n12078;
  assign n12080 = ~n12074 & n12079;
  assign n12081 = n12080 ^ x11;
  assign n12314 = n12313 ^ n12081;
  assign n12071 = n12064 ^ n11835;
  assign n12072 = ~n12065 & ~n12071;
  assign n12073 = n12072 ^ n11835;
  assign n12315 = n12314 ^ n12073;
  assign n12334 = n12333 ^ n12315;
  assign n12580 = ~n12315 & ~n12321;
  assign n12581 = ~n12325 & ~n12580;
  assign n12582 = ~n11819 & ~n12581;
  assign n12583 = ~n12315 & ~n12318;
  assign n12584 = ~n12582 & ~n12583;
  assign n12585 = ~n11816 & n12584;
  assign n12586 = n11819 & n12581;
  assign n12587 = n12315 & n12318;
  assign n12588 = ~n12586 & ~n12587;
  assign n12589 = ~n12585 & n12588;
  assign n12551 = n3829 & n4105;
  assign n12552 = x99 & n4049;
  assign n12553 = x100 & n3833;
  assign n12554 = ~n12552 & ~n12553;
  assign n12555 = x101 & n4052;
  assign n12556 = n12554 & ~n12555;
  assign n12557 = ~n12551 & n12556;
  assign n12558 = n12557 ^ x38;
  assign n12541 = n3556 & n4415;
  assign n12542 = x96 & n4420;
  assign n12543 = x97 & n4410;
  assign n12544 = ~n12542 & ~n12543;
  assign n12545 = x98 & n4614;
  assign n12546 = n12544 & ~n12545;
  assign n12547 = ~n12541 & n12546;
  assign n12548 = n12547 ^ x41;
  assign n12531 = n3054 & n5010;
  assign n12532 = x93 & n5223;
  assign n12533 = x94 & n5014;
  assign n12534 = ~n12532 & ~n12533;
  assign n12535 = x95 & n5226;
  assign n12536 = n12534 & ~n12535;
  assign n12537 = ~n12531 & n12536;
  assign n12538 = n12537 ^ x44;
  assign n12521 = n2585 & n5656;
  assign n12522 = x90 & n5895;
  assign n12523 = x91 & n5662;
  assign n12524 = ~n12522 & ~n12523;
  assign n12525 = x92 & n6111;
  assign n12526 = n12524 & ~n12525;
  assign n12527 = ~n12521 & n12526;
  assign n12528 = n12527 ^ x47;
  assign n12511 = n2164 & n6326;
  assign n12512 = x88 & n6331;
  assign n12513 = x87 & n6565;
  assign n12514 = ~n12512 & ~n12513;
  assign n12515 = x89 & n6569;
  assign n12516 = n12514 & ~n12515;
  assign n12517 = ~n12511 & n12516;
  assign n12518 = n12517 ^ x50;
  assign n12501 = n1787 & n7076;
  assign n12502 = x85 & n7080;
  assign n12503 = x84 & n7317;
  assign n12504 = ~n12502 & ~n12503;
  assign n12505 = x86 & n7319;
  assign n12506 = n12504 & ~n12505;
  assign n12507 = ~n12501 & n12506;
  assign n12508 = n12507 ^ x53;
  assign n12498 = n12222 ^ n12214;
  assign n12499 = n12260 & ~n12498;
  assign n12500 = n12499 ^ n12259;
  assign n12509 = n12508 ^ n12500;
  assign n12488 = n1445 & n7830;
  assign n12489 = x81 & n7839;
  assign n12490 = x83 & n8374;
  assign n12491 = ~n12489 & ~n12490;
  assign n12492 = x82 & n7834;
  assign n12493 = n12491 & ~n12492;
  assign n12494 = ~n12488 & n12493;
  assign n12495 = n12494 ^ x56;
  assign n12478 = ~n1141 & n8622;
  assign n12479 = x78 & n8631;
  assign n12480 = x79 & n8626;
  assign n12481 = ~n12479 & ~n12480;
  assign n12482 = x80 & n9186;
  assign n12483 = n12481 & ~n12482;
  assign n12484 = ~n12478 & n12483;
  assign n12485 = n12484 ^ x59;
  assign n12469 = n877 & n9499;
  assign n12470 = x75 & n9508;
  assign n12471 = x76 & n9503;
  assign n12472 = ~n12470 & ~n12471;
  assign n12473 = x77 & n10106;
  assign n12474 = n12472 & ~n12473;
  assign n12475 = ~n12469 & n12474;
  assign n12476 = n12475 ^ x62;
  assign n12459 = ~x8 & x72;
  assign n12460 = x73 ^ x71;
  assign n12461 = ~n10099 & n12460;
  assign n12462 = n12461 ^ x71;
  assign n12463 = ~n12459 & ~n12462;
  assign n12464 = x8 & ~x72;
  assign n12465 = ~x62 & ~x63;
  assign n12466 = ~n12464 & ~n12465;
  assign n12467 = ~n12463 & n12466;
  assign n12456 = x74 & n9798;
  assign n12457 = x73 & n10099;
  assign n12458 = ~n12456 & ~n12457;
  assign n12468 = n12467 ^ n12458;
  assign n12477 = n12476 ^ n12468;
  assign n12486 = n12485 ^ n12477;
  assign n12453 = n12245 ^ n12235;
  assign n12454 = n12236 & ~n12453;
  assign n12455 = n12454 ^ n12245;
  assign n12487 = n12486 ^ n12455;
  assign n12496 = n12495 ^ n12487;
  assign n12450 = n12257 ^ n12246;
  assign n12451 = n12258 & ~n12450;
  assign n12452 = n12451 ^ n12249;
  assign n12497 = n12496 ^ n12452;
  assign n12510 = n12509 ^ n12497;
  assign n12519 = n12518 ^ n12510;
  assign n12447 = n12261 ^ n12203;
  assign n12448 = ~n12262 & n12447;
  assign n12449 = n12448 ^ n12203;
  assign n12520 = n12519 ^ n12449;
  assign n12529 = n12528 ^ n12520;
  assign n12444 = n12271 ^ n12200;
  assign n12445 = ~n12272 & n12444;
  assign n12446 = n12445 ^ n12200;
  assign n12530 = n12529 ^ n12446;
  assign n12539 = n12538 ^ n12530;
  assign n12441 = n12281 ^ n12197;
  assign n12442 = ~n12282 & n12441;
  assign n12443 = n12442 ^ n12197;
  assign n12540 = n12539 ^ n12443;
  assign n12549 = n12548 ^ n12540;
  assign n12438 = n12283 ^ n12191;
  assign n12439 = n12284 & ~n12438;
  assign n12440 = n12439 ^ n12194;
  assign n12550 = n12549 ^ n12440;
  assign n12559 = n12558 ^ n12550;
  assign n12435 = n12293 ^ n12183;
  assign n12436 = ~n12294 & ~n12435;
  assign n12437 = n12436 ^ n12183;
  assign n12560 = n12559 ^ n12437;
  assign n12427 = n3330 & n4670;
  assign n12428 = x102 & n3500;
  assign n12429 = x103 & n3334;
  assign n12430 = ~n12428 & ~n12429;
  assign n12431 = x104 & n3502;
  assign n12432 = n12430 & ~n12431;
  assign n12433 = ~n12427 & n12432;
  assign n12434 = n12433 ^ x35;
  assign n12561 = n12560 ^ n12434;
  assign n12424 = n12295 ^ n12172;
  assign n12425 = n12296 & n12424;
  assign n12426 = n12425 ^ n12172;
  assign n12562 = n12561 ^ n12426;
  assign n12416 = n2836 & n5297;
  assign n12417 = x106 & n2840;
  assign n12418 = x105 & n2996;
  assign n12419 = ~n12417 & ~n12418;
  assign n12420 = x107 & n2998;
  assign n12421 = n12419 & ~n12420;
  assign n12422 = ~n12416 & n12421;
  assign n12423 = n12422 ^ x32;
  assign n12563 = n12562 ^ n12423;
  assign n12413 = n12297 ^ n12161;
  assign n12414 = ~n12298 & ~n12413;
  assign n12415 = n12414 ^ n12161;
  assign n12564 = n12563 ^ n12415;
  assign n12405 = n2371 & n5955;
  assign n12406 = x109 & n2377;
  assign n12407 = x108 & n2528;
  assign n12408 = ~n12406 & ~n12407;
  assign n12409 = x110 & n2531;
  assign n12410 = n12408 & ~n12409;
  assign n12411 = ~n12405 & n12410;
  assign n12412 = n12411 ^ x29;
  assign n12565 = n12564 ^ n12412;
  assign n12402 = n12299 ^ n12150;
  assign n12403 = n12300 & n12402;
  assign n12404 = n12403 ^ n12150;
  assign n12566 = n12565 ^ n12404;
  assign n12394 = n1969 & n6656;
  assign n12395 = x111 & n1978;
  assign n12396 = x113 & n2108;
  assign n12397 = ~n12395 & ~n12396;
  assign n12398 = x112 & n1973;
  assign n12399 = n12397 & ~n12398;
  assign n12400 = ~n12394 & n12399;
  assign n12401 = n12400 ^ x26;
  assign n12567 = n12566 ^ n12401;
  assign n12391 = n12301 ^ n12139;
  assign n12392 = ~n12302 & ~n12391;
  assign n12393 = n12392 ^ n12139;
  assign n12568 = n12567 ^ n12393;
  assign n12383 = n1624 & n7393;
  assign n12384 = x114 & n1742;
  assign n12385 = x115 & n1628;
  assign n12386 = ~n12384 & ~n12385;
  assign n12387 = x116 & n1744;
  assign n12388 = n12386 & ~n12387;
  assign n12389 = ~n12383 & n12388;
  assign n12390 = n12389 ^ x23;
  assign n12569 = n12568 ^ n12390;
  assign n12380 = n12303 ^ n12128;
  assign n12381 = n12304 & n12380;
  assign n12382 = n12381 ^ n12128;
  assign n12570 = n12569 ^ n12382;
  assign n12372 = n1296 & n8169;
  assign n12373 = x117 & n1403;
  assign n12374 = x118 & n1300;
  assign n12375 = ~n12373 & ~n12374;
  assign n12376 = x119 & n1406;
  assign n12377 = n12375 & ~n12376;
  assign n12378 = ~n12372 & n12377;
  assign n12379 = n12378 ^ x20;
  assign n12571 = n12570 ^ n12379;
  assign n12369 = n12305 ^ n12117;
  assign n12370 = ~n12306 & ~n12369;
  assign n12371 = n12370 ^ n12117;
  assign n12572 = n12571 ^ n12371;
  assign n12361 = n1008 & n9001;
  assign n12362 = x120 & n1101;
  assign n12363 = x121 & n1012;
  assign n12364 = ~n12362 & ~n12363;
  assign n12365 = x122 & n1104;
  assign n12366 = n12364 & ~n12365;
  assign n12367 = ~n12361 & n12366;
  assign n12368 = n12367 ^ x17;
  assign n12573 = n12572 ^ n12368;
  assign n12358 = n12307 ^ n12106;
  assign n12359 = n12308 & n12358;
  assign n12360 = n12359 ^ n12106;
  assign n12574 = n12573 ^ n12360;
  assign n12350 = n752 & n9912;
  assign n12351 = x123 & n825;
  assign n12352 = x124 & n757;
  assign n12353 = ~n12351 & ~n12352;
  assign n12354 = x125 & n828;
  assign n12355 = n12353 & ~n12354;
  assign n12356 = ~n12350 & n12355;
  assign n12357 = n12356 ^ x14;
  assign n12575 = n12574 ^ n12357;
  assign n12347 = n12309 ^ n12095;
  assign n12348 = ~n12310 & n12347;
  assign n12349 = n12348 ^ n12095;
  assign n12576 = n12575 ^ n12349;
  assign n12341 = n541 & ~n9889;
  assign n12342 = x127 & n547;
  assign n12343 = x126 & n612;
  assign n12344 = ~n12342 & ~n12343;
  assign n12345 = ~n12341 & n12344;
  assign n12346 = n12345 ^ x11;
  assign n12577 = n12576 ^ n12346;
  assign n12338 = n12311 ^ n12084;
  assign n12339 = ~n12312 & n12338;
  assign n12340 = n12339 ^ n12084;
  assign n12578 = n12577 ^ n12340;
  assign n12335 = n12081 ^ n12073;
  assign n12336 = n12314 & n12335;
  assign n12337 = n12336 ^ n12313;
  assign n12579 = n12578 ^ n12337;
  assign n12590 = n12589 ^ n12579;
  assign n12810 = n3330 & n4867;
  assign n12811 = x103 & n3500;
  assign n12812 = x104 & n3334;
  assign n12813 = ~n12811 & ~n12812;
  assign n12814 = x105 & n3502;
  assign n12815 = n12813 & ~n12814;
  assign n12816 = ~n12810 & n12815;
  assign n12817 = n12816 ^ x35;
  assign n12801 = n3829 & n4286;
  assign n12802 = x100 & n4049;
  assign n12803 = x101 & n3833;
  assign n12804 = ~n12802 & ~n12803;
  assign n12805 = x102 & n4052;
  assign n12806 = n12804 & ~n12805;
  assign n12807 = ~n12801 & n12806;
  assign n12808 = n12807 ^ x38;
  assign n12791 = n3730 & n4415;
  assign n12792 = x97 & n4420;
  assign n12793 = x98 & n4410;
  assign n12794 = ~n12792 & ~n12793;
  assign n12795 = x99 & n4614;
  assign n12796 = n12794 & ~n12795;
  assign n12797 = ~n12791 & n12796;
  assign n12798 = n12797 ^ x41;
  assign n12780 = n3209 & n5010;
  assign n12781 = x94 & n5223;
  assign n12782 = x96 & n5226;
  assign n12783 = ~n12781 & ~n12782;
  assign n12784 = x95 & n5014;
  assign n12785 = n12783 & ~n12784;
  assign n12786 = ~n12780 & n12785;
  assign n12787 = n12786 ^ x44;
  assign n12770 = n2726 & n5656;
  assign n12771 = x91 & n5895;
  assign n12772 = x93 & n6111;
  assign n12773 = ~n12771 & ~n12772;
  assign n12774 = x92 & n5662;
  assign n12775 = n12773 & ~n12774;
  assign n12776 = ~n12770 & n12775;
  assign n12777 = n12776 ^ x47;
  assign n12760 = n2292 & n6326;
  assign n12761 = x88 & n6565;
  assign n12762 = x89 & n6331;
  assign n12763 = ~n12761 & ~n12762;
  assign n12764 = x90 & n6569;
  assign n12765 = n12763 & ~n12764;
  assign n12766 = ~n12760 & n12765;
  assign n12767 = n12766 ^ x50;
  assign n12757 = n12508 ^ n12497;
  assign n12758 = n12509 & n12757;
  assign n12759 = n12758 ^ n12500;
  assign n12768 = n12767 ^ n12759;
  assign n12747 = n1903 & n7076;
  assign n12748 = x85 & n7317;
  assign n12749 = x87 & n7319;
  assign n12750 = ~n12748 & ~n12749;
  assign n12751 = x86 & n7080;
  assign n12752 = n12750 & ~n12751;
  assign n12753 = ~n12747 & n12752;
  assign n12754 = n12753 ^ x53;
  assign n12737 = n1547 & n7830;
  assign n12738 = x82 & n7839;
  assign n12739 = x84 & n8374;
  assign n12740 = ~n12738 & ~n12739;
  assign n12741 = x83 & n7834;
  assign n12742 = n12740 & ~n12741;
  assign n12743 = ~n12737 & n12742;
  assign n12744 = n12743 ^ x56;
  assign n12727 = ~x75 & n12456;
  assign n12728 = ~x74 & x75;
  assign n12729 = n9798 & n12728;
  assign n12730 = x74 ^ x73;
  assign n12731 = n10099 & n12730;
  assign n12732 = ~n12729 & ~n12731;
  assign n12733 = ~n12727 & n12732;
  assign n12724 = n12476 ^ n12467;
  assign n12725 = ~n12468 & ~n12724;
  assign n12726 = n12725 ^ n12476;
  assign n12734 = n12733 ^ n12726;
  assign n12716 = n953 & n9499;
  assign n12717 = x76 & n9508;
  assign n12718 = x77 & n9503;
  assign n12719 = ~n12717 & ~n12718;
  assign n12720 = x78 & n10106;
  assign n12721 = n12719 & ~n12720;
  assign n12722 = ~n12716 & n12721;
  assign n12723 = n12722 ^ x62;
  assign n12735 = n12734 ^ n12723;
  assign n12708 = n1230 & n8622;
  assign n12709 = x79 & n8631;
  assign n12710 = x80 & n8626;
  assign n12711 = ~n12709 & ~n12710;
  assign n12712 = x81 & n9186;
  assign n12713 = n12711 & ~n12712;
  assign n12714 = ~n12708 & n12713;
  assign n12715 = n12714 ^ x59;
  assign n12736 = n12735 ^ n12715;
  assign n12745 = n12744 ^ n12736;
  assign n12705 = n12485 ^ n12455;
  assign n12706 = ~n12486 & ~n12705;
  assign n12707 = n12706 ^ n12455;
  assign n12746 = n12745 ^ n12707;
  assign n12755 = n12754 ^ n12746;
  assign n12702 = n12495 ^ n12452;
  assign n12703 = n12496 & n12702;
  assign n12704 = n12703 ^ n12452;
  assign n12756 = n12755 ^ n12704;
  assign n12769 = n12768 ^ n12756;
  assign n12778 = n12777 ^ n12769;
  assign n12699 = n12510 ^ n12449;
  assign n12700 = ~n12519 & n12699;
  assign n12701 = n12700 ^ n12518;
  assign n12779 = n12778 ^ n12701;
  assign n12788 = n12787 ^ n12779;
  assign n12696 = n12520 ^ n12446;
  assign n12697 = ~n12529 & n12696;
  assign n12698 = n12697 ^ n12528;
  assign n12789 = n12788 ^ n12698;
  assign n12693 = n12530 ^ n12443;
  assign n12694 = ~n12539 & n12693;
  assign n12695 = n12694 ^ n12538;
  assign n12790 = n12789 ^ n12695;
  assign n12799 = n12798 ^ n12790;
  assign n12690 = n12540 ^ n12440;
  assign n12691 = ~n12549 & n12690;
  assign n12692 = n12691 ^ n12548;
  assign n12800 = n12799 ^ n12692;
  assign n12809 = n12808 ^ n12800;
  assign n12818 = n12817 ^ n12809;
  assign n12687 = n12558 ^ n12437;
  assign n12688 = n12559 & ~n12687;
  assign n12689 = n12688 ^ n12437;
  assign n12819 = n12818 ^ n12689;
  assign n12679 = n2836 & ~n5506;
  assign n12680 = x106 & n2996;
  assign n12681 = x107 & n2840;
  assign n12682 = ~n12680 & ~n12681;
  assign n12683 = x108 & n2998;
  assign n12684 = n12682 & ~n12683;
  assign n12685 = ~n12679 & n12684;
  assign n12686 = n12685 ^ x32;
  assign n12820 = n12819 ^ n12686;
  assign n12676 = n12560 ^ n12426;
  assign n12677 = ~n12561 & ~n12676;
  assign n12678 = n12677 ^ n12426;
  assign n12821 = n12820 ^ n12678;
  assign n12668 = n2371 & n6178;
  assign n12669 = x110 & n2377;
  assign n12670 = x109 & n2528;
  assign n12671 = ~n12669 & ~n12670;
  assign n12672 = x111 & n2531;
  assign n12673 = n12671 & ~n12672;
  assign n12674 = ~n12668 & n12673;
  assign n12675 = n12674 ^ x29;
  assign n12822 = n12821 ^ n12675;
  assign n12665 = n12562 ^ n12415;
  assign n12666 = n12563 & n12665;
  assign n12667 = n12666 ^ n12415;
  assign n12823 = n12822 ^ n12667;
  assign n12657 = n1969 & n6892;
  assign n12658 = x112 & n1978;
  assign n12659 = x113 & n1973;
  assign n12660 = ~n12658 & ~n12659;
  assign n12661 = x114 & n2108;
  assign n12662 = n12660 & ~n12661;
  assign n12663 = ~n12657 & n12662;
  assign n12664 = n12663 ^ x26;
  assign n12824 = n12823 ^ n12664;
  assign n12654 = n12564 ^ n12404;
  assign n12655 = ~n12565 & ~n12654;
  assign n12656 = n12655 ^ n12404;
  assign n12825 = n12824 ^ n12656;
  assign n12646 = n1624 & n7643;
  assign n12647 = x115 & n1742;
  assign n12648 = x116 & n1628;
  assign n12649 = ~n12647 & ~n12648;
  assign n12650 = x117 & n1744;
  assign n12651 = n12649 & ~n12650;
  assign n12652 = ~n12646 & n12651;
  assign n12653 = n12652 ^ x23;
  assign n12826 = n12825 ^ n12653;
  assign n12643 = n12566 ^ n12393;
  assign n12644 = n12567 & n12643;
  assign n12645 = n12644 ^ n12393;
  assign n12827 = n12826 ^ n12645;
  assign n12635 = n1296 & ~n8424;
  assign n12636 = x119 & n1300;
  assign n12637 = x118 & n1403;
  assign n12638 = ~n12636 & ~n12637;
  assign n12639 = x120 & n1406;
  assign n12640 = n12638 & ~n12639;
  assign n12641 = ~n12635 & n12640;
  assign n12642 = n12641 ^ x20;
  assign n12828 = n12827 ^ n12642;
  assign n12632 = n12568 ^ n12382;
  assign n12633 = ~n12569 & ~n12632;
  assign n12634 = n12633 ^ n12382;
  assign n12829 = n12828 ^ n12634;
  assign n12624 = n1008 & n9309;
  assign n12625 = x122 & n1012;
  assign n12626 = x121 & n1101;
  assign n12627 = ~n12625 & ~n12626;
  assign n12628 = x123 & n1104;
  assign n12629 = n12627 & ~n12628;
  assign n12630 = ~n12624 & n12629;
  assign n12631 = n12630 ^ x17;
  assign n12830 = n12829 ^ n12631;
  assign n12621 = n12570 ^ n12371;
  assign n12622 = n12571 & n12621;
  assign n12623 = n12622 ^ n12371;
  assign n12831 = n12830 ^ n12623;
  assign n12613 = n752 & ~n10174;
  assign n12614 = x124 & n825;
  assign n12615 = x126 & n828;
  assign n12616 = ~n12614 & ~n12615;
  assign n12617 = x125 & n757;
  assign n12618 = n12616 & ~n12617;
  assign n12619 = ~n12613 & n12618;
  assign n12620 = n12619 ^ x14;
  assign n12832 = n12831 ^ n12620;
  assign n12610 = n12572 ^ n12360;
  assign n12611 = ~n12573 & ~n12610;
  assign n12612 = n12611 ^ n12360;
  assign n12833 = n12832 ^ n12612;
  assign n12600 = ~x10 & n10430;
  assign n12601 = n12600 ^ n9886;
  assign n12602 = ~n543 & n12601;
  assign n12603 = x11 & n9886;
  assign n12604 = n12602 & ~n12603;
  assign n12605 = n544 ^ x10;
  assign n12606 = n540 & n12605;
  assign n12607 = x127 & n12606;
  assign n12608 = n12607 ^ x11;
  assign n12609 = ~n12604 & n12608;
  assign n12834 = n12833 ^ n12609;
  assign n12597 = n12574 ^ n12349;
  assign n12598 = n12575 & ~n12597;
  assign n12599 = n12598 ^ n12349;
  assign n12835 = n12834 ^ n12599;
  assign n12594 = n12576 ^ n12340;
  assign n12595 = n12577 & ~n12594;
  assign n12596 = n12595 ^ n12340;
  assign n12836 = n12835 ^ n12596;
  assign n12591 = n12589 ^ n12337;
  assign n12592 = n12579 & n12591;
  assign n12593 = n12592 ^ n12589;
  assign n12837 = n12836 ^ n12593;
  assign n13047 = n3330 & n5088;
  assign n13048 = x104 & n3500;
  assign n13049 = x106 & n3502;
  assign n13050 = ~n13048 & ~n13049;
  assign n13051 = x105 & n3334;
  assign n13052 = n13050 & ~n13051;
  assign n13053 = ~n13047 & n13052;
  assign n13054 = n13053 ^ x35;
  assign n13035 = n3925 & n4415;
  assign n13036 = x98 & n4420;
  assign n13037 = x100 & n4614;
  assign n13038 = ~n13036 & ~n13037;
  assign n13039 = x99 & n4410;
  assign n13040 = n13038 & ~n13039;
  assign n13041 = ~n13035 & n13040;
  assign n13042 = n13041 ^ x41;
  assign n13025 = n3388 & n5010;
  assign n13026 = x95 & n5223;
  assign n13027 = x96 & n5014;
  assign n13028 = ~n13026 & ~n13027;
  assign n13029 = x97 & n5226;
  assign n13030 = n13028 & ~n13029;
  assign n13031 = ~n13025 & n13030;
  assign n13032 = n13031 ^ x44;
  assign n13015 = n2895 & n5656;
  assign n13016 = x92 & n5895;
  assign n13017 = x93 & n5662;
  assign n13018 = ~n13016 & ~n13017;
  assign n13019 = x94 & n6111;
  assign n13020 = n13018 & ~n13019;
  assign n13021 = ~n13015 & n13020;
  assign n13022 = n13021 ^ x47;
  assign n13012 = n12769 ^ n12701;
  assign n13013 = ~n12778 & n13012;
  assign n13014 = n13013 ^ n12777;
  assign n13023 = n13022 ^ n13014;
  assign n13002 = n2447 & n6326;
  assign n13003 = x89 & n6565;
  assign n13004 = x90 & n6331;
  assign n13005 = ~n13003 & ~n13004;
  assign n13006 = x91 & n6569;
  assign n13007 = n13005 & ~n13006;
  assign n13008 = ~n13002 & n13007;
  assign n13009 = n13008 ^ x50;
  assign n12992 = n2040 & n7076;
  assign n12993 = x86 & n7317;
  assign n12994 = x87 & n7080;
  assign n12995 = ~n12993 & ~n12994;
  assign n12996 = x88 & n7319;
  assign n12997 = n12995 & ~n12996;
  assign n12998 = ~n12992 & n12997;
  assign n12999 = n12998 ^ x53;
  assign n12983 = n12726 & n12732;
  assign n12984 = ~x74 & n12457;
  assign n12985 = ~n12727 & ~n12984;
  assign n12986 = ~n12983 & n12985;
  assign n12974 = n1054 & n9499;
  assign n12975 = x77 & n9508;
  assign n12976 = x78 & n9503;
  assign n12977 = ~n12975 & ~n12976;
  assign n12978 = x79 & n10106;
  assign n12979 = n12977 & ~n12978;
  assign n12980 = ~n12974 & n12979;
  assign n12981 = n12980 ^ x62;
  assign n12969 = x76 & n9798;
  assign n12970 = x75 & n10099;
  assign n12971 = ~n12969 & ~n12970;
  assign n12972 = n12971 ^ n12458;
  assign n12973 = n12972 ^ x11;
  assign n12982 = n12981 ^ n12973;
  assign n12987 = n12986 ^ n12982;
  assign n12961 = n1345 & n8622;
  assign n12962 = x80 & n8631;
  assign n12963 = x81 & n8626;
  assign n12964 = ~n12962 & ~n12963;
  assign n12965 = x82 & n9186;
  assign n12966 = n12964 & ~n12965;
  assign n12967 = ~n12961 & n12966;
  assign n12968 = n12967 ^ x59;
  assign n12988 = n12987 ^ n12968;
  assign n12958 = n12723 ^ n12715;
  assign n12959 = n12735 & ~n12958;
  assign n12960 = n12959 ^ n12734;
  assign n12989 = n12988 ^ n12960;
  assign n12950 = n1674 & n7830;
  assign n12951 = x83 & n7839;
  assign n12952 = x85 & n8374;
  assign n12953 = ~n12951 & ~n12952;
  assign n12954 = x84 & n7834;
  assign n12955 = n12953 & ~n12954;
  assign n12956 = ~n12950 & n12955;
  assign n12957 = n12956 ^ x56;
  assign n12990 = n12989 ^ n12957;
  assign n12947 = n12736 ^ n12707;
  assign n12948 = n12745 & n12947;
  assign n12949 = n12948 ^ n12744;
  assign n12991 = n12990 ^ n12949;
  assign n13000 = n12999 ^ n12991;
  assign n12944 = n12746 ^ n12704;
  assign n12945 = ~n12755 & n12944;
  assign n12946 = n12945 ^ n12754;
  assign n13001 = n13000 ^ n12946;
  assign n13010 = n13009 ^ n13001;
  assign n12941 = n12759 ^ n12756;
  assign n12942 = n12768 & n12941;
  assign n12943 = n12942 ^ n12767;
  assign n13011 = n13010 ^ n12943;
  assign n13024 = n13023 ^ n13011;
  assign n13033 = n13032 ^ n13024;
  assign n12938 = n12779 ^ n12698;
  assign n12939 = ~n12788 & n12938;
  assign n12940 = n12939 ^ n12787;
  assign n13034 = n13033 ^ n12940;
  assign n13043 = n13042 ^ n13034;
  assign n12935 = n12798 ^ n12789;
  assign n12936 = n12790 & ~n12935;
  assign n12937 = n12936 ^ n12798;
  assign n13044 = n13043 ^ n12937;
  assign n12932 = n12808 ^ n12692;
  assign n12933 = n12800 & n12932;
  assign n12934 = n12933 ^ n12808;
  assign n13045 = n13044 ^ n12934;
  assign n12924 = n3829 & n4481;
  assign n12925 = x101 & n4049;
  assign n12926 = x103 & n4052;
  assign n12927 = ~n12925 & ~n12926;
  assign n12928 = x102 & n3833;
  assign n12929 = n12927 & ~n12928;
  assign n12930 = ~n12924 & n12929;
  assign n12931 = n12930 ^ x38;
  assign n13046 = n13045 ^ n12931;
  assign n13055 = n13054 ^ n13046;
  assign n12921 = n12817 ^ n12689;
  assign n12922 = n12818 & ~n12921;
  assign n12923 = n12922 ^ n12689;
  assign n13056 = n13055 ^ n12923;
  assign n12913 = n2836 & ~n5737;
  assign n12914 = x108 & n2840;
  assign n12915 = x107 & n2996;
  assign n12916 = ~n12914 & ~n12915;
  assign n12917 = x109 & n2998;
  assign n12918 = n12916 & ~n12917;
  assign n12919 = ~n12913 & n12918;
  assign n12920 = n12919 ^ x32;
  assign n13057 = n13056 ^ n12920;
  assign n12910 = n12819 ^ n12678;
  assign n12911 = ~n12820 & ~n12910;
  assign n12912 = n12911 ^ n12678;
  assign n13058 = n13057 ^ n12912;
  assign n12902 = n2371 & n6420;
  assign n12903 = x110 & n2528;
  assign n12904 = x112 & n2531;
  assign n12905 = ~n12903 & ~n12904;
  assign n12906 = x111 & n2377;
  assign n12907 = n12905 & ~n12906;
  assign n12908 = ~n12902 & n12907;
  assign n12909 = n12908 ^ x29;
  assign n13059 = n13058 ^ n12909;
  assign n12899 = n12821 ^ n12667;
  assign n12900 = n12822 & n12899;
  assign n12901 = n12900 ^ n12667;
  assign n13060 = n13059 ^ n12901;
  assign n12891 = n1969 & n7150;
  assign n12892 = x113 & n1978;
  assign n12893 = x114 & n1973;
  assign n12894 = ~n12892 & ~n12893;
  assign n12895 = x115 & n2108;
  assign n12896 = n12894 & ~n12895;
  assign n12897 = ~n12891 & n12896;
  assign n12898 = n12897 ^ x26;
  assign n13061 = n13060 ^ n12898;
  assign n12888 = n12823 ^ n12656;
  assign n12889 = ~n12824 & ~n12888;
  assign n12890 = n12889 ^ n12656;
  assign n13062 = n13061 ^ n12890;
  assign n12880 = n1624 & n7919;
  assign n12881 = x116 & n1742;
  assign n12882 = x117 & n1628;
  assign n12883 = ~n12881 & ~n12882;
  assign n12884 = x118 & n1744;
  assign n12885 = n12883 & ~n12884;
  assign n12886 = ~n12880 & n12885;
  assign n12887 = n12886 ^ x23;
  assign n13063 = n13062 ^ n12887;
  assign n12877 = n12825 ^ n12645;
  assign n12878 = n12826 & n12877;
  assign n12879 = n12878 ^ n12645;
  assign n13064 = n13063 ^ n12879;
  assign n12869 = n1296 & n8715;
  assign n12870 = x119 & n1403;
  assign n12871 = x121 & n1406;
  assign n12872 = ~n12870 & ~n12871;
  assign n12873 = x120 & n1300;
  assign n12874 = n12872 & ~n12873;
  assign n12875 = ~n12869 & n12874;
  assign n12876 = n12875 ^ x20;
  assign n13065 = n13064 ^ n12876;
  assign n12866 = n12827 ^ n12634;
  assign n12867 = ~n12828 & ~n12866;
  assign n12868 = n12867 ^ n12634;
  assign n13066 = n13065 ^ n12868;
  assign n12858 = n1008 & n9614;
  assign n12859 = x122 & n1101;
  assign n12860 = x123 & n1012;
  assign n12861 = ~n12859 & ~n12860;
  assign n12862 = x124 & n1104;
  assign n12863 = n12861 & ~n12862;
  assign n12864 = ~n12858 & n12863;
  assign n12865 = n12864 ^ x17;
  assign n13067 = n13066 ^ n12865;
  assign n12855 = n12829 ^ n12623;
  assign n12856 = n12830 & n12855;
  assign n12857 = n12856 ^ n12623;
  assign n13068 = n13067 ^ n12857;
  assign n12847 = n752 & ~n10447;
  assign n12848 = x125 & n825;
  assign n12849 = x126 & n757;
  assign n12850 = ~n12848 & ~n12849;
  assign n12851 = x127 & n828;
  assign n12852 = n12850 & ~n12851;
  assign n12853 = ~n12847 & n12852;
  assign n12854 = n12853 ^ x14;
  assign n13069 = n13068 ^ n12854;
  assign n12844 = n12831 ^ n12612;
  assign n12845 = ~n12832 & ~n12844;
  assign n12846 = n12845 ^ n12612;
  assign n13070 = n13069 ^ n12846;
  assign n12841 = n12833 ^ n12599;
  assign n12842 = ~n12834 & ~n12841;
  assign n12843 = n12842 ^ n12599;
  assign n13071 = n13070 ^ n12843;
  assign n12838 = n12596 ^ n12593;
  assign n12839 = ~n12836 & n12838;
  assign n12840 = n12839 ^ n12593;
  assign n13072 = n13071 ^ n12840;
  assign n13279 = n2836 & n5955;
  assign n13280 = x108 & n2996;
  assign n13281 = x109 & n2840;
  assign n13282 = ~n13280 & ~n13281;
  assign n13283 = x110 & n2998;
  assign n13284 = n13282 & ~n13283;
  assign n13285 = ~n13279 & n13284;
  assign n13286 = n13285 ^ x32;
  assign n13270 = n3330 & n5297;
  assign n13271 = x105 & n3500;
  assign n13272 = x106 & n3334;
  assign n13273 = ~n13271 & ~n13272;
  assign n13274 = x107 & n3502;
  assign n13275 = n13273 & ~n13274;
  assign n13276 = ~n13270 & n13275;
  assign n13277 = n13276 ^ x35;
  assign n13260 = n3829 & n4670;
  assign n13261 = x102 & n4049;
  assign n13262 = x104 & n4052;
  assign n13263 = ~n13261 & ~n13262;
  assign n13264 = x103 & n3833;
  assign n13265 = n13263 & ~n13264;
  assign n13266 = ~n13260 & n13265;
  assign n13267 = n13266 ^ x38;
  assign n13250 = n4105 & n4415;
  assign n13251 = x99 & n4420;
  assign n13252 = x100 & n4410;
  assign n13253 = ~n13251 & ~n13252;
  assign n13254 = x101 & n4614;
  assign n13255 = n13253 & ~n13254;
  assign n13256 = ~n13250 & n13255;
  assign n13257 = n13256 ^ x41;
  assign n13239 = n3556 & n5010;
  assign n13240 = x96 & n5223;
  assign n13241 = x98 & n5226;
  assign n13242 = ~n13240 & ~n13241;
  assign n13243 = x97 & n5014;
  assign n13244 = n13242 & ~n13243;
  assign n13245 = ~n13239 & n13244;
  assign n13246 = n13245 ^ x44;
  assign n13229 = n3054 & n5656;
  assign n13230 = x93 & n5895;
  assign n13231 = x95 & n6111;
  assign n13232 = ~n13230 & ~n13231;
  assign n13233 = x94 & n5662;
  assign n13234 = n13232 & ~n13233;
  assign n13235 = ~n13229 & n13234;
  assign n13236 = n13235 ^ x47;
  assign n13219 = n2585 & n6326;
  assign n13220 = x90 & n6565;
  assign n13221 = x92 & n6569;
  assign n13222 = ~n13220 & ~n13221;
  assign n13223 = x91 & n6331;
  assign n13224 = n13222 & ~n13223;
  assign n13225 = ~n13219 & n13224;
  assign n13226 = n13225 ^ x50;
  assign n13209 = n2164 & n7076;
  assign n13210 = x88 & n7080;
  assign n13211 = x87 & n7317;
  assign n13212 = ~n13210 & ~n13211;
  assign n13213 = x89 & n7319;
  assign n13214 = n13212 & ~n13213;
  assign n13215 = ~n13209 & n13214;
  assign n13216 = n13215 ^ x53;
  assign n13199 = n1787 & n7830;
  assign n13200 = x85 & n7834;
  assign n13201 = x84 & n7839;
  assign n13202 = ~n13200 & ~n13201;
  assign n13203 = x86 & n8374;
  assign n13204 = n13202 & ~n13203;
  assign n13205 = ~n13199 & n13204;
  assign n13206 = n13205 ^ x56;
  assign n13196 = n12987 ^ n12960;
  assign n13197 = n12988 & ~n13196;
  assign n13198 = n13197 ^ n12960;
  assign n13207 = n13206 ^ n13198;
  assign n13186 = n1445 & n8622;
  assign n13187 = x81 & n8631;
  assign n13188 = x83 & n9186;
  assign n13189 = ~n13187 & ~n13188;
  assign n13190 = x82 & n8626;
  assign n13191 = n13189 & ~n13190;
  assign n13192 = ~n13186 & n13191;
  assign n13193 = n13192 ^ x59;
  assign n13177 = ~n1141 & n9499;
  assign n13178 = x78 & n9508;
  assign n13179 = x80 & n10106;
  assign n13180 = ~n13178 & ~n13179;
  assign n13181 = x79 & n9503;
  assign n13182 = n13180 & ~n13181;
  assign n13183 = ~n13177 & n13182;
  assign n13184 = n13183 ^ x62;
  assign n13173 = x77 & n9798;
  assign n13174 = x76 & n10099;
  assign n13175 = ~n13173 & ~n13174;
  assign n13170 = n12458 ^ x11;
  assign n13171 = ~n12972 & n13170;
  assign n13172 = n13171 ^ x11;
  assign n13176 = n13175 ^ n13172;
  assign n13185 = n13184 ^ n13176;
  assign n13194 = n13193 ^ n13185;
  assign n13167 = n12986 ^ n12981;
  assign n13168 = ~n12982 & ~n13167;
  assign n13169 = n13168 ^ n12986;
  assign n13195 = n13194 ^ n13169;
  assign n13208 = n13207 ^ n13195;
  assign n13217 = n13216 ^ n13208;
  assign n13164 = n12989 ^ n12949;
  assign n13165 = n12990 & ~n13164;
  assign n13166 = n13165 ^ n12949;
  assign n13218 = n13217 ^ n13166;
  assign n13227 = n13226 ^ n13218;
  assign n13161 = n12999 ^ n12946;
  assign n13162 = n13000 & n13161;
  assign n13163 = n13162 ^ n12946;
  assign n13228 = n13227 ^ n13163;
  assign n13237 = n13236 ^ n13228;
  assign n13158 = n13009 ^ n12943;
  assign n13159 = n13010 & n13158;
  assign n13160 = n13159 ^ n12943;
  assign n13238 = n13237 ^ n13160;
  assign n13247 = n13246 ^ n13238;
  assign n13155 = n13022 ^ n13011;
  assign n13156 = n13023 & n13155;
  assign n13157 = n13156 ^ n13014;
  assign n13248 = n13247 ^ n13157;
  assign n13152 = n13032 ^ n12940;
  assign n13153 = n13033 & n13152;
  assign n13154 = n13153 ^ n12940;
  assign n13249 = n13248 ^ n13154;
  assign n13258 = n13257 ^ n13249;
  assign n13149 = n13042 ^ n12937;
  assign n13150 = n13043 & n13149;
  assign n13151 = n13150 ^ n12937;
  assign n13259 = n13258 ^ n13151;
  assign n13268 = n13267 ^ n13259;
  assign n13146 = n13044 ^ n12931;
  assign n13147 = ~n13045 & n13146;
  assign n13148 = n13147 ^ n12934;
  assign n13269 = n13268 ^ n13148;
  assign n13278 = n13277 ^ n13269;
  assign n13287 = n13286 ^ n13278;
  assign n13143 = n13054 ^ n12923;
  assign n13144 = n13055 & ~n13143;
  assign n13145 = n13144 ^ n12923;
  assign n13288 = n13287 ^ n13145;
  assign n13140 = n13056 ^ n12912;
  assign n13141 = ~n13057 & ~n13140;
  assign n13142 = n13141 ^ n12912;
  assign n13289 = n13288 ^ n13142;
  assign n13132 = n2371 & n6656;
  assign n13133 = x111 & n2528;
  assign n13134 = x113 & n2531;
  assign n13135 = ~n13133 & ~n13134;
  assign n13136 = x112 & n2377;
  assign n13137 = n13135 & ~n13136;
  assign n13138 = ~n13132 & n13137;
  assign n13139 = n13138 ^ x29;
  assign n13290 = n13289 ^ n13139;
  assign n13124 = n1969 & n7393;
  assign n13125 = x114 & n1978;
  assign n13126 = x116 & n2108;
  assign n13127 = ~n13125 & ~n13126;
  assign n13128 = x115 & n1973;
  assign n13129 = n13127 & ~n13128;
  assign n13130 = ~n13124 & n13129;
  assign n13131 = n13130 ^ x26;
  assign n13291 = n13290 ^ n13131;
  assign n13121 = n13058 ^ n12901;
  assign n13122 = n13059 & n13121;
  assign n13123 = n13122 ^ n12901;
  assign n13292 = n13291 ^ n13123;
  assign n13113 = n1624 & n8169;
  assign n13114 = x117 & n1742;
  assign n13115 = x119 & n1744;
  assign n13116 = ~n13114 & ~n13115;
  assign n13117 = x118 & n1628;
  assign n13118 = n13116 & ~n13117;
  assign n13119 = ~n13113 & n13118;
  assign n13120 = n13119 ^ x23;
  assign n13293 = n13292 ^ n13120;
  assign n13110 = n13060 ^ n12890;
  assign n13111 = ~n13061 & ~n13110;
  assign n13112 = n13111 ^ n12890;
  assign n13294 = n13293 ^ n13112;
  assign n13102 = n1296 & n9001;
  assign n13103 = x121 & n1300;
  assign n13104 = x120 & n1403;
  assign n13105 = ~n13103 & ~n13104;
  assign n13106 = x122 & n1406;
  assign n13107 = n13105 & ~n13106;
  assign n13108 = ~n13102 & n13107;
  assign n13109 = n13108 ^ x20;
  assign n13295 = n13294 ^ n13109;
  assign n13099 = n13062 ^ n12879;
  assign n13100 = n13063 & n13099;
  assign n13101 = n13100 ^ n12879;
  assign n13296 = n13295 ^ n13101;
  assign n13091 = n1008 & n9912;
  assign n13092 = x124 & n1012;
  assign n13093 = x123 & n1101;
  assign n13094 = ~n13092 & ~n13093;
  assign n13095 = x125 & n1104;
  assign n13096 = n13094 & ~n13095;
  assign n13097 = ~n13091 & n13096;
  assign n13098 = n13097 ^ x17;
  assign n13297 = n13296 ^ n13098;
  assign n13088 = n13064 ^ n12868;
  assign n13089 = ~n13065 & ~n13088;
  assign n13090 = n13089 ^ n12868;
  assign n13298 = n13297 ^ n13090;
  assign n13082 = n752 & ~n9889;
  assign n13083 = x126 & n825;
  assign n13084 = x127 & n757;
  assign n13085 = ~n13083 & ~n13084;
  assign n13086 = ~n13082 & n13085;
  assign n13087 = n13086 ^ x14;
  assign n13299 = n13298 ^ n13087;
  assign n13079 = n13066 ^ n12857;
  assign n13080 = n13067 & n13079;
  assign n13081 = n13080 ^ n12857;
  assign n13300 = n13299 ^ n13081;
  assign n13076 = n13068 ^ n12846;
  assign n13077 = ~n13069 & ~n13076;
  assign n13078 = n13077 ^ n12846;
  assign n13301 = n13300 ^ n13078;
  assign n13073 = n12843 ^ n12840;
  assign n13074 = n13071 & n13073;
  assign n13075 = n13074 ^ n12840;
  assign n13302 = n13301 ^ n13075;
  assign n13510 = n2836 & n6178;
  assign n13511 = x109 & n2996;
  assign n13512 = x110 & n2840;
  assign n13513 = ~n13511 & ~n13512;
  assign n13514 = x111 & n2998;
  assign n13515 = n13513 & ~n13514;
  assign n13516 = ~n13510 & n13515;
  assign n13517 = n13516 ^ x32;
  assign n13500 = n3330 & ~n5506;
  assign n13501 = x106 & n3500;
  assign n13502 = x107 & n3334;
  assign n13503 = ~n13501 & ~n13502;
  assign n13504 = x108 & n3502;
  assign n13505 = n13503 & ~n13504;
  assign n13506 = ~n13500 & n13505;
  assign n13507 = n13506 ^ x35;
  assign n13490 = n3829 & n4867;
  assign n13491 = x103 & n4049;
  assign n13492 = x105 & n4052;
  assign n13493 = ~n13491 & ~n13492;
  assign n13494 = x104 & n3833;
  assign n13495 = n13493 & ~n13494;
  assign n13496 = ~n13490 & n13495;
  assign n13497 = n13496 ^ x38;
  assign n13480 = n4286 & n4415;
  assign n13481 = x100 & n4420;
  assign n13482 = x102 & n4614;
  assign n13483 = ~n13481 & ~n13482;
  assign n13484 = x101 & n4410;
  assign n13485 = n13483 & ~n13484;
  assign n13486 = ~n13480 & n13485;
  assign n13487 = n13486 ^ x41;
  assign n13469 = n3730 & n5010;
  assign n13470 = x97 & n5223;
  assign n13471 = x98 & n5014;
  assign n13472 = ~n13470 & ~n13471;
  assign n13473 = x99 & n5226;
  assign n13474 = n13472 & ~n13473;
  assign n13475 = ~n13469 & n13474;
  assign n13476 = n13475 ^ x44;
  assign n13459 = n3209 & n5656;
  assign n13460 = x94 & n5895;
  assign n13461 = x96 & n6111;
  assign n13462 = ~n13460 & ~n13461;
  assign n13463 = x95 & n5662;
  assign n13464 = n13462 & ~n13463;
  assign n13465 = ~n13459 & n13464;
  assign n13466 = n13465 ^ x47;
  assign n13449 = n2726 & n6326;
  assign n13450 = x91 & n6565;
  assign n13451 = x93 & n6569;
  assign n13452 = ~n13450 & ~n13451;
  assign n13453 = x92 & n6331;
  assign n13454 = n13452 & ~n13453;
  assign n13455 = ~n13449 & n13454;
  assign n13456 = n13455 ^ x50;
  assign n13439 = n2292 & n7076;
  assign n13440 = x88 & n7317;
  assign n13441 = x89 & n7080;
  assign n13442 = ~n13440 & ~n13441;
  assign n13443 = x90 & n7319;
  assign n13444 = n13442 & ~n13443;
  assign n13445 = ~n13439 & n13444;
  assign n13446 = n13445 ^ x53;
  assign n13436 = n13206 ^ n13195;
  assign n13437 = n13207 & ~n13436;
  assign n13438 = n13437 ^ n13198;
  assign n13447 = n13446 ^ n13438;
  assign n13426 = n1903 & n7830;
  assign n13427 = x85 & n7839;
  assign n13428 = x86 & n7834;
  assign n13429 = ~n13427 & ~n13428;
  assign n13430 = x87 & n8374;
  assign n13431 = n13429 & ~n13430;
  assign n13432 = ~n13426 & n13431;
  assign n13433 = n13432 ^ x56;
  assign n13417 = n1547 & n8622;
  assign n13418 = x82 & n8631;
  assign n13419 = x84 & n9186;
  assign n13420 = ~n13418 & ~n13419;
  assign n13421 = x83 & n8626;
  assign n13422 = n13420 & ~n13421;
  assign n13423 = ~n13417 & n13422;
  assign n13424 = n13423 ^ x59;
  assign n13408 = n1230 & n9499;
  assign n13409 = x79 & n9508;
  assign n13410 = x81 & n10106;
  assign n13411 = ~n13409 & ~n13410;
  assign n13412 = x80 & n9503;
  assign n13413 = n13411 & ~n13412;
  assign n13414 = ~n13408 & n13413;
  assign n13403 = x77 ^ x76;
  assign n13404 = n10099 & n13403;
  assign n13405 = n788 & n9798;
  assign n13406 = n13405 ^ x62;
  assign n13407 = ~n13404 & n13406;
  assign n13415 = n13414 ^ n13407;
  assign n13400 = n13184 ^ n13172;
  assign n13401 = n13176 & n13400;
  assign n13402 = n13401 ^ n13184;
  assign n13416 = n13415 ^ n13402;
  assign n13425 = n13424 ^ n13416;
  assign n13434 = n13433 ^ n13425;
  assign n13397 = n13193 ^ n13169;
  assign n13398 = n13194 & ~n13397;
  assign n13399 = n13398 ^ n13169;
  assign n13435 = n13434 ^ n13399;
  assign n13448 = n13447 ^ n13435;
  assign n13457 = n13456 ^ n13448;
  assign n13394 = n13208 ^ n13166;
  assign n13395 = n13217 & ~n13394;
  assign n13396 = n13395 ^ n13216;
  assign n13458 = n13457 ^ n13396;
  assign n13467 = n13466 ^ n13458;
  assign n13391 = n13218 ^ n13163;
  assign n13392 = n13227 & ~n13391;
  assign n13393 = n13392 ^ n13226;
  assign n13468 = n13467 ^ n13393;
  assign n13477 = n13476 ^ n13468;
  assign n13388 = n13228 ^ n13160;
  assign n13389 = n13237 & ~n13388;
  assign n13390 = n13389 ^ n13236;
  assign n13478 = n13477 ^ n13390;
  assign n13385 = n13238 ^ n13157;
  assign n13386 = n13247 & ~n13385;
  assign n13387 = n13386 ^ n13246;
  assign n13479 = n13478 ^ n13387;
  assign n13488 = n13487 ^ n13479;
  assign n13382 = n13257 ^ n13154;
  assign n13383 = ~n13249 & n13382;
  assign n13384 = n13383 ^ n13257;
  assign n13489 = n13488 ^ n13384;
  assign n13498 = n13497 ^ n13489;
  assign n13379 = n13267 ^ n13151;
  assign n13380 = ~n13259 & n13379;
  assign n13381 = n13380 ^ n13267;
  assign n13499 = n13498 ^ n13381;
  assign n13508 = n13507 ^ n13499;
  assign n13376 = n13277 ^ n13148;
  assign n13377 = ~n13269 & n13376;
  assign n13378 = n13377 ^ n13277;
  assign n13509 = n13508 ^ n13378;
  assign n13518 = n13517 ^ n13509;
  assign n13373 = n13286 ^ n13145;
  assign n13374 = ~n13287 & ~n13373;
  assign n13375 = n13374 ^ n13145;
  assign n13519 = n13518 ^ n13375;
  assign n13365 = n2371 & n6892;
  assign n13366 = x112 & n2528;
  assign n13367 = x114 & n2531;
  assign n13368 = ~n13366 & ~n13367;
  assign n13369 = x113 & n2377;
  assign n13370 = n13368 & ~n13369;
  assign n13371 = ~n13365 & n13370;
  assign n13372 = n13371 ^ x29;
  assign n13520 = n13519 ^ n13372;
  assign n13362 = n13288 ^ n13139;
  assign n13363 = n13289 & n13362;
  assign n13364 = n13363 ^ n13142;
  assign n13521 = n13520 ^ n13364;
  assign n13354 = n1969 & n7643;
  assign n13355 = x115 & n1978;
  assign n13356 = x116 & n1973;
  assign n13357 = ~n13355 & ~n13356;
  assign n13358 = x117 & n2108;
  assign n13359 = n13357 & ~n13358;
  assign n13360 = ~n13354 & n13359;
  assign n13361 = n13360 ^ x26;
  assign n13522 = n13521 ^ n13361;
  assign n13346 = n1624 & ~n8424;
  assign n13347 = x119 & n1628;
  assign n13348 = x118 & n1742;
  assign n13349 = ~n13347 & ~n13348;
  assign n13350 = x120 & n1744;
  assign n13351 = n13349 & ~n13350;
  assign n13352 = ~n13346 & n13351;
  assign n13353 = n13352 ^ x23;
  assign n13523 = n13522 ^ n13353;
  assign n13343 = n13290 ^ n13123;
  assign n13344 = ~n13291 & ~n13343;
  assign n13345 = n13344 ^ n13123;
  assign n13524 = n13523 ^ n13345;
  assign n13340 = n13292 ^ n13112;
  assign n13341 = n13293 & n13340;
  assign n13342 = n13341 ^ n13112;
  assign n13525 = n13524 ^ n13342;
  assign n13332 = n1296 & n9309;
  assign n13333 = x121 & n1403;
  assign n13334 = x123 & n1406;
  assign n13335 = ~n13333 & ~n13334;
  assign n13336 = x122 & n1300;
  assign n13337 = n13335 & ~n13336;
  assign n13338 = ~n13332 & n13337;
  assign n13339 = n13338 ^ x20;
  assign n13526 = n13525 ^ n13339;
  assign n13329 = n13294 ^ n13101;
  assign n13330 = ~n13295 & ~n13329;
  assign n13331 = n13330 ^ n13101;
  assign n13527 = n13526 ^ n13331;
  assign n13321 = n1008 & ~n10174;
  assign n13322 = x125 & n1012;
  assign n13323 = x124 & n1101;
  assign n13324 = ~n13322 & ~n13323;
  assign n13325 = x126 & n1104;
  assign n13326 = n13324 & ~n13325;
  assign n13327 = ~n13321 & n13326;
  assign n13328 = n13327 ^ x17;
  assign n13528 = n13527 ^ n13328;
  assign n13312 = n607 & n10430;
  assign n13313 = x127 & n754;
  assign n13314 = x14 & ~n13313;
  assign n13315 = ~n13312 & n13314;
  assign n13316 = ~x13 & ~n13315;
  assign n13317 = x127 & n744;
  assign n13318 = ~x14 & ~n13317;
  assign n13319 = ~n13312 & n13318;
  assign n13320 = ~n13316 & ~n13319;
  assign n13529 = n13528 ^ n13320;
  assign n13309 = n13296 ^ n13090;
  assign n13310 = n13297 & n13309;
  assign n13311 = n13310 ^ n13090;
  assign n13530 = n13529 ^ n13311;
  assign n13306 = n13298 ^ n13081;
  assign n13307 = ~n13299 & ~n13306;
  assign n13308 = n13307 ^ n13081;
  assign n13531 = n13530 ^ n13308;
  assign n13303 = n13078 ^ n13075;
  assign n13304 = ~n13301 & ~n13303;
  assign n13305 = n13304 ^ n13075;
  assign n13532 = n13531 ^ n13305;
  assign n13759 = n13320 & n13528;
  assign n13760 = n13311 & n13759;
  assign n13761 = ~n13308 & ~n13760;
  assign n13762 = n13528 ^ n13311;
  assign n13763 = ~n13529 & n13762;
  assign n13764 = n13763 ^ n13311;
  assign n13765 = ~n13761 & n13764;
  assign n13766 = ~n13305 & n13765;
  assign n13767 = ~n13320 & ~n13528;
  assign n13768 = ~n13311 & n13767;
  assign n13769 = n13768 ^ n13760;
  assign n13770 = ~n13308 & n13769;
  assign n13771 = n13770 ^ n13760;
  assign n13772 = ~n13766 & ~n13771;
  assign n13773 = n13308 & ~n13768;
  assign n13774 = ~n13764 & ~n13773;
  assign n13775 = n13305 & n13774;
  assign n13776 = n13772 & ~n13775;
  assign n13743 = n1969 & n7919;
  assign n13744 = x116 & n1978;
  assign n13745 = x117 & n1973;
  assign n13746 = ~n13744 & ~n13745;
  assign n13747 = x118 & n2108;
  assign n13748 = n13746 & ~n13747;
  assign n13749 = ~n13743 & n13748;
  assign n13750 = n13749 ^ x26;
  assign n13733 = n2371 & n7150;
  assign n13734 = x114 & n2377;
  assign n13735 = x113 & n2528;
  assign n13736 = ~n13734 & ~n13735;
  assign n13737 = x115 & n2531;
  assign n13738 = n13736 & ~n13737;
  assign n13739 = ~n13733 & n13738;
  assign n13740 = n13739 ^ x29;
  assign n13723 = n2836 & n6420;
  assign n13724 = x110 & n2996;
  assign n13725 = x111 & n2840;
  assign n13726 = ~n13724 & ~n13725;
  assign n13727 = x112 & n2998;
  assign n13728 = n13726 & ~n13727;
  assign n13729 = ~n13723 & n13728;
  assign n13730 = n13729 ^ x32;
  assign n13713 = n3330 & ~n5737;
  assign n13714 = x107 & n3500;
  assign n13715 = x109 & n3502;
  assign n13716 = ~n13714 & ~n13715;
  assign n13717 = x108 & n3334;
  assign n13718 = n13716 & ~n13717;
  assign n13719 = ~n13713 & n13718;
  assign n13720 = n13719 ^ x35;
  assign n13703 = n3829 & n5088;
  assign n13704 = x104 & n4049;
  assign n13705 = x106 & n4052;
  assign n13706 = ~n13704 & ~n13705;
  assign n13707 = x105 & n3833;
  assign n13708 = n13706 & ~n13707;
  assign n13709 = ~n13703 & n13708;
  assign n13710 = n13709 ^ x38;
  assign n13693 = n4415 & n4481;
  assign n13694 = x101 & n4420;
  assign n13695 = x102 & n4410;
  assign n13696 = ~n13694 & ~n13695;
  assign n13697 = x103 & n4614;
  assign n13698 = n13696 & ~n13697;
  assign n13699 = ~n13693 & n13698;
  assign n13700 = n13699 ^ x41;
  assign n13683 = n3925 & n5010;
  assign n13684 = x98 & n5223;
  assign n13685 = x100 & n5226;
  assign n13686 = ~n13684 & ~n13685;
  assign n13687 = x99 & n5014;
  assign n13688 = n13686 & ~n13687;
  assign n13689 = ~n13683 & n13688;
  assign n13690 = n13689 ^ x44;
  assign n13673 = n3388 & n5656;
  assign n13674 = x95 & n5895;
  assign n13675 = x97 & n6111;
  assign n13676 = ~n13674 & ~n13675;
  assign n13677 = x96 & n5662;
  assign n13678 = n13676 & ~n13677;
  assign n13679 = ~n13673 & n13678;
  assign n13680 = n13679 ^ x47;
  assign n13663 = n2895 & n6326;
  assign n13664 = x92 & n6565;
  assign n13665 = x94 & n6569;
  assign n13666 = ~n13664 & ~n13665;
  assign n13667 = x93 & n6331;
  assign n13668 = n13666 & ~n13667;
  assign n13669 = ~n13663 & n13668;
  assign n13670 = n13669 ^ x50;
  assign n13653 = n2447 & n7076;
  assign n13654 = x90 & n7080;
  assign n13655 = x89 & n7317;
  assign n13656 = ~n13654 & ~n13655;
  assign n13657 = x91 & n7319;
  assign n13658 = n13656 & ~n13657;
  assign n13659 = ~n13653 & n13658;
  assign n13660 = n13659 ^ x53;
  assign n13643 = n2040 & n7830;
  assign n13644 = x86 & n7839;
  assign n13645 = x87 & n7834;
  assign n13646 = ~n13644 & ~n13645;
  assign n13647 = x88 & n8374;
  assign n13648 = n13646 & ~n13647;
  assign n13649 = ~n13643 & n13648;
  assign n13650 = n13649 ^ x56;
  assign n13633 = n1674 & n8622;
  assign n13634 = x83 & n8631;
  assign n13635 = x84 & n8626;
  assign n13636 = ~n13634 & ~n13635;
  assign n13637 = x85 & n9186;
  assign n13638 = n13636 & ~n13637;
  assign n13639 = ~n13633 & n13638;
  assign n13640 = n13639 ^ x59;
  assign n13616 = ~n13403 & n13414;
  assign n13617 = ~x76 & x77;
  assign n13618 = n10099 & ~n13617;
  assign n13619 = ~n13616 & n13618;
  assign n13620 = x63 & n788;
  assign n13621 = ~n13414 & ~n13620;
  assign n13622 = ~x77 & x78;
  assign n13623 = x63 & n13622;
  assign n13624 = ~x62 & ~n13623;
  assign n13625 = ~n13621 & n13624;
  assign n13626 = ~n13619 & ~n13625;
  assign n13627 = ~n788 & n13414;
  assign n13628 = x62 & ~x63;
  assign n13629 = ~n13622 & n13628;
  assign n13630 = ~n13627 & n13629;
  assign n13631 = n13626 & ~n13630;
  assign n13607 = n1345 & n9499;
  assign n13608 = x80 & n9508;
  assign n13609 = x81 & n9503;
  assign n13610 = ~n13608 & ~n13609;
  assign n13611 = x82 & n10106;
  assign n13612 = n13610 & ~n13611;
  assign n13613 = ~n13607 & n13612;
  assign n13614 = n13613 ^ x62;
  assign n13602 = x79 & n9798;
  assign n13603 = x78 & n10099;
  assign n13604 = ~n13602 & ~n13603;
  assign n13605 = n13604 ^ x14;
  assign n13606 = n13605 ^ n13175;
  assign n13615 = n13614 ^ n13606;
  assign n13632 = n13631 ^ n13615;
  assign n13641 = n13640 ^ n13632;
  assign n13599 = n13424 ^ n13402;
  assign n13600 = n13416 & n13599;
  assign n13601 = n13600 ^ n13424;
  assign n13642 = n13641 ^ n13601;
  assign n13651 = n13650 ^ n13642;
  assign n13596 = n13425 ^ n13399;
  assign n13597 = ~n13434 & ~n13596;
  assign n13598 = n13597 ^ n13433;
  assign n13652 = n13651 ^ n13598;
  assign n13661 = n13660 ^ n13652;
  assign n13593 = n13438 ^ n13435;
  assign n13594 = n13447 & ~n13593;
  assign n13595 = n13594 ^ n13446;
  assign n13662 = n13661 ^ n13595;
  assign n13671 = n13670 ^ n13662;
  assign n13590 = n13448 ^ n13396;
  assign n13591 = n13457 & ~n13590;
  assign n13592 = n13591 ^ n13456;
  assign n13672 = n13671 ^ n13592;
  assign n13681 = n13680 ^ n13672;
  assign n13587 = n13458 ^ n13393;
  assign n13588 = n13467 & ~n13587;
  assign n13589 = n13588 ^ n13466;
  assign n13682 = n13681 ^ n13589;
  assign n13691 = n13690 ^ n13682;
  assign n13584 = n13468 ^ n13390;
  assign n13585 = n13477 & ~n13584;
  assign n13586 = n13585 ^ n13476;
  assign n13692 = n13691 ^ n13586;
  assign n13701 = n13700 ^ n13692;
  assign n13581 = n13487 ^ n13478;
  assign n13582 = ~n13479 & n13581;
  assign n13583 = n13582 ^ n13487;
  assign n13702 = n13701 ^ n13583;
  assign n13711 = n13710 ^ n13702;
  assign n13578 = n13497 ^ n13488;
  assign n13579 = ~n13489 & n13578;
  assign n13580 = n13579 ^ n13497;
  assign n13712 = n13711 ^ n13580;
  assign n13721 = n13720 ^ n13712;
  assign n13575 = n13507 ^ n13498;
  assign n13576 = ~n13499 & n13575;
  assign n13577 = n13576 ^ n13507;
  assign n13722 = n13721 ^ n13577;
  assign n13731 = n13730 ^ n13722;
  assign n13572 = n13517 ^ n13378;
  assign n13573 = ~n13509 & n13572;
  assign n13574 = n13573 ^ n13517;
  assign n13732 = n13731 ^ n13574;
  assign n13741 = n13740 ^ n13732;
  assign n13569 = n13518 ^ n13372;
  assign n13570 = ~n13519 & ~n13569;
  assign n13571 = n13570 ^ n13375;
  assign n13742 = n13741 ^ n13571;
  assign n13751 = n13750 ^ n13742;
  assign n13566 = n13520 ^ n13361;
  assign n13567 = n13521 & n13566;
  assign n13568 = n13567 ^ n13364;
  assign n13752 = n13751 ^ n13568;
  assign n13558 = n1624 & n8715;
  assign n13559 = x119 & n1742;
  assign n13560 = x120 & n1628;
  assign n13561 = ~n13559 & ~n13560;
  assign n13562 = x121 & n1744;
  assign n13563 = n13561 & ~n13562;
  assign n13564 = ~n13558 & n13563;
  assign n13565 = n13564 ^ x23;
  assign n13753 = n13752 ^ n13565;
  assign n13555 = n13522 ^ n13345;
  assign n13556 = ~n13523 & ~n13555;
  assign n13557 = n13556 ^ n13345;
  assign n13754 = n13753 ^ n13557;
  assign n13547 = n1296 & n9614;
  assign n13548 = x123 & n1300;
  assign n13549 = x122 & n1403;
  assign n13550 = ~n13548 & ~n13549;
  assign n13551 = x124 & n1406;
  assign n13552 = n13550 & ~n13551;
  assign n13553 = ~n13547 & n13552;
  assign n13554 = n13553 ^ x20;
  assign n13755 = n13754 ^ n13554;
  assign n13544 = n13524 ^ n13339;
  assign n13545 = n13525 & n13544;
  assign n13546 = n13545 ^ n13342;
  assign n13756 = n13755 ^ n13546;
  assign n13536 = n1008 & ~n10447;
  assign n13537 = x126 & n1012;
  assign n13538 = x125 & n1101;
  assign n13539 = ~n13537 & ~n13538;
  assign n13540 = x127 & n1104;
  assign n13541 = n13539 & ~n13540;
  assign n13542 = ~n13536 & n13541;
  assign n13543 = n13542 ^ x17;
  assign n13757 = n13756 ^ n13543;
  assign n13533 = n13526 ^ n13328;
  assign n13534 = ~n13527 & ~n13533;
  assign n13535 = n13534 ^ n13331;
  assign n13758 = n13757 ^ n13535;
  assign n13777 = n13776 ^ n13758;
  assign n13994 = ~n13308 & ~n13311;
  assign n13995 = ~n13305 & ~n13994;
  assign n13996 = n13308 & n13311;
  assign n13997 = ~n13758 & ~n13767;
  assign n13998 = ~n13996 & ~n13997;
  assign n13999 = ~n13995 & n13998;
  assign n14000 = ~n13767 & n13996;
  assign n14001 = n13758 & ~n14000;
  assign n14002 = ~n13305 & ~n14001;
  assign n14003 = ~n13758 & ~n13994;
  assign n14004 = ~n13759 & ~n14003;
  assign n14005 = ~n14002 & n14004;
  assign n14006 = ~n13999 & ~n14005;
  assign n13977 = n1969 & n8169;
  assign n13978 = x117 & n1978;
  assign n13979 = x118 & n1973;
  assign n13980 = ~n13978 & ~n13979;
  assign n13981 = x119 & n2108;
  assign n13982 = n13980 & ~n13981;
  assign n13983 = ~n13977 & n13982;
  assign n13984 = n13983 ^ x26;
  assign n13968 = n2371 & n7393;
  assign n13969 = x115 & n2377;
  assign n13970 = x114 & n2528;
  assign n13971 = ~n13969 & ~n13970;
  assign n13972 = x116 & n2531;
  assign n13973 = n13971 & ~n13972;
  assign n13974 = ~n13968 & n13973;
  assign n13975 = n13974 ^ x29;
  assign n13958 = n2836 & n6656;
  assign n13959 = x111 & n2996;
  assign n13960 = x112 & n2840;
  assign n13961 = ~n13959 & ~n13960;
  assign n13962 = x113 & n2998;
  assign n13963 = n13961 & ~n13962;
  assign n13964 = ~n13958 & n13963;
  assign n13965 = n13964 ^ x32;
  assign n13947 = n3330 & n5955;
  assign n13948 = x108 & n3500;
  assign n13949 = x110 & n3502;
  assign n13950 = ~n13948 & ~n13949;
  assign n13951 = x109 & n3334;
  assign n13952 = n13950 & ~n13951;
  assign n13953 = ~n13947 & n13952;
  assign n13954 = n13953 ^ x35;
  assign n13944 = n13710 ^ n13580;
  assign n13945 = n13711 & n13944;
  assign n13946 = n13945 ^ n13580;
  assign n13955 = n13954 ^ n13946;
  assign n13935 = n3829 & n5297;
  assign n13936 = x105 & n4049;
  assign n13937 = x106 & n3833;
  assign n13938 = ~n13936 & ~n13937;
  assign n13939 = x107 & n4052;
  assign n13940 = n13938 & ~n13939;
  assign n13941 = ~n13935 & n13940;
  assign n13942 = n13941 ^ x38;
  assign n13925 = n4415 & n4670;
  assign n13926 = x102 & n4420;
  assign n13927 = x103 & n4410;
  assign n13928 = ~n13926 & ~n13927;
  assign n13929 = x104 & n4614;
  assign n13930 = n13928 & ~n13929;
  assign n13931 = ~n13925 & n13930;
  assign n13932 = n13931 ^ x41;
  assign n13914 = n4105 & n5010;
  assign n13915 = x99 & n5223;
  assign n13916 = x101 & n5226;
  assign n13917 = ~n13915 & ~n13916;
  assign n13918 = x100 & n5014;
  assign n13919 = n13917 & ~n13918;
  assign n13920 = ~n13914 & n13919;
  assign n13921 = n13920 ^ x44;
  assign n13911 = n13680 ^ n13589;
  assign n13912 = n13681 & n13911;
  assign n13913 = n13912 ^ n13589;
  assign n13922 = n13921 ^ n13913;
  assign n13901 = n3556 & n5656;
  assign n13902 = x96 & n5895;
  assign n13903 = x98 & n6111;
  assign n13904 = ~n13902 & ~n13903;
  assign n13905 = x97 & n5662;
  assign n13906 = n13904 & ~n13905;
  assign n13907 = ~n13901 & n13906;
  assign n13908 = n13907 ^ x47;
  assign n13891 = n3054 & n6326;
  assign n13892 = x93 & n6565;
  assign n13893 = x94 & n6331;
  assign n13894 = ~n13892 & ~n13893;
  assign n13895 = x95 & n6569;
  assign n13896 = n13894 & ~n13895;
  assign n13897 = ~n13891 & n13896;
  assign n13898 = n13897 ^ x50;
  assign n13881 = n2585 & n7076;
  assign n13882 = x91 & n7080;
  assign n13883 = x90 & n7317;
  assign n13884 = ~n13882 & ~n13883;
  assign n13885 = x92 & n7319;
  assign n13886 = n13884 & ~n13885;
  assign n13887 = ~n13881 & n13886;
  assign n13888 = n13887 ^ x53;
  assign n13878 = n13650 ^ n13598;
  assign n13879 = n13651 & n13878;
  assign n13880 = n13879 ^ n13598;
  assign n13889 = n13888 ^ n13880;
  assign n13868 = n2164 & n7830;
  assign n13869 = x87 & n7839;
  assign n13870 = x89 & n8374;
  assign n13871 = ~n13869 & ~n13870;
  assign n13872 = x88 & n7834;
  assign n13873 = n13871 & ~n13872;
  assign n13874 = ~n13868 & n13873;
  assign n13875 = n13874 ^ x56;
  assign n13865 = n13640 ^ n13601;
  assign n13866 = n13641 & n13865;
  assign n13867 = n13866 ^ n13601;
  assign n13876 = n13875 ^ n13867;
  assign n13855 = n1787 & n8622;
  assign n13856 = x84 & n8631;
  assign n13857 = x86 & n9186;
  assign n13858 = ~n13856 & ~n13857;
  assign n13859 = x85 & n8626;
  assign n13860 = n13858 & ~n13859;
  assign n13861 = ~n13855 & n13860;
  assign n13862 = n13861 ^ x59;
  assign n13847 = n1445 & n9499;
  assign n13848 = x81 & n9508;
  assign n13849 = x83 & n10106;
  assign n13850 = ~n13848 & ~n13849;
  assign n13851 = x82 & n9503;
  assign n13852 = n13850 & ~n13851;
  assign n13853 = ~n13847 & n13852;
  assign n13842 = n13175 ^ x14;
  assign n13843 = n13604 ^ n13175;
  assign n13844 = n13842 & ~n13843;
  assign n13845 = n13844 ^ x14;
  assign n13838 = x63 & x80;
  assign n13836 = ~x63 & n938;
  assign n13837 = n13836 ^ x79;
  assign n13839 = n13838 ^ n13837;
  assign n13840 = ~x62 & ~n13839;
  assign n13841 = n13840 ^ n13837;
  assign n13846 = n13845 ^ n13841;
  assign n13854 = n13853 ^ n13846;
  assign n13863 = n13862 ^ n13854;
  assign n13833 = n13631 ^ n13614;
  assign n13834 = ~n13615 & ~n13833;
  assign n13835 = n13834 ^ n13631;
  assign n13864 = n13863 ^ n13835;
  assign n13877 = n13876 ^ n13864;
  assign n13890 = n13889 ^ n13877;
  assign n13899 = n13898 ^ n13890;
  assign n13830 = n13660 ^ n13595;
  assign n13831 = n13661 & n13830;
  assign n13832 = n13831 ^ n13595;
  assign n13900 = n13899 ^ n13832;
  assign n13909 = n13908 ^ n13900;
  assign n13827 = n13670 ^ n13592;
  assign n13828 = n13671 & n13827;
  assign n13829 = n13828 ^ n13592;
  assign n13910 = n13909 ^ n13829;
  assign n13923 = n13922 ^ n13910;
  assign n13824 = n13690 ^ n13586;
  assign n13825 = n13691 & n13824;
  assign n13826 = n13825 ^ n13586;
  assign n13924 = n13923 ^ n13826;
  assign n13933 = n13932 ^ n13924;
  assign n13821 = n13692 ^ n13583;
  assign n13822 = ~n13701 & n13821;
  assign n13823 = n13822 ^ n13700;
  assign n13934 = n13933 ^ n13823;
  assign n13943 = n13942 ^ n13934;
  assign n13956 = n13955 ^ n13943;
  assign n13818 = n13720 ^ n13577;
  assign n13819 = n13721 & n13818;
  assign n13820 = n13819 ^ n13577;
  assign n13957 = n13956 ^ n13820;
  assign n13966 = n13965 ^ n13957;
  assign n13815 = n13730 ^ n13574;
  assign n13816 = n13731 & n13815;
  assign n13817 = n13816 ^ n13574;
  assign n13967 = n13966 ^ n13817;
  assign n13976 = n13975 ^ n13967;
  assign n13985 = n13984 ^ n13976;
  assign n13812 = n13740 ^ n13571;
  assign n13813 = n13741 & ~n13812;
  assign n13814 = n13813 ^ n13571;
  assign n13986 = n13985 ^ n13814;
  assign n13809 = n13750 ^ n13568;
  assign n13810 = ~n13751 & ~n13809;
  assign n13811 = n13810 ^ n13568;
  assign n13987 = n13986 ^ n13811;
  assign n13801 = n1624 & n9001;
  assign n13802 = x121 & n1628;
  assign n13803 = x120 & n1742;
  assign n13804 = ~n13802 & ~n13803;
  assign n13805 = x122 & n1744;
  assign n13806 = n13804 & ~n13805;
  assign n13807 = ~n13801 & n13806;
  assign n13808 = n13807 ^ x23;
  assign n13988 = n13987 ^ n13808;
  assign n13798 = n13752 ^ n13557;
  assign n13799 = n13753 & n13798;
  assign n13800 = n13799 ^ n13557;
  assign n13989 = n13988 ^ n13800;
  assign n13790 = n1296 & n9912;
  assign n13791 = x123 & n1403;
  assign n13792 = x124 & n1300;
  assign n13793 = ~n13791 & ~n13792;
  assign n13794 = x125 & n1406;
  assign n13795 = n13793 & ~n13794;
  assign n13796 = ~n13790 & n13795;
  assign n13797 = n13796 ^ x20;
  assign n13990 = n13989 ^ n13797;
  assign n13787 = n13754 ^ n13546;
  assign n13788 = ~n13755 & ~n13787;
  assign n13789 = n13788 ^ n13546;
  assign n13991 = n13990 ^ n13789;
  assign n13781 = n1008 & ~n9889;
  assign n13782 = x126 & n1101;
  assign n13783 = x127 & n1012;
  assign n13784 = ~n13782 & ~n13783;
  assign n13785 = ~n13781 & n13784;
  assign n13786 = n13785 ^ x17;
  assign n13992 = n13991 ^ n13786;
  assign n13778 = n13756 ^ n13535;
  assign n13779 = n13757 & n13778;
  assign n13780 = n13779 ^ n13535;
  assign n13993 = n13992 ^ n13780;
  assign n14007 = n14006 ^ n13993;
  assign n14224 = n13780 & n13789;
  assign n14225 = n13786 & ~n13990;
  assign n14231 = n14224 & ~n14225;
  assign n14227 = ~n13780 & ~n13789;
  assign n14228 = ~n13786 & n13990;
  assign n14232 = ~n14227 & n14228;
  assign n14233 = ~n14231 & ~n14232;
  assign n14226 = ~n14224 & n14225;
  assign n14229 = n14227 & ~n14228;
  assign n14230 = ~n14226 & ~n14229;
  assign n14234 = n14233 ^ n14230;
  assign n14235 = ~n14006 & n14234;
  assign n14236 = n14235 ^ n14233;
  assign n14237 = n13789 ^ n13780;
  assign n14238 = n13990 ^ n13786;
  assign n14239 = ~n13991 & n14238;
  assign n14240 = ~n14237 & n14239;
  assign n14241 = n14236 & ~n14240;
  assign n14213 = n834 & n10430;
  assign n14214 = x127 & n996;
  assign n14215 = x17 & ~n14214;
  assign n14216 = ~n14213 & n14215;
  assign n14217 = ~x16 & ~n14216;
  assign n14218 = x127 & n999;
  assign n14219 = ~x17 & ~n14218;
  assign n14220 = ~n14213 & n14219;
  assign n14221 = ~n14217 & ~n14220;
  assign n14204 = n1296 & ~n10174;
  assign n14205 = x124 & n1403;
  assign n14206 = x125 & n1300;
  assign n14207 = ~n14205 & ~n14206;
  assign n14208 = x126 & n1406;
  assign n14209 = n14207 & ~n14208;
  assign n14210 = ~n14204 & n14209;
  assign n14211 = n14210 ^ x20;
  assign n14194 = n1624 & n9309;
  assign n14195 = x122 & n1628;
  assign n14196 = x121 & n1742;
  assign n14197 = ~n14195 & ~n14196;
  assign n14198 = x123 & n1744;
  assign n14199 = n14197 & ~n14198;
  assign n14200 = ~n14194 & n14199;
  assign n14201 = n14200 ^ x23;
  assign n14184 = n1969 & ~n8424;
  assign n14185 = x118 & n1978;
  assign n14186 = x119 & n1973;
  assign n14187 = ~n14185 & ~n14186;
  assign n14188 = x120 & n2108;
  assign n14189 = n14187 & ~n14188;
  assign n14190 = ~n14184 & n14189;
  assign n14191 = n14190 ^ x26;
  assign n14174 = n2371 & n7643;
  assign n14175 = x115 & n2528;
  assign n14176 = x116 & n2377;
  assign n14177 = ~n14175 & ~n14176;
  assign n14178 = x117 & n2531;
  assign n14179 = n14177 & ~n14178;
  assign n14180 = ~n14174 & n14179;
  assign n14181 = n14180 ^ x29;
  assign n14164 = n2836 & n6892;
  assign n14165 = x113 & n2840;
  assign n14166 = x112 & n2996;
  assign n14167 = ~n14165 & ~n14166;
  assign n14168 = x114 & n2998;
  assign n14169 = n14167 & ~n14168;
  assign n14170 = ~n14164 & n14169;
  assign n14171 = n14170 ^ x32;
  assign n14154 = n3330 & n6178;
  assign n14155 = x109 & n3500;
  assign n14156 = x111 & n3502;
  assign n14157 = ~n14155 & ~n14156;
  assign n14158 = x110 & n3334;
  assign n14159 = n14157 & ~n14158;
  assign n14160 = ~n14154 & n14159;
  assign n14161 = n14160 ^ x35;
  assign n14144 = n3829 & ~n5506;
  assign n14145 = x106 & n4049;
  assign n14146 = x108 & n4052;
  assign n14147 = ~n14145 & ~n14146;
  assign n14148 = x107 & n3833;
  assign n14149 = n14147 & ~n14148;
  assign n14150 = ~n14144 & n14149;
  assign n14151 = n14150 ^ x38;
  assign n14134 = n4415 & n4867;
  assign n14135 = x103 & n4420;
  assign n14136 = x104 & n4410;
  assign n14137 = ~n14135 & ~n14136;
  assign n14138 = x105 & n4614;
  assign n14139 = n14137 & ~n14138;
  assign n14140 = ~n14134 & n14139;
  assign n14141 = n14140 ^ x41;
  assign n14123 = n4286 & n5010;
  assign n14124 = x100 & n5223;
  assign n14125 = x101 & n5014;
  assign n14126 = ~n14124 & ~n14125;
  assign n14127 = x102 & n5226;
  assign n14128 = n14126 & ~n14127;
  assign n14129 = ~n14123 & n14128;
  assign n14130 = n14129 ^ x44;
  assign n14113 = n3730 & n5656;
  assign n14114 = x97 & n5895;
  assign n14115 = x98 & n5662;
  assign n14116 = ~n14114 & ~n14115;
  assign n14117 = x99 & n6111;
  assign n14118 = n14116 & ~n14117;
  assign n14119 = ~n14113 & n14118;
  assign n14120 = n14119 ^ x47;
  assign n14110 = n13890 ^ n13832;
  assign n14111 = n13899 & ~n14110;
  assign n14112 = n14111 ^ n13898;
  assign n14121 = n14120 ^ n14112;
  assign n14100 = n3209 & n6326;
  assign n14101 = x94 & n6565;
  assign n14102 = x95 & n6331;
  assign n14103 = ~n14101 & ~n14102;
  assign n14104 = x96 & n6569;
  assign n14105 = n14103 & ~n14104;
  assign n14106 = ~n14100 & n14105;
  assign n14107 = n14106 ^ x50;
  assign n14090 = n2726 & n7076;
  assign n14091 = x91 & n7317;
  assign n14092 = x92 & n7080;
  assign n14093 = ~n14091 & ~n14092;
  assign n14094 = x93 & n7319;
  assign n14095 = n14093 & ~n14094;
  assign n14096 = ~n14090 & n14095;
  assign n14097 = n14096 ^ x53;
  assign n14081 = n2292 & n7830;
  assign n14082 = x88 & n7839;
  assign n14083 = x90 & n8374;
  assign n14084 = ~n14082 & ~n14083;
  assign n14085 = x89 & n7834;
  assign n14086 = n14084 & ~n14085;
  assign n14087 = ~n14081 & n14086;
  assign n14088 = n14087 ^ x56;
  assign n14071 = n1903 & n8622;
  assign n14072 = x85 & n8631;
  assign n14073 = x87 & n9186;
  assign n14074 = ~n14072 & ~n14073;
  assign n14075 = x86 & n8626;
  assign n14076 = n14074 & ~n14075;
  assign n14077 = ~n14071 & n14076;
  assign n14078 = n14077 ^ x59;
  assign n14059 = n13845 & n13853;
  assign n14060 = ~n13838 & ~n14059;
  assign n14061 = ~n13845 & ~n13853;
  assign n14062 = ~x62 & ~n14061;
  assign n14063 = ~n14060 & n14062;
  assign n14064 = ~n13837 & ~n13845;
  assign n14065 = x62 & ~n14064;
  assign n14066 = n13837 & n14059;
  assign n14067 = n14066 ^ n13853;
  assign n14068 = n14065 & ~n14067;
  assign n14069 = ~n14063 & ~n14068;
  assign n14051 = n1547 & n9499;
  assign n14052 = x82 & n9508;
  assign n14053 = x84 & n10106;
  assign n14054 = ~n14052 & ~n14053;
  assign n14055 = x83 & n9503;
  assign n14056 = n14054 & ~n14055;
  assign n14057 = ~n14051 & n14056;
  assign n14047 = n938 & n10099;
  assign n14048 = n1043 & n9798;
  assign n14049 = n14048 ^ x62;
  assign n14050 = ~n14047 & n14049;
  assign n14058 = n14057 ^ n14050;
  assign n14070 = n14069 ^ n14058;
  assign n14079 = n14078 ^ n14070;
  assign n14044 = n13854 ^ n13835;
  assign n14045 = ~n13863 & ~n14044;
  assign n14046 = n14045 ^ n13862;
  assign n14080 = n14079 ^ n14046;
  assign n14089 = n14088 ^ n14080;
  assign n14098 = n14097 ^ n14089;
  assign n14041 = n13867 ^ n13864;
  assign n14042 = n13876 & ~n14041;
  assign n14043 = n14042 ^ n13875;
  assign n14099 = n14098 ^ n14043;
  assign n14108 = n14107 ^ n14099;
  assign n14038 = n13888 ^ n13877;
  assign n14039 = n13889 & ~n14038;
  assign n14040 = n14039 ^ n13880;
  assign n14109 = n14108 ^ n14040;
  assign n14122 = n14121 ^ n14109;
  assign n14131 = n14130 ^ n14122;
  assign n14035 = n13900 ^ n13829;
  assign n14036 = n13909 & ~n14035;
  assign n14037 = n14036 ^ n13908;
  assign n14132 = n14131 ^ n14037;
  assign n14032 = n13913 ^ n13910;
  assign n14033 = n13922 & ~n14032;
  assign n14034 = n14033 ^ n13921;
  assign n14133 = n14132 ^ n14034;
  assign n14142 = n14141 ^ n14133;
  assign n14029 = n13932 ^ n13826;
  assign n14030 = ~n13924 & n14029;
  assign n14031 = n14030 ^ n13932;
  assign n14143 = n14142 ^ n14031;
  assign n14152 = n14151 ^ n14143;
  assign n14026 = n13942 ^ n13823;
  assign n14027 = ~n13934 & n14026;
  assign n14028 = n14027 ^ n13942;
  assign n14153 = n14152 ^ n14028;
  assign n14162 = n14161 ^ n14153;
  assign n14023 = n13954 ^ n13943;
  assign n14024 = n13955 & ~n14023;
  assign n14025 = n14024 ^ n13946;
  assign n14163 = n14162 ^ n14025;
  assign n14172 = n14171 ^ n14163;
  assign n14020 = n13965 ^ n13956;
  assign n14021 = ~n13957 & n14020;
  assign n14022 = n14021 ^ n13965;
  assign n14173 = n14172 ^ n14022;
  assign n14182 = n14181 ^ n14173;
  assign n14017 = n13975 ^ n13817;
  assign n14018 = ~n13967 & n14017;
  assign n14019 = n14018 ^ n13975;
  assign n14183 = n14182 ^ n14019;
  assign n14192 = n14191 ^ n14183;
  assign n14014 = n13984 ^ n13814;
  assign n14015 = ~n13985 & ~n14014;
  assign n14016 = n14015 ^ n13814;
  assign n14193 = n14192 ^ n14016;
  assign n14202 = n14201 ^ n14193;
  assign n14011 = n13986 ^ n13808;
  assign n14012 = n13987 & n14011;
  assign n14013 = n14012 ^ n13811;
  assign n14203 = n14202 ^ n14013;
  assign n14212 = n14211 ^ n14203;
  assign n14222 = n14221 ^ n14212;
  assign n14008 = n13988 ^ n13797;
  assign n14009 = ~n13989 & ~n14008;
  assign n14010 = n14009 ^ n13800;
  assign n14223 = n14222 ^ n14010;
  assign n14242 = n14241 ^ n14223;
  assign n14460 = ~n14006 & ~n14228;
  assign n14461 = n14223 & ~n14224;
  assign n14462 = ~n14225 & ~n14461;
  assign n14463 = ~n14460 & n14462;
  assign n14464 = ~n14223 & ~n14226;
  assign n14465 = ~n14006 & ~n14464;
  assign n14466 = n14223 & ~n14228;
  assign n14467 = ~n14227 & ~n14466;
  assign n14468 = ~n14465 & n14467;
  assign n14469 = ~n14463 & ~n14468;
  assign n14449 = n1296 & ~n10447;
  assign n14450 = x126 & n1300;
  assign n14451 = x125 & n1403;
  assign n14452 = ~n14450 & ~n14451;
  assign n14453 = x127 & n1406;
  assign n14454 = n14452 & ~n14453;
  assign n14455 = ~n14449 & n14454;
  assign n14456 = n14455 ^ x20;
  assign n14439 = n1624 & n9614;
  assign n14440 = x123 & n1628;
  assign n14441 = x122 & n1742;
  assign n14442 = ~n14440 & ~n14441;
  assign n14443 = x124 & n1744;
  assign n14444 = n14442 & ~n14443;
  assign n14445 = ~n14439 & n14444;
  assign n14446 = n14445 ^ x23;
  assign n14427 = n2371 & n7919;
  assign n14428 = x116 & n2528;
  assign n14429 = x117 & n2377;
  assign n14430 = ~n14428 & ~n14429;
  assign n14431 = x118 & n2531;
  assign n14432 = n14430 & ~n14431;
  assign n14433 = ~n14427 & n14432;
  assign n14434 = n14433 ^ x29;
  assign n14417 = n2836 & n7150;
  assign n14418 = x113 & n2996;
  assign n14419 = x114 & n2840;
  assign n14420 = ~n14418 & ~n14419;
  assign n14421 = x115 & n2998;
  assign n14422 = n14420 & ~n14421;
  assign n14423 = ~n14417 & n14422;
  assign n14424 = n14423 ^ x32;
  assign n14407 = n3330 & n6420;
  assign n14408 = x110 & n3500;
  assign n14409 = x112 & n3502;
  assign n14410 = ~n14408 & ~n14409;
  assign n14411 = x111 & n3334;
  assign n14412 = n14410 & ~n14411;
  assign n14413 = ~n14407 & n14412;
  assign n14414 = n14413 ^ x35;
  assign n14397 = n3829 & ~n5737;
  assign n14398 = x107 & n4049;
  assign n14399 = x108 & n3833;
  assign n14400 = ~n14398 & ~n14399;
  assign n14401 = x109 & n4052;
  assign n14402 = n14400 & ~n14401;
  assign n14403 = ~n14397 & n14402;
  assign n14404 = n14403 ^ x38;
  assign n14387 = n4415 & n5088;
  assign n14388 = x104 & n4420;
  assign n14389 = x105 & n4410;
  assign n14390 = ~n14388 & ~n14389;
  assign n14391 = x106 & n4614;
  assign n14392 = n14390 & ~n14391;
  assign n14393 = ~n14387 & n14392;
  assign n14394 = n14393 ^ x41;
  assign n14377 = n4481 & n5010;
  assign n14378 = x101 & n5223;
  assign n14379 = x103 & n5226;
  assign n14380 = ~n14378 & ~n14379;
  assign n14381 = x102 & n5014;
  assign n14382 = n14380 & ~n14381;
  assign n14383 = ~n14377 & n14382;
  assign n14384 = n14383 ^ x44;
  assign n14367 = n3925 & n5656;
  assign n14368 = x98 & n5895;
  assign n14369 = x99 & n5662;
  assign n14370 = ~n14368 & ~n14369;
  assign n14371 = x100 & n6111;
  assign n14372 = n14370 & ~n14371;
  assign n14373 = ~n14367 & n14372;
  assign n14374 = n14373 ^ x47;
  assign n14357 = n3388 & n6326;
  assign n14358 = x96 & n6331;
  assign n14359 = x95 & n6565;
  assign n14360 = ~n14358 & ~n14359;
  assign n14361 = x97 & n6569;
  assign n14362 = n14360 & ~n14361;
  assign n14363 = ~n14357 & n14362;
  assign n14364 = n14363 ^ x50;
  assign n14347 = n2895 & n7076;
  assign n14348 = x93 & n7080;
  assign n14349 = x92 & n7317;
  assign n14350 = ~n14348 & ~n14349;
  assign n14351 = x94 & n7319;
  assign n14352 = n14350 & ~n14351;
  assign n14353 = ~n14347 & n14352;
  assign n14354 = n14353 ^ x53;
  assign n14335 = n2040 & n8622;
  assign n14336 = x86 & n8631;
  assign n14337 = x87 & n8626;
  assign n14338 = ~n14336 & ~n14337;
  assign n14339 = x88 & n9186;
  assign n14340 = n14338 & ~n14339;
  assign n14341 = ~n14335 & n14340;
  assign n14342 = n14341 ^ x59;
  assign n14332 = n14078 ^ n14069;
  assign n14333 = ~n14070 & ~n14332;
  assign n14334 = n14333 ^ n14078;
  assign n14343 = n14342 ^ n14334;
  assign n14314 = ~n938 & n14057;
  assign n14315 = x79 & ~x80;
  assign n14316 = n10099 & ~n14315;
  assign n14317 = ~n14314 & n14316;
  assign n14318 = ~x80 & x81;
  assign n14319 = ~x62 & x63;
  assign n14320 = n14318 & n14319;
  assign n14321 = ~n14317 & ~n14320;
  assign n14322 = n14057 & ~n14318;
  assign n14323 = x80 & ~x81;
  assign n14324 = n13628 & ~n14323;
  assign n14325 = ~n14322 & n14324;
  assign n14326 = x63 & n14323;
  assign n14327 = ~x62 & ~n14326;
  assign n14328 = n14057 & n14327;
  assign n14329 = ~n14325 & ~n14328;
  assign n14330 = n14321 & n14329;
  assign n14305 = n1674 & n9499;
  assign n14306 = x83 & n9508;
  assign n14307 = x85 & n10106;
  assign n14308 = ~n14306 & ~n14307;
  assign n14309 = x84 & n9503;
  assign n14310 = n14308 & ~n14309;
  assign n14311 = ~n14305 & n14310;
  assign n14312 = n14311 ^ x62;
  assign n14301 = n1126 & n9798;
  assign n14302 = n1043 & n10099;
  assign n14303 = ~n14301 & ~n14302;
  assign n14304 = n14303 ^ x17;
  assign n14313 = n14312 ^ n14304;
  assign n14331 = n14330 ^ n14313;
  assign n14344 = n14343 ^ n14331;
  assign n14293 = n2447 & n7830;
  assign n14294 = x89 & n7839;
  assign n14295 = x91 & n8374;
  assign n14296 = ~n14294 & ~n14295;
  assign n14297 = x90 & n7834;
  assign n14298 = n14296 & ~n14297;
  assign n14299 = ~n14293 & n14298;
  assign n14300 = n14299 ^ x56;
  assign n14345 = n14344 ^ n14300;
  assign n14290 = n14088 ^ n14046;
  assign n14291 = ~n14080 & n14290;
  assign n14292 = n14291 ^ n14088;
  assign n14346 = n14345 ^ n14292;
  assign n14355 = n14354 ^ n14346;
  assign n14287 = n14089 ^ n14043;
  assign n14288 = n14098 & ~n14287;
  assign n14289 = n14288 ^ n14097;
  assign n14356 = n14355 ^ n14289;
  assign n14365 = n14364 ^ n14356;
  assign n14284 = n14099 ^ n14040;
  assign n14285 = n14108 & ~n14284;
  assign n14286 = n14285 ^ n14107;
  assign n14366 = n14365 ^ n14286;
  assign n14375 = n14374 ^ n14366;
  assign n14281 = n14112 ^ n14109;
  assign n14282 = n14121 & ~n14281;
  assign n14283 = n14282 ^ n14120;
  assign n14376 = n14375 ^ n14283;
  assign n14385 = n14384 ^ n14376;
  assign n14278 = n14122 ^ n14037;
  assign n14279 = n14131 & ~n14278;
  assign n14280 = n14279 ^ n14130;
  assign n14386 = n14385 ^ n14280;
  assign n14395 = n14394 ^ n14386;
  assign n14275 = n14141 ^ n14034;
  assign n14276 = ~n14133 & n14275;
  assign n14277 = n14276 ^ n14141;
  assign n14396 = n14395 ^ n14277;
  assign n14405 = n14404 ^ n14396;
  assign n14272 = n14151 ^ n14142;
  assign n14273 = ~n14143 & n14272;
  assign n14274 = n14273 ^ n14151;
  assign n14406 = n14405 ^ n14274;
  assign n14415 = n14414 ^ n14406;
  assign n14269 = n14161 ^ n14028;
  assign n14270 = ~n14153 & n14269;
  assign n14271 = n14270 ^ n14161;
  assign n14416 = n14415 ^ n14271;
  assign n14425 = n14424 ^ n14416;
  assign n14266 = n14171 ^ n14162;
  assign n14267 = ~n14163 & n14266;
  assign n14268 = n14267 ^ n14171;
  assign n14426 = n14425 ^ n14268;
  assign n14435 = n14434 ^ n14426;
  assign n14263 = n14181 ^ n14172;
  assign n14264 = ~n14173 & n14263;
  assign n14265 = n14264 ^ n14181;
  assign n14436 = n14435 ^ n14265;
  assign n14260 = n14191 ^ n14182;
  assign n14261 = ~n14183 & n14260;
  assign n14262 = n14261 ^ n14191;
  assign n14437 = n14436 ^ n14262;
  assign n14252 = n1969 & n8715;
  assign n14253 = x119 & n1978;
  assign n14254 = x120 & n1973;
  assign n14255 = ~n14253 & ~n14254;
  assign n14256 = x121 & n2108;
  assign n14257 = n14255 & ~n14256;
  assign n14258 = ~n14252 & n14257;
  assign n14259 = n14258 ^ x26;
  assign n14438 = n14437 ^ n14259;
  assign n14447 = n14446 ^ n14438;
  assign n14249 = n14201 ^ n14016;
  assign n14250 = n14193 & ~n14249;
  assign n14251 = n14250 ^ n14201;
  assign n14448 = n14447 ^ n14251;
  assign n14457 = n14456 ^ n14448;
  assign n14246 = n14211 ^ n14013;
  assign n14247 = ~n14203 & ~n14246;
  assign n14248 = n14247 ^ n14211;
  assign n14458 = n14457 ^ n14248;
  assign n14243 = n14221 ^ n14010;
  assign n14244 = n14222 & n14243;
  assign n14245 = n14244 ^ n14010;
  assign n14459 = n14458 ^ n14245;
  assign n14470 = n14469 ^ n14459;
  assign n14672 = n14245 & ~n14248;
  assign n14673 = ~n14456 & n14672;
  assign n14674 = n14448 & ~n14673;
  assign n14675 = n14456 ^ n14245;
  assign n14676 = n14456 ^ n14248;
  assign n14677 = ~n14675 & ~n14676;
  assign n14678 = n14677 ^ n14245;
  assign n14679 = ~n14674 & n14678;
  assign n14680 = ~n14469 & n14679;
  assign n14681 = ~n14245 & n14248;
  assign n14682 = n14456 & n14681;
  assign n14683 = ~n14673 & ~n14682;
  assign n14684 = ~n14457 & ~n14683;
  assign n14685 = ~n14680 & ~n14684;
  assign n14686 = ~n14448 & ~n14682;
  assign n14687 = ~n14678 & ~n14686;
  assign n14688 = n14469 & n14687;
  assign n14689 = n14685 & ~n14688;
  assign n14661 = n1624 & n9912;
  assign n14662 = x124 & n1628;
  assign n14663 = x123 & n1742;
  assign n14664 = ~n14662 & ~n14663;
  assign n14665 = x125 & n1744;
  assign n14666 = n14664 & ~n14665;
  assign n14667 = ~n14661 & n14666;
  assign n14668 = n14667 ^ x23;
  assign n14651 = n1969 & n9001;
  assign n14652 = x120 & n1978;
  assign n14653 = x121 & n1973;
  assign n14654 = ~n14652 & ~n14653;
  assign n14655 = x122 & n2108;
  assign n14656 = n14654 & ~n14655;
  assign n14657 = ~n14651 & n14656;
  assign n14658 = n14657 ^ x26;
  assign n14640 = n2371 & n8169;
  assign n14641 = x117 & n2528;
  assign n14642 = x119 & n2531;
  assign n14643 = ~n14641 & ~n14642;
  assign n14644 = x118 & n2377;
  assign n14645 = n14643 & ~n14644;
  assign n14646 = ~n14640 & n14645;
  assign n14647 = n14646 ^ x29;
  assign n14631 = n2836 & n7393;
  assign n14632 = x114 & n2996;
  assign n14633 = x115 & n2840;
  assign n14634 = ~n14632 & ~n14633;
  assign n14635 = x116 & n2998;
  assign n14636 = n14634 & ~n14635;
  assign n14637 = ~n14631 & n14636;
  assign n14638 = n14637 ^ x32;
  assign n14621 = n3330 & n6656;
  assign n14622 = x111 & n3500;
  assign n14623 = x113 & n3502;
  assign n14624 = ~n14622 & ~n14623;
  assign n14625 = x112 & n3334;
  assign n14626 = n14624 & ~n14625;
  assign n14627 = ~n14621 & n14626;
  assign n14628 = n14627 ^ x35;
  assign n14605 = n4105 & n5656;
  assign n14606 = x99 & n5895;
  assign n14607 = x101 & n6111;
  assign n14608 = ~n14606 & ~n14607;
  assign n14609 = x100 & n5662;
  assign n14610 = n14608 & ~n14609;
  assign n14611 = ~n14605 & n14610;
  assign n14612 = n14611 ^ x47;
  assign n14595 = n3556 & n6326;
  assign n14596 = x96 & n6565;
  assign n14597 = x98 & n6569;
  assign n14598 = ~n14596 & ~n14597;
  assign n14599 = x97 & n6331;
  assign n14600 = n14598 & ~n14599;
  assign n14601 = ~n14595 & n14600;
  assign n14602 = n14601 ^ x50;
  assign n14585 = n3054 & n7076;
  assign n14586 = x93 & n7317;
  assign n14587 = x94 & n7080;
  assign n14588 = ~n14586 & ~n14587;
  assign n14589 = x95 & n7319;
  assign n14590 = n14588 & ~n14589;
  assign n14591 = ~n14585 & n14590;
  assign n14592 = n14591 ^ x53;
  assign n14574 = n2585 & n7830;
  assign n14575 = x90 & n7839;
  assign n14576 = x91 & n7834;
  assign n14577 = ~n14575 & ~n14576;
  assign n14578 = x92 & n8374;
  assign n14579 = n14577 & ~n14578;
  assign n14580 = ~n14574 & n14579;
  assign n14581 = n14580 ^ x56;
  assign n14571 = n14342 ^ n14331;
  assign n14572 = n14343 & ~n14571;
  assign n14573 = n14572 ^ n14334;
  assign n14582 = n14581 ^ n14573;
  assign n14561 = n2164 & n8622;
  assign n14562 = x88 & n8626;
  assign n14563 = x89 & n9186;
  assign n14564 = ~n14562 & ~n14563;
  assign n14565 = x87 & n8631;
  assign n14566 = n14564 & ~n14565;
  assign n14567 = ~n14561 & n14566;
  assign n14568 = n14567 ^ x59;
  assign n14552 = n1787 & n9499;
  assign n14553 = x84 & n9508;
  assign n14554 = x85 & n9503;
  assign n14555 = ~n14553 & ~n14554;
  assign n14556 = x86 & n10106;
  assign n14557 = n14555 & ~n14556;
  assign n14558 = ~n14552 & n14557;
  assign n14559 = n14558 ^ x62;
  assign n14543 = x80 & n10099;
  assign n14544 = ~x17 & x81;
  assign n14545 = ~n14543 & ~n14544;
  assign n14546 = x82 & ~n10099;
  assign n14547 = n14545 & ~n14546;
  assign n14548 = x17 & ~x81;
  assign n14549 = ~n12465 & ~n14548;
  assign n14550 = ~n14547 & n14549;
  assign n14540 = x83 & n9798;
  assign n14541 = x82 & n10099;
  assign n14542 = ~n14540 & ~n14541;
  assign n14551 = n14550 ^ n14542;
  assign n14560 = n14559 ^ n14551;
  assign n14569 = n14568 ^ n14560;
  assign n14537 = n14330 ^ n14312;
  assign n14538 = n14313 & ~n14537;
  assign n14539 = n14538 ^ n14330;
  assign n14570 = n14569 ^ n14539;
  assign n14583 = n14582 ^ n14570;
  assign n14534 = n14300 ^ n14292;
  assign n14535 = n14345 & ~n14534;
  assign n14536 = n14535 ^ n14344;
  assign n14584 = n14583 ^ n14536;
  assign n14593 = n14592 ^ n14584;
  assign n14531 = n14354 ^ n14289;
  assign n14532 = ~n14355 & n14531;
  assign n14533 = n14532 ^ n14289;
  assign n14594 = n14593 ^ n14533;
  assign n14603 = n14602 ^ n14594;
  assign n14528 = n14364 ^ n14286;
  assign n14529 = ~n14365 & n14528;
  assign n14530 = n14529 ^ n14286;
  assign n14604 = n14603 ^ n14530;
  assign n14613 = n14612 ^ n14604;
  assign n14525 = n14374 ^ n14283;
  assign n14526 = ~n14375 & n14525;
  assign n14527 = n14526 ^ n14283;
  assign n14614 = n14613 ^ n14527;
  assign n14517 = n4670 & n5010;
  assign n14518 = x102 & n5223;
  assign n14519 = x103 & n5014;
  assign n14520 = ~n14518 & ~n14519;
  assign n14521 = x104 & n5226;
  assign n14522 = n14520 & ~n14521;
  assign n14523 = ~n14517 & n14522;
  assign n14524 = n14523 ^ x44;
  assign n14615 = n14614 ^ n14524;
  assign n14514 = n14384 ^ n14280;
  assign n14515 = ~n14385 & n14514;
  assign n14516 = n14515 ^ n14280;
  assign n14616 = n14615 ^ n14516;
  assign n14506 = n4415 & n5297;
  assign n14507 = x105 & n4420;
  assign n14508 = x107 & n4614;
  assign n14509 = ~n14507 & ~n14508;
  assign n14510 = x106 & n4410;
  assign n14511 = n14509 & ~n14510;
  assign n14512 = ~n14506 & n14511;
  assign n14513 = n14512 ^ x41;
  assign n14617 = n14616 ^ n14513;
  assign n14503 = n14394 ^ n14277;
  assign n14504 = ~n14395 & n14503;
  assign n14505 = n14504 ^ n14277;
  assign n14618 = n14617 ^ n14505;
  assign n14495 = n3829 & n5955;
  assign n14496 = x108 & n4049;
  assign n14497 = x109 & n3833;
  assign n14498 = ~n14496 & ~n14497;
  assign n14499 = x110 & n4052;
  assign n14500 = n14498 & ~n14499;
  assign n14501 = ~n14495 & n14500;
  assign n14502 = n14501 ^ x38;
  assign n14619 = n14618 ^ n14502;
  assign n14492 = n14404 ^ n14274;
  assign n14493 = ~n14405 & n14492;
  assign n14494 = n14493 ^ n14274;
  assign n14620 = n14619 ^ n14494;
  assign n14629 = n14628 ^ n14620;
  assign n14489 = n14406 ^ n14271;
  assign n14490 = n14415 & ~n14489;
  assign n14491 = n14490 ^ n14414;
  assign n14630 = n14629 ^ n14491;
  assign n14639 = n14638 ^ n14630;
  assign n14648 = n14647 ^ n14639;
  assign n14486 = n14424 ^ n14268;
  assign n14487 = ~n14425 & n14486;
  assign n14488 = n14487 ^ n14268;
  assign n14649 = n14648 ^ n14488;
  assign n14483 = n14434 ^ n14265;
  assign n14484 = ~n14435 & n14483;
  assign n14485 = n14484 ^ n14265;
  assign n14650 = n14649 ^ n14485;
  assign n14659 = n14658 ^ n14650;
  assign n14480 = n14436 ^ n14259;
  assign n14481 = n14437 & ~n14480;
  assign n14482 = n14481 ^ n14262;
  assign n14660 = n14659 ^ n14482;
  assign n14669 = n14668 ^ n14660;
  assign n14477 = n14446 ^ n14251;
  assign n14478 = ~n14447 & n14477;
  assign n14479 = n14478 ^ n14251;
  assign n14670 = n14669 ^ n14479;
  assign n14471 = n1296 & ~n9889;
  assign n14472 = x127 & n1300;
  assign n14473 = x126 & n1403;
  assign n14474 = ~n14472 & ~n14473;
  assign n14475 = ~n14471 & n14474;
  assign n14476 = n14475 ^ x20;
  assign n14671 = n14670 ^ n14476;
  assign n14690 = n14689 ^ n14671;
  assign n14897 = n14448 & n14456;
  assign n14898 = ~n14469 & ~n14897;
  assign n14899 = n14671 & ~n14681;
  assign n14900 = ~n14448 & ~n14456;
  assign n14901 = ~n14899 & ~n14900;
  assign n14902 = ~n14898 & n14901;
  assign n14903 = ~n14681 & n14900;
  assign n14904 = ~n14671 & ~n14903;
  assign n14905 = ~n14469 & ~n14904;
  assign n14906 = n14671 & ~n14897;
  assign n14907 = ~n14672 & ~n14906;
  assign n14908 = ~n14905 & n14907;
  assign n14909 = ~n14902 & ~n14908;
  assign n14886 = n1624 & ~n10174;
  assign n14887 = x124 & n1742;
  assign n14888 = x125 & n1628;
  assign n14889 = ~n14887 & ~n14888;
  assign n14890 = x126 & n1744;
  assign n14891 = n14889 & ~n14890;
  assign n14892 = ~n14886 & n14891;
  assign n14893 = n14892 ^ x23;
  assign n14876 = n1969 & n9309;
  assign n14877 = x121 & n1978;
  assign n14878 = x122 & n1973;
  assign n14879 = ~n14877 & ~n14878;
  assign n14880 = x123 & n2108;
  assign n14881 = n14879 & ~n14880;
  assign n14882 = ~n14876 & n14881;
  assign n14883 = n14882 ^ x26;
  assign n14866 = n2371 & ~n8424;
  assign n14867 = x118 & n2528;
  assign n14868 = x119 & n2377;
  assign n14869 = ~n14867 & ~n14868;
  assign n14870 = x120 & n2531;
  assign n14871 = n14869 & ~n14870;
  assign n14872 = ~n14866 & n14871;
  assign n14873 = n14872 ^ x29;
  assign n14856 = n2836 & n7643;
  assign n14857 = x116 & n2840;
  assign n14858 = x115 & n2996;
  assign n14859 = ~n14857 & ~n14858;
  assign n14860 = x117 & n2998;
  assign n14861 = n14859 & ~n14860;
  assign n14862 = ~n14856 & n14861;
  assign n14863 = n14862 ^ x32;
  assign n14846 = n3330 & n6892;
  assign n14847 = x112 & n3500;
  assign n14848 = x114 & n3502;
  assign n14849 = ~n14847 & ~n14848;
  assign n14850 = x113 & n3334;
  assign n14851 = n14849 & ~n14850;
  assign n14852 = ~n14846 & n14851;
  assign n14853 = n14852 ^ x35;
  assign n14836 = n3829 & n6178;
  assign n14837 = x109 & n4049;
  assign n14838 = x111 & n4052;
  assign n14839 = ~n14837 & ~n14838;
  assign n14840 = x110 & n3833;
  assign n14841 = n14839 & ~n14840;
  assign n14842 = ~n14836 & n14841;
  assign n14843 = n14842 ^ x38;
  assign n14826 = n4415 & ~n5506;
  assign n14827 = x106 & n4420;
  assign n14828 = x108 & n4614;
  assign n14829 = ~n14827 & ~n14828;
  assign n14830 = x107 & n4410;
  assign n14831 = n14829 & ~n14830;
  assign n14832 = ~n14826 & n14831;
  assign n14833 = n14832 ^ x41;
  assign n14816 = n4867 & n5010;
  assign n14817 = x103 & n5223;
  assign n14818 = x104 & n5014;
  assign n14819 = ~n14817 & ~n14818;
  assign n14820 = x105 & n5226;
  assign n14821 = n14819 & ~n14820;
  assign n14822 = ~n14816 & n14821;
  assign n14823 = n14822 ^ x44;
  assign n14803 = n3730 & n6326;
  assign n14804 = x97 & n6565;
  assign n14805 = x99 & n6569;
  assign n14806 = ~n14804 & ~n14805;
  assign n14807 = x98 & n6331;
  assign n14808 = n14806 & ~n14807;
  assign n14809 = ~n14803 & n14808;
  assign n14810 = n14809 ^ x50;
  assign n14800 = n14592 ^ n14536;
  assign n14801 = n14584 & n14800;
  assign n14802 = n14801 ^ n14592;
  assign n14811 = n14810 ^ n14802;
  assign n14790 = n3209 & n7076;
  assign n14791 = x94 & n7317;
  assign n14792 = x96 & n7319;
  assign n14793 = ~n14791 & ~n14792;
  assign n14794 = x95 & n7080;
  assign n14795 = n14793 & ~n14794;
  assign n14796 = ~n14790 & n14795;
  assign n14797 = n14796 ^ x53;
  assign n14780 = n2726 & n7830;
  assign n14781 = x91 & n7839;
  assign n14782 = x92 & n7834;
  assign n14783 = ~n14781 & ~n14782;
  assign n14784 = x93 & n8374;
  assign n14785 = n14783 & ~n14784;
  assign n14786 = ~n14780 & n14785;
  assign n14787 = n14786 ^ x56;
  assign n14777 = n14560 ^ n14539;
  assign n14778 = n14569 & n14777;
  assign n14779 = n14778 ^ n14568;
  assign n14788 = n14787 ^ n14779;
  assign n14768 = n2292 & n8622;
  assign n14769 = x88 & n8631;
  assign n14770 = x89 & n8626;
  assign n14771 = ~n14769 & ~n14770;
  assign n14772 = x90 & n9186;
  assign n14773 = n14771 & ~n14772;
  assign n14774 = ~n14768 & n14773;
  assign n14775 = n14774 ^ x59;
  assign n14758 = n1903 & n9499;
  assign n14759 = x85 & n9508;
  assign n14760 = x86 & n9503;
  assign n14761 = ~n14759 & ~n14760;
  assign n14762 = x87 & n10106;
  assign n14763 = n14761 & ~n14762;
  assign n14764 = ~n14758 & n14763;
  assign n14765 = n14764 ^ x62;
  assign n14748 = ~x83 & n14541;
  assign n14749 = x83 & ~x84;
  assign n14750 = n9798 & n14749;
  assign n14751 = ~n14748 & ~n14750;
  assign n14752 = ~x83 & x84;
  assign n14753 = n9798 & n14752;
  assign n14754 = x83 & n10099;
  assign n14755 = ~x82 & n14754;
  assign n14756 = ~n14753 & ~n14755;
  assign n14757 = n14751 & n14756;
  assign n14766 = n14765 ^ n14757;
  assign n14745 = n14559 ^ n14550;
  assign n14746 = ~n14551 & ~n14745;
  assign n14747 = n14746 ^ n14559;
  assign n14767 = n14766 ^ n14747;
  assign n14776 = n14775 ^ n14767;
  assign n14789 = n14788 ^ n14776;
  assign n14798 = n14797 ^ n14789;
  assign n14742 = n14581 ^ n14570;
  assign n14743 = n14582 & n14742;
  assign n14744 = n14743 ^ n14573;
  assign n14799 = n14798 ^ n14744;
  assign n14812 = n14811 ^ n14799;
  assign n14739 = n14602 ^ n14533;
  assign n14740 = n14594 & n14739;
  assign n14741 = n14740 ^ n14602;
  assign n14813 = n14812 ^ n14741;
  assign n14731 = n4286 & n5656;
  assign n14732 = x101 & n5662;
  assign n14733 = x100 & n5895;
  assign n14734 = ~n14732 & ~n14733;
  assign n14735 = x102 & n6111;
  assign n14736 = n14734 & ~n14735;
  assign n14737 = ~n14731 & n14736;
  assign n14738 = n14737 ^ x47;
  assign n14814 = n14813 ^ n14738;
  assign n14728 = n14612 ^ n14530;
  assign n14729 = n14604 & n14728;
  assign n14730 = n14729 ^ n14612;
  assign n14815 = n14814 ^ n14730;
  assign n14824 = n14823 ^ n14815;
  assign n14725 = n14613 ^ n14524;
  assign n14726 = ~n14614 & n14725;
  assign n14727 = n14726 ^ n14527;
  assign n14825 = n14824 ^ n14727;
  assign n14834 = n14833 ^ n14825;
  assign n14722 = n14615 ^ n14513;
  assign n14723 = ~n14616 & n14722;
  assign n14724 = n14723 ^ n14516;
  assign n14835 = n14834 ^ n14724;
  assign n14844 = n14843 ^ n14835;
  assign n14719 = n14617 ^ n14502;
  assign n14720 = ~n14618 & n14719;
  assign n14721 = n14720 ^ n14505;
  assign n14845 = n14844 ^ n14721;
  assign n14854 = n14853 ^ n14845;
  assign n14716 = n14628 ^ n14619;
  assign n14717 = n14620 & ~n14716;
  assign n14718 = n14717 ^ n14628;
  assign n14855 = n14854 ^ n14718;
  assign n14864 = n14863 ^ n14855;
  assign n14713 = n14638 ^ n14491;
  assign n14714 = n14630 & n14713;
  assign n14715 = n14714 ^ n14638;
  assign n14865 = n14864 ^ n14715;
  assign n14874 = n14873 ^ n14865;
  assign n14710 = n14639 ^ n14488;
  assign n14711 = ~n14648 & n14710;
  assign n14712 = n14711 ^ n14647;
  assign n14875 = n14874 ^ n14712;
  assign n14884 = n14883 ^ n14875;
  assign n14707 = n14658 ^ n14485;
  assign n14708 = n14650 & n14707;
  assign n14709 = n14708 ^ n14658;
  assign n14885 = n14884 ^ n14709;
  assign n14894 = n14893 ^ n14885;
  assign n14704 = n14669 ^ n14476;
  assign n14705 = ~n14670 & n14704;
  assign n14706 = n14705 ^ n14479;
  assign n14895 = n14894 ^ n14706;
  assign n14694 = n1096 & n10430;
  assign n14695 = x127 & n1283;
  assign n14696 = x20 & ~n14695;
  assign n14697 = ~n14694 & n14696;
  assign n14698 = ~x19 & ~n14697;
  assign n14699 = x127 & n1287;
  assign n14700 = ~x20 & ~n14699;
  assign n14701 = ~n14694 & n14700;
  assign n14702 = ~n14698 & ~n14701;
  assign n14691 = n14668 ^ n14659;
  assign n14692 = n14660 & ~n14691;
  assign n14693 = n14692 ^ n14668;
  assign n14703 = n14702 ^ n14693;
  assign n14896 = n14895 ^ n14703;
  assign n14910 = n14909 ^ n14896;
  assign n15097 = ~n14693 & n14702;
  assign n15102 = n14706 & n14894;
  assign n15103 = ~n15097 & n15102;
  assign n15096 = n14693 & ~n14702;
  assign n15104 = ~n14706 & ~n14894;
  assign n15105 = n15096 & ~n15104;
  assign n15106 = ~n15103 & ~n15105;
  assign n15098 = n15097 ^ n14894;
  assign n15099 = n14895 & n15098;
  assign n15100 = n15099 ^ n14706;
  assign n15101 = ~n15096 & ~n15100;
  assign n15107 = n15106 ^ n15101;
  assign n15108 = n14909 & ~n15107;
  assign n15109 = n15108 ^ n15106;
  assign n15110 = n14894 ^ n14702;
  assign n15111 = n14703 & n15110;
  assign n15112 = ~n14895 & n15111;
  assign n15113 = n15109 & ~n15112;
  assign n15086 = n1624 & ~n10447;
  assign n15087 = x126 & n1628;
  assign n15088 = x125 & n1742;
  assign n15089 = ~n15087 & ~n15088;
  assign n15090 = x127 & n1744;
  assign n15091 = n15089 & ~n15090;
  assign n15092 = ~n15086 & n15091;
  assign n15093 = n15092 ^ x23;
  assign n15076 = n1969 & n9614;
  assign n15077 = x122 & n1978;
  assign n15078 = x123 & n1973;
  assign n15079 = ~n15077 & ~n15078;
  assign n15080 = x124 & n2108;
  assign n15081 = n15079 & ~n15080;
  assign n15082 = ~n15076 & n15081;
  assign n15083 = n15082 ^ x26;
  assign n15064 = n2836 & n7919;
  assign n15065 = x116 & n2996;
  assign n15066 = x117 & n2840;
  assign n15067 = ~n15065 & ~n15066;
  assign n15068 = x118 & n2998;
  assign n15069 = n15067 & ~n15068;
  assign n15070 = ~n15064 & n15069;
  assign n15071 = n15070 ^ x32;
  assign n15054 = n3330 & n7150;
  assign n15055 = x113 & n3500;
  assign n15056 = x114 & n3334;
  assign n15057 = ~n15055 & ~n15056;
  assign n15058 = x115 & n3502;
  assign n15059 = n15057 & ~n15058;
  assign n15060 = ~n15054 & n15059;
  assign n15061 = n15060 ^ x35;
  assign n15044 = n3829 & n6420;
  assign n15045 = x110 & n4049;
  assign n15046 = x112 & n4052;
  assign n15047 = ~n15045 & ~n15046;
  assign n15048 = x111 & n3833;
  assign n15049 = n15047 & ~n15048;
  assign n15050 = ~n15044 & n15049;
  assign n15051 = n15050 ^ x38;
  assign n15034 = n4415 & ~n5737;
  assign n15035 = x107 & n4420;
  assign n15036 = x108 & n4410;
  assign n15037 = ~n15035 & ~n15036;
  assign n15038 = x109 & n4614;
  assign n15039 = n15037 & ~n15038;
  assign n15040 = ~n15034 & n15039;
  assign n15041 = n15040 ^ x41;
  assign n15024 = n5010 & n5088;
  assign n15025 = x105 & n5014;
  assign n15026 = x104 & n5223;
  assign n15027 = ~n15025 & ~n15026;
  assign n15028 = x106 & n5226;
  assign n15029 = n15027 & ~n15028;
  assign n15030 = ~n15024 & n15029;
  assign n15031 = n15030 ^ x44;
  assign n15012 = n3925 & n6326;
  assign n15013 = x98 & n6565;
  assign n15014 = x100 & n6569;
  assign n15015 = ~n15013 & ~n15014;
  assign n15016 = x99 & n6331;
  assign n15017 = n15015 & ~n15016;
  assign n15018 = ~n15012 & n15017;
  assign n15019 = n15018 ^ x50;
  assign n15009 = n14802 ^ n14799;
  assign n15010 = n14811 & ~n15009;
  assign n15011 = n15010 ^ n14810;
  assign n15020 = n15019 ^ n15011;
  assign n14999 = n3388 & n7076;
  assign n15000 = x95 & n7317;
  assign n15001 = x96 & n7080;
  assign n15002 = ~n15000 & ~n15001;
  assign n15003 = x97 & n7319;
  assign n15004 = n15002 & ~n15003;
  assign n15005 = ~n14999 & n15004;
  assign n15006 = n15005 ^ x53;
  assign n14989 = n2895 & n7830;
  assign n14990 = x92 & n7839;
  assign n14991 = x93 & n7834;
  assign n14992 = ~n14990 & ~n14991;
  assign n14993 = x94 & n8374;
  assign n14994 = n14992 & ~n14993;
  assign n14995 = ~n14989 & n14994;
  assign n14996 = n14995 ^ x56;
  assign n14979 = n2447 & n8622;
  assign n14980 = x89 & n8631;
  assign n14981 = x90 & n8626;
  assign n14982 = ~n14980 & ~n14981;
  assign n14983 = x91 & n9186;
  assign n14984 = n14982 & ~n14983;
  assign n14985 = ~n14979 & n14984;
  assign n14986 = n14985 ^ x59;
  assign n14976 = n14775 ^ n14747;
  assign n14977 = ~n14767 & n14976;
  assign n14978 = n14977 ^ n14775;
  assign n14987 = n14986 ^ n14978;
  assign n14966 = n2040 & n9499;
  assign n14967 = x86 & n9508;
  assign n14968 = x88 & n10106;
  assign n14969 = ~n14967 & ~n14968;
  assign n14970 = x87 & n9503;
  assign n14971 = n14969 & ~n14970;
  assign n14972 = ~n14966 & n14971;
  assign n14973 = n14972 ^ x62;
  assign n14962 = n1334 & n10099;
  assign n14963 = n1434 & n9798;
  assign n14964 = ~n14962 & ~n14963;
  assign n14965 = n14964 ^ x20;
  assign n14974 = n14973 ^ n14965;
  assign n14960 = n14757 & ~n14765;
  assign n14961 = n14960 ^ n14751;
  assign n14975 = n14974 ^ n14961;
  assign n14988 = n14987 ^ n14975;
  assign n14997 = n14996 ^ n14988;
  assign n14957 = n14779 ^ n14776;
  assign n14958 = n14788 & ~n14957;
  assign n14959 = n14958 ^ n14787;
  assign n14998 = n14997 ^ n14959;
  assign n15007 = n15006 ^ n14998;
  assign n14954 = n14789 ^ n14744;
  assign n14955 = n14798 & ~n14954;
  assign n14956 = n14955 ^ n14797;
  assign n15008 = n15007 ^ n14956;
  assign n15021 = n15020 ^ n15008;
  assign n14951 = n14741 ^ n14738;
  assign n14952 = n14813 & ~n14951;
  assign n14953 = n14952 ^ n14812;
  assign n15022 = n15021 ^ n14953;
  assign n14943 = n4481 & n5656;
  assign n14944 = x101 & n5895;
  assign n14945 = x103 & n6111;
  assign n14946 = ~n14944 & ~n14945;
  assign n14947 = x102 & n5662;
  assign n14948 = n14946 & ~n14947;
  assign n14949 = ~n14943 & n14948;
  assign n14950 = n14949 ^ x47;
  assign n15023 = n15022 ^ n14950;
  assign n15032 = n15031 ^ n15023;
  assign n14940 = n14823 ^ n14814;
  assign n14941 = ~n14815 & n14940;
  assign n14942 = n14941 ^ n14823;
  assign n15033 = n15032 ^ n14942;
  assign n15042 = n15041 ^ n15033;
  assign n14937 = n14833 ^ n14727;
  assign n14938 = ~n14825 & n14937;
  assign n14939 = n14938 ^ n14833;
  assign n15043 = n15042 ^ n14939;
  assign n15052 = n15051 ^ n15043;
  assign n14934 = n14843 ^ n14724;
  assign n14935 = ~n14835 & n14934;
  assign n14936 = n14935 ^ n14843;
  assign n15053 = n15052 ^ n14936;
  assign n15062 = n15061 ^ n15053;
  assign n14931 = n14853 ^ n14844;
  assign n14932 = ~n14845 & n14931;
  assign n14933 = n14932 ^ n14853;
  assign n15063 = n15062 ^ n14933;
  assign n15072 = n15071 ^ n15063;
  assign n14928 = n14863 ^ n14854;
  assign n14929 = ~n14855 & n14928;
  assign n14930 = n14929 ^ n14863;
  assign n15073 = n15072 ^ n14930;
  assign n14925 = n14873 ^ n14864;
  assign n14926 = ~n14865 & n14925;
  assign n14927 = n14926 ^ n14873;
  assign n15074 = n15073 ^ n14927;
  assign n14917 = n2371 & n8715;
  assign n14918 = x120 & n2377;
  assign n14919 = x119 & n2528;
  assign n14920 = ~n14918 & ~n14919;
  assign n14921 = x121 & n2531;
  assign n14922 = n14920 & ~n14921;
  assign n14923 = ~n14917 & n14922;
  assign n14924 = n14923 ^ x29;
  assign n15075 = n15074 ^ n14924;
  assign n15084 = n15083 ^ n15075;
  assign n14914 = n14883 ^ n14712;
  assign n14915 = ~n14875 & n14914;
  assign n14916 = n14915 ^ n14883;
  assign n15085 = n15084 ^ n14916;
  assign n15094 = n15093 ^ n15085;
  assign n14911 = n14893 ^ n14884;
  assign n14912 = ~n14885 & n14911;
  assign n14913 = n14912 ^ n14893;
  assign n15095 = n15094 ^ n14913;
  assign n15114 = n15113 ^ n15095;
  assign n15306 = n15095 & ~n15102;
  assign n15307 = ~n15097 & ~n15306;
  assign n15308 = n15095 & ~n15096;
  assign n15309 = ~n15104 & ~n15308;
  assign n15310 = ~n15307 & ~n15309;
  assign n15311 = ~n14909 & ~n15310;
  assign n15312 = ~n15095 & n15100;
  assign n15313 = n15096 & n15307;
  assign n15314 = ~n15312 & ~n15313;
  assign n15315 = ~n15311 & n15314;
  assign n15294 = n1969 & n9912;
  assign n15295 = x123 & n1978;
  assign n15296 = x125 & n2108;
  assign n15297 = ~n15295 & ~n15296;
  assign n15298 = x124 & n1973;
  assign n15299 = n15297 & ~n15298;
  assign n15300 = ~n15294 & n15299;
  assign n15301 = n15300 ^ x26;
  assign n15284 = n2371 & n9001;
  assign n15285 = x120 & n2528;
  assign n15286 = x121 & n2377;
  assign n15287 = ~n15285 & ~n15286;
  assign n15288 = x122 & n2531;
  assign n15289 = n15287 & ~n15288;
  assign n15290 = ~n15284 & n15289;
  assign n15291 = n15290 ^ x29;
  assign n15272 = n3330 & n7393;
  assign n15273 = x114 & n3500;
  assign n15274 = x116 & n3502;
  assign n15275 = ~n15273 & ~n15274;
  assign n15276 = x115 & n3334;
  assign n15277 = n15275 & ~n15276;
  assign n15278 = ~n15272 & n15277;
  assign n15279 = n15278 ^ x35;
  assign n15262 = n3829 & n6656;
  assign n15263 = x111 & n4049;
  assign n15264 = x113 & n4052;
  assign n15265 = ~n15263 & ~n15264;
  assign n15266 = x112 & n3833;
  assign n15267 = n15265 & ~n15266;
  assign n15268 = ~n15262 & n15267;
  assign n15269 = n15268 ^ x38;
  assign n15251 = n4415 & n5955;
  assign n15252 = x108 & n4420;
  assign n15253 = x110 & n4614;
  assign n15254 = ~n15252 & ~n15253;
  assign n15255 = x109 & n4410;
  assign n15256 = n15254 & ~n15255;
  assign n15257 = ~n15251 & n15256;
  assign n15258 = n15257 ^ x41;
  assign n15242 = n5010 & n5297;
  assign n15243 = x105 & n5223;
  assign n15244 = x106 & n5014;
  assign n15245 = ~n15243 & ~n15244;
  assign n15246 = x107 & n5226;
  assign n15247 = n15245 & ~n15246;
  assign n15248 = ~n15242 & n15247;
  assign n15249 = n15248 ^ x44;
  assign n15231 = n4670 & n5656;
  assign n15232 = x102 & n5895;
  assign n15233 = x103 & n5662;
  assign n15234 = ~n15232 & ~n15233;
  assign n15235 = x104 & n6111;
  assign n15236 = n15234 & ~n15235;
  assign n15237 = ~n15231 & n15236;
  assign n15238 = n15237 ^ x47;
  assign n15228 = n15019 ^ n15008;
  assign n15229 = n15020 & n15228;
  assign n15230 = n15229 ^ n15011;
  assign n15239 = n15238 ^ n15230;
  assign n15218 = n4105 & n6326;
  assign n15219 = x99 & n6565;
  assign n15220 = x100 & n6331;
  assign n15221 = ~n15219 & ~n15220;
  assign n15222 = x101 & n6569;
  assign n15223 = n15221 & ~n15222;
  assign n15224 = ~n15218 & n15223;
  assign n15225 = n15224 ^ x50;
  assign n15208 = n3556 & n7076;
  assign n15209 = x96 & n7317;
  assign n15210 = x97 & n7080;
  assign n15211 = ~n15209 & ~n15210;
  assign n15212 = x98 & n7319;
  assign n15213 = n15211 & ~n15212;
  assign n15214 = ~n15208 & n15213;
  assign n15215 = n15214 ^ x53;
  assign n15198 = n3054 & n7830;
  assign n15199 = x93 & n7839;
  assign n15200 = x95 & n8374;
  assign n15201 = ~n15199 & ~n15200;
  assign n15202 = x94 & n7834;
  assign n15203 = n15201 & ~n15202;
  assign n15204 = ~n15198 & n15203;
  assign n15205 = n15204 ^ x56;
  assign n15188 = n2585 & n8622;
  assign n15189 = x90 & n8631;
  assign n15190 = x91 & n8626;
  assign n15191 = ~n15189 & ~n15190;
  assign n15192 = x92 & n9186;
  assign n15193 = n15191 & ~n15192;
  assign n15194 = ~n15188 & n15193;
  assign n15195 = n15194 ^ x59;
  assign n15178 = n2164 & n9499;
  assign n15179 = x87 & n9508;
  assign n15180 = x89 & n10106;
  assign n15181 = ~n15179 & ~n15180;
  assign n15182 = x88 & n9503;
  assign n15183 = n15181 & ~n15182;
  assign n15184 = ~n15178 & n15183;
  assign n15185 = n15184 ^ x62;
  assign n15171 = ~x20 & x84;
  assign n15172 = ~n14754 & ~n15171;
  assign n15173 = x85 & ~n10099;
  assign n15174 = n15172 & ~n15173;
  assign n15175 = x20 & ~x84;
  assign n15176 = ~n12465 & ~n15175;
  assign n15177 = ~n15174 & n15176;
  assign n15186 = n15185 ^ n15177;
  assign n15168 = x86 & n9798;
  assign n15169 = x85 & n10099;
  assign n15170 = ~n15168 & ~n15169;
  assign n15187 = n15186 ^ n15170;
  assign n15196 = n15195 ^ n15187;
  assign n15165 = n14973 ^ n14961;
  assign n15166 = n14974 & n15165;
  assign n15167 = n15166 ^ n14961;
  assign n15197 = n15196 ^ n15167;
  assign n15206 = n15205 ^ n15197;
  assign n15162 = n14986 ^ n14975;
  assign n15163 = n14987 & n15162;
  assign n15164 = n15163 ^ n14978;
  assign n15207 = n15206 ^ n15164;
  assign n15216 = n15215 ^ n15207;
  assign n15159 = n14996 ^ n14959;
  assign n15160 = n14997 & n15159;
  assign n15161 = n15160 ^ n14959;
  assign n15217 = n15216 ^ n15161;
  assign n15226 = n15225 ^ n15217;
  assign n15156 = n15006 ^ n14956;
  assign n15157 = n15007 & n15156;
  assign n15158 = n15157 ^ n14956;
  assign n15227 = n15226 ^ n15158;
  assign n15240 = n15239 ^ n15227;
  assign n15153 = n15021 ^ n14950;
  assign n15154 = ~n15022 & n15153;
  assign n15155 = n15154 ^ n14953;
  assign n15241 = n15240 ^ n15155;
  assign n15250 = n15249 ^ n15241;
  assign n15259 = n15258 ^ n15250;
  assign n15150 = n15031 ^ n14942;
  assign n15151 = n15032 & n15150;
  assign n15152 = n15151 ^ n14942;
  assign n15260 = n15259 ^ n15152;
  assign n15147 = n15033 ^ n14939;
  assign n15148 = ~n15042 & n15147;
  assign n15149 = n15148 ^ n15041;
  assign n15261 = n15260 ^ n15149;
  assign n15270 = n15269 ^ n15261;
  assign n15144 = n15043 ^ n14936;
  assign n15145 = ~n15052 & n15144;
  assign n15146 = n15145 ^ n15051;
  assign n15271 = n15270 ^ n15146;
  assign n15280 = n15279 ^ n15271;
  assign n15141 = n15061 ^ n14933;
  assign n15142 = n15062 & n15141;
  assign n15143 = n15142 ^ n14933;
  assign n15281 = n15280 ^ n15143;
  assign n15133 = n2836 & n8169;
  assign n15134 = x117 & n2996;
  assign n15135 = x118 & n2840;
  assign n15136 = ~n15134 & ~n15135;
  assign n15137 = x119 & n2998;
  assign n15138 = n15136 & ~n15137;
  assign n15139 = ~n15133 & n15138;
  assign n15140 = n15139 ^ x32;
  assign n15282 = n15281 ^ n15140;
  assign n15130 = n15071 ^ n14930;
  assign n15131 = n15072 & n15130;
  assign n15132 = n15131 ^ n14930;
  assign n15283 = n15282 ^ n15132;
  assign n15292 = n15291 ^ n15283;
  assign n15127 = n15073 ^ n14924;
  assign n15128 = ~n15074 & n15127;
  assign n15129 = n15128 ^ n14927;
  assign n15293 = n15292 ^ n15129;
  assign n15302 = n15301 ^ n15293;
  assign n15124 = n15083 ^ n14916;
  assign n15125 = n15084 & n15124;
  assign n15126 = n15125 ^ n14916;
  assign n15303 = n15302 ^ n15126;
  assign n15118 = n1624 & ~n9889;
  assign n15119 = x127 & n1628;
  assign n15120 = x126 & n1742;
  assign n15121 = ~n15119 & ~n15120;
  assign n15122 = ~n15118 & n15121;
  assign n15123 = n15122 ^ x23;
  assign n15304 = n15303 ^ n15123;
  assign n15115 = n15085 ^ n14913;
  assign n15116 = ~n15094 & n15115;
  assign n15117 = n15116 ^ n15093;
  assign n15305 = n15304 ^ n15117;
  assign n15316 = n15315 ^ n15305;
  assign n15495 = n1398 & n10430;
  assign n15496 = x127 & n1612;
  assign n15497 = x23 & ~n15496;
  assign n15498 = ~n15495 & n15497;
  assign n15499 = ~x22 & ~n15498;
  assign n15500 = x127 & n1615;
  assign n15501 = ~x23 & ~n15500;
  assign n15502 = ~n15495 & n15501;
  assign n15503 = ~n15499 & ~n15502;
  assign n15485 = n1969 & ~n10174;
  assign n15486 = x124 & n1978;
  assign n15487 = x125 & n1973;
  assign n15488 = ~n15486 & ~n15487;
  assign n15489 = x126 & n2108;
  assign n15490 = n15488 & ~n15489;
  assign n15491 = ~n15485 & n15490;
  assign n15492 = n15491 ^ x26;
  assign n15475 = n2371 & n9309;
  assign n15476 = x121 & n2528;
  assign n15477 = x123 & n2531;
  assign n15478 = ~n15476 & ~n15477;
  assign n15479 = x122 & n2377;
  assign n15480 = n15478 & ~n15479;
  assign n15481 = ~n15475 & n15480;
  assign n15482 = n15481 ^ x29;
  assign n15465 = n2836 & ~n8424;
  assign n15466 = x118 & n2996;
  assign n15467 = x119 & n2840;
  assign n15468 = ~n15466 & ~n15467;
  assign n15469 = x120 & n2998;
  assign n15470 = n15468 & ~n15469;
  assign n15471 = ~n15465 & n15470;
  assign n15472 = n15471 ^ x32;
  assign n15455 = n3330 & n7643;
  assign n15456 = x115 & n3500;
  assign n15457 = x116 & n3334;
  assign n15458 = ~n15456 & ~n15457;
  assign n15459 = x117 & n3502;
  assign n15460 = n15458 & ~n15459;
  assign n15461 = ~n15455 & n15460;
  assign n15462 = n15461 ^ x35;
  assign n15445 = n3829 & n6892;
  assign n15446 = x112 & n4049;
  assign n15447 = x113 & n3833;
  assign n15448 = ~n15446 & ~n15447;
  assign n15449 = x114 & n4052;
  assign n15450 = n15448 & ~n15449;
  assign n15451 = ~n15445 & n15450;
  assign n15452 = n15451 ^ x38;
  assign n15435 = n4415 & n6178;
  assign n15436 = x109 & n4420;
  assign n15437 = x111 & n4614;
  assign n15438 = ~n15436 & ~n15437;
  assign n15439 = x110 & n4410;
  assign n15440 = n15438 & ~n15439;
  assign n15441 = ~n15435 & n15440;
  assign n15442 = n15441 ^ x41;
  assign n15422 = n4867 & n5656;
  assign n15423 = x103 & n5895;
  assign n15424 = x105 & n6111;
  assign n15425 = ~n15423 & ~n15424;
  assign n15426 = x104 & n5662;
  assign n15427 = n15425 & ~n15426;
  assign n15428 = ~n15422 & n15427;
  assign n15429 = n15428 ^ x47;
  assign n15419 = n15217 ^ n15158;
  assign n15420 = n15226 & ~n15419;
  assign n15421 = n15420 ^ n15225;
  assign n15430 = n15429 ^ n15421;
  assign n15409 = n4286 & n6326;
  assign n15410 = x100 & n6565;
  assign n15411 = x102 & n6569;
  assign n15412 = ~n15410 & ~n15411;
  assign n15413 = x101 & n6331;
  assign n15414 = n15412 & ~n15413;
  assign n15415 = ~n15409 & n15414;
  assign n15416 = n15415 ^ x50;
  assign n15406 = n15207 ^ n15161;
  assign n15407 = n15216 & ~n15406;
  assign n15408 = n15407 ^ n15215;
  assign n15417 = n15416 ^ n15408;
  assign n15396 = n3730 & n7076;
  assign n15397 = x97 & n7317;
  assign n15398 = x98 & n7080;
  assign n15399 = ~n15397 & ~n15398;
  assign n15400 = x99 & n7319;
  assign n15401 = n15399 & ~n15400;
  assign n15402 = ~n15396 & n15401;
  assign n15403 = n15402 ^ x53;
  assign n15393 = n15197 ^ n15164;
  assign n15394 = n15206 & ~n15393;
  assign n15395 = n15394 ^ n15205;
  assign n15404 = n15403 ^ n15395;
  assign n15383 = n3209 & n7830;
  assign n15384 = x94 & n7839;
  assign n15385 = x96 & n8374;
  assign n15386 = ~n15384 & ~n15385;
  assign n15387 = x95 & n7834;
  assign n15388 = n15386 & ~n15387;
  assign n15389 = ~n15383 & n15388;
  assign n15390 = n15389 ^ x56;
  assign n15380 = n15187 ^ n15167;
  assign n15381 = n15196 & ~n15380;
  assign n15382 = n15381 ^ n15195;
  assign n15391 = n15390 ^ n15382;
  assign n15370 = n2726 & n8622;
  assign n15371 = x91 & n8631;
  assign n15372 = x92 & n8626;
  assign n15373 = ~n15371 & ~n15372;
  assign n15374 = x93 & n9186;
  assign n15375 = n15373 & ~n15374;
  assign n15376 = ~n15370 & n15375;
  assign n15377 = n15376 ^ x59;
  assign n15367 = n15177 ^ n15170;
  assign n15368 = ~n15186 & ~n15367;
  assign n15369 = n15368 ^ n15185;
  assign n15378 = n15377 ^ n15369;
  assign n15358 = n2292 & n9499;
  assign n15359 = x88 & n9508;
  assign n15360 = x89 & n9503;
  assign n15361 = ~n15359 & ~n15360;
  assign n15362 = x90 & n10106;
  assign n15363 = n15361 & ~n15362;
  assign n15364 = ~n15358 & n15363;
  assign n15365 = n15364 ^ x62;
  assign n15355 = n1663 & n9798;
  assign n15356 = n1536 & n10099;
  assign n15357 = ~n15355 & ~n15356;
  assign n15366 = n15365 ^ n15357;
  assign n15379 = n15378 ^ n15366;
  assign n15392 = n15391 ^ n15379;
  assign n15405 = n15404 ^ n15392;
  assign n15418 = n15417 ^ n15405;
  assign n15431 = n15430 ^ n15418;
  assign n15352 = n15230 ^ n15227;
  assign n15353 = n15239 & ~n15352;
  assign n15354 = n15353 ^ n15238;
  assign n15432 = n15431 ^ n15354;
  assign n15344 = n5010 & ~n5506;
  assign n15345 = x106 & n5223;
  assign n15346 = x107 & n5014;
  assign n15347 = ~n15345 & ~n15346;
  assign n15348 = x108 & n5226;
  assign n15349 = n15347 & ~n15348;
  assign n15350 = ~n15344 & n15349;
  assign n15351 = n15350 ^ x44;
  assign n15433 = n15432 ^ n15351;
  assign n15341 = n15249 ^ n15240;
  assign n15342 = ~n15241 & n15341;
  assign n15343 = n15342 ^ n15249;
  assign n15434 = n15433 ^ n15343;
  assign n15443 = n15442 ^ n15434;
  assign n15338 = n15258 ^ n15152;
  assign n15339 = ~n15259 & n15338;
  assign n15340 = n15339 ^ n15152;
  assign n15444 = n15443 ^ n15340;
  assign n15453 = n15452 ^ n15444;
  assign n15335 = n15269 ^ n15149;
  assign n15336 = ~n15261 & n15335;
  assign n15337 = n15336 ^ n15269;
  assign n15454 = n15453 ^ n15337;
  assign n15463 = n15462 ^ n15454;
  assign n15332 = n15279 ^ n15146;
  assign n15333 = ~n15271 & n15332;
  assign n15334 = n15333 ^ n15279;
  assign n15464 = n15463 ^ n15334;
  assign n15473 = n15472 ^ n15464;
  assign n15329 = n15280 ^ n15140;
  assign n15330 = n15281 & ~n15329;
  assign n15331 = n15330 ^ n15143;
  assign n15474 = n15473 ^ n15331;
  assign n15483 = n15482 ^ n15474;
  assign n15326 = n15291 ^ n15132;
  assign n15327 = ~n15283 & n15326;
  assign n15328 = n15327 ^ n15291;
  assign n15484 = n15483 ^ n15328;
  assign n15493 = n15492 ^ n15484;
  assign n15323 = n15301 ^ n15292;
  assign n15324 = ~n15293 & n15323;
  assign n15325 = n15324 ^ n15301;
  assign n15494 = n15493 ^ n15325;
  assign n15504 = n15503 ^ n15494;
  assign n15320 = n15302 ^ n15123;
  assign n15321 = n15303 & ~n15320;
  assign n15322 = n15321 ^ n15126;
  assign n15505 = n15504 ^ n15322;
  assign n15317 = n15315 ^ n15117;
  assign n15318 = ~n15305 & ~n15317;
  assign n15319 = n15318 ^ n15315;
  assign n15506 = n15505 ^ n15319;
  assign n15686 = ~n15322 & n15504;
  assign n15687 = ~n15319 & ~n15686;
  assign n15688 = n15322 & ~n15504;
  assign n15689 = ~n15687 & ~n15688;
  assign n15675 = n1969 & ~n10447;
  assign n15676 = x125 & n1978;
  assign n15677 = x126 & n1973;
  assign n15678 = ~n15676 & ~n15677;
  assign n15679 = x127 & n2108;
  assign n15680 = n15678 & ~n15679;
  assign n15681 = ~n15675 & n15680;
  assign n15682 = n15681 ^ x26;
  assign n15665 = n2371 & n9614;
  assign n15666 = x122 & n2528;
  assign n15667 = x123 & n2377;
  assign n15668 = ~n15666 & ~n15667;
  assign n15669 = x124 & n2531;
  assign n15670 = n15668 & ~n15669;
  assign n15671 = ~n15665 & n15670;
  assign n15672 = n15671 ^ x29;
  assign n15653 = n3330 & n7919;
  assign n15654 = x116 & n3500;
  assign n15655 = x118 & n3502;
  assign n15656 = ~n15654 & ~n15655;
  assign n15657 = x117 & n3334;
  assign n15658 = n15656 & ~n15657;
  assign n15659 = ~n15653 & n15658;
  assign n15660 = n15659 ^ x35;
  assign n15643 = n3829 & n7150;
  assign n15644 = x113 & n4049;
  assign n15645 = x115 & n4052;
  assign n15646 = ~n15644 & ~n15645;
  assign n15647 = x114 & n3833;
  assign n15648 = n15646 & ~n15647;
  assign n15649 = ~n15643 & n15648;
  assign n15650 = n15649 ^ x38;
  assign n15633 = n4415 & n6420;
  assign n15634 = x110 & n4420;
  assign n15635 = x112 & n4614;
  assign n15636 = ~n15634 & ~n15635;
  assign n15637 = x111 & n4410;
  assign n15638 = n15636 & ~n15637;
  assign n15639 = ~n15633 & n15638;
  assign n15640 = n15639 ^ x41;
  assign n15619 = n4481 & n6326;
  assign n15620 = x101 & n6565;
  assign n15621 = x103 & n6569;
  assign n15622 = ~n15620 & ~n15621;
  assign n15623 = x102 & n6331;
  assign n15624 = n15622 & ~n15623;
  assign n15625 = ~n15619 & n15624;
  assign n15626 = n15625 ^ x50;
  assign n15616 = n15408 ^ n15405;
  assign n15617 = n15417 & ~n15616;
  assign n15618 = n15617 ^ n15416;
  assign n15627 = n15626 ^ n15618;
  assign n15606 = n3925 & n7076;
  assign n15607 = x98 & n7317;
  assign n15608 = x99 & n7080;
  assign n15609 = ~n15607 & ~n15608;
  assign n15610 = x100 & n7319;
  assign n15611 = n15609 & ~n15610;
  assign n15612 = ~n15606 & n15611;
  assign n15613 = n15612 ^ x53;
  assign n15603 = n15395 ^ n15392;
  assign n15604 = n15404 & ~n15603;
  assign n15605 = n15604 ^ n15403;
  assign n15614 = n15613 ^ n15605;
  assign n15591 = n2895 & n8622;
  assign n15592 = x92 & n8631;
  assign n15593 = x93 & n8626;
  assign n15594 = ~n15592 & ~n15593;
  assign n15595 = x94 & n9186;
  assign n15596 = n15594 & ~n15595;
  assign n15597 = ~n15591 & n15596;
  assign n15598 = n15597 ^ x59;
  assign n15588 = n15369 ^ n15366;
  assign n15589 = n15378 & ~n15588;
  assign n15590 = n15589 ^ n15377;
  assign n15599 = n15598 ^ n15590;
  assign n15582 = n15357 & ~n15365;
  assign n15583 = ~x86 & n15169;
  assign n15584 = ~x87 & n15168;
  assign n15585 = ~n15583 & ~n15584;
  assign n15586 = ~n15582 & n15585;
  assign n15573 = n2447 & n9499;
  assign n15574 = x89 & n9508;
  assign n15575 = x91 & n10106;
  assign n15576 = ~n15574 & ~n15575;
  assign n15577 = x90 & n9503;
  assign n15578 = n15576 & ~n15577;
  assign n15579 = ~n15573 & n15578;
  assign n15580 = n15579 ^ x62;
  assign n15569 = n1663 & n10099;
  assign n15570 = n1776 & n9798;
  assign n15571 = ~n15569 & ~n15570;
  assign n15572 = n15571 ^ x23;
  assign n15581 = n15580 ^ n15572;
  assign n15587 = n15586 ^ n15581;
  assign n15600 = n15599 ^ n15587;
  assign n15561 = n3388 & n7830;
  assign n15562 = x95 & n7839;
  assign n15563 = x96 & n7834;
  assign n15564 = ~n15562 & ~n15563;
  assign n15565 = x97 & n8374;
  assign n15566 = n15564 & ~n15565;
  assign n15567 = ~n15561 & n15566;
  assign n15568 = n15567 ^ x56;
  assign n15601 = n15600 ^ n15568;
  assign n15558 = n15382 ^ n15379;
  assign n15559 = n15391 & ~n15558;
  assign n15560 = n15559 ^ n15390;
  assign n15602 = n15601 ^ n15560;
  assign n15615 = n15614 ^ n15602;
  assign n15628 = n15627 ^ n15615;
  assign n15555 = n15421 ^ n15418;
  assign n15556 = n15430 & ~n15555;
  assign n15557 = n15556 ^ n15429;
  assign n15629 = n15628 ^ n15557;
  assign n15547 = n5088 & n5656;
  assign n15548 = x104 & n5895;
  assign n15549 = x106 & n6111;
  assign n15550 = ~n15548 & ~n15549;
  assign n15551 = x105 & n5662;
  assign n15552 = n15550 & ~n15551;
  assign n15553 = ~n15547 & n15552;
  assign n15554 = n15553 ^ x47;
  assign n15630 = n15629 ^ n15554;
  assign n15539 = n5010 & ~n5737;
  assign n15540 = x107 & n5223;
  assign n15541 = x109 & n5226;
  assign n15542 = ~n15540 & ~n15541;
  assign n15543 = x108 & n5014;
  assign n15544 = n15542 & ~n15543;
  assign n15545 = ~n15539 & n15544;
  assign n15546 = n15545 ^ x44;
  assign n15631 = n15630 ^ n15546;
  assign n15536 = n15431 ^ n15351;
  assign n15537 = n15432 & ~n15536;
  assign n15538 = n15537 ^ n15354;
  assign n15632 = n15631 ^ n15538;
  assign n15641 = n15640 ^ n15632;
  assign n15533 = n15442 ^ n15343;
  assign n15534 = ~n15434 & n15533;
  assign n15535 = n15534 ^ n15442;
  assign n15642 = n15641 ^ n15535;
  assign n15651 = n15650 ^ n15642;
  assign n15530 = n15452 ^ n15340;
  assign n15531 = ~n15444 & n15530;
  assign n15532 = n15531 ^ n15452;
  assign n15652 = n15651 ^ n15532;
  assign n15661 = n15660 ^ n15652;
  assign n15527 = n15462 ^ n15453;
  assign n15528 = ~n15454 & n15527;
  assign n15529 = n15528 ^ n15462;
  assign n15662 = n15661 ^ n15529;
  assign n15524 = n15472 ^ n15334;
  assign n15525 = ~n15464 & n15524;
  assign n15526 = n15525 ^ n15472;
  assign n15663 = n15662 ^ n15526;
  assign n15516 = n2836 & n8715;
  assign n15517 = x119 & n2996;
  assign n15518 = x120 & n2840;
  assign n15519 = ~n15517 & ~n15518;
  assign n15520 = x121 & n2998;
  assign n15521 = n15519 & ~n15520;
  assign n15522 = ~n15516 & n15521;
  assign n15523 = n15522 ^ x32;
  assign n15664 = n15663 ^ n15523;
  assign n15673 = n15672 ^ n15664;
  assign n15513 = n15482 ^ n15331;
  assign n15514 = ~n15474 & n15513;
  assign n15515 = n15514 ^ n15482;
  assign n15674 = n15673 ^ n15515;
  assign n15683 = n15682 ^ n15674;
  assign n15510 = n15492 ^ n15483;
  assign n15511 = ~n15484 & n15510;
  assign n15512 = n15511 ^ n15492;
  assign n15684 = n15683 ^ n15512;
  assign n15507 = n15503 ^ n15493;
  assign n15508 = ~n15494 & ~n15507;
  assign n15509 = n15508 ^ n15503;
  assign n15685 = n15684 ^ n15509;
  assign n15690 = n15689 ^ n15685;
  assign n15866 = ~n15509 & n15512;
  assign n15867 = ~n15674 & n15682;
  assign n15868 = ~n15866 & ~n15867;
  assign n15869 = n15868 ^ n15689;
  assign n15870 = n15512 ^ n15509;
  assign n15871 = n15674 ^ n15512;
  assign n15872 = n15683 & n15871;
  assign n15873 = n15870 & n15872;
  assign n15874 = n15873 ^ n15685;
  assign n15875 = ~n15869 & n15874;
  assign n15876 = n15682 ^ n15509;
  assign n15877 = n15872 & n15876;
  assign n15878 = ~n15875 & ~n15877;
  assign n15855 = n2371 & n9912;
  assign n15856 = x123 & n2528;
  assign n15857 = x124 & n2377;
  assign n15858 = ~n15856 & ~n15857;
  assign n15859 = x125 & n2531;
  assign n15860 = n15858 & ~n15859;
  assign n15861 = ~n15855 & n15860;
  assign n15862 = n15861 ^ x29;
  assign n15845 = n2836 & n9001;
  assign n15846 = x121 & n2840;
  assign n15847 = x120 & n2996;
  assign n15848 = ~n15846 & ~n15847;
  assign n15849 = x122 & n2998;
  assign n15850 = n15848 & ~n15849;
  assign n15851 = ~n15845 & n15850;
  assign n15852 = n15851 ^ x32;
  assign n15834 = n3330 & n8169;
  assign n15835 = x117 & n3500;
  assign n15836 = x118 & n3334;
  assign n15837 = ~n15835 & ~n15836;
  assign n15838 = x119 & n3502;
  assign n15839 = n15837 & ~n15838;
  assign n15840 = ~n15834 & n15839;
  assign n15841 = n15840 ^ x35;
  assign n15831 = n15650 ^ n15532;
  assign n15832 = n15651 & n15831;
  assign n15833 = n15832 ^ n15532;
  assign n15842 = n15841 ^ n15833;
  assign n15822 = n3829 & n7393;
  assign n15823 = x114 & n4049;
  assign n15824 = x116 & n4052;
  assign n15825 = ~n15823 & ~n15824;
  assign n15826 = x115 & n3833;
  assign n15827 = n15825 & ~n15826;
  assign n15828 = ~n15822 & n15827;
  assign n15829 = n15828 ^ x38;
  assign n15812 = n4415 & n6656;
  assign n15813 = x111 & n4420;
  assign n15814 = x113 & n4614;
  assign n15815 = ~n15813 & ~n15814;
  assign n15816 = x112 & n4410;
  assign n15817 = n15815 & ~n15816;
  assign n15818 = ~n15812 & n15817;
  assign n15819 = n15818 ^ x41;
  assign n15801 = n5010 & n5955;
  assign n15802 = x108 & n5223;
  assign n15803 = x110 & n5226;
  assign n15804 = ~n15802 & ~n15803;
  assign n15805 = x109 & n5014;
  assign n15806 = n15804 & ~n15805;
  assign n15807 = ~n15801 & n15806;
  assign n15808 = n15807 ^ x44;
  assign n15789 = n4670 & n6326;
  assign n15790 = x102 & n6565;
  assign n15791 = x103 & n6331;
  assign n15792 = ~n15790 & ~n15791;
  assign n15793 = x104 & n6569;
  assign n15794 = n15792 & ~n15793;
  assign n15795 = ~n15789 & n15794;
  assign n15796 = n15795 ^ x50;
  assign n15786 = n15613 ^ n15602;
  assign n15787 = n15614 & n15786;
  assign n15788 = n15787 ^ n15605;
  assign n15797 = n15796 ^ n15788;
  assign n15776 = n4105 & n7076;
  assign n15777 = x99 & n7317;
  assign n15778 = x100 & n7080;
  assign n15779 = ~n15777 & ~n15778;
  assign n15780 = x101 & n7319;
  assign n15781 = n15779 & ~n15780;
  assign n15782 = ~n15776 & n15781;
  assign n15783 = n15782 ^ x53;
  assign n15773 = n15600 ^ n15560;
  assign n15774 = n15601 & ~n15773;
  assign n15775 = n15774 ^ n15560;
  assign n15784 = n15783 ^ n15775;
  assign n15763 = n3556 & n7830;
  assign n15764 = x96 & n7839;
  assign n15765 = x98 & n8374;
  assign n15766 = ~n15764 & ~n15765;
  assign n15767 = x97 & n7834;
  assign n15768 = n15766 & ~n15767;
  assign n15769 = ~n15763 & n15768;
  assign n15770 = n15769 ^ x56;
  assign n15753 = n3054 & n8622;
  assign n15754 = x93 & n8631;
  assign n15755 = x95 & n9186;
  assign n15756 = ~n15754 & ~n15755;
  assign n15757 = x94 & n8626;
  assign n15758 = n15756 & ~n15757;
  assign n15759 = ~n15753 & n15758;
  assign n15760 = n15759 ^ x59;
  assign n15744 = n2585 & n9499;
  assign n15745 = x90 & n9508;
  assign n15746 = x91 & n9503;
  assign n15747 = ~n15745 & ~n15746;
  assign n15748 = x92 & n10106;
  assign n15749 = n15747 & ~n15748;
  assign n15750 = ~n15744 & n15749;
  assign n15751 = n15750 ^ x62;
  assign n15735 = x86 & n10099;
  assign n15736 = ~x23 & x87;
  assign n15737 = ~n15735 & ~n15736;
  assign n15738 = x88 & ~n10099;
  assign n15739 = n15737 & ~n15738;
  assign n15740 = x23 & ~x87;
  assign n15741 = ~n12465 & ~n15740;
  assign n15742 = ~n15739 & n15741;
  assign n15732 = x89 & n9798;
  assign n15733 = x88 & n10099;
  assign n15734 = ~n15732 & ~n15733;
  assign n15743 = n15742 ^ n15734;
  assign n15752 = n15751 ^ n15743;
  assign n15761 = n15760 ^ n15752;
  assign n15729 = n15586 ^ n15580;
  assign n15730 = n15581 & n15729;
  assign n15731 = n15730 ^ n15586;
  assign n15762 = n15761 ^ n15731;
  assign n15771 = n15770 ^ n15762;
  assign n15726 = n15598 ^ n15587;
  assign n15727 = n15599 & n15726;
  assign n15728 = n15727 ^ n15590;
  assign n15772 = n15771 ^ n15728;
  assign n15785 = n15784 ^ n15772;
  assign n15798 = n15797 ^ n15785;
  assign n15723 = n15626 ^ n15615;
  assign n15724 = n15627 & n15723;
  assign n15725 = n15724 ^ n15618;
  assign n15799 = n15798 ^ n15725;
  assign n15715 = n5297 & n5656;
  assign n15716 = x105 & n5895;
  assign n15717 = x107 & n6111;
  assign n15718 = ~n15716 & ~n15717;
  assign n15719 = x106 & n5662;
  assign n15720 = n15718 & ~n15719;
  assign n15721 = ~n15715 & n15720;
  assign n15722 = n15721 ^ x47;
  assign n15800 = n15799 ^ n15722;
  assign n15809 = n15808 ^ n15800;
  assign n15712 = n15628 ^ n15554;
  assign n15713 = ~n15629 & n15712;
  assign n15714 = n15713 ^ n15557;
  assign n15810 = n15809 ^ n15714;
  assign n15709 = n15546 ^ n15538;
  assign n15710 = ~n15631 & ~n15709;
  assign n15711 = n15710 ^ n15630;
  assign n15811 = n15810 ^ n15711;
  assign n15820 = n15819 ^ n15811;
  assign n15706 = n15632 ^ n15535;
  assign n15707 = ~n15641 & n15706;
  assign n15708 = n15707 ^ n15640;
  assign n15821 = n15820 ^ n15708;
  assign n15830 = n15829 ^ n15821;
  assign n15843 = n15842 ^ n15830;
  assign n15703 = n15660 ^ n15529;
  assign n15704 = n15661 & n15703;
  assign n15705 = n15704 ^ n15529;
  assign n15844 = n15843 ^ n15705;
  assign n15853 = n15852 ^ n15844;
  assign n15700 = n15662 ^ n15523;
  assign n15701 = ~n15663 & n15700;
  assign n15702 = n15701 ^ n15526;
  assign n15854 = n15853 ^ n15702;
  assign n15863 = n15862 ^ n15854;
  assign n15697 = n15672 ^ n15515;
  assign n15698 = n15673 & n15697;
  assign n15699 = n15698 ^ n15515;
  assign n15864 = n15863 ^ n15699;
  assign n15691 = n1969 & ~n9889;
  assign n15692 = x127 & n1973;
  assign n15693 = x126 & n1978;
  assign n15694 = ~n15692 & ~n15693;
  assign n15695 = ~n15691 & n15694;
  assign n15696 = n15695 ^ x26;
  assign n15865 = n15864 ^ n15696;
  assign n15879 = n15878 ^ n15865;
  assign n16055 = n15509 & n15674;
  assign n16056 = ~n15509 & ~n15674;
  assign n16057 = ~n15688 & ~n16056;
  assign n16058 = ~n15687 & n16057;
  assign n16059 = ~n16055 & ~n16058;
  assign n16060 = ~n15512 & ~n15682;
  assign n16061 = ~n15865 & ~n16060;
  assign n16062 = ~n16059 & ~n16061;
  assign n16063 = n15512 & n15682;
  assign n16064 = ~n15865 & ~n16055;
  assign n16065 = ~n16063 & ~n16064;
  assign n16066 = n15689 & n16065;
  assign n16067 = n16056 & ~n16060;
  assign n16068 = n15865 & ~n16063;
  assign n16069 = ~n16067 & n16068;
  assign n16070 = ~n16066 & ~n16069;
  assign n16071 = ~n16062 & n16070;
  assign n16043 = n2371 & ~n10174;
  assign n16044 = x124 & n2528;
  assign n16045 = x126 & n2531;
  assign n16046 = ~n16044 & ~n16045;
  assign n16047 = x125 & n2377;
  assign n16048 = n16046 & ~n16047;
  assign n16049 = ~n16043 & n16048;
  assign n16050 = n16049 ^ x29;
  assign n16033 = n2836 & n9309;
  assign n16034 = x121 & n2996;
  assign n16035 = x122 & n2840;
  assign n16036 = ~n16034 & ~n16035;
  assign n16037 = x123 & n2998;
  assign n16038 = n16036 & ~n16037;
  assign n16039 = ~n16033 & n16038;
  assign n16040 = n16039 ^ x32;
  assign n16021 = n3829 & n7643;
  assign n16022 = x115 & n4049;
  assign n16023 = x117 & n4052;
  assign n16024 = ~n16022 & ~n16023;
  assign n16025 = x116 & n3833;
  assign n16026 = n16024 & ~n16025;
  assign n16027 = ~n16021 & n16026;
  assign n16028 = n16027 ^ x38;
  assign n16011 = n4415 & n6892;
  assign n16012 = x112 & n4420;
  assign n16013 = x113 & n4410;
  assign n16014 = ~n16012 & ~n16013;
  assign n16015 = x114 & n4614;
  assign n16016 = n16014 & ~n16015;
  assign n16017 = ~n16011 & n16016;
  assign n16018 = n16017 ^ x41;
  assign n16001 = n5010 & n6178;
  assign n16002 = x109 & n5223;
  assign n16003 = x111 & n5226;
  assign n16004 = ~n16002 & ~n16003;
  assign n16005 = x110 & n5014;
  assign n16006 = n16004 & ~n16005;
  assign n16007 = ~n16001 & n16006;
  assign n16008 = n16007 ^ x44;
  assign n15990 = ~n5506 & n5656;
  assign n15991 = x106 & n5895;
  assign n15992 = x107 & n5662;
  assign n15993 = ~n15991 & ~n15992;
  assign n15994 = x108 & n6111;
  assign n15995 = n15993 & ~n15994;
  assign n15996 = ~n15990 & n15995;
  assign n15997 = n15996 ^ x47;
  assign n15981 = n4867 & n6326;
  assign n15982 = x103 & n6565;
  assign n15983 = x104 & n6331;
  assign n15984 = ~n15982 & ~n15983;
  assign n15985 = x105 & n6569;
  assign n15986 = n15984 & ~n15985;
  assign n15987 = ~n15981 & n15986;
  assign n15988 = n15987 ^ x50;
  assign n15970 = n4286 & n7076;
  assign n15971 = x101 & n7080;
  assign n15972 = x100 & n7317;
  assign n15973 = ~n15971 & ~n15972;
  assign n15974 = x102 & n7319;
  assign n15975 = n15973 & ~n15974;
  assign n15976 = ~n15970 & n15975;
  assign n15977 = n15976 ^ x53;
  assign n15960 = n3730 & n7830;
  assign n15961 = x97 & n7839;
  assign n15962 = x99 & n8374;
  assign n15963 = ~n15961 & ~n15962;
  assign n15964 = x98 & n7834;
  assign n15965 = n15963 & ~n15964;
  assign n15966 = ~n15960 & n15965;
  assign n15967 = n15966 ^ x56;
  assign n15951 = n3209 & n8622;
  assign n15952 = x94 & n8631;
  assign n15953 = x95 & n8626;
  assign n15954 = ~n15952 & ~n15953;
  assign n15955 = x96 & n9186;
  assign n15956 = n15954 & ~n15955;
  assign n15957 = ~n15951 & n15956;
  assign n15958 = n15957 ^ x59;
  assign n15941 = n2726 & n9499;
  assign n15942 = x91 & n9508;
  assign n15943 = x92 & n9503;
  assign n15944 = ~n15942 & ~n15943;
  assign n15945 = x93 & n10106;
  assign n15946 = n15944 & ~n15945;
  assign n15947 = ~n15941 & n15946;
  assign n15948 = n15947 ^ x62;
  assign n15931 = x89 & n10099;
  assign n15932 = ~x88 & n15931;
  assign n15933 = ~x89 & x90;
  assign n15934 = n9798 & n15933;
  assign n15935 = ~n15932 & ~n15934;
  assign n15936 = ~x89 & n15733;
  assign n15937 = x89 & ~x90;
  assign n15938 = n9798 & n15937;
  assign n15939 = ~n15936 & ~n15938;
  assign n15940 = n15935 & n15939;
  assign n15949 = n15948 ^ n15940;
  assign n15928 = n15751 ^ n15742;
  assign n15929 = ~n15743 & ~n15928;
  assign n15930 = n15929 ^ n15751;
  assign n15950 = n15949 ^ n15930;
  assign n15959 = n15958 ^ n15950;
  assign n15968 = n15967 ^ n15959;
  assign n15925 = n15752 ^ n15731;
  assign n15926 = n15761 & ~n15925;
  assign n15927 = n15926 ^ n15760;
  assign n15969 = n15968 ^ n15927;
  assign n15978 = n15977 ^ n15969;
  assign n15922 = n15762 ^ n15728;
  assign n15923 = n15771 & ~n15922;
  assign n15924 = n15923 ^ n15770;
  assign n15979 = n15978 ^ n15924;
  assign n15919 = n15775 ^ n15772;
  assign n15920 = n15784 & ~n15919;
  assign n15921 = n15920 ^ n15783;
  assign n15980 = n15979 ^ n15921;
  assign n15989 = n15988 ^ n15980;
  assign n15998 = n15997 ^ n15989;
  assign n15916 = n15788 ^ n15785;
  assign n15917 = n15797 & ~n15916;
  assign n15918 = n15917 ^ n15796;
  assign n15999 = n15998 ^ n15918;
  assign n15913 = n15798 ^ n15722;
  assign n15914 = n15799 & ~n15913;
  assign n15915 = n15914 ^ n15725;
  assign n16000 = n15999 ^ n15915;
  assign n16009 = n16008 ^ n16000;
  assign n15910 = n15808 ^ n15714;
  assign n15911 = ~n15809 & n15910;
  assign n15912 = n15911 ^ n15714;
  assign n16010 = n16009 ^ n15912;
  assign n16019 = n16018 ^ n16010;
  assign n15907 = n15819 ^ n15711;
  assign n15908 = n15811 & ~n15907;
  assign n15909 = n15908 ^ n15819;
  assign n16020 = n16019 ^ n15909;
  assign n16029 = n16028 ^ n16020;
  assign n15904 = n15829 ^ n15708;
  assign n15905 = n15821 & n15904;
  assign n15906 = n15905 ^ n15829;
  assign n16030 = n16029 ^ n15906;
  assign n15896 = n3330 & ~n8424;
  assign n15897 = x118 & n3500;
  assign n15898 = x119 & n3334;
  assign n15899 = ~n15897 & ~n15898;
  assign n15900 = x120 & n3502;
  assign n15901 = n15899 & ~n15900;
  assign n15902 = ~n15896 & n15901;
  assign n15903 = n15902 ^ x35;
  assign n16031 = n16030 ^ n15903;
  assign n15893 = n15841 ^ n15830;
  assign n15894 = n15842 & n15893;
  assign n15895 = n15894 ^ n15833;
  assign n16032 = n16031 ^ n15895;
  assign n16041 = n16040 ^ n16032;
  assign n15890 = n15852 ^ n15705;
  assign n15891 = n15844 & n15890;
  assign n15892 = n15891 ^ n15852;
  assign n16042 = n16041 ^ n15892;
  assign n16051 = n16050 ^ n16042;
  assign n15886 = n1969 & n10430;
  assign n15887 = x127 & n1978;
  assign n15888 = ~n15886 & ~n15887;
  assign n15889 = n15888 ^ x26;
  assign n16052 = n16051 ^ n15889;
  assign n15883 = n15862 ^ n15853;
  assign n15884 = n15854 & ~n15883;
  assign n15885 = n15884 ^ n15862;
  assign n16053 = n16052 ^ n15885;
  assign n15880 = n15863 ^ n15696;
  assign n15881 = ~n15864 & n15880;
  assign n15882 = n15881 ^ n15699;
  assign n16054 = n16053 ^ n15882;
  assign n16072 = n16071 ^ n16054;
  assign n16232 = ~n15882 & ~n15885;
  assign n16233 = n16071 & ~n16232;
  assign n16234 = n15882 & n15885;
  assign n16235 = n16234 ^ n15889;
  assign n16236 = n16052 & ~n16235;
  assign n16237 = n16236 ^ n16051;
  assign n16238 = n16233 & n16237;
  assign n16239 = n15889 & n16051;
  assign n16240 = n16232 & ~n16239;
  assign n16241 = ~n15889 & ~n16051;
  assign n16242 = ~n16234 & n16241;
  assign n16243 = ~n16240 & ~n16242;
  assign n16244 = ~n16071 & ~n16243;
  assign n16245 = n16051 ^ n15882;
  assign n16246 = n15889 ^ n15885;
  assign n16247 = ~n16052 & ~n16246;
  assign n16248 = ~n16245 & n16247;
  assign n16249 = ~n16244 & ~n16248;
  assign n16250 = ~n16238 & n16249;
  assign n16222 = n2371 & ~n10447;
  assign n16223 = x125 & n2528;
  assign n16224 = x126 & n2377;
  assign n16225 = ~n16223 & ~n16224;
  assign n16226 = x127 & n2531;
  assign n16227 = n16225 & ~n16226;
  assign n16228 = ~n16222 & n16227;
  assign n16229 = n16228 ^ x29;
  assign n16212 = n2836 & n9614;
  assign n16213 = x122 & n2996;
  assign n16214 = x123 & n2840;
  assign n16215 = ~n16213 & ~n16214;
  assign n16216 = x124 & n2998;
  assign n16217 = n16215 & ~n16216;
  assign n16218 = ~n16212 & n16217;
  assign n16219 = n16218 ^ x32;
  assign n16200 = n3829 & n7919;
  assign n16201 = x116 & n4049;
  assign n16202 = x118 & n4052;
  assign n16203 = ~n16201 & ~n16202;
  assign n16204 = x117 & n3833;
  assign n16205 = n16203 & ~n16204;
  assign n16206 = ~n16200 & n16205;
  assign n16207 = n16206 ^ x38;
  assign n16190 = n4415 & n7150;
  assign n16191 = x113 & n4420;
  assign n16192 = x115 & n4614;
  assign n16193 = ~n16191 & ~n16192;
  assign n16194 = x114 & n4410;
  assign n16195 = n16193 & ~n16194;
  assign n16196 = ~n16190 & n16195;
  assign n16197 = n16196 ^ x41;
  assign n16180 = n5010 & n6420;
  assign n16181 = x110 & n5223;
  assign n16182 = x112 & n5226;
  assign n16183 = ~n16181 & ~n16182;
  assign n16184 = x111 & n5014;
  assign n16185 = n16183 & ~n16184;
  assign n16186 = ~n16180 & n16185;
  assign n16187 = n16186 ^ x44;
  assign n16168 = n5088 & n6326;
  assign n16169 = x104 & n6565;
  assign n16170 = x106 & n6569;
  assign n16171 = ~n16169 & ~n16170;
  assign n16172 = x105 & n6331;
  assign n16173 = n16171 & ~n16172;
  assign n16174 = ~n16168 & n16173;
  assign n16175 = n16174 ^ x50;
  assign n16165 = n15988 ^ n15979;
  assign n16166 = ~n15980 & n16165;
  assign n16167 = n16166 ^ n15988;
  assign n16176 = n16175 ^ n16167;
  assign n16155 = n4481 & n7076;
  assign n16156 = x101 & n7317;
  assign n16157 = x103 & n7319;
  assign n16158 = ~n16156 & ~n16157;
  assign n16159 = x102 & n7080;
  assign n16160 = n16158 & ~n16159;
  assign n16161 = ~n16155 & n16160;
  assign n16162 = n16161 ^ x53;
  assign n16152 = n15969 ^ n15924;
  assign n16153 = n15978 & ~n16152;
  assign n16154 = n16153 ^ n15977;
  assign n16163 = n16162 ^ n16154;
  assign n16142 = n3925 & n7830;
  assign n16143 = x98 & n7839;
  assign n16144 = x100 & n8374;
  assign n16145 = ~n16143 & ~n16144;
  assign n16146 = x99 & n7834;
  assign n16147 = n16145 & ~n16146;
  assign n16148 = ~n16142 & n16147;
  assign n16149 = n16148 ^ x56;
  assign n16132 = n3388 & n8622;
  assign n16133 = x95 & n8631;
  assign n16134 = x96 & n8626;
  assign n16135 = ~n16133 & ~n16134;
  assign n16136 = x97 & n9186;
  assign n16137 = n16135 & ~n16136;
  assign n16138 = ~n16132 & n16137;
  assign n16139 = n16138 ^ x59;
  assign n16126 = n2024 & n10099;
  assign n16127 = n2149 & n9798;
  assign n16128 = ~n16126 & ~n16127;
  assign n16129 = n16128 ^ x26;
  assign n16124 = n15940 & ~n15948;
  assign n16125 = n16124 ^ n15939;
  assign n16130 = n16129 ^ n16125;
  assign n16116 = n2895 & n9499;
  assign n16117 = x92 & n9508;
  assign n16118 = x93 & n9503;
  assign n16119 = ~n16117 & ~n16118;
  assign n16120 = x94 & n10106;
  assign n16121 = n16119 & ~n16120;
  assign n16122 = ~n16116 & n16121;
  assign n16123 = n16122 ^ x62;
  assign n16131 = n16130 ^ n16123;
  assign n16140 = n16139 ^ n16131;
  assign n16113 = n15958 ^ n15930;
  assign n16114 = ~n15950 & n16113;
  assign n16115 = n16114 ^ n15958;
  assign n16141 = n16140 ^ n16115;
  assign n16150 = n16149 ^ n16141;
  assign n16110 = n15959 ^ n15927;
  assign n16111 = n15968 & ~n16110;
  assign n16112 = n16111 ^ n15967;
  assign n16151 = n16150 ^ n16112;
  assign n16164 = n16163 ^ n16151;
  assign n16177 = n16176 ^ n16164;
  assign n16102 = n5656 & ~n5737;
  assign n16103 = x107 & n5895;
  assign n16104 = x108 & n5662;
  assign n16105 = ~n16103 & ~n16104;
  assign n16106 = x109 & n6111;
  assign n16107 = n16105 & ~n16106;
  assign n16108 = ~n16102 & n16107;
  assign n16109 = n16108 ^ x47;
  assign n16178 = n16177 ^ n16109;
  assign n16099 = n15989 ^ n15918;
  assign n16100 = n15998 & ~n16099;
  assign n16101 = n16100 ^ n15997;
  assign n16179 = n16178 ^ n16101;
  assign n16188 = n16187 ^ n16179;
  assign n16096 = n16008 ^ n15915;
  assign n16097 = ~n16000 & n16096;
  assign n16098 = n16097 ^ n16008;
  assign n16189 = n16188 ^ n16098;
  assign n16198 = n16197 ^ n16189;
  assign n16093 = n16018 ^ n16009;
  assign n16094 = ~n16010 & n16093;
  assign n16095 = n16094 ^ n16018;
  assign n16199 = n16198 ^ n16095;
  assign n16208 = n16207 ^ n16199;
  assign n16090 = n16028 ^ n16019;
  assign n16091 = ~n16020 & n16090;
  assign n16092 = n16091 ^ n16028;
  assign n16209 = n16208 ^ n16092;
  assign n16087 = n15906 ^ n15903;
  assign n16088 = n16030 & ~n16087;
  assign n16089 = n16088 ^ n16029;
  assign n16210 = n16209 ^ n16089;
  assign n16079 = n3330 & n8715;
  assign n16080 = x119 & n3500;
  assign n16081 = x120 & n3334;
  assign n16082 = ~n16080 & ~n16081;
  assign n16083 = x121 & n3502;
  assign n16084 = n16082 & ~n16083;
  assign n16085 = ~n16079 & n16084;
  assign n16086 = n16085 ^ x35;
  assign n16211 = n16210 ^ n16086;
  assign n16220 = n16219 ^ n16211;
  assign n16076 = n16040 ^ n15895;
  assign n16077 = ~n16032 & n16076;
  assign n16078 = n16077 ^ n16040;
  assign n16221 = n16220 ^ n16078;
  assign n16230 = n16229 ^ n16221;
  assign n16073 = n16050 ^ n15892;
  assign n16074 = ~n16042 & n16073;
  assign n16075 = n16074 ^ n16050;
  assign n16231 = n16230 ^ n16075;
  assign n16251 = n16250 ^ n16231;
  assign n16418 = ~n16231 & ~n16241;
  assign n16419 = ~n16234 & ~n16418;
  assign n16420 = ~n16233 & n16419;
  assign n16421 = ~n16231 & ~n16232;
  assign n16422 = ~n16239 & ~n16421;
  assign n16423 = ~n16071 & n16422;
  assign n16424 = n16231 & ~n16237;
  assign n16425 = ~n16423 & ~n16424;
  assign n16426 = ~n16420 & n16425;
  assign n16406 = n2836 & n9912;
  assign n16407 = x123 & n2996;
  assign n16408 = x124 & n2840;
  assign n16409 = ~n16407 & ~n16408;
  assign n16410 = x125 & n2998;
  assign n16411 = n16409 & ~n16410;
  assign n16412 = ~n16406 & n16411;
  assign n16413 = n16412 ^ x32;
  assign n16396 = n3330 & n9001;
  assign n16397 = x120 & n3500;
  assign n16398 = x121 & n3334;
  assign n16399 = ~n16397 & ~n16398;
  assign n16400 = x122 & n3502;
  assign n16401 = n16399 & ~n16400;
  assign n16402 = ~n16396 & n16401;
  assign n16403 = n16402 ^ x35;
  assign n16386 = n3829 & n8169;
  assign n16387 = x117 & n4049;
  assign n16388 = x119 & n4052;
  assign n16389 = ~n16387 & ~n16388;
  assign n16390 = x118 & n3833;
  assign n16391 = n16389 & ~n16390;
  assign n16392 = ~n16386 & n16391;
  assign n16393 = n16392 ^ x38;
  assign n16376 = n4415 & n7393;
  assign n16377 = x114 & n4420;
  assign n16378 = x115 & n4410;
  assign n16379 = ~n16377 & ~n16378;
  assign n16380 = x116 & n4614;
  assign n16381 = n16379 & ~n16380;
  assign n16382 = ~n16376 & n16381;
  assign n16383 = n16382 ^ x41;
  assign n16359 = n4670 & n7076;
  assign n16360 = x102 & n7317;
  assign n16361 = x103 & n7080;
  assign n16362 = ~n16360 & ~n16361;
  assign n16363 = x104 & n7319;
  assign n16364 = n16362 & ~n16363;
  assign n16365 = ~n16359 & n16364;
  assign n16366 = n16365 ^ x53;
  assign n16349 = n4105 & n7830;
  assign n16350 = x99 & n7839;
  assign n16351 = x101 & n8374;
  assign n16352 = ~n16350 & ~n16351;
  assign n16353 = x100 & n7834;
  assign n16354 = n16352 & ~n16353;
  assign n16355 = ~n16349 & n16354;
  assign n16356 = n16355 ^ x56;
  assign n16346 = n16131 ^ n16115;
  assign n16347 = ~n16140 & n16346;
  assign n16348 = n16347 ^ n16139;
  assign n16357 = n16356 ^ n16348;
  assign n16336 = n3556 & n8622;
  assign n16337 = x96 & n8631;
  assign n16338 = x98 & n9186;
  assign n16339 = ~n16337 & ~n16338;
  assign n16340 = x97 & n8626;
  assign n16341 = n16339 & ~n16340;
  assign n16342 = ~n16336 & n16341;
  assign n16343 = n16342 ^ x59;
  assign n16327 = n3054 & n9499;
  assign n16328 = x93 & n9508;
  assign n16329 = x94 & n9503;
  assign n16330 = ~n16328 & ~n16329;
  assign n16331 = x95 & n10106;
  assign n16332 = n16330 & ~n16331;
  assign n16333 = ~n16327 & n16332;
  assign n16334 = n16333 ^ x62;
  assign n16318 = ~x26 & x90;
  assign n16319 = x91 ^ x89;
  assign n16320 = ~n10099 & n16319;
  assign n16321 = n16320 ^ x89;
  assign n16322 = ~n16318 & ~n16321;
  assign n16323 = x26 & ~x90;
  assign n16324 = ~n12465 & ~n16323;
  assign n16325 = ~n16322 & n16324;
  assign n16315 = x92 & n9798;
  assign n16316 = x91 & n10099;
  assign n16317 = ~n16315 & ~n16316;
  assign n16326 = n16325 ^ n16317;
  assign n16335 = n16334 ^ n16326;
  assign n16344 = n16343 ^ n16335;
  assign n16312 = n16129 ^ n16123;
  assign n16313 = ~n16130 & n16312;
  assign n16314 = n16313 ^ n16125;
  assign n16345 = n16344 ^ n16314;
  assign n16358 = n16357 ^ n16345;
  assign n16367 = n16366 ^ n16358;
  assign n16309 = n16149 ^ n16112;
  assign n16310 = n16150 & n16309;
  assign n16311 = n16310 ^ n16112;
  assign n16368 = n16367 ^ n16311;
  assign n16306 = n16162 ^ n16151;
  assign n16307 = n16163 & n16306;
  assign n16308 = n16307 ^ n16154;
  assign n16369 = n16368 ^ n16308;
  assign n16298 = n5297 & n6326;
  assign n16299 = x105 & n6565;
  assign n16300 = x106 & n6331;
  assign n16301 = ~n16299 & ~n16300;
  assign n16302 = x107 & n6569;
  assign n16303 = n16301 & ~n16302;
  assign n16304 = ~n16298 & n16303;
  assign n16305 = n16304 ^ x50;
  assign n16370 = n16369 ^ n16305;
  assign n16295 = n16175 ^ n16164;
  assign n16296 = n16176 & n16295;
  assign n16297 = n16296 ^ n16167;
  assign n16371 = n16370 ^ n16297;
  assign n16287 = n5656 & n5955;
  assign n16288 = x108 & n5895;
  assign n16289 = x109 & n5662;
  assign n16290 = ~n16288 & ~n16289;
  assign n16291 = x110 & n6111;
  assign n16292 = n16290 & ~n16291;
  assign n16293 = ~n16287 & n16292;
  assign n16294 = n16293 ^ x47;
  assign n16372 = n16371 ^ n16294;
  assign n16284 = n16109 ^ n16101;
  assign n16285 = ~n16178 & ~n16284;
  assign n16286 = n16285 ^ n16177;
  assign n16373 = n16372 ^ n16286;
  assign n16276 = n5010 & n6656;
  assign n16277 = x111 & n5223;
  assign n16278 = x113 & n5226;
  assign n16279 = ~n16277 & ~n16278;
  assign n16280 = x112 & n5014;
  assign n16281 = n16279 & ~n16280;
  assign n16282 = ~n16276 & n16281;
  assign n16283 = n16282 ^ x44;
  assign n16374 = n16373 ^ n16283;
  assign n16273 = n16179 ^ n16098;
  assign n16274 = ~n16188 & n16273;
  assign n16275 = n16274 ^ n16187;
  assign n16375 = n16374 ^ n16275;
  assign n16384 = n16383 ^ n16375;
  assign n16270 = n16189 ^ n16095;
  assign n16271 = ~n16198 & n16270;
  assign n16272 = n16271 ^ n16197;
  assign n16385 = n16384 ^ n16272;
  assign n16394 = n16393 ^ n16385;
  assign n16267 = n16199 ^ n16092;
  assign n16268 = ~n16208 & n16267;
  assign n16269 = n16268 ^ n16207;
  assign n16395 = n16394 ^ n16269;
  assign n16404 = n16403 ^ n16395;
  assign n16264 = n16209 ^ n16086;
  assign n16265 = ~n16210 & n16264;
  assign n16266 = n16265 ^ n16089;
  assign n16405 = n16404 ^ n16266;
  assign n16414 = n16413 ^ n16405;
  assign n16261 = n16219 ^ n16078;
  assign n16262 = n16220 & n16261;
  assign n16263 = n16262 ^ n16078;
  assign n16415 = n16414 ^ n16263;
  assign n16255 = n2371 & ~n9889;
  assign n16256 = x127 & n2377;
  assign n16257 = x126 & n2528;
  assign n16258 = ~n16256 & ~n16257;
  assign n16259 = ~n16255 & n16258;
  assign n16260 = n16259 ^ x29;
  assign n16416 = n16415 ^ n16260;
  assign n16252 = n16229 ^ n16075;
  assign n16253 = n16230 & n16252;
  assign n16254 = n16253 ^ n16075;
  assign n16417 = n16416 ^ n16254;
  assign n16427 = n16426 ^ n16417;
  assign n16588 = n2116 & n10430;
  assign n16589 = x127 & n2373;
  assign n16590 = x29 & ~n16589;
  assign n16591 = ~n16588 & n16590;
  assign n16592 = ~x28 & ~n16591;
  assign n16593 = x127 & n2374;
  assign n16594 = ~x29 & ~n16593;
  assign n16595 = ~n16588 & n16594;
  assign n16596 = ~n16592 & ~n16595;
  assign n16578 = n2836 & ~n10174;
  assign n16579 = x124 & n2996;
  assign n16580 = x125 & n2840;
  assign n16581 = ~n16579 & ~n16580;
  assign n16582 = x126 & n2998;
  assign n16583 = n16581 & ~n16582;
  assign n16584 = ~n16578 & n16583;
  assign n16585 = n16584 ^ x32;
  assign n16568 = n3330 & n9309;
  assign n16569 = x121 & n3500;
  assign n16570 = x123 & n3502;
  assign n16571 = ~n16569 & ~n16570;
  assign n16572 = x122 & n3334;
  assign n16573 = n16571 & ~n16572;
  assign n16574 = ~n16568 & n16573;
  assign n16575 = n16574 ^ x35;
  assign n16558 = n3829 & ~n8424;
  assign n16559 = x118 & n4049;
  assign n16560 = x120 & n4052;
  assign n16561 = ~n16559 & ~n16560;
  assign n16562 = x119 & n3833;
  assign n16563 = n16561 & ~n16562;
  assign n16564 = ~n16558 & n16563;
  assign n16565 = n16564 ^ x38;
  assign n16548 = n4415 & n7643;
  assign n16549 = x115 & n4420;
  assign n16550 = x117 & n4614;
  assign n16551 = ~n16549 & ~n16550;
  assign n16552 = x116 & n4410;
  assign n16553 = n16551 & ~n16552;
  assign n16554 = ~n16548 & n16553;
  assign n16555 = n16554 ^ x41;
  assign n16536 = n5656 & n6178;
  assign n16537 = x109 & n5895;
  assign n16538 = x110 & n5662;
  assign n16539 = ~n16537 & ~n16538;
  assign n16540 = x111 & n6111;
  assign n16541 = n16539 & ~n16540;
  assign n16542 = ~n16536 & n16541;
  assign n16543 = n16542 ^ x47;
  assign n16525 = ~n5506 & n6326;
  assign n16526 = x106 & n6565;
  assign n16527 = x107 & n6331;
  assign n16528 = ~n16526 & ~n16527;
  assign n16529 = x108 & n6569;
  assign n16530 = n16528 & ~n16529;
  assign n16531 = ~n16525 & n16530;
  assign n16532 = n16531 ^ x50;
  assign n16522 = n16358 ^ n16311;
  assign n16523 = n16367 & ~n16522;
  assign n16524 = n16523 ^ n16366;
  assign n16533 = n16532 ^ n16524;
  assign n16512 = n4867 & n7076;
  assign n16513 = x103 & n7317;
  assign n16514 = x105 & n7319;
  assign n16515 = ~n16513 & ~n16514;
  assign n16516 = x104 & n7080;
  assign n16517 = n16515 & ~n16516;
  assign n16518 = ~n16512 & n16517;
  assign n16519 = n16518 ^ x53;
  assign n16509 = n16348 ^ n16345;
  assign n16510 = n16357 & ~n16509;
  assign n16511 = n16510 ^ n16356;
  assign n16520 = n16519 ^ n16511;
  assign n16499 = n4286 & n7830;
  assign n16500 = x100 & n7839;
  assign n16501 = x101 & n7834;
  assign n16502 = ~n16500 & ~n16501;
  assign n16503 = x102 & n8374;
  assign n16504 = n16502 & ~n16503;
  assign n16505 = ~n16499 & n16504;
  assign n16506 = n16505 ^ x56;
  assign n16496 = n16335 ^ n16314;
  assign n16497 = n16344 & ~n16496;
  assign n16498 = n16497 ^ n16343;
  assign n16507 = n16506 ^ n16498;
  assign n16487 = n3730 & n8622;
  assign n16488 = x97 & n8631;
  assign n16489 = x99 & n9186;
  assign n16490 = ~n16488 & ~n16489;
  assign n16491 = x98 & n8626;
  assign n16492 = n16490 & ~n16491;
  assign n16493 = ~n16487 & n16492;
  assign n16494 = n16493 ^ x59;
  assign n16474 = x91 & ~x92;
  assign n16475 = n10099 & n16474;
  assign n16476 = x92 & ~x93;
  assign n16477 = n9798 & n16476;
  assign n16478 = ~n16475 & ~n16477;
  assign n16479 = ~x92 & x93;
  assign n16480 = n9798 & n16479;
  assign n16481 = x92 & n10099;
  assign n16482 = ~x91 & n16481;
  assign n16483 = ~n16480 & ~n16482;
  assign n16484 = n16478 & n16483;
  assign n16471 = n16334 ^ n16325;
  assign n16472 = ~n16326 & ~n16471;
  assign n16473 = n16472 ^ n16334;
  assign n16485 = n16484 ^ n16473;
  assign n16463 = n3209 & n9499;
  assign n16464 = x94 & n9508;
  assign n16465 = x96 & n10106;
  assign n16466 = ~n16464 & ~n16465;
  assign n16467 = x95 & n9503;
  assign n16468 = n16466 & ~n16467;
  assign n16469 = ~n16463 & n16468;
  assign n16470 = n16469 ^ x62;
  assign n16486 = n16485 ^ n16470;
  assign n16495 = n16494 ^ n16486;
  assign n16508 = n16507 ^ n16495;
  assign n16521 = n16520 ^ n16508;
  assign n16534 = n16533 ^ n16521;
  assign n16460 = n16368 ^ n16305;
  assign n16461 = n16369 & ~n16460;
  assign n16462 = n16461 ^ n16308;
  assign n16535 = n16534 ^ n16462;
  assign n16544 = n16543 ^ n16535;
  assign n16457 = n16370 ^ n16294;
  assign n16458 = n16371 & ~n16457;
  assign n16459 = n16458 ^ n16297;
  assign n16545 = n16544 ^ n16459;
  assign n16449 = n5010 & n6892;
  assign n16450 = x112 & n5223;
  assign n16451 = x114 & n5226;
  assign n16452 = ~n16450 & ~n16451;
  assign n16453 = x113 & n5014;
  assign n16454 = n16452 & ~n16453;
  assign n16455 = ~n16449 & n16454;
  assign n16456 = n16455 ^ x44;
  assign n16546 = n16545 ^ n16456;
  assign n16446 = n16372 ^ n16283;
  assign n16447 = ~n16373 & ~n16446;
  assign n16448 = n16447 ^ n16286;
  assign n16547 = n16546 ^ n16448;
  assign n16556 = n16555 ^ n16547;
  assign n16443 = n16383 ^ n16275;
  assign n16444 = n16375 & n16443;
  assign n16445 = n16444 ^ n16383;
  assign n16557 = n16556 ^ n16445;
  assign n16566 = n16565 ^ n16557;
  assign n16440 = n16393 ^ n16272;
  assign n16441 = n16385 & n16440;
  assign n16442 = n16441 ^ n16393;
  assign n16567 = n16566 ^ n16442;
  assign n16576 = n16575 ^ n16567;
  assign n16437 = n16403 ^ n16269;
  assign n16438 = n16395 & n16437;
  assign n16439 = n16438 ^ n16403;
  assign n16577 = n16576 ^ n16439;
  assign n16586 = n16585 ^ n16577;
  assign n16434 = n16413 ^ n16404;
  assign n16435 = n16405 & ~n16434;
  assign n16436 = n16435 ^ n16413;
  assign n16587 = n16586 ^ n16436;
  assign n16597 = n16596 ^ n16587;
  assign n16431 = n16414 ^ n16260;
  assign n16432 = ~n16415 & n16431;
  assign n16433 = n16432 ^ n16263;
  assign n16598 = n16597 ^ n16433;
  assign n16428 = n16426 ^ n16254;
  assign n16429 = n16417 & n16428;
  assign n16430 = n16429 ^ n16426;
  assign n16599 = n16598 ^ n16430;
  assign n16748 = n16596 ^ n16586;
  assign n16749 = n16587 & n16748;
  assign n16750 = n16749 ^ n16596;
  assign n16745 = n16585 ^ n16576;
  assign n16746 = n16577 & ~n16745;
  assign n16747 = n16746 ^ n16585;
  assign n16751 = n16750 ^ n16747;
  assign n16736 = n2836 & ~n10447;
  assign n16737 = x125 & n2996;
  assign n16738 = x126 & n2840;
  assign n16739 = ~n16737 & ~n16738;
  assign n16740 = x127 & n2998;
  assign n16741 = n16739 & ~n16740;
  assign n16742 = ~n16736 & n16741;
  assign n16743 = n16742 ^ x32;
  assign n16726 = n3330 & n9614;
  assign n16727 = x122 & n3500;
  assign n16728 = x124 & n3502;
  assign n16729 = ~n16727 & ~n16728;
  assign n16730 = x123 & n3334;
  assign n16731 = n16729 & ~n16730;
  assign n16732 = ~n16726 & n16731;
  assign n16733 = n16732 ^ x35;
  assign n16714 = n4415 & n7919;
  assign n16715 = x116 & n4420;
  assign n16716 = x118 & n4614;
  assign n16717 = ~n16715 & ~n16716;
  assign n16718 = x117 & n4410;
  assign n16719 = n16717 & ~n16718;
  assign n16720 = ~n16714 & n16719;
  assign n16721 = n16720 ^ x41;
  assign n16704 = n5010 & n7150;
  assign n16705 = x113 & n5223;
  assign n16706 = x115 & n5226;
  assign n16707 = ~n16705 & ~n16706;
  assign n16708 = x114 & n5014;
  assign n16709 = n16707 & ~n16708;
  assign n16710 = ~n16704 & n16709;
  assign n16711 = n16710 ^ x44;
  assign n16694 = n5656 & n6420;
  assign n16695 = x110 & n5895;
  assign n16696 = x111 & n5662;
  assign n16697 = ~n16695 & ~n16696;
  assign n16698 = x112 & n6111;
  assign n16699 = n16697 & ~n16698;
  assign n16700 = ~n16694 & n16699;
  assign n16701 = n16700 ^ x47;
  assign n16684 = ~n5737 & n6326;
  assign n16685 = x107 & n6565;
  assign n16686 = x108 & n6331;
  assign n16687 = ~n16685 & ~n16686;
  assign n16688 = x109 & n6569;
  assign n16689 = n16687 & ~n16688;
  assign n16690 = ~n16684 & n16689;
  assign n16691 = n16690 ^ x50;
  assign n16681 = n16524 ^ n16521;
  assign n16682 = n16533 & ~n16681;
  assign n16683 = n16682 ^ n16532;
  assign n16692 = n16691 ^ n16683;
  assign n16671 = n5088 & n7076;
  assign n16672 = x104 & n7317;
  assign n16673 = x105 & n7080;
  assign n16674 = ~n16672 & ~n16673;
  assign n16675 = x106 & n7319;
  assign n16676 = n16674 & ~n16675;
  assign n16677 = ~n16671 & n16676;
  assign n16678 = n16677 ^ x53;
  assign n16668 = n16511 ^ n16508;
  assign n16669 = n16520 & ~n16668;
  assign n16670 = n16669 ^ n16519;
  assign n16679 = n16678 ^ n16670;
  assign n16658 = n4481 & n7830;
  assign n16659 = x101 & n7839;
  assign n16660 = x103 & n8374;
  assign n16661 = ~n16659 & ~n16660;
  assign n16662 = x102 & n7834;
  assign n16663 = n16661 & ~n16662;
  assign n16664 = ~n16658 & n16663;
  assign n16665 = n16664 ^ x56;
  assign n16655 = n16498 ^ n16495;
  assign n16656 = n16507 & ~n16655;
  assign n16657 = n16656 ^ n16506;
  assign n16666 = n16665 ^ n16657;
  assign n16645 = n3925 & n8622;
  assign n16646 = x98 & n8631;
  assign n16647 = x99 & n8626;
  assign n16648 = ~n16646 & ~n16647;
  assign n16649 = x100 & n9186;
  assign n16650 = n16648 & ~n16649;
  assign n16651 = ~n16645 & n16650;
  assign n16652 = n16651 ^ x59;
  assign n16642 = n16494 ^ n16485;
  assign n16643 = ~n16486 & n16642;
  assign n16644 = n16643 ^ n16494;
  assign n16653 = n16652 ^ n16644;
  assign n16632 = n3388 & n9499;
  assign n16633 = x95 & n9508;
  assign n16634 = x96 & n9503;
  assign n16635 = ~n16633 & ~n16634;
  assign n16636 = x97 & n10106;
  assign n16637 = n16635 & ~n16636;
  assign n16638 = ~n16632 & n16637;
  assign n16639 = n16638 ^ x62;
  assign n16628 = n2433 & n10099;
  assign n16629 = n2570 & n9798;
  assign n16630 = ~n16628 & ~n16629;
  assign n16631 = n16630 ^ x29;
  assign n16640 = n16639 ^ n16631;
  assign n16626 = n16473 & n16484;
  assign n16627 = n16626 ^ n16483;
  assign n16641 = n16640 ^ n16627;
  assign n16654 = n16653 ^ n16641;
  assign n16667 = n16666 ^ n16654;
  assign n16680 = n16679 ^ n16667;
  assign n16693 = n16692 ^ n16680;
  assign n16702 = n16701 ^ n16693;
  assign n16623 = n16543 ^ n16462;
  assign n16624 = ~n16535 & n16623;
  assign n16625 = n16624 ^ n16543;
  assign n16703 = n16702 ^ n16625;
  assign n16712 = n16711 ^ n16703;
  assign n16620 = n16544 ^ n16456;
  assign n16621 = n16545 & ~n16620;
  assign n16622 = n16621 ^ n16459;
  assign n16713 = n16712 ^ n16622;
  assign n16722 = n16721 ^ n16713;
  assign n16617 = n16555 ^ n16546;
  assign n16618 = n16547 & n16617;
  assign n16619 = n16618 ^ n16555;
  assign n16723 = n16722 ^ n16619;
  assign n16614 = n16565 ^ n16556;
  assign n16615 = n16557 & ~n16614;
  assign n16616 = n16615 ^ n16565;
  assign n16724 = n16723 ^ n16616;
  assign n16606 = n3829 & n8715;
  assign n16607 = x119 & n4049;
  assign n16608 = x121 & n4052;
  assign n16609 = ~n16607 & ~n16608;
  assign n16610 = x120 & n3833;
  assign n16611 = n16609 & ~n16610;
  assign n16612 = ~n16606 & n16611;
  assign n16613 = n16612 ^ x38;
  assign n16725 = n16724 ^ n16613;
  assign n16734 = n16733 ^ n16725;
  assign n16603 = n16575 ^ n16442;
  assign n16604 = n16567 & n16603;
  assign n16605 = n16604 ^ n16575;
  assign n16735 = n16734 ^ n16605;
  assign n16744 = n16743 ^ n16735;
  assign n16752 = n16751 ^ n16744;
  assign n16600 = n16433 ^ n16430;
  assign n16601 = ~n16598 & n16600;
  assign n16602 = n16601 ^ n16430;
  assign n16753 = n16752 ^ n16602;
  assign n16902 = ~n16735 & ~n16743;
  assign n16903 = ~n16747 & n16902;
  assign n16904 = n16735 & n16743;
  assign n16905 = n16747 & n16904;
  assign n16906 = ~n16903 & ~n16905;
  assign n16907 = n16751 & ~n16906;
  assign n16908 = ~n16747 & ~n16904;
  assign n16909 = ~n16902 & ~n16908;
  assign n16912 = n16750 & ~n16909;
  assign n16913 = ~n16903 & ~n16912;
  assign n16910 = ~n16750 & n16909;
  assign n16911 = ~n16905 & ~n16910;
  assign n16914 = n16913 ^ n16911;
  assign n16915 = n16602 & n16914;
  assign n16916 = n16915 ^ n16913;
  assign n16917 = ~n16907 & n16916;
  assign n16891 = n3330 & n9912;
  assign n16892 = x123 & n3500;
  assign n16893 = x125 & n3502;
  assign n16894 = ~n16892 & ~n16893;
  assign n16895 = x124 & n3334;
  assign n16896 = n16894 & ~n16895;
  assign n16897 = ~n16891 & n16896;
  assign n16898 = n16897 ^ x35;
  assign n16881 = n3829 & n9001;
  assign n16882 = x120 & n4049;
  assign n16883 = x122 & n4052;
  assign n16884 = ~n16882 & ~n16883;
  assign n16885 = x121 & n3833;
  assign n16886 = n16884 & ~n16885;
  assign n16887 = ~n16881 & n16886;
  assign n16888 = n16887 ^ x38;
  assign n16869 = n5010 & n7393;
  assign n16870 = x114 & n5223;
  assign n16871 = x116 & n5226;
  assign n16872 = ~n16870 & ~n16871;
  assign n16873 = x115 & n5014;
  assign n16874 = n16872 & ~n16873;
  assign n16875 = ~n16869 & n16874;
  assign n16876 = n16875 ^ x44;
  assign n16859 = n5656 & n6656;
  assign n16860 = x111 & n5895;
  assign n16861 = x113 & n6111;
  assign n16862 = ~n16860 & ~n16861;
  assign n16863 = x112 & n5662;
  assign n16864 = n16862 & ~n16863;
  assign n16865 = ~n16859 & n16864;
  assign n16866 = n16865 ^ x47;
  assign n16848 = n5955 & n6326;
  assign n16849 = x108 & n6565;
  assign n16850 = x109 & n6331;
  assign n16851 = ~n16849 & ~n16850;
  assign n16852 = x110 & n6569;
  assign n16853 = n16851 & ~n16852;
  assign n16854 = ~n16848 & n16853;
  assign n16855 = n16854 ^ x50;
  assign n16845 = n16678 ^ n16667;
  assign n16846 = n16679 & ~n16845;
  assign n16847 = n16846 ^ n16670;
  assign n16856 = n16855 ^ n16847;
  assign n16835 = n5297 & n7076;
  assign n16836 = x106 & n7080;
  assign n16837 = x105 & n7317;
  assign n16838 = ~n16836 & ~n16837;
  assign n16839 = x107 & n7319;
  assign n16840 = n16838 & ~n16839;
  assign n16841 = ~n16835 & n16840;
  assign n16842 = n16841 ^ x53;
  assign n16832 = n16665 ^ n16654;
  assign n16833 = n16666 & ~n16832;
  assign n16834 = n16833 ^ n16657;
  assign n16843 = n16842 ^ n16834;
  assign n16822 = n4670 & n7830;
  assign n16823 = x103 & n7834;
  assign n16824 = x102 & n7839;
  assign n16825 = ~n16823 & ~n16824;
  assign n16826 = x104 & n8374;
  assign n16827 = n16825 & ~n16826;
  assign n16828 = ~n16822 & n16827;
  assign n16829 = n16828 ^ x56;
  assign n16812 = n4105 & n8622;
  assign n16813 = x99 & n8631;
  assign n16814 = x101 & n9186;
  assign n16815 = ~n16813 & ~n16814;
  assign n16816 = x100 & n8626;
  assign n16817 = n16815 & ~n16816;
  assign n16818 = ~n16812 & n16817;
  assign n16819 = n16818 ^ x59;
  assign n16802 = n3556 & n9499;
  assign n16803 = x97 & n9503;
  assign n16804 = x96 & n9508;
  assign n16805 = ~n16803 & ~n16804;
  assign n16806 = x98 & n10106;
  assign n16807 = n16805 & ~n16806;
  assign n16808 = ~n16802 & n16807;
  assign n16809 = n16808 ^ x62;
  assign n16795 = ~x29 & x93;
  assign n16796 = ~n16481 & ~n16795;
  assign n16797 = x94 & ~n10099;
  assign n16798 = n16796 & ~n16797;
  assign n16799 = x29 & ~x93;
  assign n16800 = ~n12465 & ~n16799;
  assign n16801 = ~n16798 & n16800;
  assign n16810 = n16809 ^ n16801;
  assign n16792 = x94 & n10099;
  assign n16793 = x95 & n9798;
  assign n16794 = ~n16792 & ~n16793;
  assign n16811 = n16810 ^ n16794;
  assign n16820 = n16819 ^ n16811;
  assign n16789 = n16639 ^ n16627;
  assign n16790 = n16640 & ~n16789;
  assign n16791 = n16790 ^ n16627;
  assign n16821 = n16820 ^ n16791;
  assign n16830 = n16829 ^ n16821;
  assign n16786 = n16652 ^ n16641;
  assign n16787 = n16653 & ~n16786;
  assign n16788 = n16787 ^ n16644;
  assign n16831 = n16830 ^ n16788;
  assign n16844 = n16843 ^ n16831;
  assign n16857 = n16856 ^ n16844;
  assign n16783 = n16691 ^ n16680;
  assign n16784 = n16692 & ~n16783;
  assign n16785 = n16784 ^ n16683;
  assign n16858 = n16857 ^ n16785;
  assign n16867 = n16866 ^ n16858;
  assign n16780 = n16701 ^ n16625;
  assign n16781 = ~n16702 & n16780;
  assign n16782 = n16781 ^ n16625;
  assign n16868 = n16867 ^ n16782;
  assign n16877 = n16876 ^ n16868;
  assign n16777 = n16711 ^ n16622;
  assign n16778 = ~n16712 & n16777;
  assign n16779 = n16778 ^ n16622;
  assign n16878 = n16877 ^ n16779;
  assign n16769 = n4415 & n8169;
  assign n16770 = x117 & n4420;
  assign n16771 = x118 & n4410;
  assign n16772 = ~n16770 & ~n16771;
  assign n16773 = x119 & n4614;
  assign n16774 = n16772 & ~n16773;
  assign n16775 = ~n16769 & n16774;
  assign n16776 = n16775 ^ x41;
  assign n16879 = n16878 ^ n16776;
  assign n16766 = n16721 ^ n16619;
  assign n16767 = ~n16722 & n16766;
  assign n16768 = n16767 ^ n16619;
  assign n16880 = n16879 ^ n16768;
  assign n16889 = n16888 ^ n16880;
  assign n16763 = n16723 ^ n16613;
  assign n16764 = n16724 & ~n16763;
  assign n16765 = n16764 ^ n16616;
  assign n16890 = n16889 ^ n16765;
  assign n16899 = n16898 ^ n16890;
  assign n16760 = n16733 ^ n16605;
  assign n16761 = ~n16734 & n16760;
  assign n16762 = n16761 ^ n16605;
  assign n16900 = n16899 ^ n16762;
  assign n16754 = n2836 & ~n9889;
  assign n16755 = x127 & n2840;
  assign n16756 = x126 & n2996;
  assign n16757 = ~n16755 & ~n16756;
  assign n16758 = ~n16754 & n16757;
  assign n16759 = n16758 ^ x32;
  assign n16901 = n16900 ^ n16759;
  assign n16918 = n16917 ^ n16901;
  assign n17067 = ~n16747 & n16750;
  assign n17068 = ~n16901 & ~n17067;
  assign n17069 = ~n16904 & ~n17068;
  assign n17070 = n16747 & ~n16750;
  assign n17071 = ~n16901 & ~n16902;
  assign n17072 = ~n17070 & ~n17071;
  assign n17073 = ~n17069 & ~n17072;
  assign n17074 = ~n16602 & ~n17073;
  assign n17075 = n16902 & ~n17068;
  assign n17076 = ~n16750 & ~n16908;
  assign n17077 = n16901 & ~n16905;
  assign n17078 = ~n17076 & n17077;
  assign n17079 = ~n17075 & ~n17078;
  assign n17080 = ~n17074 & n17079;
  assign n17054 = ~x31 & n10430;
  assign n17055 = n17054 ^ n9886;
  assign n17056 = ~n2827 & n17055;
  assign n17057 = x32 & n9886;
  assign n17058 = n17056 & ~n17057;
  assign n17059 = n2823 ^ x31;
  assign n17060 = n2835 & n17059;
  assign n17061 = x127 & n17060;
  assign n17062 = n17061 ^ x32;
  assign n17063 = ~n17058 & n17062;
  assign n17045 = n3330 & ~n10174;
  assign n17046 = x124 & n3500;
  assign n17047 = x126 & n3502;
  assign n17048 = ~n17046 & ~n17047;
  assign n17049 = x125 & n3334;
  assign n17050 = n17048 & ~n17049;
  assign n17051 = ~n17045 & n17050;
  assign n17052 = n17051 ^ x35;
  assign n17035 = n3829 & n9309;
  assign n17036 = x121 & n4049;
  assign n17037 = x122 & n3833;
  assign n17038 = ~n17036 & ~n17037;
  assign n17039 = x123 & n4052;
  assign n17040 = n17038 & ~n17039;
  assign n17041 = ~n17035 & n17040;
  assign n17042 = n17041 ^ x38;
  assign n17025 = n4415 & ~n8424;
  assign n17026 = x118 & n4420;
  assign n17027 = x120 & n4614;
  assign n17028 = ~n17026 & ~n17027;
  assign n17029 = x119 & n4410;
  assign n17030 = n17028 & ~n17029;
  assign n17031 = ~n17025 & n17030;
  assign n17032 = n17031 ^ x41;
  assign n17015 = n5010 & n7643;
  assign n17016 = x115 & n5223;
  assign n17017 = x117 & n5226;
  assign n17018 = ~n17016 & ~n17017;
  assign n17019 = x116 & n5014;
  assign n17020 = n17018 & ~n17019;
  assign n17021 = ~n17015 & n17020;
  assign n17022 = n17021 ^ x44;
  assign n17005 = n5656 & n6892;
  assign n17006 = x112 & n5895;
  assign n17007 = x114 & n6111;
  assign n17008 = ~n17006 & ~n17007;
  assign n17009 = x113 & n5662;
  assign n17010 = n17008 & ~n17009;
  assign n17011 = ~n17005 & n17010;
  assign n17012 = n17011 ^ x47;
  assign n16995 = n6178 & n6326;
  assign n16996 = x109 & n6565;
  assign n16997 = x110 & n6331;
  assign n16998 = ~n16996 & ~n16997;
  assign n16999 = x111 & n6569;
  assign n17000 = n16998 & ~n16999;
  assign n17001 = ~n16995 & n17000;
  assign n17002 = n17001 ^ x50;
  assign n16984 = ~n5506 & n7076;
  assign n16985 = x106 & n7317;
  assign n16986 = x107 & n7080;
  assign n16987 = ~n16985 & ~n16986;
  assign n16988 = x108 & n7319;
  assign n16989 = n16987 & ~n16988;
  assign n16990 = ~n16984 & n16989;
  assign n16991 = n16990 ^ x53;
  assign n16981 = n16821 ^ n16788;
  assign n16982 = ~n16830 & n16981;
  assign n16983 = n16982 ^ n16829;
  assign n16992 = n16991 ^ n16983;
  assign n16971 = n4867 & n7830;
  assign n16972 = x103 & n7839;
  assign n16973 = x105 & n8374;
  assign n16974 = ~n16972 & ~n16973;
  assign n16975 = x104 & n7834;
  assign n16976 = n16974 & ~n16975;
  assign n16977 = ~n16971 & n16976;
  assign n16978 = n16977 ^ x56;
  assign n16968 = n16811 ^ n16791;
  assign n16969 = n16820 & n16968;
  assign n16970 = n16969 ^ n16819;
  assign n16979 = n16978 ^ n16970;
  assign n16962 = n2715 & n10099;
  assign n16963 = n2881 & n9798;
  assign n16964 = ~n16962 & ~n16963;
  assign n16959 = n16801 ^ n16794;
  assign n16960 = ~n16810 & ~n16959;
  assign n16961 = n16960 ^ n16809;
  assign n16965 = n16964 ^ n16961;
  assign n16951 = n3730 & n9499;
  assign n16952 = x98 & n9503;
  assign n16953 = x97 & n9508;
  assign n16954 = ~n16952 & ~n16953;
  assign n16955 = x99 & n10106;
  assign n16956 = n16954 & ~n16955;
  assign n16957 = ~n16951 & n16956;
  assign n16958 = n16957 ^ x62;
  assign n16966 = n16965 ^ n16958;
  assign n16943 = n4286 & n8622;
  assign n16944 = x100 & n8631;
  assign n16945 = x101 & n8626;
  assign n16946 = ~n16944 & ~n16945;
  assign n16947 = x102 & n9186;
  assign n16948 = n16946 & ~n16947;
  assign n16949 = ~n16943 & n16948;
  assign n16950 = n16949 ^ x59;
  assign n16967 = n16966 ^ n16950;
  assign n16980 = n16979 ^ n16967;
  assign n16993 = n16992 ^ n16980;
  assign n16940 = n16842 ^ n16831;
  assign n16941 = n16843 & n16940;
  assign n16942 = n16941 ^ n16834;
  assign n16994 = n16993 ^ n16942;
  assign n17003 = n17002 ^ n16994;
  assign n16937 = n16855 ^ n16844;
  assign n16938 = n16856 & n16937;
  assign n16939 = n16938 ^ n16847;
  assign n17004 = n17003 ^ n16939;
  assign n17013 = n17012 ^ n17004;
  assign n16934 = n16866 ^ n16857;
  assign n16935 = n16858 & ~n16934;
  assign n16936 = n16935 ^ n16866;
  assign n17014 = n17013 ^ n16936;
  assign n17023 = n17022 ^ n17014;
  assign n16931 = n16876 ^ n16782;
  assign n16932 = n16868 & n16931;
  assign n16933 = n16932 ^ n16876;
  assign n17024 = n17023 ^ n16933;
  assign n17033 = n17032 ^ n17024;
  assign n16928 = n16877 ^ n16776;
  assign n16929 = ~n16878 & n16928;
  assign n16930 = n16929 ^ n16779;
  assign n17034 = n17033 ^ n16930;
  assign n17043 = n17042 ^ n17034;
  assign n16925 = n16888 ^ n16768;
  assign n16926 = n16880 & n16925;
  assign n16927 = n16926 ^ n16888;
  assign n17044 = n17043 ^ n16927;
  assign n17053 = n17052 ^ n17044;
  assign n17064 = n17063 ^ n17053;
  assign n16922 = n16898 ^ n16765;
  assign n16923 = n16890 & n16922;
  assign n16924 = n16923 ^ n16898;
  assign n17065 = n17064 ^ n16924;
  assign n16919 = n16899 ^ n16759;
  assign n16920 = ~n16900 & n16919;
  assign n16921 = n16920 ^ n16762;
  assign n17066 = n17065 ^ n16921;
  assign n17081 = n17080 ^ n17066;
  assign n17221 = n3330 & ~n10447;
  assign n17222 = x125 & n3500;
  assign n17223 = x126 & n3334;
  assign n17224 = ~n17222 & ~n17223;
  assign n17225 = x127 & n3502;
  assign n17226 = n17224 & ~n17225;
  assign n17227 = ~n17221 & n17226;
  assign n17228 = n17227 ^ x35;
  assign n17211 = n3829 & n9614;
  assign n17212 = x122 & n4049;
  assign n17213 = x123 & n3833;
  assign n17214 = ~n17212 & ~n17213;
  assign n17215 = x124 & n4052;
  assign n17216 = n17214 & ~n17215;
  assign n17217 = ~n17211 & n17216;
  assign n17218 = n17217 ^ x38;
  assign n17195 = n6326 & n6420;
  assign n17196 = x110 & n6565;
  assign n17197 = x111 & n6331;
  assign n17198 = ~n17196 & ~n17197;
  assign n17199 = x112 & n6569;
  assign n17200 = n17198 & ~n17199;
  assign n17201 = ~n17195 & n17200;
  assign n17202 = n17201 ^ x50;
  assign n17192 = n17002 ^ n16942;
  assign n17193 = ~n16994 & n17192;
  assign n17194 = n17193 ^ n17002;
  assign n17203 = n17202 ^ n17194;
  assign n17182 = ~n5737 & n7076;
  assign n17183 = x107 & n7317;
  assign n17184 = x109 & n7319;
  assign n17185 = ~n17183 & ~n17184;
  assign n17186 = x108 & n7080;
  assign n17187 = n17185 & ~n17186;
  assign n17188 = ~n17182 & n17187;
  assign n17189 = n17188 ^ x53;
  assign n17179 = n16991 ^ n16980;
  assign n17180 = n16992 & ~n17179;
  assign n17181 = n17180 ^ n16983;
  assign n17190 = n17189 ^ n17181;
  assign n17169 = n5088 & n7830;
  assign n17170 = x104 & n7839;
  assign n17171 = x105 & n7834;
  assign n17172 = ~n17170 & ~n17171;
  assign n17173 = x106 & n8374;
  assign n17174 = n17172 & ~n17173;
  assign n17175 = ~n17169 & n17174;
  assign n17176 = n17175 ^ x56;
  assign n17166 = n16970 ^ n16967;
  assign n17167 = n16979 & ~n17166;
  assign n17168 = n17167 ^ n16978;
  assign n17177 = n17176 ^ n17168;
  assign n17156 = n4481 & n8622;
  assign n17157 = x101 & n8631;
  assign n17158 = x102 & n8626;
  assign n17159 = ~n17157 & ~n17158;
  assign n17160 = x103 & n9186;
  assign n17161 = n17159 & ~n17160;
  assign n17162 = ~n17156 & n17161;
  assign n17163 = n17162 ^ x59;
  assign n17153 = n16958 ^ n16950;
  assign n17154 = n16966 & ~n17153;
  assign n17155 = n17154 ^ n16965;
  assign n17164 = n17163 ^ n17155;
  assign n17141 = ~x95 & n16792;
  assign n17142 = x95 & ~x96;
  assign n17143 = n9798 & n17142;
  assign n17144 = ~n17141 & ~n17143;
  assign n17145 = n16961 & n17144;
  assign n17146 = x95 & n10099;
  assign n17147 = ~x94 & n17146;
  assign n17148 = ~x95 & x96;
  assign n17149 = n9798 & n17148;
  assign n17150 = ~n17147 & ~n17149;
  assign n17151 = ~n17145 & n17150;
  assign n17132 = n3925 & n9499;
  assign n17133 = x98 & n9508;
  assign n17134 = x100 & n10106;
  assign n17135 = ~n17133 & ~n17134;
  assign n17136 = x99 & n9503;
  assign n17137 = n17135 & ~n17136;
  assign n17138 = ~n17132 & n17137;
  assign n17139 = n17138 ^ x62;
  assign n17127 = n2881 & n10099;
  assign n17128 = x97 ^ x96;
  assign n17129 = n9798 & n17128;
  assign n17130 = ~n17127 & ~n17129;
  assign n17131 = n17130 ^ x32;
  assign n17140 = n17139 ^ n17131;
  assign n17152 = n17151 ^ n17140;
  assign n17165 = n17164 ^ n17152;
  assign n17178 = n17177 ^ n17165;
  assign n17191 = n17190 ^ n17178;
  assign n17204 = n17203 ^ n17191;
  assign n17119 = n5656 & n7150;
  assign n17120 = x113 & n5895;
  assign n17121 = x114 & n5662;
  assign n17122 = ~n17120 & ~n17121;
  assign n17123 = x115 & n6111;
  assign n17124 = n17122 & ~n17123;
  assign n17125 = ~n17119 & n17124;
  assign n17126 = n17125 ^ x47;
  assign n17205 = n17204 ^ n17126;
  assign n17116 = n17012 ^ n16939;
  assign n17117 = ~n17004 & n17116;
  assign n17118 = n17117 ^ n17012;
  assign n17206 = n17205 ^ n17118;
  assign n17113 = n17022 ^ n17013;
  assign n17114 = ~n17014 & n17113;
  assign n17115 = n17114 ^ n17022;
  assign n17207 = n17206 ^ n17115;
  assign n17105 = n5010 & n7919;
  assign n17106 = x116 & n5223;
  assign n17107 = x117 & n5014;
  assign n17108 = ~n17106 & ~n17107;
  assign n17109 = x118 & n5226;
  assign n17110 = n17108 & ~n17109;
  assign n17111 = ~n17105 & n17110;
  assign n17112 = n17111 ^ x44;
  assign n17208 = n17207 ^ n17112;
  assign n17102 = n17032 ^ n17023;
  assign n17103 = ~n17024 & n17102;
  assign n17104 = n17103 ^ n17032;
  assign n17209 = n17208 ^ n17104;
  assign n17094 = n4415 & n8715;
  assign n17095 = x119 & n4420;
  assign n17096 = x121 & n4614;
  assign n17097 = ~n17095 & ~n17096;
  assign n17098 = x120 & n4410;
  assign n17099 = n17097 & ~n17098;
  assign n17100 = ~n17094 & n17099;
  assign n17101 = n17100 ^ x41;
  assign n17210 = n17209 ^ n17101;
  assign n17219 = n17218 ^ n17210;
  assign n17091 = n17042 ^ n16930;
  assign n17092 = ~n17034 & n17091;
  assign n17093 = n17092 ^ n17042;
  assign n17220 = n17219 ^ n17093;
  assign n17229 = n17228 ^ n17220;
  assign n17088 = n17052 ^ n17043;
  assign n17089 = ~n17044 & n17088;
  assign n17090 = n17089 ^ n17052;
  assign n17230 = n17229 ^ n17090;
  assign n17085 = n17053 ^ n16924;
  assign n17086 = ~n17064 & ~n17085;
  assign n17087 = n17086 ^ n17063;
  assign n17231 = n17230 ^ n17087;
  assign n17082 = n17080 ^ n16921;
  assign n17083 = n17066 & n17082;
  assign n17084 = n17083 ^ n17080;
  assign n17232 = n17231 ^ n17084;
  assign n17367 = n3330 & ~n9889;
  assign n17368 = x127 & n3334;
  assign n17369 = x126 & n3500;
  assign n17370 = ~n17368 & ~n17369;
  assign n17371 = ~n17367 & n17370;
  assign n17372 = n17371 ^ x35;
  assign n17358 = n3829 & n9912;
  assign n17359 = x123 & n4049;
  assign n17360 = x125 & n4052;
  assign n17361 = ~n17359 & ~n17360;
  assign n17362 = x124 & n3833;
  assign n17363 = n17361 & ~n17362;
  assign n17364 = ~n17358 & n17363;
  assign n17365 = n17364 ^ x38;
  assign n17348 = n4415 & n9001;
  assign n17349 = x120 & n4420;
  assign n17350 = x121 & n4410;
  assign n17351 = ~n17349 & ~n17350;
  assign n17352 = x122 & n4614;
  assign n17353 = n17351 & ~n17352;
  assign n17354 = ~n17348 & n17353;
  assign n17355 = n17354 ^ x41;
  assign n17335 = n5656 & n7393;
  assign n17336 = x114 & n5895;
  assign n17337 = x116 & n6111;
  assign n17338 = ~n17336 & ~n17337;
  assign n17339 = x115 & n5662;
  assign n17340 = n17338 & ~n17339;
  assign n17341 = ~n17335 & n17340;
  assign n17342 = n17341 ^ x47;
  assign n17325 = n6326 & n6656;
  assign n17326 = x111 & n6565;
  assign n17327 = x112 & n6331;
  assign n17328 = ~n17326 & ~n17327;
  assign n17329 = x113 & n6569;
  assign n17330 = n17328 & ~n17329;
  assign n17331 = ~n17325 & n17330;
  assign n17332 = n17331 ^ x50;
  assign n17322 = n17189 ^ n17178;
  assign n17323 = n17190 & ~n17322;
  assign n17324 = n17323 ^ n17181;
  assign n17333 = n17332 ^ n17324;
  assign n17312 = n5955 & n7076;
  assign n17313 = x108 & n7317;
  assign n17314 = x110 & n7319;
  assign n17315 = ~n17313 & ~n17314;
  assign n17316 = x109 & n7080;
  assign n17317 = n17315 & ~n17316;
  assign n17318 = ~n17312 & n17317;
  assign n17319 = n17318 ^ x53;
  assign n17309 = n17176 ^ n17165;
  assign n17310 = n17177 & ~n17309;
  assign n17311 = n17310 ^ n17168;
  assign n17320 = n17319 ^ n17311;
  assign n17299 = n5297 & n7830;
  assign n17300 = x105 & n7839;
  assign n17301 = x106 & n7834;
  assign n17302 = ~n17300 & ~n17301;
  assign n17303 = x107 & n8374;
  assign n17304 = n17302 & ~n17303;
  assign n17305 = ~n17299 & n17304;
  assign n17306 = n17305 ^ x56;
  assign n17296 = n17155 ^ n17152;
  assign n17297 = n17164 & ~n17296;
  assign n17298 = n17297 ^ n17163;
  assign n17307 = n17306 ^ n17298;
  assign n17286 = n4670 & n8622;
  assign n17287 = x102 & n8631;
  assign n17288 = x104 & n9186;
  assign n17289 = ~n17287 & ~n17288;
  assign n17290 = x103 & n8626;
  assign n17291 = n17289 & ~n17290;
  assign n17292 = ~n17286 & n17291;
  assign n17293 = n17292 ^ x59;
  assign n17276 = n4105 & n9499;
  assign n17277 = x99 & n9508;
  assign n17278 = x100 & n9503;
  assign n17279 = ~n17277 & ~n17278;
  assign n17280 = x101 & n10106;
  assign n17281 = n17279 & ~n17280;
  assign n17282 = ~n17276 & n17281;
  assign n17283 = n17282 ^ x62;
  assign n17268 = ~x32 & x96;
  assign n17269 = x97 ^ x95;
  assign n17270 = ~n10099 & n17269;
  assign n17271 = n17270 ^ x95;
  assign n17272 = ~n17268 & ~n17271;
  assign n17273 = x32 & ~x96;
  assign n17274 = ~n12465 & ~n17273;
  assign n17275 = ~n17272 & n17274;
  assign n17284 = n17283 ^ n17275;
  assign n17265 = x98 & n9798;
  assign n17266 = x97 & n10099;
  assign n17267 = ~n17265 & ~n17266;
  assign n17285 = n17284 ^ n17267;
  assign n17294 = n17293 ^ n17285;
  assign n17262 = n17151 ^ n17139;
  assign n17263 = n17140 & ~n17262;
  assign n17264 = n17263 ^ n17151;
  assign n17295 = n17294 ^ n17264;
  assign n17308 = n17307 ^ n17295;
  assign n17321 = n17320 ^ n17308;
  assign n17334 = n17333 ^ n17321;
  assign n17343 = n17342 ^ n17334;
  assign n17259 = n17202 ^ n17191;
  assign n17260 = n17203 & ~n17259;
  assign n17261 = n17260 ^ n17194;
  assign n17344 = n17343 ^ n17261;
  assign n17256 = n17126 ^ n17118;
  assign n17257 = n17205 & ~n17256;
  assign n17258 = n17257 ^ n17204;
  assign n17345 = n17344 ^ n17258;
  assign n17248 = n5010 & n8169;
  assign n17249 = x117 & n5223;
  assign n17250 = x118 & n5014;
  assign n17251 = ~n17249 & ~n17250;
  assign n17252 = x119 & n5226;
  assign n17253 = n17251 & ~n17252;
  assign n17254 = ~n17248 & n17253;
  assign n17255 = n17254 ^ x44;
  assign n17346 = n17345 ^ n17255;
  assign n17245 = n17206 ^ n17112;
  assign n17246 = n17207 & ~n17245;
  assign n17247 = n17246 ^ n17115;
  assign n17347 = n17346 ^ n17247;
  assign n17356 = n17355 ^ n17347;
  assign n17242 = n17208 ^ n17101;
  assign n17243 = n17209 & ~n17242;
  assign n17244 = n17243 ^ n17104;
  assign n17357 = n17356 ^ n17244;
  assign n17366 = n17365 ^ n17357;
  assign n17373 = n17372 ^ n17366;
  assign n17239 = n17218 ^ n17093;
  assign n17240 = ~n17219 & n17239;
  assign n17241 = n17240 ^ n17093;
  assign n17374 = n17373 ^ n17241;
  assign n17236 = n17220 ^ n17090;
  assign n17237 = n17229 & ~n17236;
  assign n17238 = n17237 ^ n17228;
  assign n17375 = n17374 ^ n17238;
  assign n17233 = n17087 ^ n17084;
  assign n17234 = n17231 & ~n17233;
  assign n17235 = n17234 ^ n17084;
  assign n17376 = n17375 ^ n17235;
  assign n17513 = n17366 & ~n17372;
  assign n17514 = n17241 ^ n17238;
  assign n17515 = ~n17366 & n17372;
  assign n17516 = n17515 ^ n17241;
  assign n17517 = n17514 & ~n17516;
  assign n17518 = n17517 ^ n17238;
  assign n17519 = ~n17513 & n17518;
  assign n17507 = n17238 & n17241;
  assign n17508 = ~n17238 & ~n17241;
  assign n17509 = n17508 ^ n17366;
  assign n17510 = ~n17373 & ~n17509;
  assign n17511 = n17510 ^ n17372;
  assign n17512 = ~n17507 & ~n17511;
  assign n17520 = n17519 ^ n17512;
  assign n17521 = ~n17235 & n17520;
  assign n17522 = n17521 ^ n17519;
  assign n17523 = n17366 ^ n17241;
  assign n17524 = ~n17514 & n17523;
  assign n17525 = n17373 & n17524;
  assign n17526 = ~n17522 & ~n17525;
  assign n17497 = n2992 & n10430;
  assign n17498 = x127 & n3317;
  assign n17499 = x35 & ~n17498;
  assign n17500 = ~n17497 & n17499;
  assign n17501 = ~x34 & ~n17500;
  assign n17502 = x127 & n3321;
  assign n17503 = ~x35 & ~n17502;
  assign n17504 = ~n17497 & n17503;
  assign n17505 = ~n17501 & ~n17504;
  assign n17487 = n3829 & ~n10174;
  assign n17488 = x124 & n4049;
  assign n17489 = x126 & n4052;
  assign n17490 = ~n17488 & ~n17489;
  assign n17491 = x125 & n3833;
  assign n17492 = n17490 & ~n17491;
  assign n17493 = ~n17487 & n17492;
  assign n17494 = n17493 ^ x38;
  assign n17477 = n4415 & n9309;
  assign n17478 = x121 & n4420;
  assign n17479 = x123 & n4614;
  assign n17480 = ~n17478 & ~n17479;
  assign n17481 = x122 & n4410;
  assign n17482 = n17480 & ~n17481;
  assign n17483 = ~n17477 & n17482;
  assign n17484 = n17483 ^ x41;
  assign n17465 = n5656 & n7643;
  assign n17466 = x115 & n5895;
  assign n17467 = x117 & n6111;
  assign n17468 = ~n17466 & ~n17467;
  assign n17469 = x116 & n5662;
  assign n17470 = n17468 & ~n17469;
  assign n17471 = ~n17465 & n17470;
  assign n17472 = n17471 ^ x47;
  assign n17454 = n6326 & n6892;
  assign n17455 = x112 & n6565;
  assign n17456 = x113 & n6331;
  assign n17457 = ~n17455 & ~n17456;
  assign n17458 = x114 & n6569;
  assign n17459 = n17457 & ~n17458;
  assign n17460 = ~n17454 & n17459;
  assign n17461 = n17460 ^ x50;
  assign n17451 = n17319 ^ n17308;
  assign n17452 = n17320 & n17451;
  assign n17453 = n17452 ^ n17311;
  assign n17462 = n17461 ^ n17453;
  assign n17441 = n6178 & n7076;
  assign n17442 = x110 & n7080;
  assign n17443 = x109 & n7317;
  assign n17444 = ~n17442 & ~n17443;
  assign n17445 = x111 & n7319;
  assign n17446 = n17444 & ~n17445;
  assign n17447 = ~n17441 & n17446;
  assign n17448 = n17447 ^ x53;
  assign n17438 = n17298 ^ n17295;
  assign n17439 = n17307 & n17438;
  assign n17440 = n17439 ^ n17306;
  assign n17449 = n17448 ^ n17440;
  assign n17428 = ~n5506 & n7830;
  assign n17429 = x106 & n7839;
  assign n17430 = x107 & n7834;
  assign n17431 = ~n17429 & ~n17430;
  assign n17432 = x108 & n8374;
  assign n17433 = n17431 & ~n17432;
  assign n17434 = ~n17428 & n17433;
  assign n17435 = n17434 ^ x56;
  assign n17425 = n17285 ^ n17264;
  assign n17426 = n17294 & n17425;
  assign n17427 = n17426 ^ n17293;
  assign n17436 = n17435 ^ n17427;
  assign n17416 = n4867 & n8622;
  assign n17417 = x103 & n8631;
  assign n17418 = x104 & n8626;
  assign n17419 = ~n17417 & ~n17418;
  assign n17420 = x105 & n9186;
  assign n17421 = n17419 & ~n17420;
  assign n17422 = ~n17416 & n17421;
  assign n17423 = n17422 ^ x59;
  assign n17411 = n3198 & n10099;
  assign n17412 = n3373 & n9798;
  assign n17413 = ~n17411 & ~n17412;
  assign n17408 = n17275 ^ n17267;
  assign n17409 = ~n17284 & ~n17408;
  assign n17410 = n17409 ^ n17283;
  assign n17414 = n17413 ^ n17410;
  assign n17400 = n4286 & n9499;
  assign n17401 = x100 & n9508;
  assign n17402 = x102 & n10106;
  assign n17403 = ~n17401 & ~n17402;
  assign n17404 = x101 & n9503;
  assign n17405 = n17403 & ~n17404;
  assign n17406 = ~n17400 & n17405;
  assign n17407 = n17406 ^ x62;
  assign n17415 = n17414 ^ n17407;
  assign n17424 = n17423 ^ n17415;
  assign n17437 = n17436 ^ n17424;
  assign n17450 = n17449 ^ n17437;
  assign n17463 = n17462 ^ n17450;
  assign n17397 = n17324 ^ n17321;
  assign n17398 = n17333 & n17397;
  assign n17399 = n17398 ^ n17332;
  assign n17464 = n17463 ^ n17399;
  assign n17473 = n17472 ^ n17464;
  assign n17394 = n17342 ^ n17261;
  assign n17395 = n17343 & n17394;
  assign n17396 = n17395 ^ n17261;
  assign n17474 = n17473 ^ n17396;
  assign n17386 = n5010 & ~n8424;
  assign n17387 = x118 & n5223;
  assign n17388 = x120 & n5226;
  assign n17389 = ~n17387 & ~n17388;
  assign n17390 = x119 & n5014;
  assign n17391 = n17389 & ~n17390;
  assign n17392 = ~n17386 & n17391;
  assign n17393 = n17392 ^ x44;
  assign n17475 = n17474 ^ n17393;
  assign n17383 = n17344 ^ n17255;
  assign n17384 = ~n17345 & n17383;
  assign n17385 = n17384 ^ n17258;
  assign n17476 = n17475 ^ n17385;
  assign n17485 = n17484 ^ n17476;
  assign n17380 = n17355 ^ n17247;
  assign n17381 = n17347 & n17380;
  assign n17382 = n17381 ^ n17355;
  assign n17486 = n17485 ^ n17382;
  assign n17495 = n17494 ^ n17486;
  assign n17377 = n17365 ^ n17356;
  assign n17378 = n17357 & ~n17377;
  assign n17379 = n17378 ^ n17365;
  assign n17496 = n17495 ^ n17379;
  assign n17506 = n17505 ^ n17496;
  assign n17527 = n17526 ^ n17506;
  assign n17661 = n17506 & ~n17507;
  assign n17662 = ~n17513 & ~n17661;
  assign n17663 = n17506 & ~n17515;
  assign n17664 = ~n17508 & ~n17663;
  assign n17665 = ~n17662 & ~n17664;
  assign n17666 = n17235 & ~n17665;
  assign n17667 = ~n17506 & n17511;
  assign n17668 = n17507 & n17664;
  assign n17669 = ~n17667 & ~n17668;
  assign n17670 = ~n17666 & n17669;
  assign n17650 = n3829 & ~n10447;
  assign n17651 = x125 & n4049;
  assign n17652 = x127 & n4052;
  assign n17653 = ~n17651 & ~n17652;
  assign n17654 = x126 & n3833;
  assign n17655 = n17653 & ~n17654;
  assign n17656 = ~n17650 & n17655;
  assign n17657 = n17656 ^ x38;
  assign n17640 = n4415 & n9614;
  assign n17641 = x122 & n4420;
  assign n17642 = x123 & n4410;
  assign n17643 = ~n17641 & ~n17642;
  assign n17644 = x124 & n4614;
  assign n17645 = n17643 & ~n17644;
  assign n17646 = ~n17640 & n17645;
  assign n17647 = n17646 ^ x41;
  assign n17630 = n5010 & n8715;
  assign n17631 = x119 & n5223;
  assign n17632 = x121 & n5226;
  assign n17633 = ~n17631 & ~n17632;
  assign n17634 = x120 & n5014;
  assign n17635 = n17633 & ~n17634;
  assign n17636 = ~n17630 & n17635;
  assign n17637 = n17636 ^ x44;
  assign n17616 = n6420 & n7076;
  assign n17617 = x111 & n7080;
  assign n17618 = x110 & n7317;
  assign n17619 = ~n17617 & ~n17618;
  assign n17620 = x112 & n7319;
  assign n17621 = n17619 & ~n17620;
  assign n17622 = ~n17616 & n17621;
  assign n17623 = n17622 ^ x53;
  assign n17606 = ~n5737 & n7830;
  assign n17607 = x107 & n7839;
  assign n17608 = x109 & n8374;
  assign n17609 = ~n17607 & ~n17608;
  assign n17610 = x108 & n7834;
  assign n17611 = n17609 & ~n17610;
  assign n17612 = ~n17606 & n17611;
  assign n17613 = n17612 ^ x56;
  assign n17603 = n17435 ^ n17424;
  assign n17604 = n17436 & ~n17603;
  assign n17605 = n17604 ^ n17427;
  assign n17614 = n17613 ^ n17605;
  assign n17593 = n5088 & n8622;
  assign n17594 = x104 & n8631;
  assign n17595 = x106 & n9186;
  assign n17596 = ~n17594 & ~n17595;
  assign n17597 = x105 & n8626;
  assign n17598 = n17596 & ~n17597;
  assign n17599 = ~n17593 & n17598;
  assign n17600 = n17599 ^ x59;
  assign n17590 = n17423 ^ n17414;
  assign n17591 = ~n17415 & n17590;
  assign n17592 = n17591 ^ n17423;
  assign n17601 = n17600 ^ n17592;
  assign n17578 = ~x98 & n17266;
  assign n17579 = x98 & ~x99;
  assign n17580 = n9798 & n17579;
  assign n17581 = ~n17578 & ~n17580;
  assign n17582 = n17410 & n17581;
  assign n17583 = x98 & n10099;
  assign n17584 = ~x97 & n17583;
  assign n17585 = ~x98 & x99;
  assign n17586 = n9798 & n17585;
  assign n17587 = ~n17584 & ~n17586;
  assign n17588 = ~n17582 & n17587;
  assign n17569 = n4481 & n9499;
  assign n17570 = x101 & n9508;
  assign n17571 = x103 & n10106;
  assign n17572 = ~n17570 & ~n17571;
  assign n17573 = x102 & n9503;
  assign n17574 = n17572 & ~n17573;
  assign n17575 = ~n17569 & n17574;
  assign n17576 = n17575 ^ x62;
  assign n17565 = n3373 & n10099;
  assign n17566 = n3538 & n9798;
  assign n17567 = ~n17565 & ~n17566;
  assign n17568 = n17567 ^ x35;
  assign n17577 = n17576 ^ n17568;
  assign n17589 = n17588 ^ n17577;
  assign n17602 = n17601 ^ n17589;
  assign n17615 = n17614 ^ n17602;
  assign n17624 = n17623 ^ n17615;
  assign n17562 = n17440 ^ n17437;
  assign n17563 = n17449 & ~n17562;
  assign n17564 = n17563 ^ n17448;
  assign n17625 = n17624 ^ n17564;
  assign n17559 = n17453 ^ n17450;
  assign n17560 = n17462 & ~n17559;
  assign n17561 = n17560 ^ n17461;
  assign n17626 = n17625 ^ n17561;
  assign n17551 = n6326 & n7150;
  assign n17552 = x113 & n6565;
  assign n17553 = x115 & n6569;
  assign n17554 = ~n17552 & ~n17553;
  assign n17555 = x114 & n6331;
  assign n17556 = n17554 & ~n17555;
  assign n17557 = ~n17551 & n17556;
  assign n17558 = n17557 ^ x50;
  assign n17627 = n17626 ^ n17558;
  assign n17543 = n5656 & n7919;
  assign n17544 = x116 & n5895;
  assign n17545 = x117 & n5662;
  assign n17546 = ~n17544 & ~n17545;
  assign n17547 = x118 & n6111;
  assign n17548 = n17546 & ~n17547;
  assign n17549 = ~n17543 & n17548;
  assign n17550 = n17549 ^ x47;
  assign n17628 = n17627 ^ n17550;
  assign n17540 = n17472 ^ n17463;
  assign n17541 = ~n17464 & n17540;
  assign n17542 = n17541 ^ n17472;
  assign n17629 = n17628 ^ n17542;
  assign n17638 = n17637 ^ n17629;
  assign n17537 = n17473 ^ n17393;
  assign n17538 = n17474 & ~n17537;
  assign n17539 = n17538 ^ n17396;
  assign n17639 = n17638 ^ n17539;
  assign n17648 = n17647 ^ n17639;
  assign n17534 = n17484 ^ n17385;
  assign n17535 = ~n17476 & n17534;
  assign n17536 = n17535 ^ n17484;
  assign n17649 = n17648 ^ n17536;
  assign n17658 = n17657 ^ n17649;
  assign n17531 = n17494 ^ n17485;
  assign n17532 = ~n17486 & n17531;
  assign n17533 = n17532 ^ n17494;
  assign n17659 = n17658 ^ n17533;
  assign n17528 = n17505 ^ n17495;
  assign n17529 = ~n17496 & ~n17528;
  assign n17530 = n17529 ^ n17505;
  assign n17660 = n17659 ^ n17530;
  assign n17671 = n17670 ^ n17660;
  assign n17789 = n4415 & n9912;
  assign n17790 = x123 & n4420;
  assign n17791 = x124 & n4410;
  assign n17792 = ~n17790 & ~n17791;
  assign n17793 = x125 & n4614;
  assign n17794 = n17792 & ~n17793;
  assign n17795 = ~n17789 & n17794;
  assign n17796 = n17795 ^ x41;
  assign n17779 = n5010 & n9001;
  assign n17780 = x120 & n5223;
  assign n17781 = x121 & n5014;
  assign n17782 = ~n17780 & ~n17781;
  assign n17783 = x122 & n5226;
  assign n17784 = n17782 & ~n17783;
  assign n17785 = ~n17779 & n17784;
  assign n17786 = n17785 ^ x44;
  assign n17766 = n6326 & n7393;
  assign n17767 = x114 & n6565;
  assign n17768 = x116 & n6569;
  assign n17769 = ~n17767 & ~n17768;
  assign n17770 = x115 & n6331;
  assign n17771 = n17769 & ~n17770;
  assign n17772 = ~n17766 & n17771;
  assign n17773 = n17772 ^ x50;
  assign n17763 = n17623 ^ n17564;
  assign n17764 = ~n17624 & n17763;
  assign n17765 = n17764 ^ n17564;
  assign n17774 = n17773 ^ n17765;
  assign n17753 = n6656 & n7076;
  assign n17754 = x111 & n7317;
  assign n17755 = x112 & n7080;
  assign n17756 = ~n17754 & ~n17755;
  assign n17757 = x113 & n7319;
  assign n17758 = n17756 & ~n17757;
  assign n17759 = ~n17753 & n17758;
  assign n17760 = n17759 ^ x53;
  assign n17750 = n17613 ^ n17602;
  assign n17751 = n17614 & ~n17750;
  assign n17752 = n17751 ^ n17605;
  assign n17761 = n17760 ^ n17752;
  assign n17740 = n5955 & n7830;
  assign n17741 = x108 & n7839;
  assign n17742 = x110 & n8374;
  assign n17743 = ~n17741 & ~n17742;
  assign n17744 = x109 & n7834;
  assign n17745 = n17743 & ~n17744;
  assign n17746 = ~n17740 & n17745;
  assign n17747 = n17746 ^ x56;
  assign n17737 = n17600 ^ n17589;
  assign n17738 = n17601 & ~n17737;
  assign n17739 = n17738 ^ n17592;
  assign n17748 = n17747 ^ n17739;
  assign n17727 = n5297 & n8622;
  assign n17728 = x105 & n8631;
  assign n17729 = x106 & n8626;
  assign n17730 = ~n17728 & ~n17729;
  assign n17731 = x107 & n9186;
  assign n17732 = n17730 & ~n17731;
  assign n17733 = ~n17727 & n17732;
  assign n17734 = n17733 ^ x59;
  assign n17724 = n17588 ^ n17576;
  assign n17725 = n17577 & ~n17724;
  assign n17726 = n17725 ^ n17588;
  assign n17735 = n17734 ^ n17726;
  assign n17715 = n4670 & n9499;
  assign n17716 = x102 & n9508;
  assign n17717 = x103 & n9503;
  assign n17718 = ~n17716 & ~n17717;
  assign n17719 = x104 & n10106;
  assign n17720 = n17718 & ~n17719;
  assign n17721 = ~n17715 & n17720;
  assign n17722 = n17721 ^ x62;
  assign n17707 = ~x35 & x99;
  assign n17708 = n3539 & ~n10099;
  assign n17709 = n17708 ^ x98;
  assign n17710 = ~n17707 & ~n17709;
  assign n17711 = x35 & ~x99;
  assign n17712 = ~n12465 & ~n17711;
  assign n17713 = ~n17710 & n17712;
  assign n17704 = x101 & n9798;
  assign n17705 = x100 & n10099;
  assign n17706 = ~n17704 & ~n17705;
  assign n17714 = n17713 ^ n17706;
  assign n17723 = n17722 ^ n17714;
  assign n17736 = n17735 ^ n17723;
  assign n17749 = n17748 ^ n17736;
  assign n17762 = n17761 ^ n17749;
  assign n17775 = n17774 ^ n17762;
  assign n17701 = n17625 ^ n17558;
  assign n17702 = n17626 & ~n17701;
  assign n17703 = n17702 ^ n17561;
  assign n17776 = n17775 ^ n17703;
  assign n17693 = n5656 & n8169;
  assign n17694 = x117 & n5895;
  assign n17695 = x118 & n5662;
  assign n17696 = ~n17694 & ~n17695;
  assign n17697 = x119 & n6111;
  assign n17698 = n17696 & ~n17697;
  assign n17699 = ~n17693 & n17698;
  assign n17700 = n17699 ^ x47;
  assign n17777 = n17776 ^ n17700;
  assign n17690 = n17550 ^ n17542;
  assign n17691 = n17628 & ~n17690;
  assign n17692 = n17691 ^ n17627;
  assign n17778 = n17777 ^ n17692;
  assign n17787 = n17786 ^ n17778;
  assign n17687 = n17637 ^ n17539;
  assign n17688 = ~n17638 & n17687;
  assign n17689 = n17688 ^ n17539;
  assign n17788 = n17787 ^ n17689;
  assign n17797 = n17796 ^ n17788;
  assign n17684 = n17647 ^ n17536;
  assign n17685 = ~n17648 & n17684;
  assign n17686 = n17685 ^ n17536;
  assign n17798 = n17797 ^ n17686;
  assign n17678 = n3829 & ~n9889;
  assign n17679 = x126 & n4049;
  assign n17680 = x127 & n3833;
  assign n17681 = ~n17679 & ~n17680;
  assign n17682 = ~n17678 & n17681;
  assign n17683 = n17682 ^ x38;
  assign n17799 = n17798 ^ n17683;
  assign n17675 = n17657 ^ n17533;
  assign n17676 = ~n17658 & n17675;
  assign n17677 = n17676 ^ n17533;
  assign n17800 = n17799 ^ n17677;
  assign n17672 = n17670 ^ n17530;
  assign n17673 = n17660 & n17672;
  assign n17674 = n17673 ^ n17670;
  assign n17801 = n17800 ^ n17674;
  assign n17921 = n3496 & n10430;
  assign n17922 = x127 & n3816;
  assign n17923 = x38 & ~n17922;
  assign n17924 = ~n17921 & n17923;
  assign n17925 = ~x37 & ~n17924;
  assign n17926 = x127 & n3820;
  assign n17927 = ~x38 & ~n17926;
  assign n17928 = ~n17921 & n17927;
  assign n17929 = ~n17925 & ~n17928;
  assign n17911 = n4415 & ~n10174;
  assign n17912 = x124 & n4420;
  assign n17913 = x125 & n4410;
  assign n17914 = ~n17912 & ~n17913;
  assign n17915 = x126 & n4614;
  assign n17916 = n17914 & ~n17915;
  assign n17917 = ~n17911 & n17916;
  assign n17918 = n17917 ^ x41;
  assign n17901 = n5010 & n9309;
  assign n17902 = x121 & n5223;
  assign n17903 = x122 & n5014;
  assign n17904 = ~n17902 & ~n17903;
  assign n17905 = x123 & n5226;
  assign n17906 = n17904 & ~n17905;
  assign n17907 = ~n17901 & n17906;
  assign n17908 = n17907 ^ x44;
  assign n17888 = n6326 & n7643;
  assign n17889 = x115 & n6565;
  assign n17890 = x117 & n6569;
  assign n17891 = ~n17889 & ~n17890;
  assign n17892 = x116 & n6331;
  assign n17893 = n17891 & ~n17892;
  assign n17894 = ~n17888 & n17893;
  assign n17895 = n17894 ^ x50;
  assign n17879 = n6892 & n7076;
  assign n17880 = x112 & n7317;
  assign n17881 = x113 & n7080;
  assign n17882 = ~n17880 & ~n17881;
  assign n17883 = x114 & n7319;
  assign n17884 = n17882 & ~n17883;
  assign n17885 = ~n17879 & n17884;
  assign n17886 = n17885 ^ x53;
  assign n17868 = n6178 & n7830;
  assign n17869 = x109 & n7839;
  assign n17870 = x110 & n7834;
  assign n17871 = ~n17869 & ~n17870;
  assign n17872 = x111 & n8374;
  assign n17873 = n17871 & ~n17872;
  assign n17874 = ~n17868 & n17873;
  assign n17875 = n17874 ^ x56;
  assign n17865 = n17734 ^ n17723;
  assign n17866 = ~n17735 & ~n17865;
  assign n17867 = n17866 ^ n17726;
  assign n17876 = n17875 ^ n17867;
  assign n17855 = ~n5506 & n8622;
  assign n17856 = x107 & n8626;
  assign n17857 = x106 & n8631;
  assign n17858 = ~n17856 & ~n17857;
  assign n17859 = x108 & n9186;
  assign n17860 = n17858 & ~n17859;
  assign n17861 = ~n17855 & n17860;
  assign n17862 = n17861 ^ x59;
  assign n17845 = ~x102 & n17704;
  assign n17846 = ~x101 & n17705;
  assign n17847 = ~n17845 & ~n17846;
  assign n17848 = ~x101 & x102;
  assign n17849 = n9798 & n17848;
  assign n17850 = ~x100 & x101;
  assign n17851 = n10099 & n17850;
  assign n17852 = ~n17849 & ~n17851;
  assign n17853 = n17847 & n17852;
  assign n17842 = n17722 ^ n17713;
  assign n17843 = ~n17714 & ~n17842;
  assign n17844 = n17843 ^ n17722;
  assign n17854 = n17853 ^ n17844;
  assign n17863 = n17862 ^ n17854;
  assign n17834 = n4867 & n9499;
  assign n17835 = x104 & n9503;
  assign n17836 = x103 & n9508;
  assign n17837 = ~n17835 & ~n17836;
  assign n17838 = x105 & n10106;
  assign n17839 = n17837 & ~n17838;
  assign n17840 = ~n17834 & n17839;
  assign n17841 = n17840 ^ x62;
  assign n17864 = n17863 ^ n17841;
  assign n17877 = n17876 ^ n17864;
  assign n17831 = n17747 ^ n17736;
  assign n17832 = n17748 & n17831;
  assign n17833 = n17832 ^ n17739;
  assign n17878 = n17877 ^ n17833;
  assign n17887 = n17886 ^ n17878;
  assign n17896 = n17895 ^ n17887;
  assign n17828 = n17752 ^ n17749;
  assign n17829 = n17761 & n17828;
  assign n17830 = n17829 ^ n17760;
  assign n17897 = n17896 ^ n17830;
  assign n17825 = n17765 ^ n17762;
  assign n17826 = n17774 & n17825;
  assign n17827 = n17826 ^ n17773;
  assign n17898 = n17897 ^ n17827;
  assign n17817 = n5656 & ~n8424;
  assign n17818 = x118 & n5895;
  assign n17819 = x119 & n5662;
  assign n17820 = ~n17818 & ~n17819;
  assign n17821 = x120 & n6111;
  assign n17822 = n17820 & ~n17821;
  assign n17823 = ~n17817 & n17822;
  assign n17824 = n17823 ^ x47;
  assign n17899 = n17898 ^ n17824;
  assign n17814 = n17775 ^ n17700;
  assign n17815 = ~n17776 & n17814;
  assign n17816 = n17815 ^ n17703;
  assign n17900 = n17899 ^ n17816;
  assign n17909 = n17908 ^ n17900;
  assign n17811 = n17786 ^ n17692;
  assign n17812 = n17778 & n17811;
  assign n17813 = n17812 ^ n17786;
  assign n17910 = n17909 ^ n17813;
  assign n17919 = n17918 ^ n17910;
  assign n17808 = n17796 ^ n17689;
  assign n17809 = n17788 & n17808;
  assign n17810 = n17809 ^ n17796;
  assign n17920 = n17919 ^ n17810;
  assign n17930 = n17929 ^ n17920;
  assign n17805 = n17797 ^ n17683;
  assign n17806 = ~n17798 & n17805;
  assign n17807 = n17806 ^ n17686;
  assign n17931 = n17930 ^ n17807;
  assign n17802 = n17677 ^ n17674;
  assign n17803 = n17800 & ~n17802;
  assign n17804 = n17803 ^ n17674;
  assign n17932 = n17931 ^ n17804;
  assign n18045 = ~n17807 & ~n17930;
  assign n18046 = ~n17804 & ~n18045;
  assign n18047 = n17807 & n17930;
  assign n18048 = ~n18046 & ~n18047;
  assign n18029 = n6326 & n7919;
  assign n18030 = x116 & n6565;
  assign n18031 = x118 & n6569;
  assign n18032 = ~n18030 & ~n18031;
  assign n18033 = x117 & n6331;
  assign n18034 = n18032 & ~n18033;
  assign n18035 = ~n18029 & n18034;
  assign n18036 = n18035 ^ x50;
  assign n18026 = n17887 ^ n17830;
  assign n18027 = ~n17896 & n18026;
  assign n18028 = n18027 ^ n17895;
  assign n18037 = n18036 ^ n18028;
  assign n18016 = n7076 & n7150;
  assign n18017 = x113 & n7317;
  assign n18018 = x114 & n7080;
  assign n18019 = ~n18017 & ~n18018;
  assign n18020 = x115 & n7319;
  assign n18021 = n18019 & ~n18020;
  assign n18022 = ~n18016 & n18021;
  assign n18023 = n18022 ^ x53;
  assign n18013 = n17886 ^ n17833;
  assign n18014 = n17878 & n18013;
  assign n18015 = n18014 ^ n17886;
  assign n18024 = n18023 ^ n18015;
  assign n18003 = n6420 & n7830;
  assign n18004 = x110 & n7839;
  assign n18005 = x111 & n7834;
  assign n18006 = ~n18004 & ~n18005;
  assign n18007 = x112 & n8374;
  assign n18008 = n18006 & ~n18007;
  assign n18009 = ~n18003 & n18008;
  assign n18010 = n18009 ^ x56;
  assign n18000 = n17867 ^ n17864;
  assign n18001 = ~n17876 & n18000;
  assign n18002 = n18001 ^ n17875;
  assign n18011 = n18010 ^ n18002;
  assign n17990 = ~n5737 & n8622;
  assign n17991 = x107 & n8631;
  assign n17992 = x109 & n9186;
  assign n17993 = ~n17991 & ~n17992;
  assign n17994 = x108 & n8626;
  assign n17995 = n17993 & ~n17994;
  assign n17996 = ~n17990 & n17995;
  assign n17997 = n17996 ^ x59;
  assign n17987 = n17854 ^ n17841;
  assign n17988 = n17863 & ~n17987;
  assign n17989 = n17988 ^ n17862;
  assign n17998 = n17997 ^ n17989;
  assign n17977 = n5088 & n9499;
  assign n17978 = x104 & n9508;
  assign n17979 = x106 & n10106;
  assign n17980 = ~n17978 & ~n17979;
  assign n17981 = x105 & n9503;
  assign n17982 = n17980 & ~n17981;
  assign n17983 = ~n17977 & n17982;
  assign n17984 = n17983 ^ x62;
  assign n17972 = x103 & n9798;
  assign n17973 = x102 & n10099;
  assign n17974 = ~n17972 & ~n17973;
  assign n17975 = n17974 ^ n17706;
  assign n17976 = n17975 ^ x38;
  assign n17985 = n17984 ^ n17976;
  assign n17970 = n17844 & n17853;
  assign n17971 = n17970 ^ n17847;
  assign n17986 = n17985 ^ n17971;
  assign n17999 = n17998 ^ n17986;
  assign n18012 = n18011 ^ n17999;
  assign n18025 = n18024 ^ n18012;
  assign n18038 = n18037 ^ n18025;
  assign n17962 = n5656 & n8715;
  assign n17963 = x119 & n5895;
  assign n17964 = x120 & n5662;
  assign n17965 = ~n17963 & ~n17964;
  assign n17966 = x121 & n6111;
  assign n17967 = n17965 & ~n17966;
  assign n17968 = ~n17962 & n17967;
  assign n17969 = n17968 ^ x47;
  assign n18039 = n18038 ^ n17969;
  assign n17959 = n17827 ^ n17824;
  assign n17960 = ~n17898 & ~n17959;
  assign n17961 = n17960 ^ n17897;
  assign n18040 = n18039 ^ n17961;
  assign n17956 = n17908 ^ n17816;
  assign n17957 = n17900 & n17956;
  assign n17958 = n17957 ^ n17908;
  assign n18041 = n18040 ^ n17958;
  assign n17948 = n5010 & n9614;
  assign n17949 = x122 & n5223;
  assign n17950 = x123 & n5014;
  assign n17951 = ~n17949 & ~n17950;
  assign n17952 = x124 & n5226;
  assign n17953 = n17951 & ~n17952;
  assign n17954 = ~n17948 & n17953;
  assign n17955 = n17954 ^ x44;
  assign n18042 = n18041 ^ n17955;
  assign n17945 = n17929 ^ n17919;
  assign n17946 = n17920 & n17945;
  assign n17947 = n17946 ^ n17929;
  assign n18043 = n18042 ^ n17947;
  assign n17936 = n4415 & ~n10447;
  assign n17937 = x125 & n4420;
  assign n17938 = x127 & n4614;
  assign n17939 = ~n17937 & ~n17938;
  assign n17940 = x126 & n4410;
  assign n17941 = n17939 & ~n17940;
  assign n17942 = ~n17936 & n17941;
  assign n17943 = n17942 ^ x41;
  assign n17933 = n17918 ^ n17813;
  assign n17934 = n17910 & n17933;
  assign n17935 = n17934 ^ n17918;
  assign n17944 = n17943 ^ n17935;
  assign n18044 = n18043 ^ n17944;
  assign n18049 = n18048 ^ n18044;
  assign n18156 = n17935 & n17943;
  assign n18155 = ~n17935 & ~n17943;
  assign n18157 = n18156 ^ n18155;
  assign n18158 = ~n18042 & n18157;
  assign n18159 = n18158 ^ n18156;
  assign n18160 = n18043 & n18159;
  assign n18165 = ~n18042 & n18155;
  assign n18166 = ~n17947 & ~n18165;
  assign n18167 = n18042 ^ n17935;
  assign n18168 = ~n17944 & n18167;
  assign n18169 = n18168 ^ n18042;
  assign n18170 = ~n18166 & ~n18169;
  assign n18161 = n18156 ^ n18042;
  assign n18162 = ~n18043 & ~n18161;
  assign n18163 = n18162 ^ n17947;
  assign n18164 = ~n18155 & ~n18163;
  assign n18171 = n18170 ^ n18164;
  assign n18172 = ~n18048 & n18171;
  assign n18173 = n18172 ^ n18170;
  assign n18174 = ~n18160 & ~n18173;
  assign n18143 = n5010 & n9912;
  assign n18144 = x123 & n5223;
  assign n18145 = x124 & n5014;
  assign n18146 = ~n18144 & ~n18145;
  assign n18147 = x125 & n5226;
  assign n18148 = n18146 & ~n18147;
  assign n18149 = ~n18143 & n18148;
  assign n18150 = n18149 ^ x44;
  assign n18133 = n5656 & n9001;
  assign n18134 = x120 & n5895;
  assign n18135 = x122 & n6111;
  assign n18136 = ~n18134 & ~n18135;
  assign n18137 = x121 & n5662;
  assign n18138 = n18136 & ~n18137;
  assign n18139 = ~n18133 & n18138;
  assign n18140 = n18139 ^ x47;
  assign n18123 = n6326 & n8169;
  assign n18124 = x117 & n6565;
  assign n18125 = x118 & n6331;
  assign n18126 = ~n18124 & ~n18125;
  assign n18127 = x119 & n6569;
  assign n18128 = n18126 & ~n18127;
  assign n18129 = ~n18123 & n18128;
  assign n18130 = n18129 ^ x50;
  assign n18113 = n7076 & n7393;
  assign n18114 = x114 & n7317;
  assign n18115 = x115 & n7080;
  assign n18116 = ~n18114 & ~n18115;
  assign n18117 = x116 & n7319;
  assign n18118 = n18116 & ~n18117;
  assign n18119 = ~n18113 & n18118;
  assign n18120 = n18119 ^ x53;
  assign n18110 = n18010 ^ n17999;
  assign n18111 = n18011 & n18110;
  assign n18112 = n18111 ^ n18002;
  assign n18121 = n18120 ^ n18112;
  assign n18100 = n6656 & n7830;
  assign n18101 = x111 & n7839;
  assign n18102 = x113 & n8374;
  assign n18103 = ~n18101 & ~n18102;
  assign n18104 = x112 & n7834;
  assign n18105 = n18103 & ~n18104;
  assign n18106 = ~n18100 & n18105;
  assign n18107 = n18106 ^ x56;
  assign n18097 = n17997 ^ n17986;
  assign n18098 = n17998 & n18097;
  assign n18099 = n18098 ^ n17989;
  assign n18108 = n18107 ^ n18099;
  assign n18087 = n5955 & n8622;
  assign n18088 = x108 & n8631;
  assign n18089 = x109 & n8626;
  assign n18090 = ~n18088 & ~n18089;
  assign n18091 = x110 & n9186;
  assign n18092 = n18090 & ~n18091;
  assign n18093 = ~n18087 & n18092;
  assign n18094 = n18093 ^ x59;
  assign n18078 = n5297 & n9499;
  assign n18079 = x105 & n9508;
  assign n18080 = x107 & n10106;
  assign n18081 = ~n18079 & ~n18080;
  assign n18082 = x106 & n9503;
  assign n18083 = n18081 & ~n18082;
  assign n18084 = ~n18078 & n18083;
  assign n18085 = n18084 ^ x62;
  assign n18074 = x104 & n9798;
  assign n18075 = x103 & n10099;
  assign n18076 = ~n18074 & ~n18075;
  assign n18071 = n17706 ^ x38;
  assign n18072 = ~n17975 & n18071;
  assign n18073 = n18072 ^ x38;
  assign n18077 = n18076 ^ n18073;
  assign n18086 = n18085 ^ n18077;
  assign n18095 = n18094 ^ n18086;
  assign n18068 = n17984 ^ n17971;
  assign n18069 = ~n17985 & ~n18068;
  assign n18070 = n18069 ^ n17971;
  assign n18096 = n18095 ^ n18070;
  assign n18109 = n18108 ^ n18096;
  assign n18122 = n18121 ^ n18109;
  assign n18131 = n18130 ^ n18122;
  assign n18065 = n18023 ^ n18012;
  assign n18066 = n18024 & n18065;
  assign n18067 = n18066 ^ n18015;
  assign n18132 = n18131 ^ n18067;
  assign n18141 = n18140 ^ n18132;
  assign n18062 = n18036 ^ n18025;
  assign n18063 = n18037 & n18062;
  assign n18064 = n18063 ^ n18028;
  assign n18142 = n18141 ^ n18064;
  assign n18151 = n18150 ^ n18142;
  assign n18059 = n17969 ^ n17961;
  assign n18060 = ~n18039 & n18059;
  assign n18061 = n18060 ^ n18038;
  assign n18152 = n18151 ^ n18061;
  assign n18056 = n18040 ^ n17955;
  assign n18057 = n18041 & ~n18056;
  assign n18058 = n18057 ^ n17958;
  assign n18153 = n18152 ^ n18058;
  assign n18050 = n4415 & ~n9889;
  assign n18051 = x126 & n4420;
  assign n18052 = x127 & n4410;
  assign n18053 = ~n18051 & ~n18052;
  assign n18054 = ~n18050 & n18053;
  assign n18055 = n18054 ^ x41;
  assign n18154 = n18153 ^ n18055;
  assign n18175 = n18174 ^ n18154;
  assign n18278 = ~n18047 & ~n18156;
  assign n18279 = ~n18046 & n18278;
  assign n18280 = ~n18155 & ~n18279;
  assign n18281 = n17947 & ~n18042;
  assign n18282 = ~n18154 & ~n18281;
  assign n18283 = ~n18280 & ~n18282;
  assign n18284 = ~n17947 & n18042;
  assign n18285 = ~n18154 & ~n18155;
  assign n18286 = ~n18284 & ~n18285;
  assign n18287 = n18048 & n18286;
  assign n18288 = n18154 & n18163;
  assign n18289 = ~n18287 & ~n18288;
  assign n18290 = ~n18283 & n18289;
  assign n18271 = n4415 & n10430;
  assign n18272 = x127 & n4420;
  assign n18273 = ~n18271 & ~n18272;
  assign n18274 = n18273 ^ x41;
  assign n18268 = n18142 ^ n18061;
  assign n18269 = n18151 & n18268;
  assign n18270 = n18269 ^ n18150;
  assign n18275 = n18274 ^ n18270;
  assign n18259 = n5010 & ~n10174;
  assign n18260 = x125 & n5014;
  assign n18261 = x124 & n5223;
  assign n18262 = ~n18260 & ~n18261;
  assign n18263 = x126 & n5226;
  assign n18264 = n18262 & ~n18263;
  assign n18265 = ~n18259 & n18264;
  assign n18266 = n18265 ^ x44;
  assign n18246 = n6326 & ~n8424;
  assign n18247 = x118 & n6565;
  assign n18248 = x119 & n6331;
  assign n18249 = ~n18247 & ~n18248;
  assign n18250 = x120 & n6569;
  assign n18251 = n18249 & ~n18250;
  assign n18252 = ~n18246 & n18251;
  assign n18253 = n18252 ^ x50;
  assign n18243 = n18120 ^ n18109;
  assign n18244 = n18121 & ~n18243;
  assign n18245 = n18244 ^ n18112;
  assign n18254 = n18253 ^ n18245;
  assign n18233 = n7076 & n7643;
  assign n18234 = x115 & n7317;
  assign n18235 = x116 & n7080;
  assign n18236 = ~n18234 & ~n18235;
  assign n18237 = x117 & n7319;
  assign n18238 = n18236 & ~n18237;
  assign n18239 = ~n18233 & n18238;
  assign n18240 = n18239 ^ x53;
  assign n18230 = n18099 ^ n18096;
  assign n18231 = n18108 & ~n18230;
  assign n18232 = n18231 ^ n18107;
  assign n18241 = n18240 ^ n18232;
  assign n18220 = n6892 & n7830;
  assign n18221 = x112 & n7839;
  assign n18222 = x114 & n8374;
  assign n18223 = ~n18221 & ~n18222;
  assign n18224 = x113 & n7834;
  assign n18225 = n18223 & ~n18224;
  assign n18226 = ~n18220 & n18225;
  assign n18227 = n18226 ^ x56;
  assign n18217 = n18094 ^ n18070;
  assign n18218 = n18095 & ~n18217;
  assign n18219 = n18218 ^ n18070;
  assign n18228 = n18227 ^ n18219;
  assign n18208 = n6178 & n8622;
  assign n18209 = x109 & n8631;
  assign n18210 = x110 & n8626;
  assign n18211 = ~n18209 & ~n18210;
  assign n18212 = x111 & n9186;
  assign n18213 = n18211 & ~n18212;
  assign n18214 = ~n18208 & n18213;
  assign n18215 = n18214 ^ x59;
  assign n18203 = x105 & n9798;
  assign n18204 = x104 & n10099;
  assign n18205 = ~n18203 & ~n18204;
  assign n18201 = n18085 ^ n18073;
  assign n18202 = ~n18077 & ~n18201;
  assign n18206 = n18205 ^ n18202;
  assign n18193 = ~n5506 & n9499;
  assign n18194 = x106 & n9508;
  assign n18195 = x108 & n10106;
  assign n18196 = ~n18194 & ~n18195;
  assign n18197 = x107 & n9503;
  assign n18198 = n18196 & ~n18197;
  assign n18199 = ~n18193 & n18198;
  assign n18200 = n18199 ^ x62;
  assign n18207 = n18206 ^ n18200;
  assign n18216 = n18215 ^ n18207;
  assign n18229 = n18228 ^ n18216;
  assign n18242 = n18241 ^ n18229;
  assign n18255 = n18254 ^ n18242;
  assign n18190 = n18122 ^ n18067;
  assign n18191 = n18131 & ~n18190;
  assign n18192 = n18191 ^ n18130;
  assign n18256 = n18255 ^ n18192;
  assign n18182 = n5656 & n9309;
  assign n18183 = x121 & n5895;
  assign n18184 = x123 & n6111;
  assign n18185 = ~n18183 & ~n18184;
  assign n18186 = x122 & n5662;
  assign n18187 = n18185 & ~n18186;
  assign n18188 = ~n18182 & n18187;
  assign n18189 = n18188 ^ x47;
  assign n18257 = n18256 ^ n18189;
  assign n18179 = n18132 ^ n18064;
  assign n18180 = n18141 & ~n18179;
  assign n18181 = n18180 ^ n18140;
  assign n18258 = n18257 ^ n18181;
  assign n18267 = n18266 ^ n18258;
  assign n18276 = n18275 ^ n18267;
  assign n18176 = n18152 ^ n18055;
  assign n18177 = ~n18153 & n18176;
  assign n18178 = n18177 ^ n18058;
  assign n18277 = n18276 ^ n18178;
  assign n18291 = n18290 ^ n18277;
  assign n18388 = n18274 ^ n18267;
  assign n18389 = n18275 & n18388;
  assign n18390 = n18389 ^ n18270;
  assign n18391 = n18178 & n18390;
  assign n18392 = ~n18267 & n18274;
  assign n18393 = n18270 & n18392;
  assign n18394 = ~n18391 & ~n18393;
  assign n18395 = n18290 & ~n18394;
  assign n18396 = n18178 & n18393;
  assign n18397 = n18267 & ~n18274;
  assign n18398 = ~n18270 & n18397;
  assign n18399 = ~n18178 & n18398;
  assign n18400 = ~n18396 & ~n18399;
  assign n18401 = ~n18395 & n18400;
  assign n18402 = n18178 & ~n18398;
  assign n18403 = ~n18390 & ~n18402;
  assign n18404 = ~n18290 & n18403;
  assign n18405 = n18401 & ~n18404;
  assign n18378 = n5010 & ~n10447;
  assign n18379 = x125 & n5223;
  assign n18380 = x127 & n5226;
  assign n18381 = ~n18379 & ~n18380;
  assign n18382 = x126 & n5014;
  assign n18383 = n18381 & ~n18382;
  assign n18384 = ~n18378 & n18383;
  assign n18385 = n18384 ^ x44;
  assign n18368 = n5656 & n9614;
  assign n18369 = x122 & n5895;
  assign n18370 = x124 & n6111;
  assign n18371 = ~n18369 & ~n18370;
  assign n18372 = x123 & n5662;
  assign n18373 = n18371 & ~n18372;
  assign n18374 = ~n18368 & n18373;
  assign n18375 = n18374 ^ x47;
  assign n18358 = n6326 & n8715;
  assign n18359 = x120 & n6331;
  assign n18360 = x119 & n6565;
  assign n18361 = ~n18359 & ~n18360;
  assign n18362 = x121 & n6569;
  assign n18363 = n18361 & ~n18362;
  assign n18364 = ~n18358 & n18363;
  assign n18365 = n18364 ^ x50;
  assign n18355 = n18253 ^ n18242;
  assign n18356 = n18254 & n18355;
  assign n18357 = n18356 ^ n18245;
  assign n18366 = n18365 ^ n18357;
  assign n18345 = n7076 & n7919;
  assign n18346 = x116 & n7317;
  assign n18347 = x118 & n7319;
  assign n18348 = ~n18346 & ~n18347;
  assign n18349 = x117 & n7080;
  assign n18350 = n18348 & ~n18349;
  assign n18351 = ~n18345 & n18350;
  assign n18352 = n18351 ^ x53;
  assign n18342 = n18232 ^ n18229;
  assign n18343 = n18241 & n18342;
  assign n18344 = n18343 ^ n18240;
  assign n18353 = n18352 ^ n18344;
  assign n18332 = n7150 & n7830;
  assign n18333 = x113 & n7839;
  assign n18334 = x115 & n8374;
  assign n18335 = ~n18333 & ~n18334;
  assign n18336 = x114 & n7834;
  assign n18337 = n18335 & ~n18336;
  assign n18338 = ~n18332 & n18337;
  assign n18339 = n18338 ^ x56;
  assign n18322 = n6420 & n8622;
  assign n18323 = x110 & n8631;
  assign n18324 = x111 & n8626;
  assign n18325 = ~n18323 & ~n18324;
  assign n18326 = x112 & n9186;
  assign n18327 = n18325 & ~n18326;
  assign n18328 = ~n18322 & n18327;
  assign n18329 = n18328 ^ x59;
  assign n18312 = ~n5737 & n9499;
  assign n18313 = x107 & n9508;
  assign n18314 = x109 & n10106;
  assign n18315 = ~n18313 & ~n18314;
  assign n18316 = x108 & n9503;
  assign n18317 = n18315 & ~n18316;
  assign n18318 = ~n18312 & n18317;
  assign n18319 = n18318 ^ x62;
  assign n18309 = n18205 ^ n18076;
  assign n18310 = n18202 & ~n18309;
  assign n18311 = n18310 ^ n18076;
  assign n18320 = n18319 ^ n18311;
  assign n18304 = x106 & n9798;
  assign n18305 = x105 & n10099;
  assign n18306 = ~n18304 & ~n18305;
  assign n18307 = n18306 ^ n18076;
  assign n18308 = n18307 ^ x41;
  assign n18321 = n18320 ^ n18308;
  assign n18330 = n18329 ^ n18321;
  assign n18301 = n18215 ^ n18206;
  assign n18302 = ~n18207 & n18301;
  assign n18303 = n18302 ^ n18215;
  assign n18331 = n18330 ^ n18303;
  assign n18340 = n18339 ^ n18331;
  assign n18298 = n18219 ^ n18216;
  assign n18299 = ~n18228 & n18298;
  assign n18300 = n18299 ^ n18227;
  assign n18341 = n18340 ^ n18300;
  assign n18354 = n18353 ^ n18341;
  assign n18367 = n18366 ^ n18354;
  assign n18376 = n18375 ^ n18367;
  assign n18295 = n18255 ^ n18189;
  assign n18296 = ~n18256 & n18295;
  assign n18297 = n18296 ^ n18192;
  assign n18377 = n18376 ^ n18297;
  assign n18386 = n18385 ^ n18377;
  assign n18292 = n18266 ^ n18181;
  assign n18293 = n18258 & n18292;
  assign n18294 = n18293 ^ n18266;
  assign n18387 = n18386 ^ n18294;
  assign n18406 = n18405 ^ n18387;
  assign n18503 = ~n18387 & ~n18403;
  assign n18504 = ~n18396 & ~n18503;
  assign n18505 = ~n18290 & n18504;
  assign n18506 = n18387 & n18394;
  assign n18507 = ~n18399 & ~n18506;
  assign n18508 = ~n18505 & n18507;
  assign n18490 = n5656 & n9912;
  assign n18491 = x123 & n5895;
  assign n18492 = x124 & n5662;
  assign n18493 = ~n18491 & ~n18492;
  assign n18494 = x125 & n6111;
  assign n18495 = n18493 & ~n18494;
  assign n18496 = ~n18490 & n18495;
  assign n18497 = n18496 ^ x47;
  assign n18487 = n18365 ^ n18354;
  assign n18488 = n18366 & n18487;
  assign n18489 = n18488 ^ n18357;
  assign n18498 = n18497 ^ n18489;
  assign n18475 = n7076 & n8169;
  assign n18476 = x117 & n7317;
  assign n18477 = x118 & n7080;
  assign n18478 = ~n18476 & ~n18477;
  assign n18479 = x119 & n7319;
  assign n18480 = n18478 & ~n18479;
  assign n18481 = ~n18475 & n18480;
  assign n18482 = n18481 ^ x53;
  assign n18465 = n7393 & n7830;
  assign n18466 = x114 & n7839;
  assign n18467 = x115 & n7834;
  assign n18468 = ~n18466 & ~n18467;
  assign n18469 = x116 & n8374;
  assign n18470 = n18468 & ~n18469;
  assign n18471 = ~n18465 & n18470;
  assign n18472 = n18471 ^ x56;
  assign n18462 = n18329 ^ n18303;
  assign n18463 = n18330 & n18462;
  assign n18464 = n18463 ^ n18303;
  assign n18473 = n18472 ^ n18464;
  assign n18452 = n6656 & n8622;
  assign n18453 = x111 & n8631;
  assign n18454 = x112 & n8626;
  assign n18455 = ~n18453 & ~n18454;
  assign n18456 = x113 & n9186;
  assign n18457 = n18455 & ~n18456;
  assign n18458 = ~n18452 & n18457;
  assign n18459 = n18458 ^ x59;
  assign n18449 = n18319 ^ n18308;
  assign n18450 = ~n18320 & ~n18449;
  assign n18451 = n18450 ^ n18311;
  assign n18460 = n18459 ^ n18451;
  assign n18440 = n5955 & n9499;
  assign n18441 = x109 & n9503;
  assign n18442 = x108 & n9508;
  assign n18443 = ~n18441 & ~n18442;
  assign n18444 = x110 & n10106;
  assign n18445 = n18443 & ~n18444;
  assign n18446 = ~n18440 & n18445;
  assign n18447 = n18446 ^ x62;
  assign n18436 = x107 & n9798;
  assign n18437 = x106 & n10099;
  assign n18438 = ~n18436 & ~n18437;
  assign n18433 = n18076 ^ x41;
  assign n18434 = ~n18307 & n18433;
  assign n18435 = n18434 ^ x41;
  assign n18439 = n18438 ^ n18435;
  assign n18448 = n18447 ^ n18439;
  assign n18461 = n18460 ^ n18448;
  assign n18474 = n18473 ^ n18461;
  assign n18483 = n18482 ^ n18474;
  assign n18430 = n18339 ^ n18300;
  assign n18431 = n18340 & n18430;
  assign n18432 = n18431 ^ n18300;
  assign n18484 = n18483 ^ n18432;
  assign n18427 = n18352 ^ n18341;
  assign n18428 = n18353 & n18427;
  assign n18429 = n18428 ^ n18344;
  assign n18485 = n18484 ^ n18429;
  assign n18419 = n6326 & n9001;
  assign n18420 = x120 & n6565;
  assign n18421 = x121 & n6331;
  assign n18422 = ~n18420 & ~n18421;
  assign n18423 = x122 & n6569;
  assign n18424 = n18422 & ~n18423;
  assign n18425 = ~n18419 & n18424;
  assign n18426 = n18425 ^ x50;
  assign n18486 = n18485 ^ n18426;
  assign n18499 = n18498 ^ n18486;
  assign n18416 = n18375 ^ n18297;
  assign n18417 = n18376 & n18416;
  assign n18418 = n18417 ^ n18297;
  assign n18500 = n18499 ^ n18418;
  assign n18410 = n5010 & ~n9889;
  assign n18411 = x127 & n5014;
  assign n18412 = x126 & n5223;
  assign n18413 = ~n18411 & ~n18412;
  assign n18414 = ~n18410 & n18413;
  assign n18415 = n18414 ^ x44;
  assign n18501 = n18500 ^ n18415;
  assign n18407 = n18385 ^ n18294;
  assign n18408 = n18386 & n18407;
  assign n18409 = n18408 ^ n18294;
  assign n18502 = n18501 ^ n18409;
  assign n18509 = n18508 ^ n18502;
  assign n18607 = ~n18409 & ~n18501;
  assign n18608 = n18507 & ~n18607;
  assign n18609 = ~n18505 & n18608;
  assign n18610 = n18409 & n18501;
  assign n18611 = ~n18609 & ~n18610;
  assign n18595 = n4611 & n10430;
  assign n18596 = x127 & n4998;
  assign n18597 = x44 & ~n18596;
  assign n18598 = ~n18595 & n18597;
  assign n18599 = ~x43 & ~n18598;
  assign n18600 = x127 & n5001;
  assign n18601 = ~x44 & ~n18600;
  assign n18602 = ~n18595 & n18601;
  assign n18603 = ~n18599 & ~n18602;
  assign n18592 = n18489 ^ n18486;
  assign n18593 = n18498 & ~n18592;
  assign n18594 = n18593 ^ n18497;
  assign n18604 = n18603 ^ n18594;
  assign n18582 = n5656 & ~n10174;
  assign n18583 = x124 & n5895;
  assign n18584 = x126 & n6111;
  assign n18585 = ~n18583 & ~n18584;
  assign n18586 = x125 & n5662;
  assign n18587 = n18585 & ~n18586;
  assign n18588 = ~n18582 & n18587;
  assign n18589 = n18588 ^ x47;
  assign n18572 = n6326 & n9309;
  assign n18573 = x121 & n6565;
  assign n18574 = x122 & n6331;
  assign n18575 = ~n18573 & ~n18574;
  assign n18576 = x123 & n6569;
  assign n18577 = n18575 & ~n18576;
  assign n18578 = ~n18572 & n18577;
  assign n18579 = n18578 ^ x50;
  assign n18562 = n7076 & ~n8424;
  assign n18563 = x118 & n7317;
  assign n18564 = x119 & n7080;
  assign n18565 = ~n18563 & ~n18564;
  assign n18566 = x120 & n7319;
  assign n18567 = n18565 & ~n18566;
  assign n18568 = ~n18562 & n18567;
  assign n18569 = n18568 ^ x53;
  assign n18552 = n7643 & n7830;
  assign n18553 = x115 & n7839;
  assign n18554 = x116 & n7834;
  assign n18555 = ~n18553 & ~n18554;
  assign n18556 = x117 & n8374;
  assign n18557 = n18555 & ~n18556;
  assign n18558 = ~n18552 & n18557;
  assign n18559 = n18558 ^ x56;
  assign n18543 = n6892 & n8622;
  assign n18544 = x112 & n8631;
  assign n18545 = x113 & n8626;
  assign n18546 = ~n18544 & ~n18545;
  assign n18547 = x114 & n9186;
  assign n18548 = n18546 & ~n18547;
  assign n18549 = ~n18543 & n18548;
  assign n18550 = n18549 ^ x59;
  assign n18534 = n6178 & n9499;
  assign n18535 = x109 & n9508;
  assign n18536 = x111 & n10106;
  assign n18537 = ~n18535 & ~n18536;
  assign n18538 = x110 & n9503;
  assign n18539 = n18537 & ~n18538;
  assign n18540 = ~n18534 & n18539;
  assign n18528 = x107 ^ x106;
  assign n18529 = n10099 & n18528;
  assign n18530 = x108 ^ x107;
  assign n18531 = n9798 & n18530;
  assign n18532 = n18531 ^ x62;
  assign n18533 = ~n18529 & n18532;
  assign n18541 = n18540 ^ n18533;
  assign n18525 = n18447 ^ n18435;
  assign n18526 = n18439 & n18525;
  assign n18527 = n18526 ^ n18447;
  assign n18542 = n18541 ^ n18527;
  assign n18551 = n18550 ^ n18542;
  assign n18560 = n18559 ^ n18551;
  assign n18522 = n18451 ^ n18448;
  assign n18523 = ~n18460 & ~n18522;
  assign n18524 = n18523 ^ n18459;
  assign n18561 = n18560 ^ n18524;
  assign n18570 = n18569 ^ n18561;
  assign n18519 = n18464 ^ n18461;
  assign n18520 = n18473 & ~n18519;
  assign n18521 = n18520 ^ n18472;
  assign n18571 = n18570 ^ n18521;
  assign n18580 = n18579 ^ n18571;
  assign n18516 = n18474 ^ n18432;
  assign n18517 = n18483 & ~n18516;
  assign n18518 = n18517 ^ n18482;
  assign n18581 = n18580 ^ n18518;
  assign n18590 = n18589 ^ n18581;
  assign n18513 = n18484 ^ n18426;
  assign n18514 = n18485 & ~n18513;
  assign n18515 = n18514 ^ n18429;
  assign n18591 = n18590 ^ n18515;
  assign n18605 = n18604 ^ n18591;
  assign n18510 = n18499 ^ n18415;
  assign n18511 = n18500 & ~n18510;
  assign n18512 = n18511 ^ n18418;
  assign n18606 = n18605 ^ n18512;
  assign n18612 = n18611 ^ n18606;
  assign n18706 = n18591 ^ n18512;
  assign n18707 = n18594 ^ n18591;
  assign n18708 = n18706 & n18707;
  assign n18709 = n18604 & n18708;
  assign n18717 = n18706 ^ n18594;
  assign n18718 = n18717 ^ n18603;
  assign n18719 = n18718 ^ n18709;
  assign n18720 = ~n18611 & n18719;
  assign n18710 = n18512 & n18594;
  assign n18711 = n18603 ^ n18591;
  assign n18712 = ~n18512 & ~n18594;
  assign n18713 = n18712 ^ n18591;
  assign n18714 = n18711 & ~n18713;
  assign n18715 = n18714 ^ n18603;
  assign n18716 = ~n18710 & n18715;
  assign n18721 = n18720 ^ n18716;
  assign n18722 = ~n18709 & ~n18721;
  assign n18696 = n5656 & ~n10447;
  assign n18697 = x125 & n5895;
  assign n18698 = x126 & n5662;
  assign n18699 = ~n18697 & ~n18698;
  assign n18700 = x127 & n6111;
  assign n18701 = n18699 & ~n18700;
  assign n18702 = ~n18696 & n18701;
  assign n18703 = n18702 ^ x47;
  assign n18686 = n6326 & n9614;
  assign n18687 = x122 & n6565;
  assign n18688 = x123 & n6331;
  assign n18689 = ~n18687 & ~n18688;
  assign n18690 = x124 & n6569;
  assign n18691 = n18689 & ~n18690;
  assign n18692 = ~n18686 & n18691;
  assign n18693 = n18692 ^ x50;
  assign n18676 = n7076 & n8715;
  assign n18677 = x119 & n7317;
  assign n18678 = x120 & n7080;
  assign n18679 = ~n18677 & ~n18678;
  assign n18680 = x121 & n7319;
  assign n18681 = n18679 & ~n18680;
  assign n18682 = ~n18676 & n18681;
  assign n18683 = n18682 ^ x53;
  assign n18673 = n18561 ^ n18521;
  assign n18674 = ~n18570 & n18673;
  assign n18675 = n18674 ^ n18569;
  assign n18684 = n18683 ^ n18675;
  assign n18661 = n7150 & n8622;
  assign n18662 = x113 & n8631;
  assign n18663 = x114 & n8626;
  assign n18664 = ~n18662 & ~n18663;
  assign n18665 = x115 & n9186;
  assign n18666 = n18664 & ~n18665;
  assign n18667 = ~n18661 & n18666;
  assign n18668 = n18667 ^ x59;
  assign n18658 = n18550 ^ n18527;
  assign n18659 = n18542 & n18658;
  assign n18660 = n18659 ^ n18550;
  assign n18669 = n18668 ^ n18660;
  assign n18644 = ~n5072 & n18540;
  assign n18645 = ~n5070 & n13628;
  assign n18646 = ~n18644 & n18645;
  assign n18647 = x63 & n5070;
  assign n18648 = ~x62 & ~n18647;
  assign n18649 = n18540 & n18648;
  assign n18650 = ~n18646 & ~n18649;
  assign n18651 = ~n4853 & n18540;
  assign n18652 = ~n4855 & n10099;
  assign n18653 = ~n18651 & n18652;
  assign n18654 = n5072 & n14319;
  assign n18655 = ~n18653 & ~n18654;
  assign n18656 = n18650 & n18655;
  assign n18635 = n6420 & n9499;
  assign n18636 = x110 & n9508;
  assign n18637 = x112 & n10106;
  assign n18638 = ~n18636 & ~n18637;
  assign n18639 = x111 & n9503;
  assign n18640 = n18638 & ~n18639;
  assign n18641 = ~n18635 & n18640;
  assign n18642 = n18641 ^ x62;
  assign n18630 = x109 & n9798;
  assign n18631 = x108 & n10099;
  assign n18632 = ~n18630 & ~n18631;
  assign n18633 = n18632 ^ n18438;
  assign n18634 = n18633 ^ x44;
  assign n18643 = n18642 ^ n18634;
  assign n18657 = n18656 ^ n18643;
  assign n18670 = n18669 ^ n18657;
  assign n18622 = n7830 & n7919;
  assign n18623 = x116 & n7839;
  assign n18624 = x117 & n7834;
  assign n18625 = ~n18623 & ~n18624;
  assign n18626 = x118 & n8374;
  assign n18627 = n18625 & ~n18626;
  assign n18628 = ~n18622 & n18627;
  assign n18629 = n18628 ^ x56;
  assign n18671 = n18670 ^ n18629;
  assign n18619 = n18551 ^ n18524;
  assign n18620 = ~n18560 & n18619;
  assign n18621 = n18620 ^ n18559;
  assign n18672 = n18671 ^ n18621;
  assign n18685 = n18684 ^ n18672;
  assign n18694 = n18693 ^ n18685;
  assign n18616 = n18571 ^ n18518;
  assign n18617 = ~n18580 & n18616;
  assign n18618 = n18617 ^ n18579;
  assign n18695 = n18694 ^ n18618;
  assign n18704 = n18703 ^ n18695;
  assign n18613 = n18581 ^ n18515;
  assign n18614 = ~n18590 & n18613;
  assign n18615 = n18614 ^ n18589;
  assign n18705 = n18704 ^ n18615;
  assign n18723 = n18722 ^ n18705;
  assign n18807 = n18611 & ~n18710;
  assign n18808 = ~n18591 & ~n18603;
  assign n18809 = n18705 & ~n18808;
  assign n18810 = ~n18712 & ~n18809;
  assign n18811 = ~n18807 & n18810;
  assign n18812 = n18591 & n18603;
  assign n18813 = n18705 & ~n18710;
  assign n18814 = ~n18812 & ~n18813;
  assign n18815 = ~n18611 & n18814;
  assign n18816 = ~n18705 & ~n18715;
  assign n18817 = ~n18815 & ~n18816;
  assign n18818 = ~n18811 & n18817;
  assign n18798 = n5656 & ~n9889;
  assign n18799 = x126 & n5895;
  assign n18800 = x127 & n5662;
  assign n18801 = ~n18799 & ~n18800;
  assign n18802 = ~n18798 & n18801;
  assign n18803 = n18802 ^ x47;
  assign n18788 = n6326 & n9912;
  assign n18789 = x123 & n6565;
  assign n18790 = x124 & n6331;
  assign n18791 = ~n18789 & ~n18790;
  assign n18792 = x125 & n6569;
  assign n18793 = n18791 & ~n18792;
  assign n18794 = ~n18788 & n18793;
  assign n18795 = n18794 ^ x50;
  assign n18778 = n7076 & n9001;
  assign n18779 = x120 & n7317;
  assign n18780 = x121 & n7080;
  assign n18781 = ~n18779 & ~n18780;
  assign n18782 = x122 & n7319;
  assign n18783 = n18781 & ~n18782;
  assign n18784 = ~n18778 & n18783;
  assign n18785 = n18784 ^ x53;
  assign n18768 = n7830 & n8169;
  assign n18769 = x117 & n7839;
  assign n18770 = x118 & n7834;
  assign n18771 = ~n18769 & ~n18770;
  assign n18772 = x119 & n8374;
  assign n18773 = n18771 & ~n18772;
  assign n18774 = ~n18768 & n18773;
  assign n18775 = n18774 ^ x56;
  assign n18758 = n7393 & n8622;
  assign n18759 = x114 & n8631;
  assign n18760 = x116 & n9186;
  assign n18761 = ~n18759 & ~n18760;
  assign n18762 = x115 & n8626;
  assign n18763 = n18761 & ~n18762;
  assign n18764 = ~n18758 & n18763;
  assign n18765 = n18764 ^ x59;
  assign n18748 = n6656 & n9499;
  assign n18749 = x111 & n9508;
  assign n18750 = x112 & n9503;
  assign n18751 = ~n18749 & ~n18750;
  assign n18752 = x113 & n10106;
  assign n18753 = n18751 & ~n18752;
  assign n18754 = ~n18748 & n18753;
  assign n18755 = n18754 ^ x62;
  assign n18745 = n18438 ^ x44;
  assign n18746 = ~n18633 & n18745;
  assign n18747 = n18746 ^ x44;
  assign n18756 = n18755 ^ n18747;
  assign n18742 = x110 & n9798;
  assign n18743 = x109 & n10099;
  assign n18744 = ~n18742 & ~n18743;
  assign n18757 = n18756 ^ n18744;
  assign n18766 = n18765 ^ n18757;
  assign n18739 = n18656 ^ n18642;
  assign n18740 = ~n18643 & ~n18739;
  assign n18741 = n18740 ^ n18656;
  assign n18767 = n18766 ^ n18741;
  assign n18776 = n18775 ^ n18767;
  assign n18736 = n18668 ^ n18657;
  assign n18737 = n18669 & n18736;
  assign n18738 = n18737 ^ n18660;
  assign n18777 = n18776 ^ n18738;
  assign n18786 = n18785 ^ n18777;
  assign n18733 = n18670 ^ n18621;
  assign n18734 = n18671 & ~n18733;
  assign n18735 = n18734 ^ n18621;
  assign n18787 = n18786 ^ n18735;
  assign n18796 = n18795 ^ n18787;
  assign n18730 = n18683 ^ n18672;
  assign n18731 = n18684 & n18730;
  assign n18732 = n18731 ^ n18675;
  assign n18797 = n18796 ^ n18732;
  assign n18804 = n18803 ^ n18797;
  assign n18727 = n18693 ^ n18618;
  assign n18728 = n18694 & n18727;
  assign n18729 = n18728 ^ n18618;
  assign n18805 = n18804 ^ n18729;
  assign n18724 = n18703 ^ n18615;
  assign n18725 = n18704 & n18724;
  assign n18726 = n18725 ^ n18615;
  assign n18806 = n18805 ^ n18726;
  assign n18819 = n18818 ^ n18806;
  assign n18899 = ~n18797 & ~n18803;
  assign n18900 = n18726 & n18729;
  assign n18912 = n18899 & ~n18900;
  assign n18902 = ~n18726 & ~n18729;
  assign n18904 = n18797 & n18803;
  assign n18913 = n18902 & ~n18904;
  assign n18914 = ~n18912 & ~n18913;
  assign n18906 = n18797 ^ n18729;
  assign n18907 = ~n18804 & ~n18906;
  assign n18908 = n18729 ^ n18726;
  assign n18909 = n18907 & ~n18908;
  assign n18901 = n18900 ^ n18899;
  assign n18903 = n18902 ^ n18901;
  assign n18905 = n18904 ^ n18903;
  assign n18910 = n18909 ^ n18905;
  assign n18911 = ~n18818 & n18910;
  assign n18915 = n18914 ^ n18911;
  assign n18916 = n18803 ^ n18726;
  assign n18917 = n18907 & ~n18916;
  assign n18918 = n18915 & ~n18917;
  assign n18888 = n5218 & n10430;
  assign n18889 = x127 & n5658;
  assign n18890 = x47 & ~n18889;
  assign n18891 = ~n18888 & n18890;
  assign n18892 = ~x46 & ~n18891;
  assign n18893 = x127 & n5659;
  assign n18894 = ~x47 & ~n18893;
  assign n18895 = ~n18888 & n18894;
  assign n18896 = ~n18892 & ~n18895;
  assign n18878 = n6326 & ~n10174;
  assign n18879 = x124 & n6565;
  assign n18880 = x126 & n6569;
  assign n18881 = ~n18879 & ~n18880;
  assign n18882 = x125 & n6331;
  assign n18883 = n18881 & ~n18882;
  assign n18884 = ~n18878 & n18883;
  assign n18885 = n18884 ^ x50;
  assign n18868 = n7076 & n9309;
  assign n18869 = x121 & n7317;
  assign n18870 = x122 & n7080;
  assign n18871 = ~n18869 & ~n18870;
  assign n18872 = x123 & n7319;
  assign n18873 = n18871 & ~n18872;
  assign n18874 = ~n18868 & n18873;
  assign n18875 = n18874 ^ x53;
  assign n18858 = n7830 & ~n8424;
  assign n18859 = x118 & n7839;
  assign n18860 = x119 & n7834;
  assign n18861 = ~n18859 & ~n18860;
  assign n18862 = x120 & n8374;
  assign n18863 = n18861 & ~n18862;
  assign n18864 = ~n18858 & n18863;
  assign n18865 = n18864 ^ x56;
  assign n18855 = n18757 ^ n18741;
  assign n18856 = ~n18766 & ~n18855;
  assign n18857 = n18856 ^ n18765;
  assign n18866 = n18865 ^ n18857;
  assign n18845 = n7643 & n8622;
  assign n18846 = x115 & n8631;
  assign n18847 = x117 & n9186;
  assign n18848 = ~n18846 & ~n18847;
  assign n18849 = x116 & n8626;
  assign n18850 = n18848 & ~n18849;
  assign n18851 = ~n18845 & n18850;
  assign n18852 = n18851 ^ x59;
  assign n18837 = n6892 & n9499;
  assign n18838 = x112 & n9508;
  assign n18839 = x113 & n9503;
  assign n18840 = ~n18838 & ~n18839;
  assign n18841 = x114 & n10106;
  assign n18842 = n18840 & ~n18841;
  assign n18843 = ~n18837 & n18842;
  assign n18844 = n18843 ^ x62;
  assign n18853 = n18852 ^ n18844;
  assign n18832 = n5954 & n10099;
  assign n18833 = x111 ^ x110;
  assign n18834 = n9798 & n18833;
  assign n18835 = ~n18832 & ~n18834;
  assign n18829 = n18747 ^ n18744;
  assign n18830 = n18756 & n18829;
  assign n18831 = n18830 ^ n18755;
  assign n18836 = n18835 ^ n18831;
  assign n18854 = n18853 ^ n18836;
  assign n18867 = n18866 ^ n18854;
  assign n18876 = n18875 ^ n18867;
  assign n18826 = n18767 ^ n18738;
  assign n18827 = n18776 & ~n18826;
  assign n18828 = n18827 ^ n18775;
  assign n18877 = n18876 ^ n18828;
  assign n18886 = n18885 ^ n18877;
  assign n18823 = n18777 ^ n18735;
  assign n18824 = n18786 & ~n18823;
  assign n18825 = n18824 ^ n18785;
  assign n18887 = n18886 ^ n18825;
  assign n18897 = n18896 ^ n18887;
  assign n18820 = n18787 ^ n18732;
  assign n18821 = n18796 & ~n18820;
  assign n18822 = n18821 ^ n18795;
  assign n18898 = n18897 ^ n18822;
  assign n18919 = n18918 ^ n18898;
  assign n19001 = n18818 & ~n18900;
  assign n19002 = n18898 & ~n18904;
  assign n19003 = ~n18902 & ~n19002;
  assign n19004 = ~n19001 & n19003;
  assign n19005 = ~n18898 & ~n18913;
  assign n19006 = n18818 & ~n19005;
  assign n19007 = n18898 & ~n18900;
  assign n19008 = ~n18899 & ~n19007;
  assign n19009 = ~n19006 & n19008;
  assign n19010 = ~n19004 & ~n19009;
  assign n18996 = n18887 ^ n18822;
  assign n18997 = ~n18897 & ~n18996;
  assign n18998 = n18997 ^ n18896;
  assign n18993 = n18877 ^ n18825;
  assign n18994 = n18886 & ~n18993;
  assign n18995 = n18994 ^ n18885;
  assign n18999 = n18998 ^ n18995;
  assign n18984 = n6326 & ~n10447;
  assign n18985 = x125 & n6565;
  assign n18986 = x126 & n6331;
  assign n18987 = ~n18985 & ~n18986;
  assign n18988 = x127 & n6569;
  assign n18989 = n18987 & ~n18988;
  assign n18990 = ~n18984 & n18989;
  assign n18991 = n18990 ^ x50;
  assign n18974 = n7076 & n9614;
  assign n18975 = x122 & n7317;
  assign n18976 = x124 & n7319;
  assign n18977 = ~n18975 & ~n18976;
  assign n18978 = x123 & n7080;
  assign n18979 = n18977 & ~n18978;
  assign n18980 = ~n18974 & n18979;
  assign n18981 = n18980 ^ x53;
  assign n18962 = n7919 & n8622;
  assign n18963 = x116 & n8631;
  assign n18964 = x118 & n9186;
  assign n18965 = ~n18963 & ~n18964;
  assign n18966 = x117 & n8626;
  assign n18967 = n18965 & ~n18966;
  assign n18968 = ~n18962 & n18967;
  assign n18969 = n18968 ^ x59;
  assign n18959 = n18844 ^ n18836;
  assign n18960 = n18853 & ~n18959;
  assign n18961 = n18960 ^ n18852;
  assign n18970 = n18969 ^ n18961;
  assign n18947 = ~x110 & n18743;
  assign n18948 = x110 & ~x111;
  assign n18949 = n9798 & n18948;
  assign n18950 = ~n18947 & ~n18949;
  assign n18951 = n18831 & n18950;
  assign n18952 = x110 & n10099;
  assign n18953 = ~x109 & n18952;
  assign n18954 = ~x110 & x111;
  assign n18955 = n9798 & n18954;
  assign n18956 = ~n18953 & ~n18955;
  assign n18957 = ~n18951 & n18956;
  assign n18938 = n7150 & n9499;
  assign n18939 = x113 & n9508;
  assign n18940 = x114 & n9503;
  assign n18941 = ~n18939 & ~n18940;
  assign n18942 = x115 & n10106;
  assign n18943 = n18941 & ~n18942;
  assign n18944 = ~n18938 & n18943;
  assign n18945 = n18944 ^ x62;
  assign n18934 = n10099 & n18833;
  assign n18935 = n5939 & n9798;
  assign n18936 = ~n18934 & ~n18935;
  assign n18937 = n18936 ^ x47;
  assign n18946 = n18945 ^ n18937;
  assign n18958 = n18957 ^ n18946;
  assign n18971 = n18970 ^ n18958;
  assign n18926 = n7830 & n8715;
  assign n18927 = x119 & n7839;
  assign n18928 = x121 & n8374;
  assign n18929 = ~n18927 & ~n18928;
  assign n18930 = x120 & n7834;
  assign n18931 = n18929 & ~n18930;
  assign n18932 = ~n18926 & n18931;
  assign n18933 = n18932 ^ x56;
  assign n18972 = n18971 ^ n18933;
  assign n18923 = n18865 ^ n18854;
  assign n18924 = n18866 & ~n18923;
  assign n18925 = n18924 ^ n18857;
  assign n18973 = n18972 ^ n18925;
  assign n18982 = n18981 ^ n18973;
  assign n18920 = n18867 ^ n18828;
  assign n18921 = n18876 & ~n18920;
  assign n18922 = n18921 ^ n18875;
  assign n18983 = n18982 ^ n18922;
  assign n18992 = n18991 ^ n18983;
  assign n19000 = n18999 ^ n18992;
  assign n19011 = n19010 ^ n19000;
  assign n19083 = ~n18983 & ~n18991;
  assign n19084 = ~n19010 & ~n19083;
  assign n19085 = n18983 & n18991;
  assign n19086 = n19085 ^ n18995;
  assign n19087 = ~n18999 & ~n19086;
  assign n19088 = n19087 ^ n18998;
  assign n19089 = n19084 & ~n19088;
  assign n19090 = n18995 & ~n18998;
  assign n19091 = n19083 & ~n19090;
  assign n19092 = ~n18995 & n18998;
  assign n19093 = ~n19085 & n19092;
  assign n19094 = ~n19091 & ~n19093;
  assign n19095 = n19010 & ~n19094;
  assign n19096 = n18995 ^ n18991;
  assign n19097 = ~n18992 & ~n19096;
  assign n19098 = n18999 & n19097;
  assign n19099 = ~n19095 & ~n19098;
  assign n19100 = ~n19089 & n19099;
  assign n19071 = n7076 & n9912;
  assign n19072 = x123 & n7317;
  assign n19073 = x125 & n7319;
  assign n19074 = ~n19072 & ~n19073;
  assign n19075 = x124 & n7080;
  assign n19076 = n19074 & ~n19075;
  assign n19077 = ~n19071 & n19076;
  assign n19078 = n19077 ^ x53;
  assign n19068 = n18933 ^ n18925;
  assign n19069 = n18972 & ~n19068;
  assign n19070 = n19069 ^ n18971;
  assign n19079 = n19078 ^ n19070;
  assign n19058 = n7830 & n9001;
  assign n19059 = x120 & n7839;
  assign n19060 = x121 & n7834;
  assign n19061 = ~n19059 & ~n19060;
  assign n19062 = x122 & n8374;
  assign n19063 = n19061 & ~n19062;
  assign n19064 = ~n19058 & n19063;
  assign n19065 = n19064 ^ x56;
  assign n19055 = n18969 ^ n18958;
  assign n19056 = n18970 & ~n19055;
  assign n19057 = n19056 ^ n18961;
  assign n19066 = n19065 ^ n19057;
  assign n19045 = n8169 & n8622;
  assign n19046 = x118 & n8626;
  assign n19047 = x117 & n8631;
  assign n19048 = ~n19046 & ~n19047;
  assign n19049 = x119 & n9186;
  assign n19050 = n19048 & ~n19049;
  assign n19051 = ~n19045 & n19050;
  assign n19052 = n19051 ^ x59;
  assign n19036 = n7393 & n9499;
  assign n19037 = x114 & n9508;
  assign n19038 = x115 & n9503;
  assign n19039 = ~n19037 & ~n19038;
  assign n19040 = x116 & n10106;
  assign n19041 = n19039 & ~n19040;
  assign n19042 = ~n19036 & n19041;
  assign n19043 = n19042 ^ x62;
  assign n19027 = ~x47 & x111;
  assign n19028 = x112 ^ x110;
  assign n19029 = ~n10099 & n19028;
  assign n19030 = n19029 ^ x110;
  assign n19031 = ~n19027 & ~n19030;
  assign n19032 = x47 & ~x111;
  assign n19033 = ~n12465 & ~n19032;
  assign n19034 = ~n19031 & n19033;
  assign n19024 = x113 & n9798;
  assign n19025 = x112 & n10099;
  assign n19026 = ~n19024 & ~n19025;
  assign n19035 = n19034 ^ n19026;
  assign n19044 = n19043 ^ n19035;
  assign n19053 = n19052 ^ n19044;
  assign n19021 = n18957 ^ n18945;
  assign n19022 = n18946 & ~n19021;
  assign n19023 = n19022 ^ n18957;
  assign n19054 = n19053 ^ n19023;
  assign n19067 = n19066 ^ n19054;
  assign n19080 = n19079 ^ n19067;
  assign n19018 = n18981 ^ n18922;
  assign n19019 = ~n18982 & n19018;
  assign n19020 = n19019 ^ n18922;
  assign n19081 = n19080 ^ n19020;
  assign n19012 = n6326 & ~n9889;
  assign n19013 = x127 & n6331;
  assign n19014 = x126 & n6565;
  assign n19015 = ~n19013 & ~n19014;
  assign n19016 = ~n19012 & n19015;
  assign n19017 = n19016 ^ x50;
  assign n19082 = n19081 ^ n19017;
  assign n19101 = n19100 ^ n19082;
  assign n19172 = ~n19082 & ~n19092;
  assign n19173 = ~n19085 & ~n19172;
  assign n19174 = ~n19084 & n19173;
  assign n19175 = ~n19082 & ~n19083;
  assign n19176 = ~n19090 & ~n19175;
  assign n19177 = n19010 & n19176;
  assign n19178 = n19082 & n19088;
  assign n19179 = ~n19177 & ~n19178;
  assign n19180 = ~n19174 & n19179;
  assign n19160 = n7076 & ~n10174;
  assign n19161 = x124 & n7317;
  assign n19162 = x125 & n7080;
  assign n19163 = ~n19161 & ~n19162;
  assign n19164 = x126 & n7319;
  assign n19165 = n19163 & ~n19164;
  assign n19166 = ~n19160 & n19165;
  assign n19167 = n19166 ^ x53;
  assign n19157 = n19065 ^ n19054;
  assign n19158 = n19066 & n19157;
  assign n19159 = n19158 ^ n19057;
  assign n19168 = n19167 ^ n19159;
  assign n19147 = n7830 & n9309;
  assign n19148 = x121 & n7839;
  assign n19149 = x123 & n8374;
  assign n19150 = ~n19148 & ~n19149;
  assign n19151 = x122 & n7834;
  assign n19152 = n19150 & ~n19151;
  assign n19153 = ~n19147 & n19152;
  assign n19154 = n19153 ^ x56;
  assign n19138 = ~n8424 & n8622;
  assign n19139 = x118 & n8631;
  assign n19140 = x119 & n8626;
  assign n19141 = ~n19139 & ~n19140;
  assign n19142 = x120 & n9186;
  assign n19143 = n19141 & ~n19142;
  assign n19144 = ~n19138 & n19143;
  assign n19145 = n19144 ^ x59;
  assign n19129 = n7643 & n9499;
  assign n19130 = x115 & n9508;
  assign n19131 = x117 & n10106;
  assign n19132 = ~n19130 & ~n19131;
  assign n19133 = x116 & n9503;
  assign n19134 = n19132 & ~n19133;
  assign n19135 = ~n19129 & n19134;
  assign n19124 = x113 ^ x112;
  assign n19125 = n10099 & n19124;
  assign n19126 = n6409 & n9798;
  assign n19127 = n19126 ^ x62;
  assign n19128 = ~n19125 & n19127;
  assign n19136 = n19135 ^ n19128;
  assign n19121 = n19043 ^ n19034;
  assign n19122 = ~n19035 & ~n19121;
  assign n19123 = n19122 ^ n19043;
  assign n19137 = n19136 ^ n19123;
  assign n19146 = n19145 ^ n19137;
  assign n19155 = n19154 ^ n19146;
  assign n19118 = n19052 ^ n19023;
  assign n19119 = ~n19053 & ~n19118;
  assign n19120 = n19119 ^ n19023;
  assign n19156 = n19155 ^ n19120;
  assign n19169 = n19168 ^ n19156;
  assign n19115 = n19080 ^ n19017;
  assign n19116 = ~n19081 & n19115;
  assign n19117 = n19116 ^ n19020;
  assign n19170 = n19169 ^ n19117;
  assign n19105 = n5900 & n10430;
  assign n19106 = x127 & n6322;
  assign n19107 = x50 & ~n19106;
  assign n19108 = ~n19105 & n19107;
  assign n19109 = ~x49 & ~n19108;
  assign n19110 = x127 & n6328;
  assign n19111 = ~x50 & ~n19110;
  assign n19112 = ~n19105 & n19111;
  assign n19113 = ~n19109 & ~n19112;
  assign n19102 = n19070 ^ n19067;
  assign n19103 = n19079 & n19102;
  assign n19104 = n19103 ^ n19078;
  assign n19114 = n19113 ^ n19104;
  assign n19171 = n19170 ^ n19114;
  assign n19181 = n19180 ^ n19171;
  assign n19253 = n19104 & ~n19113;
  assign n19254 = ~n19180 & ~n19253;
  assign n19255 = ~n19104 & n19113;
  assign n19256 = n19255 ^ n19169;
  assign n19257 = n19170 & n19256;
  assign n19258 = n19257 ^ n19117;
  assign n19259 = n19254 & ~n19258;
  assign n19260 = ~n19117 & ~n19169;
  assign n19261 = n19253 & ~n19260;
  assign n19262 = n19117 & n19169;
  assign n19263 = ~n19255 & n19262;
  assign n19264 = ~n19261 & ~n19263;
  assign n19265 = n19180 & ~n19264;
  assign n19266 = n19117 ^ n19113;
  assign n19267 = n19114 & n19266;
  assign n19268 = ~n19170 & n19267;
  assign n19269 = ~n19265 & ~n19268;
  assign n19270 = ~n19259 & n19269;
  assign n19243 = n7076 & ~n10447;
  assign n19244 = x125 & n7317;
  assign n19245 = x126 & n7080;
  assign n19246 = ~n19244 & ~n19245;
  assign n19247 = x127 & n7319;
  assign n19248 = n19246 & ~n19247;
  assign n19249 = ~n19243 & n19248;
  assign n19250 = n19249 ^ x53;
  assign n19233 = n7830 & n9614;
  assign n19234 = x122 & n7839;
  assign n19235 = x123 & n7834;
  assign n19236 = ~n19234 & ~n19235;
  assign n19237 = x124 & n8374;
  assign n19238 = n19236 & ~n19237;
  assign n19239 = ~n19233 & n19238;
  assign n19240 = n19239 ^ x56;
  assign n19223 = n8622 & n8715;
  assign n19224 = x120 & n8626;
  assign n19225 = x119 & n8631;
  assign n19226 = ~n19224 & ~n19225;
  assign n19227 = x121 & n9186;
  assign n19228 = n19226 & ~n19227;
  assign n19229 = ~n19223 & n19228;
  assign n19230 = n19229 ^ x59;
  assign n19220 = n19145 ^ n19123;
  assign n19221 = n19137 & n19220;
  assign n19222 = n19221 ^ n19145;
  assign n19231 = n19230 ^ n19222;
  assign n19202 = x113 & ~x114;
  assign n19203 = n19135 & ~n19202;
  assign n19204 = ~x113 & x114;
  assign n19205 = n13628 & ~n19204;
  assign n19206 = ~n19203 & n19205;
  assign n19207 = x63 & n19204;
  assign n19208 = ~x62 & ~n19207;
  assign n19209 = n19135 & n19208;
  assign n19210 = ~n19206 & ~n19209;
  assign n19211 = x112 & ~x113;
  assign n19212 = n19135 & ~n19211;
  assign n19213 = ~x112 & x113;
  assign n19214 = n10099 & ~n19213;
  assign n19215 = ~n19212 & n19214;
  assign n19216 = n14319 & n19202;
  assign n19217 = ~n19215 & ~n19216;
  assign n19218 = n19210 & n19217;
  assign n19193 = n7919 & n9499;
  assign n19194 = x116 & n9508;
  assign n19195 = x118 & n10106;
  assign n19196 = ~n19194 & ~n19195;
  assign n19197 = x117 & n9503;
  assign n19198 = n19196 & ~n19197;
  assign n19199 = ~n19193 & n19198;
  assign n19200 = n19199 ^ x62;
  assign n19188 = x115 & n9798;
  assign n19189 = x114 & n10099;
  assign n19190 = ~n19188 & ~n19189;
  assign n19191 = n19190 ^ x50;
  assign n19192 = n19191 ^ n19026;
  assign n19201 = n19200 ^ n19192;
  assign n19219 = n19218 ^ n19201;
  assign n19232 = n19231 ^ n19219;
  assign n19241 = n19240 ^ n19232;
  assign n19185 = n19146 ^ n19120;
  assign n19186 = ~n19155 & ~n19185;
  assign n19187 = n19186 ^ n19154;
  assign n19242 = n19241 ^ n19187;
  assign n19251 = n19250 ^ n19242;
  assign n19182 = n19159 ^ n19156;
  assign n19183 = n19168 & ~n19182;
  assign n19184 = n19183 ^ n19167;
  assign n19252 = n19251 ^ n19184;
  assign n19271 = n19270 ^ n19252;
  assign n19330 = n19252 & ~n19262;
  assign n19331 = ~n19255 & ~n19330;
  assign n19332 = ~n19254 & n19331;
  assign n19333 = n19252 & ~n19253;
  assign n19334 = ~n19260 & ~n19333;
  assign n19335 = n19180 & n19334;
  assign n19336 = ~n19252 & n19258;
  assign n19337 = ~n19335 & ~n19336;
  assign n19338 = ~n19332 & n19337;
  assign n19317 = n7830 & n9912;
  assign n19318 = x123 & n7839;
  assign n19319 = x124 & n7834;
  assign n19320 = ~n19318 & ~n19319;
  assign n19321 = x125 & n8374;
  assign n19322 = n19320 & ~n19321;
  assign n19323 = ~n19317 & n19322;
  assign n19324 = n19323 ^ x56;
  assign n19314 = n19230 ^ n19219;
  assign n19315 = n19231 & n19314;
  assign n19316 = n19315 ^ n19222;
  assign n19325 = n19324 ^ n19316;
  assign n19304 = n8622 & n9001;
  assign n19305 = x120 & n8631;
  assign n19306 = x121 & n8626;
  assign n19307 = ~n19305 & ~n19306;
  assign n19308 = x122 & n9186;
  assign n19309 = n19307 & ~n19308;
  assign n19310 = ~n19304 & n19309;
  assign n19311 = n19310 ^ x59;
  assign n19294 = n8169 & n9499;
  assign n19295 = x117 & n9508;
  assign n19296 = x118 & n9503;
  assign n19297 = ~n19295 & ~n19296;
  assign n19298 = x119 & n10106;
  assign n19299 = n19297 & ~n19298;
  assign n19300 = ~n19294 & n19299;
  assign n19301 = n19300 ^ x62;
  assign n19290 = n19026 ^ x50;
  assign n19291 = n19190 ^ n19026;
  assign n19292 = n19290 & ~n19291;
  assign n19293 = n19292 ^ x50;
  assign n19302 = n19301 ^ n19293;
  assign n19287 = x115 & n10099;
  assign n19288 = x116 & n9798;
  assign n19289 = ~n19287 & ~n19288;
  assign n19303 = n19302 ^ n19289;
  assign n19312 = n19311 ^ n19303;
  assign n19284 = n19218 ^ n19200;
  assign n19285 = ~n19201 & ~n19284;
  assign n19286 = n19285 ^ n19218;
  assign n19313 = n19312 ^ n19286;
  assign n19326 = n19325 ^ n19313;
  assign n19281 = n19240 ^ n19187;
  assign n19282 = n19241 & n19281;
  assign n19283 = n19282 ^ n19187;
  assign n19327 = n19326 ^ n19283;
  assign n19275 = n7076 & ~n9889;
  assign n19276 = x127 & n7080;
  assign n19277 = x126 & n7317;
  assign n19278 = ~n19276 & ~n19277;
  assign n19279 = ~n19275 & n19278;
  assign n19280 = n19279 ^ x53;
  assign n19328 = n19327 ^ n19280;
  assign n19272 = n19250 ^ n19184;
  assign n19273 = n19251 & n19272;
  assign n19274 = n19273 ^ n19184;
  assign n19329 = n19328 ^ n19274;
  assign n19339 = n19338 ^ n19329;
  assign n19403 = ~n19274 & ~n19328;
  assign n19404 = ~n19338 & ~n19403;
  assign n19405 = n19274 & n19328;
  assign n19406 = ~n19404 & ~n19405;
  assign n19391 = n6561 & n10430;
  assign n19392 = x127 & n7066;
  assign n19393 = x53 & ~n19392;
  assign n19394 = ~n19391 & n19393;
  assign n19395 = ~x52 & ~n19394;
  assign n19396 = x127 & n7070;
  assign n19397 = ~x53 & ~n19396;
  assign n19398 = ~n19391 & n19397;
  assign n19399 = ~n19395 & ~n19398;
  assign n19382 = n7830 & ~n10174;
  assign n19383 = x124 & n7839;
  assign n19384 = x126 & n8374;
  assign n19385 = ~n19383 & ~n19384;
  assign n19386 = x125 & n7834;
  assign n19387 = n19385 & ~n19386;
  assign n19388 = ~n19382 & n19387;
  assign n19389 = n19388 ^ x56;
  assign n19371 = n8622 & n9309;
  assign n19372 = x121 & n8631;
  assign n19373 = x122 & n8626;
  assign n19374 = ~n19372 & ~n19373;
  assign n19375 = x123 & n9186;
  assign n19376 = n19374 & ~n19375;
  assign n19377 = ~n19371 & n19376;
  assign n19378 = n19377 ^ x59;
  assign n19363 = ~n8424 & n9499;
  assign n19364 = x118 & n9508;
  assign n19365 = x119 & n9503;
  assign n19366 = ~n19364 & ~n19365;
  assign n19367 = x120 & n10106;
  assign n19368 = n19366 & ~n19367;
  assign n19369 = ~n19363 & n19368;
  assign n19370 = n19369 ^ x62;
  assign n19379 = n19378 ^ n19370;
  assign n19352 = ~x116 & n19287;
  assign n19353 = x116 & ~x117;
  assign n19354 = n9798 & n19353;
  assign n19355 = ~n19352 & ~n19354;
  assign n19356 = x116 & n10099;
  assign n19357 = ~x115 & n19356;
  assign n19358 = ~x116 & x117;
  assign n19359 = n9798 & n19358;
  assign n19360 = ~n19357 & ~n19359;
  assign n19361 = n19355 & n19360;
  assign n19349 = n19293 ^ n19289;
  assign n19350 = n19302 & n19349;
  assign n19351 = n19350 ^ n19301;
  assign n19362 = n19361 ^ n19351;
  assign n19380 = n19379 ^ n19362;
  assign n19346 = n19303 ^ n19286;
  assign n19347 = ~n19312 & ~n19346;
  assign n19348 = n19347 ^ n19311;
  assign n19381 = n19380 ^ n19348;
  assign n19390 = n19389 ^ n19381;
  assign n19400 = n19399 ^ n19390;
  assign n19343 = n19316 ^ n19313;
  assign n19344 = n19325 & ~n19343;
  assign n19345 = n19344 ^ n19324;
  assign n19401 = n19400 ^ n19345;
  assign n19340 = n19326 ^ n19280;
  assign n19341 = n19327 & ~n19340;
  assign n19342 = n19341 ^ n19283;
  assign n19402 = n19401 ^ n19342;
  assign n19407 = n19406 ^ n19402;
  assign n19455 = n19342 & ~n19401;
  assign n19456 = ~n19405 & ~n19455;
  assign n19457 = ~n19404 & n19456;
  assign n19458 = ~n19342 & n19401;
  assign n19459 = ~n19457 & ~n19458;
  assign n19450 = n19390 ^ n19345;
  assign n19451 = ~n19400 & ~n19450;
  assign n19452 = n19451 ^ n19399;
  assign n19447 = n19389 ^ n19348;
  assign n19448 = ~n19381 & n19447;
  assign n19449 = n19448 ^ n19389;
  assign n19453 = n19452 ^ n19449;
  assign n19436 = n8622 & n9614;
  assign n19437 = x122 & n8631;
  assign n19438 = x123 & n8626;
  assign n19439 = ~n19437 & ~n19438;
  assign n19440 = x124 & n9186;
  assign n19441 = n19439 & ~n19440;
  assign n19442 = ~n19436 & n19441;
  assign n19443 = n19442 ^ x59;
  assign n19433 = n19370 ^ n19362;
  assign n19434 = n19379 & ~n19433;
  assign n19435 = n19434 ^ n19378;
  assign n19444 = n19443 ^ n19435;
  assign n19423 = n8715 & n9499;
  assign n19424 = x119 & n9508;
  assign n19425 = x120 & n9503;
  assign n19426 = ~n19424 & ~n19425;
  assign n19427 = x121 & n10106;
  assign n19428 = n19426 & ~n19427;
  assign n19429 = ~n19423 & n19428;
  assign n19430 = n19429 ^ x62;
  assign n19418 = x117 ^ x116;
  assign n19419 = n10099 & n19418;
  assign n19420 = n7378 & n9798;
  assign n19421 = ~n19419 & ~n19420;
  assign n19422 = n19421 ^ x53;
  assign n19431 = n19430 ^ n19422;
  assign n19416 = n19351 & n19361;
  assign n19417 = n19416 ^ n19360;
  assign n19432 = n19431 ^ n19417;
  assign n19445 = n19444 ^ n19432;
  assign n19408 = n7830 & ~n10447;
  assign n19409 = x125 & n7839;
  assign n19410 = x127 & n8374;
  assign n19411 = ~n19409 & ~n19410;
  assign n19412 = x126 & n7834;
  assign n19413 = n19411 & ~n19412;
  assign n19414 = ~n19408 & n19413;
  assign n19415 = n19414 ^ x56;
  assign n19446 = n19445 ^ n19415;
  assign n19454 = n19453 ^ n19446;
  assign n19460 = n19459 ^ n19454;
  assign n19506 = ~n19415 & ~n19445;
  assign n19507 = n19459 & ~n19506;
  assign n19508 = ~n19449 & n19452;
  assign n19509 = n19415 & n19445;
  assign n19510 = ~n19508 & n19509;
  assign n19511 = n19449 & ~n19452;
  assign n19512 = ~n19510 & ~n19511;
  assign n19513 = n19507 & ~n19512;
  assign n19514 = n19506 & ~n19511;
  assign n19515 = ~n19508 & ~n19514;
  assign n19516 = ~n19509 & ~n19515;
  assign n19517 = ~n19459 & n19516;
  assign n19518 = ~n19510 & ~n19514;
  assign n19519 = n19453 & ~n19518;
  assign n19520 = ~n19517 & ~n19519;
  assign n19521 = ~n19513 & n19520;
  assign n19494 = n8622 & n9912;
  assign n19495 = x123 & n8631;
  assign n19496 = x125 & n9186;
  assign n19497 = ~n19495 & ~n19496;
  assign n19498 = x124 & n8626;
  assign n19499 = n19497 & ~n19498;
  assign n19500 = ~n19494 & n19499;
  assign n19501 = n19500 ^ x59;
  assign n19491 = n19430 ^ n19417;
  assign n19492 = n19431 & ~n19491;
  assign n19493 = n19492 ^ n19417;
  assign n19502 = n19501 ^ n19493;
  assign n19482 = n9001 & n9499;
  assign n19483 = x120 & n9508;
  assign n19484 = x121 & n9503;
  assign n19485 = ~n19483 & ~n19484;
  assign n19486 = x122 & n10106;
  assign n19487 = n19485 & ~n19486;
  assign n19488 = ~n19482 & n19487;
  assign n19489 = n19488 ^ x62;
  assign n19473 = ~x53 & x117;
  assign n19474 = x118 ^ x116;
  assign n19475 = ~n10099 & n19474;
  assign n19476 = n19475 ^ x116;
  assign n19477 = ~n19473 & ~n19476;
  assign n19478 = x53 & ~x117;
  assign n19479 = ~n12465 & ~n19478;
  assign n19480 = ~n19477 & n19479;
  assign n19470 = x119 & n9798;
  assign n19471 = x118 & n10099;
  assign n19472 = ~n19470 & ~n19471;
  assign n19481 = n19480 ^ n19472;
  assign n19490 = n19489 ^ n19481;
  assign n19503 = n19502 ^ n19490;
  assign n19467 = n19443 ^ n19432;
  assign n19468 = n19444 & ~n19467;
  assign n19469 = n19468 ^ n19435;
  assign n19504 = n19503 ^ n19469;
  assign n19461 = n7830 & ~n9889;
  assign n19462 = x126 & n7839;
  assign n19463 = x127 & n7834;
  assign n19464 = ~n19462 & ~n19463;
  assign n19465 = ~n19461 & n19464;
  assign n19466 = n19465 ^ x56;
  assign n19505 = n19504 ^ n19466;
  assign n19522 = n19521 ^ n19505;
  assign n19565 = ~n19505 & ~n19508;
  assign n19566 = ~n19509 & ~n19565;
  assign n19567 = ~n19507 & n19566;
  assign n19568 = ~n19505 & ~n19506;
  assign n19569 = ~n19511 & ~n19568;
  assign n19570 = ~n19459 & n19569;
  assign n19571 = n19505 & n19512;
  assign n19572 = ~n19570 & ~n19571;
  assign n19573 = ~n19567 & n19572;
  assign n19554 = n8622 & ~n10174;
  assign n19555 = x124 & n8631;
  assign n19556 = x125 & n8626;
  assign n19557 = ~n19555 & ~n19556;
  assign n19558 = x126 & n9186;
  assign n19559 = n19557 & ~n19558;
  assign n19560 = ~n19554 & n19559;
  assign n19561 = n19560 ^ x59;
  assign n19544 = n9309 & n9499;
  assign n19545 = x121 & n9508;
  assign n19546 = x123 & n10106;
  assign n19547 = ~n19545 & ~n19546;
  assign n19548 = x122 & n9503;
  assign n19549 = n19547 & ~n19548;
  assign n19550 = ~n19544 & n19549;
  assign n19551 = n19550 ^ x62;
  assign n19537 = ~x120 & n19470;
  assign n19538 = n7627 & n10099;
  assign n19539 = ~n19537 & ~n19538;
  assign n19540 = n7625 & n10099;
  assign n19541 = n7900 & n9798;
  assign n19542 = ~n19540 & ~n19541;
  assign n19543 = n19539 & n19542;
  assign n19552 = n19551 ^ n19543;
  assign n19534 = n19489 ^ n19480;
  assign n19535 = ~n19481 & ~n19534;
  assign n19536 = n19535 ^ n19489;
  assign n19553 = n19552 ^ n19536;
  assign n19562 = n19561 ^ n19553;
  assign n19531 = n19503 ^ n19466;
  assign n19532 = ~n19504 & n19531;
  assign n19533 = n19532 ^ n19469;
  assign n19563 = n19562 ^ n19533;
  assign n19526 = n7830 & n10430;
  assign n19527 = x127 & n7839;
  assign n19528 = ~n19526 & ~n19527;
  assign n19529 = n19528 ^ x56;
  assign n19523 = n19501 ^ n19490;
  assign n19524 = ~n19502 & ~n19523;
  assign n19525 = n19524 ^ n19493;
  assign n19530 = n19529 ^ n19525;
  assign n19564 = n19563 ^ n19530;
  assign n19574 = n19573 ^ n19564;
  assign n19605 = n19525 & ~n19529;
  assign n19606 = n19573 & ~n19605;
  assign n19607 = ~n19525 & n19529;
  assign n19608 = n19607 ^ n19562;
  assign n19609 = n19563 & ~n19608;
  assign n19610 = n19609 ^ n19533;
  assign n19611 = n19606 & n19610;
  assign n19612 = n19562 ^ n19529;
  assign n19613 = n19530 & n19612;
  assign n19614 = n19613 ^ n19562;
  assign n19615 = ~n19533 & ~n19614;
  assign n19616 = ~n19562 & n19605;
  assign n19617 = ~n19615 & ~n19616;
  assign n19618 = ~n19573 & ~n19617;
  assign n19619 = n19607 ^ n19605;
  assign n19620 = n19562 & n19619;
  assign n19621 = n19620 ^ n19605;
  assign n19622 = ~n19563 & n19621;
  assign n19623 = ~n19618 & ~n19622;
  assign n19624 = ~n19611 & n19623;
  assign n19595 = n8622 & ~n10447;
  assign n19596 = x125 & n8631;
  assign n19597 = x127 & n9186;
  assign n19598 = ~n19596 & ~n19597;
  assign n19599 = x126 & n8626;
  assign n19600 = n19598 & ~n19599;
  assign n19601 = ~n19595 & n19600;
  assign n19602 = n19601 ^ x59;
  assign n19592 = n19561 ^ n19536;
  assign n19593 = ~n19553 & n19592;
  assign n19594 = n19593 ^ n19561;
  assign n19603 = n19602 ^ n19594;
  assign n19582 = n9499 & n9614;
  assign n19583 = x122 & n9508;
  assign n19584 = x123 & n9503;
  assign n19585 = ~n19583 & ~n19584;
  assign n19586 = x124 & n10106;
  assign n19587 = n19585 & ~n19586;
  assign n19588 = ~n19582 & n19587;
  assign n19589 = n19588 ^ x62;
  assign n19577 = x121 & n9798;
  assign n19578 = x120 & n10099;
  assign n19579 = ~n19577 & ~n19578;
  assign n19580 = n19579 ^ x56;
  assign n19581 = n19580 ^ n19472;
  assign n19590 = n19589 ^ n19581;
  assign n19575 = n19543 & ~n19551;
  assign n19576 = n19575 ^ n19542;
  assign n19591 = n19590 ^ n19576;
  assign n19604 = n19603 ^ n19591;
  assign n19625 = n19624 ^ n19604;
  assign n19658 = ~n19533 & ~n19562;
  assign n19659 = n19604 & ~n19658;
  assign n19660 = ~n19607 & ~n19659;
  assign n19661 = ~n19606 & n19660;
  assign n19662 = n19533 & n19562;
  assign n19663 = n19604 & ~n19605;
  assign n19664 = ~n19662 & ~n19663;
  assign n19665 = ~n19573 & n19664;
  assign n19666 = ~n19604 & ~n19610;
  assign n19667 = ~n19665 & ~n19666;
  assign n19668 = ~n19661 & n19667;
  assign n19650 = n8622 & ~n9889;
  assign n19651 = x127 & n8626;
  assign n19652 = x126 & n8631;
  assign n19653 = ~n19651 & ~n19652;
  assign n19654 = ~n19650 & n19653;
  assign n19655 = n19654 ^ x59;
  assign n19639 = n9499 & n9912;
  assign n19640 = x123 & n9508;
  assign n19641 = x124 & n9503;
  assign n19642 = ~n19640 & ~n19641;
  assign n19643 = x125 & n10106;
  assign n19644 = n19642 & ~n19643;
  assign n19645 = ~n19639 & n19644;
  assign n19646 = n19645 ^ x62;
  assign n19635 = n19472 ^ x56;
  assign n19636 = n19579 ^ n19472;
  assign n19637 = n19635 & ~n19636;
  assign n19638 = n19637 ^ x56;
  assign n19647 = n19646 ^ n19638;
  assign n19632 = x122 & n9798;
  assign n19633 = x121 & n10099;
  assign n19634 = ~n19632 & ~n19633;
  assign n19648 = n19647 ^ n19634;
  assign n19629 = n19589 ^ n19576;
  assign n19630 = ~n19590 & n19629;
  assign n19631 = n19630 ^ n19576;
  assign n19649 = n19648 ^ n19631;
  assign n19656 = n19655 ^ n19649;
  assign n19626 = n19602 ^ n19591;
  assign n19627 = n19603 & ~n19626;
  assign n19628 = n19627 ^ n19594;
  assign n19657 = n19656 ^ n19628;
  assign n19669 = n19668 ^ n19657;
  assign n19699 = n8622 & n10430;
  assign n19700 = x127 & n8631;
  assign n19701 = ~n19699 & ~n19700;
  assign n19702 = n19701 ^ x59;
  assign n19696 = n19655 ^ n19631;
  assign n19697 = n19649 & n19696;
  assign n19698 = n19697 ^ n19655;
  assign n19703 = n19702 ^ n19698;
  assign n19684 = ~x122 & n19633;
  assign n19685 = x122 & ~x123;
  assign n19686 = n9798 & n19685;
  assign n19687 = ~n19684 & ~n19686;
  assign n19688 = x122 & n10099;
  assign n19689 = ~x121 & n19688;
  assign n19690 = ~x122 & x123;
  assign n19691 = n9798 & n19690;
  assign n19692 = ~n19689 & ~n19691;
  assign n19693 = n19687 & n19692;
  assign n19681 = n19638 ^ n19634;
  assign n19682 = n19647 & n19681;
  assign n19683 = n19682 ^ n19646;
  assign n19694 = n19693 ^ n19683;
  assign n19673 = n9499 & ~n10174;
  assign n19674 = x124 & n9508;
  assign n19675 = x125 & n9503;
  assign n19676 = ~n19674 & ~n19675;
  assign n19677 = x126 & n10106;
  assign n19678 = n19676 & ~n19677;
  assign n19679 = ~n19673 & n19678;
  assign n19680 = n19679 ^ x62;
  assign n19695 = n19694 ^ n19680;
  assign n19704 = n19703 ^ n19695;
  assign n19670 = n19668 ^ n19628;
  assign n19671 = n19657 & n19670;
  assign n19672 = n19671 ^ n19668;
  assign n19705 = n19704 ^ n19672;
  assign n19723 = n19698 & n19702;
  assign n19724 = ~n19680 & ~n19694;
  assign n19725 = n19723 & ~n19724;
  assign n19726 = ~n19698 & ~n19702;
  assign n19727 = n19680 & n19694;
  assign n19728 = n19726 & ~n19727;
  assign n19729 = ~n19725 & ~n19728;
  assign n19730 = ~n19695 & ~n19729;
  assign n19733 = ~n19726 & n19727;
  assign n19734 = ~n19725 & ~n19733;
  assign n19731 = ~n19723 & n19724;
  assign n19732 = ~n19728 & ~n19731;
  assign n19735 = n19734 ^ n19732;
  assign n19736 = ~n19672 & n19735;
  assign n19737 = n19736 ^ n19734;
  assign n19738 = ~n19730 & n19737;
  assign n19713 = n9499 & ~n10447;
  assign n19714 = x125 & n9508;
  assign n19715 = x127 & n10106;
  assign n19716 = ~n19714 & ~n19715;
  assign n19717 = x126 & n9503;
  assign n19718 = n19716 & ~n19717;
  assign n19719 = ~n19713 & n19718;
  assign n19720 = n19719 ^ x62;
  assign n19708 = n8724 & n10099;
  assign n19709 = x124 ^ x123;
  assign n19710 = n9798 & n19709;
  assign n19711 = ~n19708 & ~n19710;
  assign n19712 = n19711 ^ x59;
  assign n19721 = n19720 ^ n19712;
  assign n19706 = n19683 & n19693;
  assign n19707 = n19706 ^ n19692;
  assign n19722 = n19721 ^ n19707;
  assign n19739 = n19738 ^ n19722;
  assign n19763 = n19722 & ~n19726;
  assign n19764 = ~n19727 & ~n19763;
  assign n19765 = ~n19722 & ~n19723;
  assign n19766 = ~n19731 & ~n19765;
  assign n19767 = ~n19764 & n19766;
  assign n19768 = ~n19672 & ~n19767;
  assign n19769 = n19724 & ~n19763;
  assign n19770 = ~n19733 & n19765;
  assign n19771 = ~n19769 & ~n19770;
  assign n19772 = ~n19768 & n19771;
  assign n19754 = n9499 & ~n9889;
  assign n19755 = x127 & n9503;
  assign n19756 = x126 & n9508;
  assign n19757 = ~n19755 & ~n19756;
  assign n19758 = ~n19754 & n19757;
  assign n19759 = n19758 ^ x62;
  assign n19746 = ~x59 & x123;
  assign n19747 = x124 ^ x122;
  assign n19748 = ~n10099 & n19747;
  assign n19749 = n19748 ^ x122;
  assign n19750 = ~n19746 & ~n19749;
  assign n19751 = x59 & ~x123;
  assign n19752 = ~n12465 & ~n19751;
  assign n19753 = ~n19750 & n19752;
  assign n19760 = n19759 ^ n19753;
  assign n19743 = x124 & n10099;
  assign n19744 = x125 & n9798;
  assign n19745 = ~n19743 & ~n19744;
  assign n19761 = n19760 ^ n19745;
  assign n19740 = n19720 ^ n19707;
  assign n19741 = n19721 & ~n19740;
  assign n19742 = n19741 ^ n19707;
  assign n19762 = n19761 ^ n19742;
  assign n19773 = n19772 ^ n19762;
  assign n19788 = n19742 & ~n19761;
  assign n19789 = n19771 & ~n19788;
  assign n19790 = ~n19768 & n19789;
  assign n19791 = ~n19742 & n19761;
  assign n19792 = ~n19790 & ~n19791;
  assign n19783 = n9499 & n10430;
  assign n19784 = x127 & n9508;
  assign n19785 = ~n19783 & ~n19784;
  assign n19777 = n9911 & n10099;
  assign n19778 = x126 ^ x125;
  assign n19779 = ~x62 & ~n19778;
  assign n19780 = ~n19777 & ~n19779;
  assign n19781 = ~x63 & n19778;
  assign n19782 = n19780 & ~n19781;
  assign n19786 = n19785 ^ n19782;
  assign n19774 = n19753 ^ n19745;
  assign n19775 = ~n19760 & ~n19774;
  assign n19776 = n19775 ^ n19759;
  assign n19787 = n19786 ^ n19776;
  assign n19793 = n19792 ^ n19787;
  assign n19804 = n19785 ^ x126;
  assign n19805 = n19778 & ~n19804;
  assign n19806 = x63 & n19805;
  assign n19807 = n19806 ^ n19785;
  assign n19808 = ~x62 & n19807;
  assign n19809 = ~n9288 & n19785;
  assign n19810 = ~n9286 & n10099;
  assign n19811 = ~n19809 & n19810;
  assign n19812 = ~n9595 & n19785;
  assign n19813 = ~n9597 & n13628;
  assign n19814 = ~n19812 & n19813;
  assign n19815 = ~n19811 & ~n19814;
  assign n19816 = ~n19808 & n19815;
  assign n19797 = x126 ^ x124;
  assign n19798 = n10099 & n19797;
  assign n19799 = x127 ^ x125;
  assign n19800 = ~x63 & n19799;
  assign n19801 = ~n19798 & ~n19800;
  assign n19802 = ~x62 & ~n19799;
  assign n19803 = n19801 & ~n19802;
  assign n19817 = n19816 ^ n19803;
  assign n19794 = n19792 ^ n19776;
  assign n19795 = n19787 & ~n19794;
  assign n19796 = n19795 ^ n19792;
  assign n19818 = n19817 ^ n19796;
  assign n19822 = x124 & x126;
  assign n19823 = x127 & ~n19822;
  assign n19824 = ~x125 & ~x127;
  assign n19825 = ~x62 & ~n19824;
  assign n19826 = ~n19823 & ~n19825;
  assign n19827 = x63 & ~n19826;
  assign n19828 = n9887 & n19743;
  assign n19829 = x125 & x127;
  assign n19830 = n13628 & n19829;
  assign n19831 = ~n19828 & ~n19830;
  assign n19832 = ~n19827 & n19831;
  assign n19819 = n19816 ^ n19796;
  assign n19820 = n19817 & n19819;
  assign n19821 = n19820 ^ n19796;
  assign n19833 = n19832 ^ n19821;
  assign y0 = n129;
  assign y1 = n132;
  assign y2 = n145;
  assign y3 = n170;
  assign y4 = ~n194;
  assign y5 = n241;
  assign y6 = ~n282;
  assign y7 = n340;
  assign y8 = ~n394;
  assign y9 = ~n445;
  assign y10 = n498;
  assign y11 = ~n574;
  assign y12 = n636;
  assign y13 = ~n700;
  assign y14 = ~n780;
  assign y15 = ~n855;
  assign y16 = n934;
  assign y17 = n1035;
  assign y18 = n1122;
  assign y19 = ~n1211;
  assign y20 = ~n1325;
  assign y21 = ~n1426;
  assign y22 = n1528;
  assign y23 = ~n1655;
  assign y24 = n1768;
  assign y25 = ~n1883;
  assign y26 = ~n2020;
  assign y27 = ~n2145;
  assign y28 = ~n2273;
  assign y29 = n2425;
  assign y30 = n2566;
  assign y31 = n2707;
  assign y32 = n2873;
  assign y33 = ~n3028;
  assign y34 = n3189;
  assign y35 = ~n3369;
  assign y36 = n3534;
  assign y37 = n3704;
  assign y38 = n3903;
  assign y39 = ~n4084;
  assign y40 = n4266;
  assign y41 = ~n4461;
  assign y42 = n4650;
  assign y43 = ~n4845;
  assign y44 = n5066;
  assign y45 = n5273;
  assign y46 = ~n5484;
  assign y47 = n5717;
  assign y48 = n5935;
  assign y49 = n6156;
  assign y50 = n6401;
  assign y51 = n6634;
  assign y52 = ~n6872;
  assign y53 = n7130;
  assign y54 = ~n7374;
  assign y55 = n7621;
  assign y56 = n7890;
  assign y57 = ~n8162;
  assign y58 = ~n8423;
  assign y59 = ~n8714;
  assign y60 = n8989;
  assign y61 = ~n9276;
  assign y62 = n9581;
  assign y63 = ~n9875;
  assign y64 = ~n10164;
  assign y65 = n10440;
  assign y66 = ~n10712;
  assign y67 = n10989;
  assign y68 = ~n11270;
  assign y69 = ~n11549;
  assign y70 = n11813;
  assign y71 = ~n12070;
  assign y72 = n12334;
  assign y73 = n12590;
  assign y74 = ~n12837;
  assign y75 = n13072;
  assign y76 = ~n13302;
  assign y77 = ~n13532;
  assign y78 = ~n13777;
  assign y79 = ~n14007;
  assign y80 = ~n14242;
  assign y81 = n14470;
  assign y82 = n14690;
  assign y83 = ~n14910;
  assign y84 = n15114;
  assign y85 = n15316;
  assign y86 = ~n15506;
  assign y87 = n15690;
  assign y88 = n15879;
  assign y89 = ~n16072;
  assign y90 = n16251;
  assign y91 = n16427;
  assign y92 = ~n16599;
  assign y93 = n16753;
  assign y94 = n16918;
  assign y95 = n17081;
  assign y96 = n17232;
  assign y97 = n17376;
  assign y98 = n17527;
  assign y99 = ~n17671;
  assign y100 = ~n17801;
  assign y101 = n17932;
  assign y102 = ~n18049;
  assign y103 = n18175;
  assign y104 = n18291;
  assign y105 = n18406;
  assign y106 = ~n18509;
  assign y107 = n18612;
  assign y108 = n18723;
  assign y109 = n18819;
  assign y110 = n18919;
  assign y111 = ~n19011;
  assign y112 = n19101;
  assign y113 = n19181;
  assign y114 = n19271;
  assign y115 = n19339;
  assign y116 = ~n19407;
  assign y117 = n19460;
  assign y118 = n19522;
  assign y119 = n19574;
  assign y120 = ~n19625;
  assign y121 = n19669;
  assign y122 = ~n19705;
  assign y123 = ~n19739;
  assign y124 = n19773;
  assign y125 = ~n19793;
  assign y126 = ~n19818;
  assign y127 = n19833;
endmodule
