module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63;
  wire n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628;
  assign n129 = x105 ^ x58;
  assign n130 = x96 ^ x32;
  assign n131 = n129 & ~n130;
  assign n132 = x82 ^ x0;
  assign n133 = x72 ^ x8;
  assign n134 = ~n132 & n133;
  assign n135 = x65 ^ x16;
  assign n136 = x120 ^ x24;
  assign n137 = ~n135 & ~n136;
  assign n138 = n134 & n137;
  assign n139 = n131 & n138;
  assign n140 = n132 & ~n133;
  assign n141 = ~n135 & n136;
  assign n142 = n140 & n141;
  assign n143 = n135 & n136;
  assign n144 = ~n132 & ~n133;
  assign n145 = n143 & n144;
  assign n146 = ~n142 & ~n145;
  assign n147 = n131 & ~n146;
  assign n148 = ~n129 & ~n130;
  assign n149 = n132 & n133;
  assign n150 = n135 & ~n136;
  assign n151 = n149 & n150;
  assign n152 = n144 & n150;
  assign n153 = ~n151 & ~n152;
  assign n154 = n148 & ~n153;
  assign n155 = ~n147 & ~n154;
  assign n156 = n129 & n130;
  assign n157 = n145 & n156;
  assign n158 = n134 & n150;
  assign n159 = n137 & n140;
  assign n160 = ~n158 & ~n159;
  assign n161 = n148 & ~n160;
  assign n162 = n137 & n144;
  assign n163 = n140 & n150;
  assign n164 = ~n162 & ~n163;
  assign n165 = n131 & ~n164;
  assign n166 = ~n161 & ~n165;
  assign n167 = ~n157 & n166;
  assign n168 = n143 & n149;
  assign n169 = n131 & n168;
  assign n170 = ~n129 & n130;
  assign n171 = ~n164 & n170;
  assign n172 = ~n169 & ~n171;
  assign n173 = n134 & n143;
  assign n174 = n140 & n143;
  assign n175 = ~n173 & ~n174;
  assign n176 = n170 & ~n175;
  assign n177 = n141 & n144;
  assign n178 = n170 & n177;
  assign n179 = n148 & n173;
  assign n180 = ~n178 & ~n179;
  assign n181 = n134 & n141;
  assign n182 = n137 & n149;
  assign n183 = ~n181 & ~n182;
  assign n184 = n131 & ~n183;
  assign n185 = n141 & n149;
  assign n186 = ~n138 & ~n151;
  assign n187 = ~n185 & n186;
  assign n188 = n170 & ~n187;
  assign n189 = ~n184 & ~n188;
  assign n190 = ~n148 & ~n156;
  assign n191 = ~n174 & ~n181;
  assign n192 = ~n142 & n191;
  assign n193 = ~n190 & ~n192;
  assign n194 = n153 & ~n158;
  assign n195 = ~n182 & n194;
  assign n196 = n156 & ~n195;
  assign n197 = ~n193 & ~n196;
  assign n198 = n189 & n197;
  assign n199 = n180 & n198;
  assign n200 = ~n176 & n199;
  assign n201 = n172 & n200;
  assign n202 = n167 & n201;
  assign n203 = n155 & n202;
  assign n204 = ~n139 & n203;
  assign n205 = n204 ^ x27;
  assign n206 = n205 ^ x113;
  assign n207 = x85 ^ x2;
  assign n208 = x67 ^ x28;
  assign n209 = ~n207 & n208;
  assign n210 = x91 ^ x60;
  assign n211 = x102 ^ x52;
  assign n212 = x100 ^ x36;
  assign n213 = x117 ^ x44;
  assign n214 = n212 & ~n213;
  assign n215 = ~n211 & n214;
  assign n216 = ~n210 & n215;
  assign n217 = n209 & n216;
  assign n218 = ~n207 & ~n208;
  assign n219 = ~n212 & n213;
  assign n220 = ~n210 & n211;
  assign n221 = n219 & n220;
  assign n222 = n210 & n212;
  assign n223 = ~n211 & n213;
  assign n224 = n222 & n223;
  assign n225 = ~n221 & ~n224;
  assign n226 = n218 & ~n225;
  assign n227 = ~n217 & ~n226;
  assign n228 = n207 & ~n208;
  assign n229 = ~n213 & n222;
  assign n230 = ~n211 & n229;
  assign n231 = n228 & n230;
  assign n232 = n207 & n208;
  assign n233 = n224 & n232;
  assign n234 = n213 & n222;
  assign n235 = n211 & n234;
  assign n236 = ~n212 & ~n213;
  assign n237 = n211 & n236;
  assign n238 = n210 & n237;
  assign n239 = ~n235 & ~n238;
  assign n240 = n218 & ~n239;
  assign n241 = ~n233 & ~n240;
  assign n242 = ~n231 & n241;
  assign n243 = n209 & n221;
  assign n244 = ~n212 & n223;
  assign n245 = ~n210 & n244;
  assign n246 = ~n216 & ~n245;
  assign n247 = n232 & ~n246;
  assign n248 = ~n243 & ~n247;
  assign n249 = n214 & n220;
  assign n250 = n232 & n249;
  assign n251 = n216 & n218;
  assign n252 = ~n250 & ~n251;
  assign n253 = ~n211 & n236;
  assign n254 = ~n210 & n253;
  assign n255 = n212 & n220;
  assign n256 = n213 & n255;
  assign n257 = ~n238 & ~n256;
  assign n258 = ~n254 & n257;
  assign n259 = ~n230 & n258;
  assign n260 = n232 & ~n259;
  assign n261 = n211 & n229;
  assign n262 = n212 & n223;
  assign n263 = ~n210 & n262;
  assign n264 = ~n261 & ~n263;
  assign n265 = n211 & n219;
  assign n266 = n210 & n265;
  assign n267 = n210 & n244;
  assign n268 = ~n254 & ~n267;
  assign n269 = ~n224 & n268;
  assign n270 = ~n266 & n269;
  assign n271 = n264 & n270;
  assign n272 = n209 & ~n271;
  assign n273 = n210 & n253;
  assign n274 = ~n249 & ~n273;
  assign n275 = ~n266 & n274;
  assign n276 = n275 ^ n207;
  assign n277 = n276 ^ n275;
  assign n278 = n220 & n236;
  assign n279 = ~n263 & ~n278;
  assign n280 = ~n235 & n279;
  assign n281 = ~n267 & n274;
  assign n282 = n280 & n281;
  assign n283 = ~n256 & n282;
  assign n284 = n283 ^ n275;
  assign n285 = n277 & n284;
  assign n286 = n285 ^ n275;
  assign n287 = ~n208 & ~n286;
  assign n288 = ~n272 & ~n287;
  assign n289 = ~n260 & n288;
  assign n290 = n252 & n289;
  assign n291 = n248 & n290;
  assign n292 = n242 & n291;
  assign n293 = n227 & n292;
  assign n294 = n293 ^ x1;
  assign n295 = n294 ^ x123;
  assign n296 = ~n206 & n295;
  assign n297 = x124 ^ x4;
  assign n298 = x83 ^ x30;
  assign n299 = ~n297 & n298;
  assign n300 = x84 ^ x62;
  assign n301 = x78 ^ x38;
  assign n302 = n300 & ~n301;
  assign n303 = x126 ^ x46;
  assign n304 = x101 ^ x54;
  assign n305 = ~n303 & n304;
  assign n306 = n302 & n305;
  assign n307 = n300 & n301;
  assign n308 = ~n303 & ~n304;
  assign n309 = n307 & n308;
  assign n310 = ~n306 & ~n309;
  assign n311 = n299 & ~n310;
  assign n312 = n297 & ~n298;
  assign n313 = n303 ^ n300;
  assign n314 = n313 ^ n301;
  assign n315 = n314 ^ n300;
  assign n316 = n315 ^ n304;
  assign n317 = n316 ^ n301;
  assign n318 = n301 ^ n300;
  assign n319 = n304 ^ n300;
  assign n320 = n319 ^ n300;
  assign n321 = n318 & n320;
  assign n322 = n321 ^ n300;
  assign n323 = ~n317 & ~n322;
  assign n324 = n323 ^ n314;
  assign n325 = n312 & n324;
  assign n326 = n298 ^ n297;
  assign n327 = ~n300 & n301;
  assign n328 = n308 & n327;
  assign n329 = n303 & n304;
  assign n330 = ~n300 & ~n301;
  assign n331 = n329 & n330;
  assign n332 = ~n328 & ~n331;
  assign n333 = ~n326 & ~n332;
  assign n334 = n297 & n298;
  assign n335 = n302 & n308;
  assign n336 = n302 & n329;
  assign n337 = n303 & ~n304;
  assign n338 = n327 & n337;
  assign n339 = n302 & n337;
  assign n340 = n305 & n307;
  assign n341 = ~n339 & ~n340;
  assign n342 = ~n338 & n341;
  assign n343 = ~n336 & n342;
  assign n344 = ~n335 & n343;
  assign n345 = n334 & ~n344;
  assign n346 = n327 & n329;
  assign n347 = n330 & n337;
  assign n348 = n305 & n327;
  assign n349 = ~n347 & ~n348;
  assign n350 = ~n346 & n349;
  assign n351 = ~n328 & n350;
  assign n352 = ~n336 & n351;
  assign n353 = n299 & ~n352;
  assign n354 = ~n297 & ~n298;
  assign n355 = n307 & n329;
  assign n356 = ~n335 & ~n355;
  assign n357 = ~n339 & n356;
  assign n358 = n349 & n357;
  assign n359 = ~n340 & n358;
  assign n360 = n354 & ~n359;
  assign n361 = ~n353 & ~n360;
  assign n362 = ~n345 & n361;
  assign n363 = ~n333 & n362;
  assign n364 = ~n325 & n363;
  assign n365 = ~n311 & n364;
  assign n366 = n305 & n330;
  assign n367 = n366 ^ n297;
  assign n368 = n367 ^ n366;
  assign n369 = n366 ^ n331;
  assign n370 = ~n368 & n369;
  assign n371 = n370 ^ n366;
  assign n372 = n298 & n371;
  assign n373 = n365 & ~n372;
  assign n374 = n373 ^ x35;
  assign n375 = n374 ^ x99;
  assign n376 = x110 ^ x36;
  assign n377 = x92 ^ x62;
  assign n378 = ~n376 & ~n377;
  assign n379 = x86 ^ x4;
  assign n380 = x68 ^ x20;
  assign n381 = n379 & n380;
  assign n382 = x93 ^ x28;
  assign n383 = x116 ^ x12;
  assign n384 = ~n382 & ~n383;
  assign n385 = n381 & n384;
  assign n386 = n378 & n385;
  assign n387 = ~n376 & n377;
  assign n388 = n382 & n383;
  assign n389 = ~n379 & n380;
  assign n390 = n388 & n389;
  assign n391 = n382 & ~n383;
  assign n392 = n381 & n391;
  assign n393 = ~n390 & ~n392;
  assign n394 = ~n379 & ~n380;
  assign n395 = n384 & n394;
  assign n396 = n379 & ~n380;
  assign n397 = ~n382 & n383;
  assign n398 = n396 & n397;
  assign n399 = ~n395 & ~n398;
  assign n400 = n393 & n399;
  assign n401 = n387 & ~n400;
  assign n402 = ~n386 & ~n401;
  assign n403 = n378 & n398;
  assign n404 = n384 & n396;
  assign n405 = n384 & n389;
  assign n406 = ~n404 & ~n405;
  assign n407 = n387 & ~n406;
  assign n408 = ~n403 & ~n407;
  assign n409 = n388 & n396;
  assign n410 = n391 & n394;
  assign n411 = ~n409 & ~n410;
  assign n412 = n377 & ~n411;
  assign n413 = n389 & n391;
  assign n414 = ~n392 & ~n413;
  assign n415 = n381 & n388;
  assign n416 = n388 & n394;
  assign n417 = ~n415 & ~n416;
  assign n418 = n414 & n417;
  assign n419 = n378 & ~n418;
  assign n420 = n376 & n377;
  assign n421 = n391 & n396;
  assign n422 = ~n413 & ~n421;
  assign n423 = ~n404 & n422;
  assign n424 = n420 & ~n423;
  assign n425 = ~n419 & ~n424;
  assign n426 = ~n412 & n425;
  assign n427 = n377 ^ n376;
  assign n428 = n389 & n397;
  assign n429 = n428 ^ n377;
  assign n430 = n429 ^ n428;
  assign n431 = n394 & n397;
  assign n432 = n381 & n397;
  assign n433 = ~n431 & ~n432;
  assign n434 = ~n390 & n433;
  assign n435 = ~n415 & n434;
  assign n436 = n411 & n435;
  assign n437 = n406 & n436;
  assign n438 = n437 ^ n428;
  assign n439 = n438 ^ n428;
  assign n440 = ~n430 & ~n439;
  assign n441 = n440 ^ n428;
  assign n442 = n427 & n441;
  assign n443 = n442 ^ n428;
  assign n444 = n426 & ~n443;
  assign n445 = n408 & n444;
  assign n446 = n431 ^ n420;
  assign n447 = n431 ^ n378;
  assign n448 = n447 ^ n378;
  assign n449 = n432 ^ n378;
  assign n450 = ~n448 & ~n449;
  assign n451 = n450 ^ n378;
  assign n452 = n446 & n451;
  assign n453 = n452 ^ n420;
  assign n454 = n445 & ~n453;
  assign n455 = n402 & n454;
  assign n456 = n455 ^ x43;
  assign n457 = n456 ^ x80;
  assign n458 = n375 & n457;
  assign n459 = x104 ^ x60;
  assign n460 = x122 ^ x34;
  assign n461 = n459 & ~n460;
  assign n462 = x99 ^ x18;
  assign n463 = x90 ^ x10;
  assign n464 = n462 & n463;
  assign n465 = x81 ^ x2;
  assign n466 = x64 ^ x26;
  assign n467 = n465 & ~n466;
  assign n468 = n464 & n467;
  assign n469 = n461 & n468;
  assign n470 = n459 & n460;
  assign n471 = n465 & n466;
  assign n472 = ~n462 & n463;
  assign n473 = n471 & n472;
  assign n474 = n470 & n473;
  assign n475 = ~n469 & ~n474;
  assign n476 = ~n465 & ~n466;
  assign n477 = n462 & ~n463;
  assign n478 = n476 & n477;
  assign n479 = ~n465 & n466;
  assign n480 = n464 & n479;
  assign n481 = ~n478 & ~n480;
  assign n482 = n459 & ~n481;
  assign n483 = n472 & n476;
  assign n484 = n471 & n477;
  assign n485 = n467 & n477;
  assign n486 = ~n462 & ~n463;
  assign n487 = n471 & n486;
  assign n488 = ~n485 & ~n487;
  assign n489 = ~n484 & n488;
  assign n490 = ~n483 & n489;
  assign n491 = n461 & ~n490;
  assign n492 = n467 & n472;
  assign n493 = n464 & n471;
  assign n494 = n467 & n486;
  assign n495 = ~n493 & ~n494;
  assign n496 = ~n484 & n495;
  assign n497 = ~n492 & n496;
  assign n498 = n470 & ~n497;
  assign n499 = ~n491 & ~n498;
  assign n500 = ~n482 & n499;
  assign n501 = ~n459 & ~n460;
  assign n502 = ~n484 & ~n494;
  assign n503 = ~n473 & n502;
  assign n504 = n472 & n479;
  assign n505 = n479 & n486;
  assign n506 = n464 & n476;
  assign n507 = ~n505 & ~n506;
  assign n508 = ~n504 & n507;
  assign n509 = n503 & n508;
  assign n510 = n481 & n509;
  assign n511 = n501 & n510;
  assign n512 = ~n459 & n460;
  assign n513 = n476 & n486;
  assign n514 = ~n485 & n509;
  assign n515 = ~n513 & n514;
  assign n516 = n512 & ~n515;
  assign n517 = ~n511 & ~n516;
  assign n518 = n500 & n517;
  assign n519 = n475 & n518;
  assign n520 = n513 ^ n460;
  assign n521 = n520 ^ n513;
  assign n522 = n513 ^ n504;
  assign n523 = ~n521 & n522;
  assign n524 = n523 ^ n513;
  assign n525 = n459 & n524;
  assign n526 = n519 & ~n525;
  assign n527 = n526 ^ x51;
  assign n528 = n527 ^ x81;
  assign n529 = x114 ^ x56;
  assign n530 = x123 ^ x40;
  assign n531 = n529 & n530;
  assign n532 = x97 ^ x48;
  assign n533 = x112 ^ x32;
  assign n534 = n532 & ~n533;
  assign n535 = n531 & n534;
  assign n536 = x73 ^ x6;
  assign n537 = x80 ^ x24;
  assign n538 = ~n536 & n537;
  assign n539 = ~n532 & ~n533;
  assign n540 = ~n529 & ~n530;
  assign n541 = n539 & n540;
  assign n542 = n538 & n541;
  assign n543 = n536 & n537;
  assign n544 = n532 & n533;
  assign n545 = n529 & ~n530;
  assign n546 = n544 & n545;
  assign n547 = n543 & n546;
  assign n548 = ~n542 & ~n547;
  assign n549 = n538 & n546;
  assign n550 = ~n536 & ~n537;
  assign n551 = ~n532 & n533;
  assign n552 = ~n529 & n530;
  assign n553 = n551 & n552;
  assign n554 = n550 & n553;
  assign n555 = ~n549 & ~n554;
  assign n556 = n544 & n552;
  assign n557 = n538 & n556;
  assign n558 = n531 & n539;
  assign n559 = n543 & n558;
  assign n560 = ~n557 & ~n559;
  assign n561 = n539 & n545;
  assign n562 = n543 & n561;
  assign n563 = n536 & ~n537;
  assign n564 = n540 & n551;
  assign n565 = ~n541 & ~n564;
  assign n566 = n563 & ~n565;
  assign n567 = n537 ^ n536;
  assign n568 = n534 & n540;
  assign n569 = ~n567 & n568;
  assign n570 = ~n561 & ~n564;
  assign n571 = n534 & n545;
  assign n572 = n531 & n544;
  assign n573 = ~n558 & ~n572;
  assign n574 = ~n571 & n573;
  assign n575 = n570 & n574;
  assign n576 = n550 & ~n575;
  assign n577 = ~n569 & ~n576;
  assign n578 = n534 & n552;
  assign n579 = ~n553 & ~n556;
  assign n580 = ~n578 & n579;
  assign n581 = n543 & ~n580;
  assign n582 = n545 & n551;
  assign n583 = n539 & n552;
  assign n584 = n540 & n544;
  assign n585 = ~n583 & ~n584;
  assign n586 = ~n553 & n585;
  assign n587 = ~n582 & n586;
  assign n588 = n538 & ~n587;
  assign n589 = ~n578 & ~n584;
  assign n590 = n533 ^ n532;
  assign n591 = n590 ^ n532;
  assign n592 = n532 ^ n530;
  assign n593 = n591 & n592;
  assign n594 = n593 ^ n532;
  assign n595 = n529 & n594;
  assign n596 = n589 & ~n595;
  assign n597 = n563 & ~n596;
  assign n598 = ~n588 & ~n597;
  assign n599 = ~n581 & n598;
  assign n600 = n577 & n599;
  assign n601 = ~n566 & n600;
  assign n602 = ~n562 & n601;
  assign n603 = n560 & n602;
  assign n604 = n555 & n603;
  assign n605 = n548 & n604;
  assign n606 = ~n535 & n605;
  assign n607 = n606 ^ x59;
  assign n608 = n607 ^ x90;
  assign n609 = n528 & ~n608;
  assign n610 = n458 & n609;
  assign n611 = n296 & n610;
  assign n612 = ~n375 & n457;
  assign n613 = n528 & n608;
  assign n614 = n612 & n613;
  assign n615 = n296 & n614;
  assign n616 = n206 & ~n295;
  assign n617 = n609 & n612;
  assign n618 = n616 & n617;
  assign n619 = ~n615 & ~n618;
  assign n620 = ~n611 & n619;
  assign n621 = n614 & n616;
  assign n622 = ~n528 & n608;
  assign n623 = n458 & n622;
  assign n624 = n616 & n623;
  assign n625 = n206 & n295;
  assign n626 = n610 & n625;
  assign n627 = ~n624 & ~n626;
  assign n628 = ~n621 & n627;
  assign n629 = n296 & n623;
  assign n630 = ~n206 & ~n295;
  assign n631 = n612 & n622;
  assign n632 = n375 & ~n457;
  assign n633 = n622 & n632;
  assign n634 = ~n631 & ~n633;
  assign n635 = n630 & ~n634;
  assign n636 = ~n629 & ~n635;
  assign n637 = ~n375 & ~n457;
  assign n638 = n613 & n637;
  assign n639 = n458 & n613;
  assign n640 = ~n638 & ~n639;
  assign n641 = n630 & ~n640;
  assign n642 = ~n528 & ~n608;
  assign n643 = n458 & n642;
  assign n644 = n612 & n642;
  assign n645 = ~n643 & ~n644;
  assign n646 = n296 & ~n645;
  assign n647 = ~n641 & ~n646;
  assign n648 = n609 & n632;
  assign n649 = ~n644 & ~n648;
  assign n650 = n616 & ~n649;
  assign n651 = n295 ^ n206;
  assign n652 = n632 & n642;
  assign n653 = n622 & n637;
  assign n654 = n613 & n632;
  assign n655 = ~n653 & ~n654;
  assign n656 = ~n652 & n655;
  assign n657 = n651 & ~n656;
  assign n658 = n630 & n652;
  assign n659 = n609 & n637;
  assign n660 = ~n643 & ~n659;
  assign n661 = n625 & ~n660;
  assign n662 = ~n658 & ~n661;
  assign n663 = n637 & n642;
  assign n664 = ~n610 & ~n659;
  assign n665 = ~n663 & n664;
  assign n666 = n630 & ~n665;
  assign n667 = ~n614 & ~n663;
  assign n668 = ~n638 & n667;
  assign n669 = ~n633 & n668;
  assign n670 = ~n644 & n669;
  assign n671 = n625 & ~n670;
  assign n672 = ~n666 & ~n671;
  assign n673 = n662 & n672;
  assign n674 = ~n657 & n673;
  assign n675 = ~n650 & n674;
  assign n676 = n647 & n675;
  assign n677 = n636 & n676;
  assign n678 = n628 & n677;
  assign n679 = n620 & n678;
  assign n680 = n679 ^ x4;
  assign n681 = n680 ^ x100;
  assign n682 = ~n468 & ~n478;
  assign n683 = ~n505 & n682;
  assign n684 = n477 & n479;
  assign n685 = ~n506 & ~n684;
  assign n686 = n495 & n685;
  assign n687 = n683 & n686;
  assign n688 = ~n473 & n687;
  assign n689 = n512 & n688;
  assign n690 = n496 & n685;
  assign n691 = n461 & ~n690;
  assign n692 = ~n689 & ~n691;
  assign n693 = ~n480 & n683;
  assign n694 = ~n485 & n693;
  assign n695 = n470 & ~n694;
  assign n696 = n466 ^ n462;
  assign n697 = n696 ^ n463;
  assign n698 = n697 ^ n466;
  assign n699 = n466 ^ n465;
  assign n700 = n699 ^ n465;
  assign n701 = n465 ^ n463;
  assign n702 = n701 ^ n465;
  assign n703 = n700 & ~n702;
  assign n704 = n703 ^ n465;
  assign n705 = n698 & n704;
  assign n706 = n705 ^ n696;
  assign n707 = n706 ^ n483;
  assign n708 = n707 ^ n483;
  assign n709 = n483 ^ n460;
  assign n710 = n709 ^ n483;
  assign n711 = n708 & ~n710;
  assign n712 = n711 ^ n483;
  assign n713 = ~n459 & n712;
  assign n714 = n713 ^ n483;
  assign n715 = ~n695 & ~n714;
  assign n716 = n692 & n715;
  assign n717 = n475 & n716;
  assign n718 = ~n525 & n717;
  assign n719 = n718 ^ x37;
  assign n720 = n719 ^ x102;
  assign n721 = n232 & n266;
  assign n722 = n242 & ~n721;
  assign n723 = n218 & n230;
  assign n724 = ~n249 & n270;
  assign n725 = ~n245 & n724;
  assign n726 = ~n256 & n725;
  assign n727 = n228 & ~n726;
  assign n728 = ~n723 & ~n727;
  assign n729 = n208 ^ n207;
  assign n730 = n261 & ~n729;
  assign n731 = ~n256 & ~n278;
  assign n732 = ~n267 & n731;
  assign n733 = n232 & ~n732;
  assign n734 = n246 & ~n273;
  assign n735 = ~n263 & n734;
  assign n736 = n218 & ~n735;
  assign n737 = ~n209 & ~n736;
  assign n738 = n218 & ~n246;
  assign n739 = ~n266 & ~n273;
  assign n740 = ~n229 & n739;
  assign n741 = ~n738 & n740;
  assign n742 = n279 & n741;
  assign n743 = ~n256 & n742;
  assign n744 = ~n737 & ~n743;
  assign n745 = ~n733 & ~n744;
  assign n746 = ~n730 & n745;
  assign n747 = n728 & n746;
  assign n748 = n248 & n747;
  assign n749 = n722 & n748;
  assign n750 = n749 ^ x63;
  assign n751 = n750 ^ x84;
  assign n752 = n720 & n751;
  assign n753 = x121 ^ x26;
  assign n754 = x66 ^ x0;
  assign n755 = n753 & ~n754;
  assign n756 = x98 ^ x58;
  assign n757 = x89 ^ x50;
  assign n758 = ~n756 & n757;
  assign n759 = x88 ^ x42;
  assign n760 = x107 ^ x34;
  assign n761 = ~n759 & ~n760;
  assign n762 = n758 & n761;
  assign n763 = n755 & n762;
  assign n764 = n753 & n754;
  assign n765 = n759 & n760;
  assign n766 = n758 & n765;
  assign n767 = n764 & n766;
  assign n768 = ~n753 & n754;
  assign n769 = n759 & ~n760;
  assign n770 = n758 & n769;
  assign n771 = n756 & n757;
  assign n772 = n761 & n771;
  assign n773 = ~n759 & n760;
  assign n774 = n756 & ~n757;
  assign n775 = n773 & n774;
  assign n776 = ~n772 & ~n775;
  assign n777 = ~n770 & n776;
  assign n778 = n768 & ~n777;
  assign n779 = ~n767 & ~n778;
  assign n780 = ~n763 & n779;
  assign n781 = n754 ^ n753;
  assign n782 = n761 & n774;
  assign n783 = ~n781 & n782;
  assign n784 = n766 & n768;
  assign n785 = ~n783 & ~n784;
  assign n786 = ~n756 & ~n757;
  assign n787 = n761 & n786;
  assign n788 = n764 & n787;
  assign n789 = ~n753 & ~n754;
  assign n790 = n766 & n789;
  assign n791 = n765 & n771;
  assign n792 = n769 & n774;
  assign n793 = ~n791 & ~n792;
  assign n794 = n755 & ~n793;
  assign n795 = ~n790 & ~n794;
  assign n796 = ~n788 & n795;
  assign n797 = n765 & n786;
  assign n798 = n764 & n797;
  assign n799 = n769 & n786;
  assign n800 = n768 & n799;
  assign n801 = ~n798 & ~n800;
  assign n802 = n768 & n791;
  assign n803 = n758 & n773;
  assign n804 = n773 & n786;
  assign n805 = ~n803 & ~n804;
  assign n806 = n755 & ~n805;
  assign n807 = ~n802 & ~n806;
  assign n808 = ~n770 & ~n782;
  assign n809 = n755 & ~n808;
  assign n810 = n789 & ~n805;
  assign n811 = ~n809 & ~n810;
  assign n812 = ~n792 & ~n804;
  assign n813 = n768 & ~n812;
  assign n814 = n769 & n771;
  assign n815 = n765 & n774;
  assign n816 = ~n814 & ~n815;
  assign n817 = ~n762 & n816;
  assign n818 = ~n781 & ~n817;
  assign n819 = ~n813 & ~n818;
  assign n820 = n811 & n819;
  assign n821 = n807 & n820;
  assign n822 = n771 & n773;
  assign n823 = n822 ^ n799;
  assign n824 = n823 ^ n822;
  assign n825 = n822 ^ n754;
  assign n826 = n825 ^ n822;
  assign n827 = n824 & ~n826;
  assign n828 = n827 ^ n822;
  assign n829 = n781 & n828;
  assign n830 = n829 ^ n822;
  assign n831 = n821 & ~n830;
  assign n832 = n801 & n831;
  assign n833 = n796 & n832;
  assign n834 = n785 & n833;
  assign n835 = n780 & n834;
  assign n836 = n835 ^ x5;
  assign n837 = n836 ^ x78;
  assign n838 = x94 ^ x56;
  assign n839 = x108 ^ x38;
  assign n840 = n838 & n839;
  assign n841 = x125 ^ x14;
  assign n842 = x77 ^ x30;
  assign n843 = x76 ^ x22;
  assign n844 = x118 ^ x6;
  assign n845 = ~n843 & ~n844;
  assign n846 = ~n842 & n845;
  assign n847 = ~n841 & n846;
  assign n848 = ~n842 & n843;
  assign n849 = ~n841 & n848;
  assign n850 = n844 & n849;
  assign n851 = ~n847 & ~n850;
  assign n852 = n840 & ~n851;
  assign n853 = n838 & ~n839;
  assign n854 = n841 & n842;
  assign n855 = n843 & n854;
  assign n856 = n844 & n855;
  assign n857 = n845 & n854;
  assign n858 = ~n856 & ~n857;
  assign n859 = n853 & ~n858;
  assign n860 = ~n838 & n839;
  assign n861 = n841 & n848;
  assign n862 = n844 & n861;
  assign n863 = n841 & n846;
  assign n864 = ~n862 & ~n863;
  assign n865 = n860 & ~n864;
  assign n866 = ~n859 & ~n865;
  assign n867 = ~n838 & ~n839;
  assign n868 = ~n843 & n844;
  assign n869 = ~n842 & n868;
  assign n870 = n867 & n869;
  assign n871 = ~n840 & ~n867;
  assign n872 = ~n844 & n849;
  assign n873 = ~n863 & ~n872;
  assign n874 = ~n871 & ~n873;
  assign n875 = ~n870 & ~n874;
  assign n876 = ~n841 & n842;
  assign n877 = n843 & n876;
  assign n878 = n853 & n877;
  assign n879 = ~n844 & n861;
  assign n880 = ~n850 & ~n879;
  assign n881 = n860 & ~n880;
  assign n882 = ~n844 & n855;
  assign n883 = n854 & n868;
  assign n884 = ~n882 & ~n883;
  assign n885 = n845 & n876;
  assign n886 = n844 & n877;
  assign n887 = ~n885 & ~n886;
  assign n888 = n884 & n887;
  assign n889 = n867 & ~n888;
  assign n890 = ~n853 & ~n889;
  assign n891 = n841 & n869;
  assign n892 = ~n872 & ~n891;
  assign n893 = ~n862 & n892;
  assign n894 = ~n867 & ~n885;
  assign n895 = ~n888 & ~n894;
  assign n896 = n893 & ~n895;
  assign n897 = ~n890 & ~n896;
  assign n898 = n868 & n876;
  assign n900 = ~n879 & n884;
  assign n899 = n858 & ~n885;
  assign n901 = n900 ^ n899;
  assign n902 = n899 ^ n860;
  assign n903 = n902 ^ n860;
  assign n904 = n860 ^ n840;
  assign n905 = n903 & ~n904;
  assign n906 = n905 ^ n860;
  assign n907 = n901 & n906;
  assign n908 = n907 ^ n900;
  assign n909 = ~n898 & n908;
  assign n910 = n839 & ~n909;
  assign n911 = ~n897 & ~n910;
  assign n912 = ~n881 & n911;
  assign n913 = ~n878 & n912;
  assign n914 = n875 & n913;
  assign n915 = n866 & n914;
  assign n916 = ~n852 & n915;
  assign n917 = n916 ^ x29;
  assign n918 = n917 ^ x85;
  assign n919 = ~n564 & ~n583;
  assign n920 = ~n567 & ~n919;
  assign n921 = n574 & n580;
  assign n922 = n538 & ~n921;
  assign n923 = ~n568 & n589;
  assign n924 = n923 ^ n537;
  assign n925 = n924 ^ n923;
  assign n926 = ~n553 & ~n568;
  assign n927 = ~n558 & n926;
  assign n928 = ~n535 & n927;
  assign n929 = ~n582 & n928;
  assign n930 = n929 ^ n923;
  assign n931 = ~n925 & n930;
  assign n932 = n931 ^ n923;
  assign n933 = n536 & ~n932;
  assign n934 = ~n922 & ~n933;
  assign n935 = ~n920 & n934;
  assign n936 = n531 & n590;
  assign n937 = ~n571 & ~n936;
  assign n938 = ~n556 & n937;
  assign n939 = ~n546 & n938;
  assign n940 = n939 ^ n572;
  assign n941 = n940 ^ n572;
  assign n942 = n572 ^ n537;
  assign n943 = n942 ^ n572;
  assign n944 = ~n941 & ~n943;
  assign n945 = n944 ^ n572;
  assign n946 = ~n536 & n945;
  assign n947 = n946 ^ n572;
  assign n948 = n935 & ~n947;
  assign n949 = ~n566 & n948;
  assign n950 = ~n562 & n949;
  assign n951 = n555 & n950;
  assign n952 = n548 & n951;
  assign n953 = n952 ^ x13;
  assign n954 = n953 ^ x108;
  assign n955 = n299 & n355;
  assign n956 = n334 & n346;
  assign n957 = ~n955 & ~n956;
  assign n958 = n297 & n331;
  assign n959 = n312 & ~n350;
  assign n960 = ~n958 & ~n959;
  assign n961 = n299 & n340;
  assign n962 = n308 & n330;
  assign n963 = ~n328 & ~n962;
  assign n964 = n334 & ~n963;
  assign n965 = ~n961 & ~n964;
  assign n966 = ~n338 & ~n347;
  assign n967 = ~n328 & ~n366;
  assign n968 = n966 & n967;
  assign n969 = n354 & ~n968;
  assign n970 = ~n309 & n357;
  assign n971 = n312 & ~n970;
  assign n972 = n306 & n334;
  assign n973 = n307 & n337;
  assign n974 = n335 & n354;
  assign n975 = ~n973 & ~n974;
  assign n976 = ~n972 & n975;
  assign n977 = ~n336 & n976;
  assign n978 = ~n340 & n977;
  assign n979 = ~n326 & ~n978;
  assign n980 = n335 & ~n970;
  assign n981 = n966 & ~n980;
  assign n982 = ~n346 & n981;
  assign n983 = n299 & ~n982;
  assign n984 = ~n979 & ~n983;
  assign n985 = ~n971 & n984;
  assign n986 = ~n969 & n985;
  assign n987 = n965 & n986;
  assign n988 = n960 & n987;
  assign n989 = n957 & n988;
  assign n990 = ~n311 & n989;
  assign n991 = n990 ^ x21;
  assign n992 = n991 ^ x91;
  assign n993 = ~n954 & n992;
  assign n994 = ~n918 & n993;
  assign n995 = n837 & n994;
  assign n996 = ~n837 & ~n918;
  assign n997 = n954 & n996;
  assign n998 = n992 & n997;
  assign n999 = ~n995 & ~n998;
  assign n1000 = n752 & ~n999;
  assign n1001 = n720 & ~n751;
  assign n1002 = n837 & n954;
  assign n1003 = ~n918 & n1002;
  assign n1004 = ~n992 & n1003;
  assign n1005 = ~n954 & n996;
  assign n1006 = ~n992 & n1005;
  assign n1007 = ~n1004 & ~n1006;
  assign n1008 = n1001 & ~n1007;
  assign n1009 = ~n1000 & ~n1008;
  assign n1010 = n752 & n1004;
  assign n1011 = ~n720 & ~n751;
  assign n1012 = ~n752 & ~n1011;
  assign n1013 = n1006 & ~n1012;
  assign n1014 = ~n918 & ~n954;
  assign n1015 = n837 & n1014;
  assign n1016 = ~n992 & n1015;
  assign n1017 = n999 & ~n1016;
  assign n1018 = n1011 & ~n1017;
  assign n1019 = ~n720 & n751;
  assign n1020 = n993 & n996;
  assign n1021 = n1019 & n1020;
  assign n1022 = n918 & n954;
  assign n1023 = ~n837 & n1022;
  assign n1024 = n992 & n1023;
  assign n1025 = n918 & ~n992;
  assign n1026 = n1002 & n1025;
  assign n1027 = ~n1024 & ~n1026;
  assign n1028 = n1011 & ~n1027;
  assign n1029 = ~n1021 & ~n1028;
  assign n1030 = n918 & n993;
  assign n1031 = ~n837 & n1030;
  assign n1032 = ~n1004 & ~n1031;
  assign n1033 = n1011 & ~n1032;
  assign n1034 = ~n992 & n997;
  assign n1035 = n992 & n1003;
  assign n1036 = n837 & n1030;
  assign n1037 = ~n1035 & ~n1036;
  assign n1038 = ~n1025 & n1037;
  assign n1039 = ~n1034 & n1038;
  assign n1040 = n1019 & ~n1039;
  assign n1041 = ~n1033 & ~n1040;
  assign n1042 = ~n1016 & ~n1020;
  assign n1043 = n1001 & ~n1042;
  assign n1051 = n918 & n1002;
  assign n1052 = n992 & n1051;
  assign n1046 = ~n954 & n1025;
  assign n1053 = ~n837 & n1046;
  assign n1044 = n954 & n1025;
  assign n1045 = ~n837 & n1044;
  assign n1054 = ~n1036 & ~n1045;
  assign n1055 = ~n1053 & n1054;
  assign n1056 = ~n1052 & n1055;
  assign n1047 = n837 & n1046;
  assign n1048 = ~n1045 & ~n1047;
  assign n1049 = ~n1031 & n1048;
  assign n1050 = ~n1024 & n1049;
  assign n1057 = n1056 ^ n1050;
  assign n1058 = n1056 ^ n751;
  assign n1059 = n1058 ^ n1056;
  assign n1060 = n1057 & n1059;
  assign n1061 = n1060 ^ n1056;
  assign n1062 = n720 & ~n1061;
  assign n1063 = ~n1043 & ~n1062;
  assign n1064 = n1041 & n1063;
  assign n1065 = n1029 & n1064;
  assign n1066 = ~n1018 & n1065;
  assign n1067 = ~n1013 & n1066;
  assign n1068 = ~n1010 & n1067;
  assign n1069 = n1009 & n1068;
  assign n1070 = n1069 ^ x30;
  assign n1071 = n1070 ^ x126;
  assign n1072 = n681 & n1071;
  assign n1073 = ~n871 & n885;
  assign n1074 = ~n841 & n869;
  assign n1075 = ~n879 & ~n1074;
  assign n1076 = ~n849 & n1075;
  assign n1077 = n853 & ~n1076;
  assign n1078 = ~n1073 & ~n1077;
  assign n1079 = n858 & ~n883;
  assign n1080 = n867 & ~n1079;
  assign n1081 = ~n844 & n877;
  assign n1082 = ~n855 & ~n1081;
  assign n1083 = n840 & ~n1082;
  assign n1084 = ~n863 & ~n891;
  assign n1085 = n840 & ~n1084;
  assign n1086 = ~n886 & n1079;
  assign n1087 = n853 & ~n1086;
  assign n1088 = ~n1085 & ~n1087;
  assign n1089 = n867 & ~n1076;
  assign n1090 = n843 ^ n842;
  assign n1091 = n1090 ^ n841;
  assign n1092 = n1091 ^ n841;
  assign n1093 = n844 & n1092;
  assign n1094 = n842 & n1093;
  assign n1095 = n1094 ^ n1091;
  assign n1096 = n860 & ~n1095;
  assign n1097 = ~n1089 & ~n1096;
  assign n1098 = n1088 & n1097;
  assign n1099 = ~n852 & n1098;
  assign n1100 = ~n1083 & n1099;
  assign n1101 = ~n1080 & n1100;
  assign n1102 = n1078 & n1101;
  assign n1103 = n1102 ^ x11;
  assign n1104 = n1103 ^ x82;
  assign n1105 = ~n772 & n816;
  assign n1106 = n768 & ~n1105;
  assign n1107 = ~n775 & ~n792;
  assign n1108 = ~n822 & n1107;
  assign n1109 = ~n781 & ~n1108;
  assign n1110 = n759 ^ n756;
  assign n1111 = n1110 ^ n760;
  assign n1112 = n1111 ^ n757;
  assign n1113 = n760 ^ n757;
  assign n1114 = n760 ^ n756;
  assign n1115 = n1114 ^ n760;
  assign n1116 = n1113 & n1115;
  assign n1117 = n1116 ^ n760;
  assign n1118 = n1112 & ~n1117;
  assign n1119 = n1118 ^ n760;
  assign n1120 = n755 & ~n1119;
  assign n1121 = ~n787 & n805;
  assign n1122 = ~n799 & n1121;
  assign n1123 = n768 & ~n1122;
  assign n1125 = ~n770 & ~n797;
  assign n1124 = ~n782 & ~n799;
  assign n1126 = n1125 ^ n1124;
  assign n1127 = n1124 ^ n789;
  assign n1128 = n1127 ^ n789;
  assign n1129 = n789 ^ n764;
  assign n1130 = ~n1128 & ~n1129;
  assign n1131 = n1130 ^ n789;
  assign n1132 = n1126 & ~n1131;
  assign n1133 = n1132 ^ n1125;
  assign n1134 = ~n766 & n1133;
  assign n1135 = ~n762 & n1134;
  assign n1136 = ~n781 & ~n1135;
  assign n1137 = ~n1123 & ~n1136;
  assign n1138 = ~n1120 & n1137;
  assign n1139 = ~n1109 & n1138;
  assign n1140 = ~n1106 & n1139;
  assign n1141 = n791 ^ n754;
  assign n1142 = n1141 ^ n791;
  assign n1143 = n815 ^ n791;
  assign n1144 = ~n1142 & n1143;
  assign n1145 = n1144 ^ n791;
  assign n1146 = ~n781 & n1145;
  assign n1147 = n1140 & ~n1146;
  assign n1148 = n807 & n1147;
  assign n1149 = n1148 ^ x3;
  assign n1150 = n1149 ^ x73;
  assign n1151 = ~n1104 & n1150;
  assign n1152 = n374 ^ x114;
  assign n1153 = ~n567 & n582;
  assign n1154 = ~n571 & n586;
  assign n1155 = ~n578 & n1154;
  assign n1156 = n543 & ~n1155;
  assign n1157 = ~n1153 & ~n1156;
  assign n1158 = ~n546 & ~n561;
  assign n1159 = ~n535 & n1158;
  assign n1160 = n550 & ~n1159;
  assign n1161 = ~n584 & ~n595;
  assign n1162 = ~n561 & n1161;
  assign n1163 = n538 & ~n1162;
  assign n1164 = ~n1160 & ~n1163;
  assign n1165 = n550 & ~n926;
  assign n1166 = n580 & ~n1165;
  assign n1167 = ~n564 & n1166;
  assign n1168 = n1167 ^ n563;
  assign n1169 = ~n546 & n574;
  assign n1170 = n1169 ^ n1167;
  assign n1171 = n1170 ^ n1169;
  assign n1172 = ~n556 & n926;
  assign n1173 = ~n578 & n1172;
  assign n1174 = n550 & ~n1173;
  assign n1175 = n1174 ^ n1169;
  assign n1176 = ~n1171 & n1175;
  assign n1177 = n1176 ^ n1169;
  assign n1178 = ~n1168 & n1177;
  assign n1179 = n1178 ^ n563;
  assign n1180 = n1164 & ~n1179;
  assign n1181 = n1157 & n1180;
  assign n1182 = n560 & n1181;
  assign n1183 = n548 & n1182;
  assign n1184 = n1183 ^ x61;
  assign n1185 = n1184 ^ x96;
  assign n1186 = ~n1152 & ~n1185;
  assign n1187 = n232 & n256;
  assign n1188 = n209 & ~n281;
  assign n1189 = ~n1187 & ~n1188;
  assign n1190 = n245 & ~n729;
  assign n1191 = ~n263 & n740;
  assign n1192 = n232 & ~n1191;
  assign n1193 = ~n1190 & ~n1192;
  assign n1194 = n218 & ~n731;
  assign n1195 = ~n254 & n280;
  assign n1196 = n209 & ~n1195;
  assign n1197 = ~n224 & ~n238;
  assign n1198 = ~n266 & n1197;
  assign n1199 = ~n228 & n1198;
  assign n1200 = ~n230 & n1199;
  assign n1201 = n213 ^ n212;
  assign n1202 = n1201 ^ n212;
  assign n1203 = n212 ^ n210;
  assign n1204 = n1203 ^ n213;
  assign n1205 = n1204 ^ n212;
  assign n1206 = n1205 ^ n212;
  assign n1207 = ~n1202 & n1206;
  assign n1208 = n1207 ^ n212;
  assign n1209 = ~n211 & ~n1208;
  assign n1210 = n1209 ^ n1204;
  assign n1211 = n228 & n1210;
  assign n1212 = ~n218 & ~n1211;
  assign n1213 = ~n1200 & ~n1212;
  assign n1214 = ~n1196 & ~n1213;
  assign n1215 = ~n1194 & n1214;
  assign n1216 = n1193 & n1215;
  assign n1217 = n252 & n1216;
  assign n1218 = n1189 & n1217;
  assign n1219 = ~n243 & n1218;
  assign n1220 = n1219 ^ x19;
  assign n1221 = n1220 ^ x120;
  assign n1222 = n1186 & n1221;
  assign n1223 = n1151 & n1222;
  assign n1224 = n1152 & ~n1185;
  assign n1225 = n205 ^ x121;
  assign n1226 = n1104 & n1150;
  assign n1227 = ~n1225 & n1226;
  assign n1228 = ~n1104 & ~n1150;
  assign n1229 = n1221 & n1225;
  assign n1230 = n1228 & n1229;
  assign n1231 = ~n1227 & ~n1230;
  assign n1232 = n1224 & ~n1231;
  assign n1233 = ~n1223 & ~n1232;
  assign n1234 = ~n1152 & n1185;
  assign n1235 = ~n1221 & ~n1225;
  assign n1236 = n1150 & n1235;
  assign n1237 = n1225 & n1226;
  assign n1238 = n1229 ^ n1225;
  assign n1239 = ~n1228 & ~n1238;
  assign n1240 = n1239 ^ n1225;
  assign n1241 = ~n1237 & n1240;
  assign n1242 = ~n1236 & n1241;
  assign n1243 = n1234 & n1242;
  assign n1244 = n1151 & n1235;
  assign n1245 = n1104 & ~n1150;
  assign n1246 = n1225 ^ n1221;
  assign n1247 = n1245 & n1246;
  assign n1248 = ~n1221 & n1228;
  assign n1249 = ~n1221 & n1225;
  assign n1250 = n1226 & n1249;
  assign n1251 = ~n1248 & ~n1250;
  assign n1252 = ~n1247 & n1251;
  assign n1253 = ~n1244 & n1252;
  assign n1254 = n1186 & ~n1253;
  assign n1255 = ~n1243 & ~n1254;
  assign n1256 = n1226 & n1229;
  assign n1257 = n1104 & n1235;
  assign n1258 = n1151 & n1246;
  assign n1259 = n1228 & n1235;
  assign n1260 = ~n1258 & ~n1259;
  assign n1261 = ~n1257 & n1260;
  assign n1262 = ~n1256 & n1261;
  assign n1263 = n1224 & ~n1262;
  assign n1264 = n1152 & n1185;
  assign n1265 = n1221 & ~n1225;
  assign n1266 = n1245 & n1265;
  assign n1267 = n1150 ^ n1104;
  assign n1268 = n1229 & ~n1267;
  assign n1269 = ~n1266 & ~n1268;
  assign n1270 = n1251 & n1269;
  assign n1271 = ~n1236 & n1270;
  assign n1272 = n1264 & ~n1271;
  assign n1273 = ~n1263 & ~n1272;
  assign n1274 = n1255 & n1273;
  assign n1275 = n1233 & n1274;
  assign n1276 = n1275 ^ x54;
  assign n1277 = n1276 ^ x77;
  assign n1278 = n404 & ~n427;
  assign n1279 = ~n385 & ~n428;
  assign n1280 = n378 & ~n1279;
  assign n1281 = ~n1278 & ~n1280;
  assign n1282 = ~n376 & n410;
  assign n1283 = ~n405 & n422;
  assign n1284 = ~n398 & n1283;
  assign n1285 = n434 & n1284;
  assign n1286 = n387 & ~n1285;
  assign n1287 = ~n394 & n414;
  assign n1288 = ~n396 & n1287;
  assign n1289 = ~n378 & n1288;
  assign n1290 = n413 & n420;
  assign n1291 = ~n409 & ~n1290;
  assign n1292 = n393 & ~n416;
  assign n1293 = n1291 & n1292;
  assign n1294 = ~n427 & ~n1293;
  assign n1295 = ~n1289 & n1294;
  assign n1296 = ~n385 & ~n395;
  assign n1297 = ~n431 & n1296;
  assign n1298 = n420 & ~n1297;
  assign n1299 = n376 & ~n377;
  assign n1300 = n417 & n1284;
  assign n1301 = ~n410 & n1300;
  assign n1302 = ~n432 & n1301;
  assign n1303 = n1299 & ~n1302;
  assign n1304 = ~n1298 & ~n1303;
  assign n1305 = ~n1295 & n1304;
  assign n1306 = ~n1286 & n1305;
  assign n1307 = ~n1282 & n1306;
  assign n1308 = n1281 & n1307;
  assign n1309 = n1308 ^ x33;
  assign n1310 = n1309 ^ x88;
  assign n1311 = n607 ^ x97;
  assign n1312 = ~n1310 & n1311;
  assign n1313 = ~n787 & ~n797;
  assign n1314 = n755 & ~n1313;
  assign n1315 = n796 & ~n1314;
  assign n1316 = ~n781 & n799;
  assign n1317 = n768 & ~n1313;
  assign n1318 = ~n1316 & ~n1317;
  assign n1319 = n789 & ~n808;
  assign n1320 = ~n804 & ~n814;
  assign n1321 = n755 & ~n1320;
  assign n1322 = n776 & ~n815;
  assign n1323 = ~n803 & n1322;
  assign n1324 = ~n781 & ~n1323;
  assign n1325 = ~n1321 & ~n1324;
  assign n1326 = ~n1319 & n1325;
  assign n1327 = ~n782 & ~n803;
  assign n1328 = ~n791 & n1327;
  assign n1329 = n1328 ^ n822;
  assign n1330 = n1329 ^ n822;
  assign n1331 = n826 & ~n1330;
  assign n1332 = n1331 ^ n822;
  assign n1333 = ~n753 & n1332;
  assign n1334 = n1333 ^ n822;
  assign n1335 = n1326 & ~n1334;
  assign n1336 = n780 & n1335;
  assign n1337 = n1318 & n1336;
  assign n1338 = n1315 & n1337;
  assign n1339 = n1338 ^ x17;
  assign n1340 = n1339 ^ x122;
  assign n1341 = n294 ^ x74;
  assign n1342 = n1340 & n1341;
  assign n1343 = ~n331 & ~n340;
  assign n1344 = n312 & ~n1343;
  assign n1345 = ~n326 & n973;
  assign n1346 = ~n309 & n341;
  assign n1347 = n299 & ~n1346;
  assign n1348 = ~n348 & ~n962;
  assign n1349 = n966 & n1348;
  assign n1350 = n1349 ^ n326;
  assign n1351 = n1350 ^ n1349;
  assign n1352 = n334 & n347;
  assign n1353 = n967 & ~n1352;
  assign n1354 = ~n346 & n1353;
  assign n1355 = ~n335 & n1354;
  assign n1356 = n1355 ^ n1349;
  assign n1357 = ~n1351 & n1356;
  assign n1358 = n1357 ^ n1349;
  assign n1359 = ~n1347 & n1358;
  assign n1360 = ~n372 & n1359;
  assign n1361 = ~n1345 & n1360;
  assign n1362 = ~n1344 & n1361;
  assign n1365 = ~n309 & ~n336;
  assign n1363 = ~n306 & ~n355;
  assign n1364 = ~n339 & n1363;
  assign n1366 = n1365 ^ n1364;
  assign n1367 = n1366 ^ n1365;
  assign n1368 = n1365 ^ n298;
  assign n1369 = n1368 ^ n1365;
  assign n1370 = ~n1367 & ~n1369;
  assign n1371 = n1370 ^ n1365;
  assign n1372 = ~n297 & ~n1371;
  assign n1373 = n1372 ^ n1365;
  assign n1374 = n1362 & n1373;
  assign n1375 = n1374 ^ x9;
  assign n1376 = n1375 ^ x64;
  assign n1377 = n853 & n861;
  assign n1378 = n840 & ~n884;
  assign n1379 = ~n1377 & ~n1378;
  assign n1380 = ~n858 & n867;
  assign n1381 = ~n871 & n877;
  assign n1382 = ~n898 & ~n1081;
  assign n1383 = n853 & ~n1382;
  assign n1384 = ~n882 & ~n891;
  assign n1385 = ~n898 & n1384;
  assign n1386 = ~n847 & n1385;
  assign n1387 = n860 & ~n1386;
  assign n1388 = ~n1383 & ~n1387;
  assign n1389 = n839 ^ n838;
  assign n1391 = n892 & ~n1074;
  assign n1392 = ~n847 & n1391;
  assign n1390 = n893 & ~n1074;
  assign n1393 = n1392 ^ n1390;
  assign n1394 = n1392 ^ n839;
  assign n1395 = n1394 ^ n1392;
  assign n1396 = n1393 & ~n1395;
  assign n1397 = n1396 ^ n1392;
  assign n1398 = ~n1389 & ~n1397;
  assign n1399 = n1388 & ~n1398;
  assign n1400 = n866 & n1399;
  assign n1401 = ~n1381 & n1400;
  assign n1402 = ~n1380 & n1401;
  assign n1403 = n1379 & n1402;
  assign n1404 = n887 ^ n839;
  assign n1405 = n1404 ^ n887;
  assign n1406 = n887 ^ n851;
  assign n1407 = ~n1405 & n1406;
  assign n1408 = n1407 ^ n887;
  assign n1409 = n1389 & ~n1408;
  assign n1410 = n1403 & ~n1409;
  assign n1411 = n1410 ^ x25;
  assign n1412 = n1411 ^ x112;
  assign n1413 = ~n1376 & n1412;
  assign n1414 = n1342 & n1413;
  assign n1415 = n1312 & n1414;
  assign n1416 = n1310 & n1311;
  assign n1417 = ~n1376 & ~n1412;
  assign n1418 = n1340 & ~n1341;
  assign n1419 = n1417 & n1418;
  assign n1420 = ~n1340 & n1341;
  assign n1421 = n1376 & ~n1412;
  assign n1422 = n1420 & n1421;
  assign n1423 = ~n1419 & ~n1422;
  assign n1424 = n1416 & ~n1423;
  assign n1425 = ~n1415 & ~n1424;
  assign n1426 = ~n1310 & ~n1311;
  assign n1427 = n1414 & n1426;
  assign n1428 = ~n1340 & ~n1341;
  assign n1429 = n1417 & n1428;
  assign n1430 = n1416 & n1429;
  assign n1431 = ~n1427 & ~n1430;
  assign n1432 = n1376 & n1412;
  assign n1433 = n1420 & n1432;
  assign n1434 = n1416 & n1433;
  assign n1435 = n1421 & n1428;
  assign n1436 = n1312 & n1435;
  assign n1437 = ~n1434 & ~n1436;
  assign n1438 = n1310 & ~n1311;
  assign n1439 = n1413 & n1420;
  assign n1440 = n1428 & n1432;
  assign n1441 = ~n1439 & ~n1440;
  assign n1442 = n1438 & ~n1441;
  assign n1443 = n1437 & ~n1442;
  assign n1444 = n1413 & n1428;
  assign n1445 = n1416 & n1444;
  assign n1446 = n1418 & n1432;
  assign n1447 = n1312 & n1446;
  assign n1448 = ~n1445 & ~n1447;
  assign n1449 = n1422 & n1438;
  assign n1450 = n1417 & n1420;
  assign n1451 = n1312 & n1450;
  assign n1452 = ~n1449 & ~n1451;
  assign n1453 = n1342 & n1432;
  assign n1454 = n1342 & n1417;
  assign n1455 = ~n1453 & ~n1454;
  assign n1456 = n1416 & ~n1455;
  assign n1457 = ~n1433 & ~n1446;
  assign n1458 = n1342 & n1421;
  assign n1459 = ~n1419 & ~n1458;
  assign n1460 = n1457 & n1459;
  assign n1461 = n1438 & ~n1460;
  assign n1462 = ~n1456 & ~n1461;
  assign n1463 = n1413 & n1418;
  assign n1464 = ~n1439 & ~n1463;
  assign n1465 = ~n1458 & n1464;
  assign n1466 = ~n1440 & n1465;
  assign n1467 = n1466 ^ n1311;
  assign n1468 = n1467 ^ n1466;
  assign n1469 = n1341 ^ n1340;
  assign n1470 = n1469 ^ n1412;
  assign n1471 = n1470 ^ n1376;
  assign n1472 = n1471 ^ n1341;
  assign n1473 = n1472 ^ n1412;
  assign n1474 = n1376 ^ n1341;
  assign n1475 = n1412 ^ n1376;
  assign n1476 = ~n1474 & n1475;
  assign n1477 = n1476 ^ n1376;
  assign n1478 = n1473 & ~n1477;
  assign n1479 = n1478 ^ n1470;
  assign n1480 = ~n1435 & ~n1479;
  assign n1481 = n1480 ^ n1466;
  assign n1482 = ~n1468 & n1481;
  assign n1483 = n1482 ^ n1466;
  assign n1484 = ~n1310 & ~n1483;
  assign n1485 = n1462 & ~n1484;
  assign n1486 = n1452 & n1485;
  assign n1487 = n1429 ^ n1311;
  assign n1488 = n1487 ^ n1429;
  assign n1489 = n1418 & n1421;
  assign n1490 = n1489 ^ n1429;
  assign n1491 = n1488 & n1490;
  assign n1492 = n1491 ^ n1429;
  assign n1493 = n1310 & n1492;
  assign n1494 = n1486 & ~n1493;
  assign n1495 = n1448 & n1494;
  assign n1496 = n1443 & n1495;
  assign n1497 = n1431 & n1496;
  assign n1498 = n1425 & n1497;
  assign n1499 = n1498 ^ x38;
  assign n1500 = n1499 ^ x117;
  assign n1501 = ~n1277 & ~n1500;
  assign n1502 = n512 & n513;
  assign n1503 = ~n468 & ~n504;
  assign n1504 = ~n483 & n1503;
  assign n1505 = n501 & ~n1504;
  assign n1506 = ~n1502 & ~n1505;
  assign n1507 = ~n489 & n501;
  assign n1508 = n470 & n515;
  assign n1509 = ~n1507 & ~n1508;
  assign n1510 = n461 & ~n509;
  assign n1511 = ~n493 & n503;
  assign n1512 = ~n492 & n1511;
  assign n1513 = n512 & ~n1512;
  assign n1514 = ~n1510 & ~n1513;
  assign n1515 = n1509 & n1514;
  assign n1516 = n481 & n1515;
  assign n1517 = n1506 & n1516;
  assign n1518 = n1517 ^ x57;
  assign n1519 = n1518 ^ x86;
  assign n1520 = ~n146 & n170;
  assign n1521 = n131 & ~n192;
  assign n1522 = ~n1520 & ~n1521;
  assign n1523 = n131 & n158;
  assign n1524 = ~n138 & n191;
  assign n1525 = n148 & ~n1524;
  assign n1526 = ~n1523 & ~n1525;
  assign n1527 = n153 & ~n162;
  assign n1528 = n170 & ~n1527;
  assign n1529 = ~n152 & ~n159;
  assign n1530 = n186 & n1529;
  assign n1531 = n156 & ~n1530;
  assign n1532 = ~n1528 & ~n1531;
  assign n1533 = ~n168 & ~n177;
  assign n1534 = n1533 ^ n148;
  assign n1535 = n1533 ^ n156;
  assign n1536 = n1535 ^ n156;
  assign n1537 = n163 ^ n156;
  assign n1538 = n1536 & ~n1537;
  assign n1539 = n1538 ^ n156;
  assign n1540 = ~n1534 & n1539;
  assign n1541 = n1540 ^ n148;
  assign n1542 = n1532 & ~n1541;
  assign n1543 = ~n173 & ~n185;
  assign n1544 = n1543 ^ n182;
  assign n1545 = n1544 ^ n182;
  assign n1546 = n182 ^ n129;
  assign n1547 = n1546 ^ n182;
  assign n1548 = ~n1545 & n1547;
  assign n1549 = n1548 ^ n182;
  assign n1550 = ~n130 & n1549;
  assign n1551 = n1550 ^ n182;
  assign n1552 = n1542 & ~n1551;
  assign n1553 = ~n176 & n1552;
  assign n1554 = n167 & n1553;
  assign n1555 = n1526 & n1554;
  assign n1556 = n1522 & n1555;
  assign n1557 = n1556 ^ x39;
  assign n1558 = n1557 ^ x100;
  assign n1559 = n1519 & ~n1558;
  assign n1560 = ~n339 & n1365;
  assign n1561 = n334 & ~n1560;
  assign n1562 = ~n338 & n967;
  assign n1563 = ~n339 & n1562;
  assign n1564 = n299 & ~n1563;
  assign n1565 = ~n1561 & ~n1564;
  assign n1566 = n324 & n354;
  assign n1567 = ~n340 & n1348;
  assign n1568 = n297 & ~n1567;
  assign n1569 = n332 & n1364;
  assign n1570 = n312 & ~n1569;
  assign n1571 = ~n1568 & ~n1570;
  assign n1572 = ~n1566 & n1571;
  assign n1573 = n1565 & n1572;
  assign n1574 = n957 & n1573;
  assign n1575 = ~n311 & n1574;
  assign n1576 = ~n372 & n1575;
  assign n1577 = n1576 ^ x7;
  assign n1578 = n1577 ^ x110;
  assign n1579 = n764 & n770;
  assign n1580 = n755 & ~n776;
  assign n1581 = ~n1579 & ~n1580;
  assign n1582 = ~n781 & n791;
  assign n1583 = n753 & n803;
  assign n1584 = ~n1582 & ~n1583;
  assign n1585 = ~n804 & n1107;
  assign n1586 = n789 & ~n1585;
  assign n1587 = ~n762 & n1322;
  assign n1588 = n768 & ~n1587;
  assign n1589 = ~n1586 & ~n1588;
  assign n1590 = n1584 & n1589;
  assign n1591 = n1581 & n1590;
  assign n1592 = ~n830 & n1591;
  assign n1593 = n801 & n1592;
  assign n1594 = n785 & n1593;
  assign n1595 = n1318 & n1594;
  assign n1596 = n1315 & n1595;
  assign n1597 = n1596 ^ x23;
  assign n1598 = n1597 ^ x68;
  assign n1599 = ~n1578 & n1598;
  assign n1600 = ~n406 & ~n427;
  assign n1601 = n378 & ~n417;
  assign n1602 = ~n1600 & ~n1601;
  assign n1603 = n378 & n432;
  assign n1604 = n410 & ~n427;
  assign n1605 = ~n1603 & ~n1604;
  assign n1606 = n420 & ~n1292;
  assign n1607 = ~n415 & n422;
  assign n1608 = ~n428 & n1607;
  assign n1609 = n387 & ~n1608;
  assign n1610 = n383 ^ n380;
  assign n1611 = n382 ^ n379;
  assign n1612 = n1611 ^ n380;
  assign n1613 = n1612 ^ n380;
  assign n1614 = n1610 & ~n1613;
  assign n1615 = ~n379 & n1614;
  assign n1616 = n1615 ^ n1612;
  assign n1617 = n1299 & ~n1616;
  assign n1618 = ~n1609 & ~n1617;
  assign n1619 = ~n1606 & n1618;
  assign n1620 = n1605 & n1619;
  assign n1621 = ~n453 & n1620;
  assign n1622 = n402 & n1621;
  assign n1623 = n1602 & n1622;
  assign n1624 = n1623 ^ x31;
  assign n1625 = n1624 ^ x69;
  assign n1626 = n550 & ~n585;
  assign n1627 = n538 & ~n937;
  assign n1628 = ~n1626 & ~n1627;
  assign n1629 = n536 & n556;
  assign n1630 = ~n567 & n578;
  assign n1631 = ~n1629 & ~n1630;
  assign n1632 = ~n541 & ~n584;
  assign n1633 = n543 & ~n1632;
  assign n1634 = ~n578 & n919;
  assign n1635 = n538 & ~n1634;
  assign n1636 = n570 & n937;
  assign n1637 = ~n558 & n1636;
  assign n1638 = ~n568 & n1637;
  assign n1639 = n563 & ~n1638;
  assign n1640 = ~n1635 & ~n1639;
  assign n1641 = ~n571 & n1158;
  assign n1642 = n1641 ^ n582;
  assign n1643 = n1641 ^ n550;
  assign n1644 = n1643 ^ n550;
  assign n1645 = n550 ^ n543;
  assign n1646 = n1644 & ~n1645;
  assign n1647 = n1646 ^ n550;
  assign n1648 = ~n1642 & n1647;
  assign n1649 = n1648 ^ n582;
  assign n1650 = ~n572 & ~n1649;
  assign n1651 = ~n567 & ~n1650;
  assign n1652 = n1640 & ~n1651;
  assign n1653 = ~n562 & n1652;
  assign n1654 = n560 & n1653;
  assign n1655 = ~n1633 & n1654;
  assign n1656 = n1631 & n1655;
  assign n1657 = n1628 & n1656;
  assign n1658 = n555 & n1657;
  assign n1659 = n1658 ^ x15;
  assign n1660 = n1659 ^ x117;
  assign n1661 = ~n1625 & n1660;
  assign n1662 = n1599 & n1661;
  assign n1663 = n1559 & n1662;
  assign n1664 = ~n1519 & ~n1558;
  assign n1665 = ~n1578 & ~n1598;
  assign n1666 = n1625 & n1660;
  assign n1667 = n1665 & n1666;
  assign n1668 = n1664 & n1667;
  assign n1669 = ~n1663 & ~n1668;
  assign n1670 = n1599 & n1666;
  assign n1671 = n1578 & n1598;
  assign n1672 = n1625 & ~n1660;
  assign n1673 = n1671 & n1672;
  assign n1674 = ~n1670 & ~n1673;
  assign n1675 = n1559 & ~n1674;
  assign n1676 = n1661 & n1671;
  assign n1677 = n1559 & n1676;
  assign n1678 = ~n1625 & ~n1660;
  assign n1679 = n1665 & n1678;
  assign n1680 = n1664 & n1679;
  assign n1681 = n1578 & ~n1598;
  assign n1682 = n1678 & n1681;
  assign n1683 = n1559 & n1682;
  assign n1684 = ~n1680 & ~n1683;
  assign n1685 = ~n1519 & n1558;
  assign n1686 = n1666 & n1671;
  assign n1687 = ~n1667 & ~n1686;
  assign n1688 = n1685 & ~n1687;
  assign n1689 = ~n1559 & ~n1685;
  assign n1690 = n1661 & n1681;
  assign n1691 = n1599 & n1678;
  assign n1692 = ~n1690 & ~n1691;
  assign n1693 = n1689 & ~n1692;
  assign n1694 = ~n1682 & ~n1690;
  assign n1695 = ~n1662 & n1694;
  assign n1696 = n1685 & ~n1695;
  assign n1697 = ~n1693 & ~n1696;
  assign n1698 = n1519 & n1558;
  assign n1699 = n1672 & n1681;
  assign n1700 = ~n1670 & ~n1699;
  assign n1701 = n1698 & ~n1700;
  assign n1702 = n1661 & n1665;
  assign n1703 = n1599 & n1672;
  assign n1704 = ~n1699 & ~n1703;
  assign n1705 = ~n1702 & n1704;
  assign n1706 = n1559 & ~n1705;
  assign n1707 = ~n1701 & ~n1706;
  assign n1710 = n1665 & n1672;
  assign n1714 = ~n1673 & ~n1710;
  assign n1708 = n1666 & n1681;
  assign n1709 = n1671 & n1678;
  assign n1711 = ~n1686 & ~n1710;
  assign n1712 = ~n1709 & n1711;
  assign n1713 = ~n1708 & n1712;
  assign n1715 = n1714 ^ n1713;
  assign n1716 = n1715 ^ n1714;
  assign n1717 = n1714 ^ n1519;
  assign n1718 = n1717 ^ n1714;
  assign n1719 = ~n1716 & ~n1718;
  assign n1720 = n1719 ^ n1714;
  assign n1721 = ~n1558 & ~n1720;
  assign n1722 = n1721 ^ n1714;
  assign n1723 = n1707 & n1722;
  assign n1724 = n1697 & n1723;
  assign n1725 = ~n1688 & n1724;
  assign n1726 = n1684 & n1725;
  assign n1727 = ~n1677 & n1726;
  assign n1728 = ~n1675 & n1727;
  assign n1729 = n1669 & n1728;
  assign n1730 = n1709 ^ n1519;
  assign n1731 = n1730 ^ n1709;
  assign n1732 = ~n1676 & ~n1702;
  assign n1733 = n1732 ^ n1709;
  assign n1734 = n1731 & ~n1733;
  assign n1735 = n1734 ^ n1709;
  assign n1736 = n1558 & n1735;
  assign n1737 = n1729 & ~n1736;
  assign n1738 = n1737 ^ x46;
  assign n1739 = n1738 ^ x102;
  assign n1740 = n917 ^ x126;
  assign n1741 = n1149 ^ x77;
  assign n1742 = ~n1740 & ~n1741;
  assign n1743 = n719 ^ x92;
  assign n1744 = n1184 ^ x83;
  assign n1745 = ~n1743 & ~n1744;
  assign n1746 = ~n376 & n421;
  assign n1747 = ~n432 & n1292;
  assign n1748 = n387 & ~n1747;
  assign n1749 = ~n1746 & ~n1748;
  assign n1750 = ~n385 & n411;
  assign n1751 = n417 & n1750;
  assign n1752 = n420 & ~n1751;
  assign n1753 = n400 & n433;
  assign n1754 = ~n413 & n1753;
  assign n1755 = ~n410 & n1754;
  assign n1756 = n1299 & ~n1755;
  assign n1757 = ~n1752 & ~n1756;
  assign n1758 = n1749 & n1757;
  assign n1759 = n428 ^ n393;
  assign n1760 = n1759 ^ n428;
  assign n1761 = n428 ^ n376;
  assign n1762 = n1761 ^ n428;
  assign n1763 = ~n1760 & ~n1762;
  assign n1764 = n1763 ^ n428;
  assign n1765 = ~n377 & n1764;
  assign n1766 = n1765 ^ n428;
  assign n1767 = n1758 & ~n1766;
  assign n1768 = n408 & n1767;
  assign n1769 = n1602 & n1768;
  assign n1770 = n1769 ^ x45;
  assign n1771 = n1770 ^ x109;
  assign n1772 = n131 & n177;
  assign n1773 = ~n157 & ~n1772;
  assign n1774 = n170 & n181;
  assign n1775 = n145 & n148;
  assign n1776 = ~n1774 & ~n1775;
  assign n1777 = ~n151 & ~n163;
  assign n1778 = ~n185 & n1777;
  assign n1779 = n131 & ~n1778;
  assign n1781 = n160 & n186;
  assign n1780 = n164 & n1529;
  assign n1782 = n1781 ^ n1780;
  assign n1783 = n130 ^ n129;
  assign n1784 = n1783 ^ n129;
  assign n1785 = n1780 ^ n129;
  assign n1786 = ~n1784 & ~n1785;
  assign n1787 = n1786 ^ n129;
  assign n1788 = n1782 & ~n1787;
  assign n1789 = n1788 ^ n1781;
  assign n1790 = n1543 & n1789;
  assign n1791 = ~n142 & n1790;
  assign n1792 = n1791 ^ n129;
  assign n1793 = n1792 ^ n1791;
  assign n1794 = ~n168 & ~n182;
  assign n1795 = n1794 ^ n1791;
  assign n1796 = n1795 ^ n1791;
  assign n1797 = ~n1793 & ~n1796;
  assign n1798 = n1797 ^ n1791;
  assign n1799 = ~n130 & ~n1798;
  assign n1800 = n1799 ^ n1791;
  assign n1801 = ~n1779 & n1800;
  assign n1802 = n1776 & n1801;
  assign n1803 = n1773 & n1802;
  assign n1804 = n155 & n1803;
  assign n1805 = n1526 & n1804;
  assign n1806 = ~n139 & n1805;
  assign n1807 = n1806 ^ x53;
  assign n1808 = n1807 ^ x94;
  assign n1809 = n1771 & ~n1808;
  assign n1810 = n1745 & n1809;
  assign n1811 = n1742 & n1810;
  assign n1812 = ~n1740 & n1741;
  assign n1813 = ~n1771 & ~n1808;
  assign n1814 = n1745 & n1813;
  assign n1815 = n1743 & ~n1744;
  assign n1816 = n1809 & n1815;
  assign n1817 = ~n1814 & ~n1816;
  assign n1818 = n1812 & ~n1817;
  assign n1819 = ~n1811 & ~n1818;
  assign n1820 = n1813 & n1815;
  assign n1821 = ~n1743 & n1744;
  assign n1822 = n1809 & n1821;
  assign n1823 = ~n1820 & ~n1822;
  assign n1824 = n1812 & ~n1823;
  assign n1825 = n1740 & ~n1741;
  assign n1826 = ~n1771 & n1808;
  assign n1827 = n1815 & n1826;
  assign n1828 = n1771 & n1808;
  assign n1829 = n1745 & n1828;
  assign n1830 = ~n1827 & ~n1829;
  assign n1831 = n1817 & n1830;
  assign n1832 = n1825 & ~n1831;
  assign n1833 = ~n1824 & ~n1832;
  assign n1834 = n1740 & n1741;
  assign n1835 = n1743 & n1744;
  assign n1836 = n1809 & n1835;
  assign n1837 = n1821 & n1826;
  assign n1838 = n1828 & n1835;
  assign n1839 = ~n1822 & ~n1838;
  assign n1840 = ~n1837 & n1839;
  assign n1841 = ~n1836 & n1840;
  assign n1842 = n1834 & ~n1841;
  assign n1843 = n1815 & n1828;
  assign n1844 = ~n1814 & ~n1843;
  assign n1845 = ~n1827 & n1844;
  assign n1846 = n1742 & ~n1845;
  assign n1847 = n1821 & n1828;
  assign n1848 = n1826 & n1835;
  assign n1849 = ~n1847 & ~n1848;
  assign n1850 = n1812 & ~n1849;
  assign n1851 = n1813 & n1821;
  assign n1852 = ~n1837 & ~n1851;
  assign n1853 = n1742 & ~n1852;
  assign n1854 = n1745 & n1826;
  assign n1855 = ~n1820 & ~n1829;
  assign n1856 = ~n1854 & n1855;
  assign n1857 = n1834 & ~n1856;
  assign n1858 = ~n1812 & ~n1825;
  assign n1859 = n1812 & n1836;
  assign n1860 = ~n1836 & ~n1838;
  assign n1861 = ~n1825 & n1860;
  assign n1862 = n1813 & n1835;
  assign n1863 = ~n1838 & n1852;
  assign n1864 = ~n1862 & n1863;
  assign n1865 = ~n1861 & ~n1864;
  assign n1866 = ~n1859 & ~n1865;
  assign n1867 = ~n1858 & ~n1866;
  assign n1868 = ~n1857 & ~n1867;
  assign n1869 = ~n1853 & n1868;
  assign n1870 = n1741 ^ n1740;
  assign n1871 = n1827 ^ n1741;
  assign n1872 = n1871 ^ n1827;
  assign n1873 = ~n1836 & ~n1862;
  assign n1874 = n1873 ^ n1827;
  assign n1875 = ~n1872 & ~n1874;
  assign n1876 = n1875 ^ n1827;
  assign n1877 = ~n1870 & n1876;
  assign n1878 = n1869 & ~n1877;
  assign n1879 = ~n1850 & n1878;
  assign n1880 = ~n1846 & n1879;
  assign n1881 = ~n1842 & n1880;
  assign n1882 = n1833 & n1881;
  assign n1883 = n1819 & n1882;
  assign n1884 = n1883 ^ x62;
  assign n1885 = n1884 ^ x91;
  assign n1886 = n1739 & n1885;
  assign n1887 = n1501 & n1886;
  assign n1888 = ~n1739 & ~n1885;
  assign n1889 = n1501 & n1888;
  assign n1890 = ~n1277 & n1500;
  assign n1891 = ~n1739 & n1885;
  assign n1892 = n1890 & n1891;
  assign n1893 = n1277 & ~n1500;
  assign n1894 = n1886 & n1893;
  assign n1895 = ~n1892 & ~n1894;
  assign n1896 = n1891 & n1893;
  assign n1897 = n1277 & n1500;
  assign n1898 = n1739 & ~n1885;
  assign n1899 = n1897 & n1898;
  assign n1900 = ~n1896 & ~n1899;
  assign n1901 = n1895 & n1900;
  assign n1902 = ~n1889 & n1901;
  assign n1903 = ~n1887 & n1902;
  assign n1904 = n1072 & ~n1903;
  assign n1905 = ~n681 & n1071;
  assign n1906 = n1890 & n1898;
  assign n1907 = n1501 & n1891;
  assign n1908 = n1891 & n1897;
  assign n1909 = ~n1887 & ~n1908;
  assign n1910 = ~n1907 & n1909;
  assign n1911 = n1888 & n1890;
  assign n1912 = n1893 & n1898;
  assign n1913 = ~n1911 & ~n1912;
  assign n1914 = n1910 & n1913;
  assign n1915 = ~n1906 & n1914;
  assign n1916 = n1905 & ~n1915;
  assign n1917 = ~n681 & ~n1071;
  assign n1918 = n1886 & n1890;
  assign n1919 = n1501 & n1898;
  assign n1920 = n1888 & n1897;
  assign n1921 = ~n1919 & ~n1920;
  assign n1922 = n1895 & n1921;
  assign n1923 = ~n1918 & n1922;
  assign n1924 = n1913 & n1923;
  assign n1925 = ~n1896 & n1924;
  assign n1926 = n1917 & ~n1925;
  assign n1927 = ~n1916 & ~n1926;
  assign n1928 = ~n1904 & n1927;
  assign n1929 = n1500 ^ n1277;
  assign n1930 = n1929 ^ n1885;
  assign n1931 = n1930 ^ n1500;
  assign n1932 = n1931 ^ n1739;
  assign n1933 = n1932 ^ n1885;
  assign n1934 = n1739 ^ n1500;
  assign n1935 = n1934 ^ n1500;
  assign n1936 = n1885 ^ n1500;
  assign n1937 = ~n1935 & n1936;
  assign n1938 = n1937 ^ n1500;
  assign n1939 = n1933 & n1938;
  assign n1940 = n1939 ^ n1930;
  assign n1941 = n1940 ^ n1921;
  assign n1942 = n1941 ^ n1921;
  assign n1943 = n1921 ^ n681;
  assign n1944 = n1943 ^ n1921;
  assign n1945 = n1942 & n1944;
  assign n1946 = n1945 ^ n1921;
  assign n1947 = ~n1071 & ~n1946;
  assign n1948 = n1947 ^ n1921;
  assign n1949 = n1928 & n1948;
  assign n1950 = n1949 ^ n374;
  assign n1951 = n1950 ^ x82;
  assign n1952 = n836 ^ x116;
  assign n1953 = n1624 ^ x75;
  assign n1954 = ~n1952 & n1953;
  assign n1955 = n461 & ~n706;
  assign n1956 = n501 & ~n690;
  assign n1957 = ~n1955 & ~n1956;
  assign n1958 = n470 & ~n688;
  assign n1959 = ~n473 & n694;
  assign n1960 = ~n483 & n1959;
  assign n1961 = n512 & ~n1960;
  assign n1962 = ~n1958 & ~n1961;
  assign n1963 = n1957 & n1962;
  assign n1964 = n1506 & n1963;
  assign n1965 = n1964 ^ x55;
  assign n1966 = n1965 ^ x93;
  assign n1967 = n1557 ^ x70;
  assign n1968 = ~n1966 & ~n1967;
  assign n1969 = ~n864 & n867;
  assign n1970 = n892 & n1082;
  assign n1971 = n884 & n1970;
  assign n1972 = n853 & ~n1971;
  assign n1973 = ~n1969 & ~n1972;
  assign n1974 = n858 & n1390;
  assign n1975 = n860 & ~n1974;
  assign n1976 = n1079 & ~n1081;
  assign n1977 = ~n867 & n1976;
  assign n1978 = ~n857 & ~n898;
  assign n1979 = n887 & n1978;
  assign n1980 = ~n840 & n1979;
  assign n1981 = ~n1977 & ~n1980;
  assign n1982 = n1075 & ~n1981;
  assign n1983 = ~n871 & ~n1982;
  assign n1984 = ~n1975 & ~n1983;
  assign n1985 = n1973 & n1984;
  assign n1986 = ~n1409 & n1985;
  assign n1987 = ~n852 & n1986;
  assign n1988 = n1987 ^ x47;
  assign n1989 = n1988 ^ x118;
  assign n1990 = n750 ^ x76;
  assign n1991 = ~n1989 & n1990;
  assign n1992 = n1968 & n1991;
  assign n1993 = n1966 & n1967;
  assign n1994 = n1991 & n1993;
  assign n1995 = ~n1992 & ~n1994;
  assign n1996 = n1954 & ~n1995;
  assign n1997 = n1952 & n1953;
  assign n1998 = n1989 & n1990;
  assign n1999 = n1968 & n1998;
  assign n2000 = ~n1966 & n1967;
  assign n2001 = n1991 & n2000;
  assign n2002 = ~n1999 & ~n2001;
  assign n2003 = n1997 & ~n2002;
  assign n2004 = ~n1996 & ~n2003;
  assign n2005 = ~n1989 & ~n1990;
  assign n2006 = n1968 & n2005;
  assign n2007 = n1997 & n2006;
  assign n2008 = n1989 & ~n1990;
  assign n2009 = n1968 & n2008;
  assign n2010 = n1954 & n2009;
  assign n2011 = ~n2007 & ~n2010;
  assign n2012 = n1966 & ~n1967;
  assign n2013 = n1998 & n2012;
  assign n2014 = ~n1994 & ~n2013;
  assign n2015 = n1997 & ~n2014;
  assign n2016 = n1952 & ~n1953;
  assign n2017 = ~n1997 & ~n2016;
  assign n2018 = n2000 & n2005;
  assign n2019 = n2005 & n2012;
  assign n2020 = ~n2018 & ~n2019;
  assign n2021 = ~n2017 & ~n2020;
  assign n2022 = ~n2015 & ~n2021;
  assign n2023 = ~n1952 & ~n1953;
  assign n2024 = n1967 ^ n1966;
  assign n2025 = n2024 ^ n1990;
  assign n2026 = n2025 ^ n1967;
  assign n2027 = n2026 ^ n1989;
  assign n2028 = n2027 ^ n1990;
  assign n2029 = n1990 ^ n1967;
  assign n2030 = n1989 ^ n1967;
  assign n2031 = n2030 ^ n1967;
  assign n2032 = n2029 & ~n2031;
  assign n2033 = n2032 ^ n1967;
  assign n2034 = n2028 & n2033;
  assign n2035 = n2034 ^ n2025;
  assign n2036 = n2023 & n2035;
  assign n2037 = n1998 & n2000;
  assign n2038 = ~n2013 & ~n2037;
  assign n2039 = n1993 & n2005;
  assign n2040 = ~n2006 & ~n2039;
  assign n2041 = n2038 & n2040;
  assign n2042 = n1954 & ~n2041;
  assign n2043 = ~n2009 & n2038;
  assign n2044 = ~n2039 & n2043;
  assign n2045 = ~n2001 & n2044;
  assign n2046 = ~n1992 & n2045;
  assign n2047 = n2016 & ~n2046;
  assign n2048 = ~n2042 & ~n2047;
  assign n2049 = ~n2036 & n2048;
  assign n2050 = n2022 & n2049;
  assign n2051 = n2011 & n2050;
  assign n2052 = n2004 & n2051;
  assign n2053 = n1993 & n2008;
  assign n2054 = n2053 ^ n1952;
  assign n2055 = n2054 ^ n2053;
  assign n2056 = n2000 & n2008;
  assign n2057 = n2056 ^ n2053;
  assign n2058 = n2055 & n2057;
  assign n2059 = n2058 ^ n2053;
  assign n2060 = n1953 & n2059;
  assign n2061 = n2052 & ~n2060;
  assign n2062 = n2061 ^ x6;
  assign n2063 = n2062 ^ x114;
  assign n2064 = n1685 & n1708;
  assign n2065 = n1698 & ~n1704;
  assign n2066 = n1664 & ~n1714;
  assign n2067 = ~n2065 & ~n2066;
  assign n2068 = ~n1691 & ~n1708;
  assign n2069 = ~n1710 & n2068;
  assign n2070 = n1559 & ~n2069;
  assign n2071 = ~n1679 & ~n1682;
  assign n2072 = ~n1703 & n2071;
  assign n2073 = n1685 & ~n2072;
  assign n2074 = ~n2070 & ~n2073;
  assign n2075 = n2067 & n2074;
  assign n2076 = n1664 & n1709;
  assign n2077 = n1698 & n1702;
  assign n2078 = n1558 ^ n1519;
  assign n2079 = ~n1695 & ~n2078;
  assign n2080 = ~n2077 & ~n2079;
  assign n2081 = ~n2076 & n2080;
  assign n2082 = ~n1670 & ~n1686;
  assign n2083 = n2082 ^ n1689;
  assign n2084 = n2083 ^ n2082;
  assign n2085 = ~n1702 & ~n1709;
  assign n2086 = n2085 ^ n2082;
  assign n2087 = ~n2084 & n2086;
  assign n2088 = n2087 ^ n2082;
  assign n2089 = n2081 & n2088;
  assign n2090 = n2075 & n2089;
  assign n2091 = ~n1688 & n2090;
  assign n2092 = ~n1677 & n2091;
  assign n2093 = ~n2064 & n2092;
  assign n2094 = ~n1675 & n2093;
  assign n2095 = n2094 ^ x24;
  assign n2096 = n2095 ^ x121;
  assign n2097 = n2063 & ~n2096;
  assign n2098 = n1151 & n1249;
  assign n2099 = ~n1150 & n1246;
  assign n2100 = n1224 & n2099;
  assign n2101 = n1225 & n1245;
  assign n2102 = ~n1151 & n1235;
  assign n2103 = ~n2101 & ~n2102;
  assign n2104 = n1186 & ~n2103;
  assign n2105 = ~n2100 & ~n2104;
  assign n2106 = n1151 & n1225;
  assign n2107 = n1246 ^ n1245;
  assign n2108 = n2107 ^ n1246;
  assign n2109 = n1246 ^ n1229;
  assign n2110 = ~n2108 & n2109;
  assign n2111 = n2110 ^ n1246;
  assign n2112 = ~n2106 & ~n2111;
  assign n2113 = ~n1236 & n2112;
  assign n2114 = n2113 ^ n1152;
  assign n2115 = n2114 ^ n2113;
  assign n2116 = n1225 ^ n1104;
  assign n2117 = n2116 ^ n1221;
  assign n2118 = n2117 ^ n1104;
  assign n2119 = n2118 ^ n1150;
  assign n2120 = n2119 ^ n1221;
  assign n2121 = n1221 ^ n1104;
  assign n2122 = n1267 ^ n1104;
  assign n2123 = ~n2121 & ~n2122;
  assign n2124 = n2123 ^ n1104;
  assign n2125 = ~n2120 & n2124;
  assign n2126 = n2125 ^ n2117;
  assign n2127 = n2126 ^ n2113;
  assign n2128 = n2115 & ~n2127;
  assign n2129 = n2128 ^ n2113;
  assign n2130 = n1185 & ~n2129;
  assign n2131 = n2105 & ~n2130;
  assign n2132 = ~n2098 & n2131;
  assign n2133 = n1233 & n2132;
  assign n2134 = n2133 ^ x56;
  assign n2135 = n2134 ^ x90;
  assign n2136 = n1001 & n1026;
  assign n2137 = n1011 & n1047;
  assign n2138 = ~n2136 & ~n2137;
  assign n2139 = ~n1024 & ~n1045;
  assign n2140 = n1011 & ~n2139;
  assign n2141 = n999 & n1042;
  assign n2142 = n752 & ~n2141;
  assign n2143 = ~n1024 & ~n1053;
  assign n2144 = n720 & ~n2143;
  assign n2145 = ~n2142 & ~n2144;
  assign n2146 = ~n995 & ~n1034;
  assign n2147 = ~n1016 & n2146;
  assign n2148 = ~n1031 & n2147;
  assign n2149 = n1011 & ~n2148;
  assign n2150 = ~n998 & ~n1035;
  assign n2151 = n1055 & n2150;
  assign n2152 = n1019 & ~n2151;
  assign n2153 = n1001 & ~n1037;
  assign n2154 = n1007 & ~n1031;
  assign n2155 = n1012 & ~n2154;
  assign n2156 = ~n2153 & ~n2155;
  assign n2157 = n1052 ^ n752;
  assign n2158 = n1052 ^ n1011;
  assign n2159 = n2158 ^ n1011;
  assign n2160 = n1047 ^ n1011;
  assign n2161 = ~n2159 & ~n2160;
  assign n2162 = n2161 ^ n1011;
  assign n2163 = n2157 & n2162;
  assign n2164 = n2163 ^ n752;
  assign n2165 = n2156 & ~n2164;
  assign n2166 = ~n2152 & n2165;
  assign n2167 = ~n2149 & n2166;
  assign n2168 = n2145 & n2167;
  assign n2169 = ~n2140 & n2168;
  assign n2170 = n2138 & n2169;
  assign n2171 = n2170 ^ x32;
  assign n2172 = n2171 ^ x88;
  assign n2173 = ~n2135 & n2172;
  assign n2174 = n1416 & n1450;
  assign n2175 = ~n1435 & ~n1458;
  assign n2176 = n1438 & ~n2175;
  assign n2177 = ~n2174 & ~n2176;
  assign n2178 = ~n1414 & ~n1446;
  assign n2179 = n1438 & ~n2178;
  assign n2180 = ~n1433 & ~n1440;
  assign n2181 = n1426 & ~n2180;
  assign n2182 = ~n2179 & ~n2181;
  assign n2183 = n1438 & n1453;
  assign n2184 = n1416 & n1440;
  assign n2185 = ~n2183 & ~n2184;
  assign n2186 = n1310 & n1433;
  assign n2187 = n1438 & n1450;
  assign n2188 = ~n2186 & ~n2187;
  assign n2189 = n1312 & n1479;
  assign n2190 = n1459 & ~n1463;
  assign n2191 = n1416 & ~n2190;
  assign n2192 = ~n1429 & ~n1454;
  assign n2193 = ~n1453 & n2192;
  assign n2194 = n1464 & ~n1489;
  assign n2195 = n2193 & n2194;
  assign n2196 = n1426 & ~n2195;
  assign n2197 = ~n2191 & ~n2196;
  assign n2198 = ~n2189 & n2197;
  assign n2199 = n2188 & n2198;
  assign n2200 = ~n1415 & n2199;
  assign n2201 = n2185 & n2200;
  assign n2202 = ~n1493 & n2201;
  assign n2203 = n1448 & n2202;
  assign n2204 = n2182 & n2203;
  assign n2205 = n2177 & n2204;
  assign n2206 = n2205 ^ x48;
  assign n2207 = n2206 ^ x73;
  assign n2208 = n1816 & n1834;
  assign n2209 = n1812 & n1862;
  assign n2210 = ~n2208 & ~n2209;
  assign n2211 = n1825 & ~n1873;
  assign n2212 = n2210 & ~n2211;
  assign n2213 = n1834 & n1854;
  assign n2214 = n1825 & n1827;
  assign n2215 = ~n2213 & ~n2214;
  assign n2216 = n1742 & ~n1839;
  assign n2217 = ~n1810 & ~n1848;
  assign n2218 = ~n1837 & n2217;
  assign n2219 = n1825 & ~n2218;
  assign n2220 = ~n2216 & ~n2219;
  assign n2221 = n1834 & n1843;
  assign n2222 = ~n1851 & ~n1854;
  assign n2223 = ~n1836 & n2222;
  assign n2224 = n1812 & ~n2223;
  assign n2225 = ~n1855 & ~n1858;
  assign n2226 = ~n1847 & ~n1851;
  assign n2227 = n1839 & n2226;
  assign n2228 = n1834 & ~n2227;
  assign n2229 = ~n1820 & n1844;
  assign n2230 = ~n1854 & n2229;
  assign n2231 = n1742 & ~n2230;
  assign n2232 = ~n2228 & ~n2231;
  assign n2233 = ~n2225 & n2232;
  assign n2234 = ~n2224 & n2233;
  assign n2235 = ~n2221 & n2234;
  assign n2236 = n2220 & n2235;
  assign n2237 = n2215 & n2236;
  assign n2238 = n2212 & n2237;
  assign n2239 = ~n1877 & n2238;
  assign n2240 = ~n1850 & n2239;
  assign n2241 = n2240 ^ x40;
  assign n2242 = n2241 ^ x99;
  assign n2243 = ~n2207 & n2242;
  assign n2244 = n2173 & n2243;
  assign n2245 = n2097 & n2244;
  assign n2246 = ~n2063 & n2096;
  assign n2247 = n2207 & ~n2242;
  assign n2248 = n2173 & n2247;
  assign n2249 = n2246 & n2248;
  assign n2250 = n2135 & ~n2172;
  assign n2251 = ~n2207 & ~n2242;
  assign n2252 = n2250 & n2251;
  assign n2253 = n2097 & n2252;
  assign n2254 = ~n2249 & ~n2253;
  assign n2255 = n2135 & n2172;
  assign n2256 = n2247 & n2255;
  assign n2257 = n2097 & n2256;
  assign n2258 = n2207 & n2242;
  assign n2259 = n2255 & n2258;
  assign n2260 = n2250 & n2258;
  assign n2261 = ~n2259 & ~n2260;
  assign n2262 = ~n2135 & ~n2172;
  assign n2263 = n2247 & n2262;
  assign n2264 = n2173 & n2251;
  assign n2265 = ~n2263 & ~n2264;
  assign n2266 = n2261 & n2265;
  assign n2267 = n2063 & ~n2266;
  assign n2268 = n2247 & n2250;
  assign n2269 = n2251 & n2255;
  assign n2270 = ~n2268 & ~n2269;
  assign n2271 = ~n2260 & n2270;
  assign n2272 = ~n2256 & n2271;
  assign n2273 = n2246 & ~n2272;
  assign n2274 = n2063 & n2096;
  assign n2275 = n2243 & n2255;
  assign n2276 = n2173 & n2258;
  assign n2277 = n2251 & n2262;
  assign n2278 = ~n2276 & ~n2277;
  assign n2279 = ~n2275 & n2278;
  assign n2280 = ~n2252 & n2279;
  assign n2281 = n2274 & ~n2280;
  assign n2282 = n2243 & n2250;
  assign n2283 = n2282 ^ n2063;
  assign n2286 = n2243 & n2262;
  assign n2287 = ~n2276 & ~n2286;
  assign n2284 = n2242 & n2255;
  assign n2285 = ~n2268 & ~n2284;
  assign n2288 = n2287 ^ n2285;
  assign n2289 = n2287 ^ n2096;
  assign n2290 = n2289 ^ n2287;
  assign n2291 = n2288 & ~n2290;
  assign n2292 = n2291 ^ n2287;
  assign n2293 = n2292 ^ n2282;
  assign n2294 = n2283 & ~n2293;
  assign n2295 = n2294 ^ n2291;
  assign n2296 = n2295 ^ n2287;
  assign n2297 = n2296 ^ n2063;
  assign n2298 = ~n2282 & ~n2297;
  assign n2299 = n2298 ^ n2282;
  assign n2300 = n2299 ^ n2063;
  assign n2301 = ~n2281 & ~n2300;
  assign n2302 = ~n2273 & n2301;
  assign n2303 = ~n2267 & n2302;
  assign n2304 = ~n2063 & ~n2096;
  assign n2305 = n2304 ^ n2248;
  assign n2306 = n2248 ^ n2097;
  assign n2307 = n2306 ^ n2097;
  assign n2308 = n2258 & n2262;
  assign n2309 = n2265 & ~n2308;
  assign n2310 = n2309 ^ n2097;
  assign n2311 = ~n2307 & n2310;
  assign n2312 = n2311 ^ n2097;
  assign n2313 = n2305 & n2312;
  assign n2314 = n2313 ^ n2304;
  assign n2315 = n2303 & ~n2314;
  assign n2316 = ~n2257 & n2315;
  assign n2317 = n2254 & n2316;
  assign n2318 = ~n2245 & n2317;
  assign n2319 = n2318 ^ n1184;
  assign n2320 = n2319 ^ x64;
  assign n2321 = n1951 & ~n2320;
  assign n2322 = n2134 ^ x70;
  assign n2323 = n1499 ^ x84;
  assign n2324 = ~n2322 & ~n2323;
  assign n2325 = n2062 ^ x94;
  assign n2326 = n1070 ^ x116;
  assign n2327 = ~n2325 & n2326;
  assign n2328 = n296 & n652;
  assign n2329 = n617 & n630;
  assign n2330 = ~n2328 & ~n2329;
  assign n2331 = n630 & ~n649;
  assign n2332 = ~n643 & ~n648;
  assign n2333 = n616 & ~n2332;
  assign n2334 = n617 & n625;
  assign n2335 = n634 & n640;
  assign n2336 = n625 & ~n2335;
  assign n2337 = n625 & n648;
  assign n2338 = ~n631 & ~n654;
  assign n2339 = ~n639 & n2338;
  assign n2340 = n630 & ~n2339;
  assign n2341 = ~n2337 & ~n2340;
  assign n2342 = n662 & n2341;
  assign n2343 = ~n2336 & n2342;
  assign n2344 = ~n623 & ~n633;
  assign n2345 = n667 ^ n640;
  assign n2346 = n667 ^ n616;
  assign n2347 = n2346 ^ n616;
  assign n2348 = n616 ^ n296;
  assign n2349 = n2347 & ~n2348;
  assign n2350 = n2349 ^ n616;
  assign n2351 = n2345 & n2350;
  assign n2352 = n2351 ^ n640;
  assign n2353 = n2344 & n2352;
  assign n2354 = n651 & ~n2353;
  assign n2355 = n2343 & ~n2354;
  assign n2356 = ~n2334 & n2355;
  assign n2357 = ~n2333 & n2356;
  assign n2358 = ~n2331 & n2357;
  assign n2359 = n620 & n2358;
  assign n2360 = n2330 & n2359;
  assign n2361 = ~n659 & n2360;
  assign n2362 = n2361 ^ x22;
  assign n2363 = n2362 ^ x83;
  assign n2364 = n1577 ^ x65;
  assign n2365 = n1411 ^ x72;
  assign n2366 = n2364 & n2365;
  assign n2367 = n1309 ^ x104;
  assign n2368 = n218 & n267;
  assign n2369 = ~n230 & n279;
  assign n2370 = ~n729 & ~n2369;
  assign n2371 = n225 & n264;
  assign n2372 = n274 & n2371;
  assign n2373 = ~n245 & n2372;
  assign n2374 = n228 & ~n2373;
  assign n2375 = ~n235 & ~n254;
  assign n2376 = n2375 ^ n207;
  assign n2377 = n2376 ^ n2375;
  assign n2378 = n257 & ~n261;
  assign n2379 = n2378 ^ n2375;
  assign n2380 = ~n2377 & n2379;
  assign n2381 = n2380 ^ n2375;
  assign n2382 = n208 & ~n2381;
  assign n2383 = ~n2374 & ~n2382;
  assign n2384 = ~n2370 & n2383;
  assign n2385 = ~n2368 & n2384;
  assign n2386 = n722 & n2385;
  assign n2387 = n227 & n2386;
  assign n2388 = n1189 & n2387;
  assign n2389 = ~n243 & n2388;
  assign n2390 = n2389 ^ x41;
  assign n2391 = n2390 ^ x115;
  assign n2392 = ~n2367 & ~n2391;
  assign n2393 = n1518 ^ x106;
  assign n2394 = n156 & n168;
  assign n2395 = ~n174 & ~n185;
  assign n2396 = ~n190 & ~n2395;
  assign n2397 = ~n2394 & ~n2396;
  assign n2398 = n131 & ~n160;
  assign n2399 = ~n151 & ~n158;
  assign n2400 = n170 & ~n2399;
  assign n2401 = n160 & ~n162;
  assign n2402 = ~n182 & n2401;
  assign n2403 = ~n148 & n2402;
  assign n2404 = ~n156 & ~n159;
  assign n2405 = ~n2402 & ~n2404;
  assign n2406 = ~n177 & ~n2405;
  assign n2407 = n186 & n2406;
  assign n2408 = ~n2403 & ~n2407;
  assign n2409 = ~n190 & n2408;
  assign n2410 = ~n2400 & ~n2409;
  assign n2411 = ~n2398 & n2410;
  assign n2412 = n2397 & n2411;
  assign n2413 = n1776 & n2412;
  assign n2414 = n180 & n2413;
  assign n2415 = n1773 & n2414;
  assign n2416 = n172 & n2415;
  assign n2417 = n1522 & n2416;
  assign n2418 = ~n139 & n2417;
  assign n2419 = n2418 ^ x49;
  assign n2420 = n2419 ^ x89;
  assign n2421 = ~n2393 & n2420;
  assign n2422 = n2392 & n2421;
  assign n2423 = n2393 & ~n2420;
  assign n2424 = n2392 & n2423;
  assign n2425 = ~n2422 & ~n2424;
  assign n2426 = n2366 & ~n2425;
  assign n2427 = n2364 & ~n2365;
  assign n2428 = n2367 & n2391;
  assign n2429 = ~n2393 & ~n2420;
  assign n2430 = n2428 & n2429;
  assign n2431 = n2427 & n2430;
  assign n2432 = n2421 & n2428;
  assign n2433 = n2366 & n2432;
  assign n2434 = ~n2364 & ~n2365;
  assign n2435 = n2422 & n2434;
  assign n2436 = ~n2364 & n2365;
  assign n2437 = n2393 & n2420;
  assign n2438 = n2392 & n2437;
  assign n2439 = n2367 & ~n2391;
  assign n2440 = n2423 & n2439;
  assign n2441 = ~n2438 & ~n2440;
  assign n2442 = n2436 & ~n2441;
  assign n2443 = ~n2435 & ~n2442;
  assign n2444 = ~n2367 & n2391;
  assign n2445 = n2423 & n2444;
  assign n2446 = n2366 & n2445;
  assign n2447 = n2365 ^ n2364;
  assign n2448 = n2424 ^ n2365;
  assign n2449 = n2448 ^ n2424;
  assign n2450 = n2421 & n2439;
  assign n2451 = ~n2422 & ~n2450;
  assign n2452 = n2451 ^ n2424;
  assign n2453 = n2449 & ~n2452;
  assign n2454 = n2453 ^ n2424;
  assign n2455 = n2447 & n2454;
  assign n2456 = ~n2446 & ~n2455;
  assign n2457 = n2437 & n2444;
  assign n2458 = n2436 & n2457;
  assign n2459 = n2364 & n2450;
  assign n2460 = n2429 & n2444;
  assign n2461 = n2366 & n2460;
  assign n2462 = ~n2459 & ~n2461;
  assign n2463 = n2392 & n2429;
  assign n2464 = n2429 & n2439;
  assign n2465 = ~n2463 & ~n2464;
  assign n2466 = ~n2432 & n2465;
  assign n2467 = n2434 & ~n2466;
  assign n2468 = n2428 & n2437;
  assign n2469 = ~n2430 & ~n2463;
  assign n2470 = ~n2468 & n2469;
  assign n2471 = n2436 & ~n2470;
  assign n2472 = ~n2467 & ~n2471;
  assign n2473 = n2421 & n2444;
  assign n2474 = ~n2445 & ~n2473;
  assign n2475 = n2441 & ~n2457;
  assign n2476 = n2474 & n2475;
  assign n2477 = n2427 & ~n2476;
  assign n2478 = n2437 & n2439;
  assign n2482 = n2423 & n2428;
  assign n2483 = ~n2478 & ~n2482;
  assign n2479 = ~n2457 & ~n2478;
  assign n2480 = ~n2445 & n2479;
  assign n2481 = ~n2468 & n2480;
  assign n2484 = n2483 ^ n2481;
  assign n2485 = n2483 ^ n2365;
  assign n2486 = n2485 ^ n2483;
  assign n2487 = n2484 & ~n2486;
  assign n2488 = n2487 ^ n2483;
  assign n2489 = ~n2447 & ~n2488;
  assign n2490 = ~n2477 & ~n2489;
  assign n2491 = n2472 & n2490;
  assign n2492 = n2462 & n2491;
  assign n2493 = ~n2458 & n2492;
  assign n2494 = n2456 & n2493;
  assign n2495 = n2443 & n2494;
  assign n2496 = ~n2433 & n2495;
  assign n2497 = ~n2431 & n2496;
  assign n2498 = ~n2426 & n2497;
  assign n2499 = n2498 ^ x14;
  assign n2500 = n2499 ^ x101;
  assign n2501 = ~n2363 & ~n2500;
  assign n2502 = n2327 & n2501;
  assign n2503 = n2324 & n2502;
  assign n2504 = ~n2322 & n2323;
  assign n2505 = n2325 & n2326;
  assign n2506 = ~n2363 & n2500;
  assign n2507 = n2505 & n2506;
  assign n2508 = n2363 & n2500;
  assign n2509 = n2505 & n2508;
  assign n2510 = ~n2507 & ~n2509;
  assign n2511 = n2504 & ~n2510;
  assign n2512 = n2327 & n2508;
  assign n2513 = n2323 & n2512;
  assign n2514 = n2322 & n2323;
  assign n2515 = n2363 & ~n2500;
  assign n2516 = n2327 & n2515;
  assign n2517 = n2514 & n2516;
  assign n2518 = ~n2513 & ~n2517;
  assign n2519 = n2502 & n2504;
  assign n2520 = n2323 ^ n2322;
  assign n2521 = n2327 & n2506;
  assign n2522 = n2505 & n2515;
  assign n2523 = ~n2521 & ~n2522;
  assign n2524 = ~n2520 & ~n2523;
  assign n2525 = ~n2519 & ~n2524;
  assign n2526 = n2518 & n2525;
  assign n2527 = n2501 & n2505;
  assign n2528 = n2324 & n2527;
  assign n2529 = n2322 & ~n2323;
  assign n2530 = n2325 & ~n2326;
  assign n2531 = n2506 & n2530;
  assign n2532 = ~n2325 & ~n2326;
  assign n2533 = n2508 & n2532;
  assign n2534 = ~n2531 & ~n2533;
  assign n2535 = n2508 & n2530;
  assign n2536 = n2515 & n2532;
  assign n2537 = ~n2535 & ~n2536;
  assign n2538 = n2534 & n2537;
  assign n2539 = n2529 & ~n2538;
  assign n2540 = n2506 & n2532;
  assign n2541 = ~n2535 & ~n2540;
  assign n2542 = n2514 & ~n2541;
  assign n2543 = n2504 & n2540;
  assign n2544 = n2324 & ~n2534;
  assign n2545 = ~n2502 & ~n2522;
  assign n2546 = n2529 & ~n2545;
  assign n2547 = ~n2544 & ~n2546;
  assign n2548 = ~n2543 & n2547;
  assign n2549 = n2324 & ~n2537;
  assign n2550 = ~n2509 & ~n2527;
  assign n2551 = n2529 & ~n2550;
  assign n2552 = ~n2549 & ~n2551;
  assign n2553 = n2501 & n2530;
  assign n2554 = n2501 & n2532;
  assign n2555 = ~n2553 & ~n2554;
  assign n2556 = n2514 & ~n2555;
  assign n2557 = n2515 & n2530;
  assign n2558 = ~n2531 & ~n2536;
  assign n2559 = ~n2557 & n2558;
  assign n2560 = n2504 & ~n2559;
  assign n2561 = ~n2556 & ~n2560;
  assign n2562 = n2552 & n2561;
  assign n2563 = n2548 & n2562;
  assign n2564 = ~n2542 & n2563;
  assign n2565 = ~n2539 & n2564;
  assign n2566 = ~n2528 & n2565;
  assign n2567 = n2526 & n2566;
  assign n2568 = ~n2511 & n2567;
  assign n2569 = ~n2503 & n2568;
  assign n2570 = n2569 ^ n1103;
  assign n2571 = n2570 ^ x115;
  assign n2572 = n1438 & n1463;
  assign n2573 = ~n1444 & n1460;
  assign n2574 = ~n1454 & n2573;
  assign n2575 = n1312 & ~n2574;
  assign n2576 = ~n2572 & ~n2575;
  assign n2577 = n1416 & ~n2178;
  assign n2578 = n1438 & n1454;
  assign n2579 = ~n1422 & ~n2578;
  assign n2580 = ~n1429 & n2579;
  assign n2581 = ~n1489 & n2580;
  assign n2582 = ~n1450 & n2581;
  assign n2583 = n2582 ^ n1426;
  assign n2584 = n1441 & n2178;
  assign n2585 = n2584 ^ n2582;
  assign n2586 = n2585 ^ n2584;
  assign n2587 = n1438 & ~n2192;
  assign n2588 = n2587 ^ n2584;
  assign n2589 = ~n2586 & n2588;
  assign n2590 = n2589 ^ n2584;
  assign n2591 = ~n2583 & n2590;
  assign n2592 = n2591 ^ n1426;
  assign n2593 = ~n2577 & ~n2592;
  assign n2594 = n2576 & n2593;
  assign n2595 = ~n1430 & n2594;
  assign n2596 = n2185 & n2595;
  assign n2597 = n1443 & n2596;
  assign n2598 = n1425 & n2597;
  assign n2599 = n2177 & n2598;
  assign n2600 = n2599 ^ x26;
  assign n2601 = n2600 ^ x97;
  assign n2602 = n1810 & n1834;
  assign n2603 = n2215 & ~n2602;
  assign n2604 = n1825 & n1847;
  assign n2605 = n1812 & n1837;
  assign n2606 = ~n2604 & ~n2605;
  assign n2607 = n1744 ^ n1743;
  assign n2608 = n2607 ^ n1808;
  assign n2609 = n2608 ^ n1771;
  assign n2610 = n2609 ^ n1744;
  assign n2611 = n2610 ^ n1808;
  assign n2612 = n1808 ^ n1771;
  assign n2613 = n1771 ^ n1744;
  assign n2614 = n2612 & ~n2613;
  assign n2615 = n2614 ^ n1771;
  assign n2616 = ~n2611 & n2615;
  assign n2617 = n2616 ^ n2608;
  assign n2618 = ~n1827 & ~n2617;
  assign n2619 = ~n1836 & n2618;
  assign n2620 = n1742 & ~n2619;
  assign n2621 = ~n1820 & n1864;
  assign n2622 = n1834 & ~n2621;
  assign n2623 = ~n1810 & n1844;
  assign n2624 = ~n1812 & n2623;
  assign n2625 = ~n1822 & ~n1843;
  assign n2626 = ~n1854 & n2625;
  assign n2627 = ~n1825 & n2626;
  assign n2628 = ~n2624 & ~n2627;
  assign n2629 = ~n1816 & ~n2628;
  assign n2630 = ~n1858 & ~n2629;
  assign n2631 = ~n2622 & ~n2630;
  assign n2632 = ~n2620 & n2631;
  assign n2633 = n2606 & n2632;
  assign n2634 = n2212 & n2633;
  assign n2635 = n2603 & n2634;
  assign n2636 = ~n1850 & n2635;
  assign n2637 = n2636 ^ x0;
  assign n2638 = n2637 ^ x107;
  assign n2639 = n2601 & n2638;
  assign n2640 = n2008 & n2012;
  assign n2641 = n2023 & n2640;
  assign n2642 = n2004 & ~n2641;
  assign n2643 = n1997 & n2009;
  assign n2644 = n1997 & n2039;
  assign n2645 = n1954 & n2640;
  assign n2646 = ~n2644 & ~n2645;
  assign n2647 = ~n2643 & n2646;
  assign n2648 = n1991 & n2012;
  assign n2649 = n2023 & n2648;
  assign n2650 = n2011 & ~n2649;
  assign n2651 = ~n1952 & n2018;
  assign n2652 = n2023 & ~n2045;
  assign n2653 = ~n2651 & ~n2652;
  assign n2654 = n2016 & n2035;
  assign n2655 = ~n2013 & ~n2053;
  assign n2656 = ~n2648 & n2655;
  assign n2657 = n1997 & ~n2656;
  assign n2658 = ~n1999 & ~n2039;
  assign n2659 = ~n2056 & n2658;
  assign n2660 = n1954 & ~n2659;
  assign n2661 = ~n2657 & ~n2660;
  assign n2662 = ~n2654 & n2661;
  assign n2663 = n2653 & n2662;
  assign n2664 = n2650 & n2663;
  assign n2665 = n2647 & n2664;
  assign n2666 = n2642 & n2665;
  assign n2667 = n2666 ^ x34;
  assign n2668 = n2667 ^ x112;
  assign n2669 = n1229 & n1234;
  assign n2670 = n1151 & n2669;
  assign n2671 = ~n1231 & n1264;
  assign n2672 = ~n2670 & ~n2671;
  assign n2673 = ~n2098 & ~n2099;
  assign n2674 = n1264 & ~n2673;
  assign n2675 = n1261 & ~n2101;
  assign n2676 = n1234 & ~n2675;
  assign n2677 = ~n2674 & ~n2676;
  assign n2678 = ~n1185 & n2129;
  assign n2679 = n2677 & ~n2678;
  assign n2680 = n2672 & n2679;
  assign n2681 = n2680 ^ x50;
  assign n2682 = n2681 ^ x65;
  assign n2683 = ~n2668 & n2682;
  assign n2684 = n2422 & n2427;
  assign n2685 = ~n2432 & ~n2460;
  assign n2686 = n2436 & ~n2685;
  assign n2687 = ~n2684 & ~n2686;
  assign n2688 = ~n2431 & n2687;
  assign n2689 = n2436 & n2450;
  assign n2690 = n2434 & ~n2474;
  assign n2691 = ~n2689 & ~n2690;
  assign n2692 = n2427 & ~n2685;
  assign n2693 = ~n2450 & ~n2464;
  assign n2694 = n2474 & n2693;
  assign n2695 = ~n2468 & n2694;
  assign n2696 = n2366 & ~n2695;
  assign n2697 = ~n2692 & ~n2696;
  assign n2698 = ~n2430 & ~n2464;
  assign n2699 = n2434 & ~n2698;
  assign n2700 = n2424 & n2434;
  assign n2701 = ~n2427 & ~n2434;
  assign n2702 = ~n2479 & ~n2701;
  assign n2703 = ~n2700 & ~n2702;
  assign n2704 = n2427 & n2440;
  assign n2705 = ~n2468 & ~n2482;
  assign n2706 = n2465 & n2705;
  assign n2707 = n2436 & ~n2706;
  assign n2708 = ~n2704 & ~n2707;
  assign n2709 = n2703 & n2708;
  assign n2710 = ~n2699 & n2709;
  assign n2711 = n2697 & n2710;
  assign n2712 = n2691 & n2711;
  assign n2713 = n2688 & n2712;
  assign n2714 = ~n2426 & n2713;
  assign n2715 = ~n2438 & n2714;
  assign n2716 = n2715 ^ x58;
  assign n2717 = n2716 ^ x74;
  assign n2718 = n720 & n1052;
  assign n2719 = n752 & n1036;
  assign n2720 = ~n2718 & ~n2719;
  assign n2721 = ~n1012 & n1053;
  assign n2722 = n992 ^ n954;
  assign n2723 = n954 ^ n837;
  assign n2724 = n2723 ^ n992;
  assign n2725 = n2724 ^ n954;
  assign n2726 = n2722 & ~n2725;
  assign n2727 = n2726 ^ n954;
  assign n2728 = ~n918 & ~n2727;
  assign n2729 = n2728 ^ n2724;
  assign n2730 = n1019 & n2729;
  assign n2731 = n999 & ~n1045;
  assign n2732 = n1001 & ~n2731;
  assign n2733 = ~n1004 & ~n1011;
  assign n2734 = ~n1016 & n2150;
  assign n2735 = ~n2733 & ~n2734;
  assign n2736 = ~n1010 & ~n2735;
  assign n2737 = ~n1034 & n2736;
  assign n2738 = ~n1012 & ~n2737;
  assign n2739 = ~n2732 & ~n2738;
  assign n2740 = ~n2730 & n2739;
  assign n2741 = ~n2721 & n2740;
  assign n2742 = n2720 & n2741;
  assign n2743 = n1031 ^ n995;
  assign n2744 = n2743 ^ n1031;
  assign n2745 = n1031 ^ n751;
  assign n2746 = n2745 ^ n1031;
  assign n2747 = n2744 & n2746;
  assign n2748 = n2747 ^ n1031;
  assign n2749 = ~n720 & n2748;
  assign n2750 = n2749 ^ n1031;
  assign n2751 = n2742 & ~n2750;
  assign n2752 = n1009 & n2751;
  assign n2753 = n2138 & n2752;
  assign n2754 = n1029 & n2753;
  assign n2755 = n2754 ^ x42;
  assign n2756 = n2755 ^ x64;
  assign n2757 = ~n2717 & n2756;
  assign n2758 = n2683 & n2757;
  assign n2759 = n2639 & n2758;
  assign n2760 = n2601 & ~n2638;
  assign n2761 = n2717 & ~n2756;
  assign n2762 = n2683 & n2761;
  assign n2763 = n2668 & ~n2682;
  assign n2764 = n2761 & n2763;
  assign n2765 = ~n2762 & ~n2764;
  assign n2766 = n2760 & ~n2765;
  assign n2767 = ~n2601 & ~n2638;
  assign n2768 = ~n2668 & ~n2682;
  assign n2769 = n2761 & n2768;
  assign n2770 = n2668 & n2682;
  assign n2771 = n2761 & n2770;
  assign n2772 = ~n2769 & ~n2771;
  assign n2773 = n2767 & ~n2772;
  assign n2774 = ~n2766 & ~n2773;
  assign n2775 = n2757 & n2763;
  assign n2776 = ~n2717 & ~n2756;
  assign n2777 = n2768 & n2776;
  assign n2778 = ~n2775 & ~n2777;
  assign n2779 = n2639 & ~n2778;
  assign n2780 = ~n2601 & n2638;
  assign n2781 = ~n2762 & ~n2771;
  assign n2782 = n2780 & ~n2781;
  assign n2783 = ~n2779 & ~n2782;
  assign n2784 = ~n2760 & ~n2780;
  assign n2785 = n2717 & n2756;
  assign n2786 = n2770 & n2785;
  assign n2787 = n2763 & n2785;
  assign n2788 = ~n2786 & ~n2787;
  assign n2789 = ~n2784 & ~n2788;
  assign n2790 = n2768 & n2785;
  assign n2791 = n2772 & ~n2790;
  assign n2792 = ~n2762 & n2791;
  assign n2793 = n2639 & ~n2792;
  assign n2794 = n2757 & n2770;
  assign n2795 = n2683 & n2776;
  assign n2796 = ~n2775 & ~n2795;
  assign n2797 = ~n2758 & n2796;
  assign n2798 = ~n2794 & n2797;
  assign n2799 = n2767 & ~n2798;
  assign n2800 = ~n2793 & ~n2799;
  assign n2801 = n2638 ^ n2601;
  assign n2805 = n2763 & n2776;
  assign n2802 = n2757 & n2768;
  assign n2808 = n2683 & n2785;
  assign n2809 = ~n2802 & ~n2808;
  assign n2810 = ~n2795 & n2809;
  assign n2811 = ~n2805 & n2810;
  assign n2803 = n2770 & n2776;
  assign n2804 = ~n2802 & ~n2803;
  assign n2806 = ~n2777 & ~n2805;
  assign n2807 = n2804 & n2806;
  assign n2812 = n2811 ^ n2807;
  assign n2813 = n2811 ^ n2638;
  assign n2814 = n2813 ^ n2811;
  assign n2815 = n2812 & n2814;
  assign n2816 = n2815 ^ n2811;
  assign n2817 = n2801 & ~n2816;
  assign n2818 = n2800 & ~n2817;
  assign n2819 = ~n2789 & n2818;
  assign n2820 = n2783 & n2819;
  assign n2821 = n2774 & n2820;
  assign n2822 = n2794 ^ n2638;
  assign n2823 = n2822 ^ n2794;
  assign n2824 = ~n2764 & ~n2790;
  assign n2825 = n2824 ^ n2794;
  assign n2826 = ~n2823 & ~n2825;
  assign n2827 = n2826 ^ n2794;
  assign n2828 = ~n2801 & n2827;
  assign n2829 = n2821 & ~n2828;
  assign n2830 = ~n2759 & n2829;
  assign n2831 = n2830 ^ n1149;
  assign n2832 = n2831 ^ x106;
  assign n2833 = ~n638 & ~n653;
  assign n2834 = n625 & ~n2833;
  assign n2835 = n296 & ~n640;
  assign n2836 = ~n643 & n2338;
  assign n2837 = ~n663 & n2836;
  assign n2838 = n625 & ~n2837;
  assign n2839 = ~n633 & ~n659;
  assign n2840 = n640 & n2839;
  assign n2841 = n616 & ~n2840;
  assign n2842 = ~n2838 & ~n2841;
  assign n2843 = n644 & n651;
  assign n2844 = ~n648 & ~n654;
  assign n2845 = n296 & ~n2844;
  assign n2846 = n655 & n660;
  assign n2847 = ~n610 & n2846;
  assign n2848 = n630 & ~n2847;
  assign n2849 = ~n2845 & ~n2848;
  assign n2850 = ~n2843 & n2849;
  assign n2851 = n2842 & n2850;
  assign n2852 = n628 & n2851;
  assign n2853 = ~n2835 & n2852;
  assign n2854 = n652 ^ n295;
  assign n2855 = n2854 ^ n652;
  assign n2856 = n663 ^ n652;
  assign n2857 = n2855 & n2856;
  assign n2858 = n2857 ^ n652;
  assign n2859 = n651 & n2858;
  assign n2860 = n2853 & ~n2859;
  assign n2861 = n636 & n2860;
  assign n2862 = ~n2834 & n2861;
  assign n2863 = ~n2334 & n2862;
  assign n2864 = n2330 & n2863;
  assign n2865 = n2864 ^ x2;
  assign n2866 = n2865 ^ x124;
  assign n2867 = ~n1676 & ~n1691;
  assign n2868 = ~n1679 & n2867;
  assign n2869 = n1685 & ~n2868;
  assign n2870 = n1559 & ~n1712;
  assign n2871 = ~n2869 & ~n2870;
  assign n2872 = ~n1686 & n1695;
  assign n2873 = n1664 & ~n2872;
  assign n2874 = n1689 & ~n1704;
  assign n2875 = ~n1662 & n2068;
  assign n2876 = ~n1679 & n2875;
  assign n2877 = n1698 & ~n2876;
  assign n2878 = ~n2874 & ~n2877;
  assign n2879 = n1685 ^ n1667;
  assign n2880 = n1667 ^ n1559;
  assign n2881 = n2880 ^ n1559;
  assign n2882 = n1714 ^ n1559;
  assign n2883 = ~n2881 & n2882;
  assign n2884 = n2883 ^ n1559;
  assign n2885 = n2879 & n2884;
  assign n2886 = n2885 ^ n1685;
  assign n2887 = n2878 & ~n2886;
  assign n2888 = ~n2873 & n2887;
  assign n2889 = n2871 & n2888;
  assign n2890 = n1684 & n2889;
  assign n2891 = ~n2064 & n2890;
  assign n2892 = ~n1675 & n2891;
  assign n2893 = n1669 & n2892;
  assign n2894 = ~n1736 & n2893;
  assign n2895 = n2894 ^ x28;
  assign n2896 = n2895 ^ x110;
  assign n2897 = ~n2866 & n2896;
  assign n2898 = n1186 & ~n1242;
  assign n2899 = n1151 & ~n1225;
  assign n2900 = n1252 & ~n2899;
  assign n2901 = n1234 & ~n2900;
  assign n2902 = ~n2898 & ~n2901;
  assign n2903 = n1224 & n1271;
  assign n2904 = ~n1262 & n1264;
  assign n2905 = ~n2903 & ~n2904;
  assign n2906 = n2902 & n2905;
  assign n2907 = n2672 & n2906;
  assign n2908 = n2907 ^ x36;
  assign n2909 = n2908 ^ x76;
  assign n2910 = ~n2366 & ~n2434;
  assign n2911 = ~n2705 & ~n2910;
  assign n2912 = ~n2693 & ~n2701;
  assign n2913 = ~n2911 & ~n2912;
  assign n2914 = n2434 & n2438;
  assign n2915 = n2436 & n2445;
  assign n2916 = ~n2914 & ~n2915;
  assign n2917 = ~n2457 & n2465;
  assign n2918 = n2366 & ~n2917;
  assign n2919 = ~n2424 & ~n2468;
  assign n2920 = n2479 & n2919;
  assign n2921 = n2427 & ~n2920;
  assign n2922 = ~n2918 & ~n2921;
  assign n2923 = n2916 & n2922;
  assign n2924 = n2913 & n2923;
  assign n2925 = n2691 & n2924;
  assign n2926 = n2443 & n2925;
  assign n2927 = n2436 & n2479;
  assign n2928 = n2927 ^ n2436;
  assign n2929 = n2926 & ~n2928;
  assign n2930 = n2688 & n2929;
  assign n2931 = ~n2433 & n2930;
  assign n2932 = ~n2426 & n2931;
  assign n2933 = n2932 ^ x60;
  assign n2934 = n2933 ^ x67;
  assign n2935 = ~n2909 & n2934;
  assign n2936 = n1426 & n1444;
  assign n2937 = n1416 & n1446;
  assign n2938 = n1310 & ~n2194;
  assign n2939 = n1423 & n2192;
  assign n2940 = n1416 & n1454;
  assign n2941 = ~n1426 & ~n2940;
  assign n2942 = ~n2939 & ~n2941;
  assign n2943 = n1457 & n2193;
  assign n2944 = ~n1463 & n2943;
  assign n2945 = n1312 & ~n2944;
  assign n2946 = ~n2942 & ~n2945;
  assign n2947 = ~n2938 & n2946;
  assign n2948 = ~n2937 & n2947;
  assign n2949 = ~n2936 & n2948;
  assign n2950 = n1431 & n2949;
  assign n2951 = n2182 & n2950;
  assign n2952 = n1452 & n2951;
  assign n2953 = n1437 & n2952;
  assign n2954 = n2177 & n2953;
  assign n2955 = n2954 ^ x52;
  assign n2956 = n2955 ^ x78;
  assign n2957 = ~n1024 & ~n1052;
  assign n2958 = n752 & ~n2957;
  assign n2959 = n1048 & ~n1053;
  assign n2960 = n1001 & ~n2959;
  assign n2961 = ~n2958 & ~n2960;
  assign n2962 = ~n1012 & n1026;
  assign n2963 = n1007 & ~n1034;
  assign n2964 = n1019 & ~n2963;
  assign n2965 = n752 & ~n2147;
  assign n2966 = ~n1020 & n2733;
  assign n2967 = n2150 & n2966;
  assign n2968 = n1001 & ~n2967;
  assign n2969 = ~n2965 & ~n2968;
  assign n2970 = ~n995 & n1037;
  assign n2971 = n1011 & ~n2970;
  assign n2972 = ~n1036 & n1048;
  assign n2973 = ~n1024 & n2972;
  assign n2974 = n1019 & ~n2973;
  assign n2975 = ~n2971 & ~n2974;
  assign n2976 = ~n1013 & n2975;
  assign n2977 = n2969 & n2976;
  assign n2978 = ~n2964 & n2977;
  assign n2979 = ~n2962 & n2978;
  assign n2980 = n2961 & n2979;
  assign n2981 = ~n2137 & n2980;
  assign n2982 = ~n2750 & n2981;
  assign n2983 = ~n2140 & n2982;
  assign n2984 = n2983 ^ x44;
  assign n2985 = n2984 ^ x93;
  assign n2986 = n2956 & ~n2985;
  assign n2987 = n2935 & n2986;
  assign n2988 = n2897 & n2987;
  assign n2989 = n2866 & ~n2896;
  assign n2990 = n2987 & n2989;
  assign n2991 = n2866 & n2896;
  assign n2992 = ~n2956 & n2985;
  assign n2993 = ~n2909 & ~n2934;
  assign n2994 = n2992 & n2993;
  assign n2995 = n2991 & n2994;
  assign n2996 = ~n2990 & ~n2995;
  assign n2997 = n2909 & n2934;
  assign n2998 = ~n2956 & ~n2985;
  assign n2999 = n2997 & n2998;
  assign n3000 = n2956 & n2985;
  assign n3001 = n2935 & n3000;
  assign n3002 = ~n2999 & ~n3001;
  assign n3003 = n2989 & ~n3002;
  assign n3004 = n2993 & n3000;
  assign n3005 = n2909 & ~n2934;
  assign n3006 = n2998 & n3005;
  assign n3007 = n3000 & n3005;
  assign n3008 = ~n3006 & ~n3007;
  assign n3009 = ~n3004 & n3008;
  assign n3010 = n2991 & ~n3009;
  assign n3011 = ~n2897 & ~n2989;
  assign n3012 = n2992 & n2997;
  assign n3013 = n2986 & n3005;
  assign n3014 = n3008 & ~n3013;
  assign n3015 = ~n2989 & n3014;
  assign n3016 = n2993 & n2998;
  assign n3017 = ~n3004 & ~n3013;
  assign n3018 = ~n3016 & n3017;
  assign n3019 = ~n2897 & n3018;
  assign n3020 = ~n3015 & ~n3019;
  assign n3021 = ~n3012 & ~n3020;
  assign n3022 = ~n3011 & ~n3021;
  assign n3023 = ~n3010 & ~n3022;
  assign n3024 = n2997 & n3000;
  assign n3025 = n2935 & n2992;
  assign n3026 = ~n3024 & ~n3025;
  assign n3027 = n2897 & ~n3026;
  assign n3028 = ~n2866 & ~n2896;
  assign n3029 = n2935 & n2998;
  assign n3030 = ~n2999 & ~n3029;
  assign n3031 = n2986 & n2997;
  assign n3032 = ~n3001 & ~n3031;
  assign n3033 = n3030 & n3032;
  assign n3034 = n3028 & ~n3033;
  assign n3035 = n2986 & n2993;
  assign n3038 = ~n2994 & ~n3007;
  assign n3039 = ~n3035 & n3038;
  assign n3036 = ~n3031 & ~n3035;
  assign n3037 = ~n3029 & n3036;
  assign n3040 = n3039 ^ n3037;
  assign n3041 = n2896 ^ n2866;
  assign n3042 = n3037 ^ n2896;
  assign n3043 = n3041 & n3042;
  assign n3044 = n3043 ^ n2896;
  assign n3045 = n3040 & n3044;
  assign n3046 = n3045 ^ n3039;
  assign n3047 = ~n3025 & n3046;
  assign n3048 = n3011 & ~n3047;
  assign n3049 = ~n3034 & ~n3048;
  assign n3050 = ~n3027 & n3049;
  assign n3051 = n3023 & n3050;
  assign n3052 = ~n3003 & n3051;
  assign n3053 = n2996 & n3052;
  assign n3054 = ~n2988 & n3053;
  assign n3055 = n3016 ^ n2896;
  assign n3056 = n3055 ^ n3016;
  assign n3057 = n2992 & n3005;
  assign n3058 = n3057 ^ n3016;
  assign n3059 = ~n3056 & n3058;
  assign n3060 = n3059 ^ n3016;
  assign n3061 = n3041 & n3060;
  assign n3062 = n3054 & ~n3061;
  assign n3063 = n3062 ^ n1220;
  assign n3064 = n3063 ^ x88;
  assign n3065 = ~n2832 & n3064;
  assign n3066 = ~n2571 & n3065;
  assign n3067 = n2832 ^ n2571;
  assign n3068 = n2171 ^ x72;
  assign n3069 = n2716 ^ x81;
  assign n3070 = ~n3068 & ~n3069;
  assign n3071 = n2095 ^ x96;
  assign n3072 = ~n2017 & n2640;
  assign n3073 = n1993 & n1998;
  assign n3074 = ~n1999 & ~n3073;
  assign n3075 = ~n2648 & n3074;
  assign n3076 = ~n1994 & n3075;
  assign n3077 = n1997 & ~n3076;
  assign n3078 = ~n1954 & ~n2016;
  assign n3079 = ~n2001 & n2014;
  assign n3080 = ~n2016 & n3079;
  assign n3081 = ~n1994 & ~n2009;
  assign n3082 = n2002 & n3081;
  assign n3083 = ~n1954 & n3082;
  assign n3084 = ~n3080 & ~n3083;
  assign n3085 = n2020 & ~n3084;
  assign n3086 = ~n3078 & ~n3085;
  assign n3087 = ~n3077 & ~n3086;
  assign n3088 = ~n3072 & n3087;
  assign n3089 = ~n1992 & ~n3073;
  assign n3090 = n2041 & n3089;
  assign n3091 = ~n2056 & n3090;
  assign n3092 = n3091 ^ n2053;
  assign n3093 = ~n2055 & ~n3092;
  assign n3094 = n3093 ^ n2053;
  assign n3095 = ~n1953 & n3094;
  assign n3096 = n3088 & ~n3095;
  assign n3097 = n2646 & n3096;
  assign n3098 = n2650 & n3097;
  assign n3099 = ~n2060 & n3098;
  assign n3100 = n3099 ^ x8;
  assign n3101 = n3100 ^ x113;
  assign n3102 = ~n3071 & ~n3101;
  assign n3103 = ~n639 & n2332;
  assign n3104 = n667 & n3103;
  assign n3105 = n634 & n3104;
  assign n3106 = n630 & ~n3105;
  assign n3108 = n660 & n2339;
  assign n3107 = n649 & n2344;
  assign n3109 = n3108 ^ n3107;
  assign n3110 = n3109 ^ n3108;
  assign n3111 = n3108 ^ n295;
  assign n3112 = n3111 ^ n3108;
  assign n3113 = ~n3110 & n3112;
  assign n3114 = n3113 ^ n3108;
  assign n3115 = ~n651 & ~n3114;
  assign n3116 = n3115 ^ n3108;
  assign n3117 = ~n3106 & n3116;
  assign n3118 = n619 & n3117;
  assign n3119 = ~n2859 & n3118;
  assign n3120 = n627 & n3119;
  assign n3121 = ~n2834 & n3120;
  assign n3122 = ~n2334 & n3121;
  assign n3123 = n2330 & n3122;
  assign n3124 = n3123 ^ x16;
  assign n3125 = n3124 ^ x106;
  assign n3126 = n2637 ^ x123;
  assign n3127 = ~n3125 & ~n3126;
  assign n3128 = n3102 & n3127;
  assign n3129 = n3070 & n3128;
  assign n3130 = n3069 ^ n3068;
  assign n3131 = n3128 ^ n3069;
  assign n3132 = n3131 ^ n3128;
  assign n3133 = n3071 & ~n3101;
  assign n3134 = n3125 & n3126;
  assign n3135 = n3133 & n3134;
  assign n3136 = n3071 & n3101;
  assign n3137 = n3127 & n3136;
  assign n3138 = ~n3135 & ~n3137;
  assign n3139 = n3138 ^ n3128;
  assign n3140 = ~n3132 & ~n3139;
  assign n3141 = n3140 ^ n3128;
  assign n3142 = ~n3130 & n3141;
  assign n3143 = ~n3129 & ~n3142;
  assign n3144 = n3068 & ~n3069;
  assign n3145 = ~n3125 & n3126;
  assign n3146 = n3133 & n3145;
  assign n3147 = n3125 & ~n3126;
  assign n3148 = n3133 & n3147;
  assign n3149 = ~n3146 & ~n3148;
  assign n3150 = n3144 & ~n3149;
  assign n3151 = ~n3068 & n3069;
  assign n3152 = n3136 & n3145;
  assign n3153 = n3136 & n3147;
  assign n3154 = ~n3152 & ~n3153;
  assign n3155 = n3151 & ~n3154;
  assign n3156 = ~n3150 & ~n3155;
  assign n3157 = n3127 & n3133;
  assign n3158 = n3151 & n3157;
  assign n3159 = ~n3071 & n3101;
  assign n3160 = n3134 & n3159;
  assign n3161 = ~n3128 & ~n3160;
  assign n3162 = n3144 & ~n3161;
  assign n3163 = ~n3158 & ~n3162;
  assign n3164 = n3068 & n3069;
  assign n3165 = ~n3154 & n3164;
  assign n3166 = n3102 & n3134;
  assign n3167 = n3127 & n3159;
  assign n3168 = ~n3166 & ~n3167;
  assign n3169 = n3151 & ~n3168;
  assign n3170 = ~n3165 & ~n3169;
  assign n3171 = n3102 & n3147;
  assign n3172 = ~n3135 & ~n3171;
  assign n3173 = n3151 & ~n3172;
  assign n3174 = n3134 & n3136;
  assign n3175 = n3168 & ~n3174;
  assign n3176 = n3144 & ~n3175;
  assign n3177 = ~n3173 & ~n3176;
  assign n3178 = n3102 & n3145;
  assign n3179 = n3138 & ~n3178;
  assign n3180 = n3164 & ~n3179;
  assign n3181 = n3145 & n3159;
  assign n3182 = ~n3171 & ~n3181;
  assign n3183 = ~n3070 & ~n3164;
  assign n3184 = n3147 & n3159;
  assign n3185 = ~n3181 & ~n3184;
  assign n3186 = ~n3178 & n3185;
  assign n3187 = ~n3164 & n3186;
  assign n3188 = ~n3183 & ~n3187;
  assign n3189 = ~n3182 & n3188;
  assign n3190 = ~n3146 & ~n3188;
  assign n3191 = ~n3153 & n3190;
  assign n3192 = n3070 & ~n3191;
  assign n3193 = ~n3189 & ~n3192;
  assign n3194 = ~n3180 & n3193;
  assign n3195 = n3177 & n3194;
  assign n3196 = n3170 & n3195;
  assign n3197 = n3160 ^ n3069;
  assign n3198 = n3197 ^ n3160;
  assign n3199 = n3160 ^ n3137;
  assign n3200 = ~n3198 & n3199;
  assign n3201 = n3200 ^ n3160;
  assign n3202 = n3130 & n3201;
  assign n3203 = n3196 & ~n3202;
  assign n3204 = n3163 & n3203;
  assign n3205 = n3156 & n3204;
  assign n3206 = n3143 & n3205;
  assign n3207 = n3206 ^ n205;
  assign n3208 = n3207 ^ x89;
  assign n3209 = ~n3067 & n3208;
  assign n3210 = n2571 & ~n3208;
  assign n3211 = n3064 & n3210;
  assign n3212 = ~n3209 & ~n3211;
  assign n3213 = ~n3066 & n3212;
  assign n3214 = n2832 & ~n3064;
  assign n3215 = ~n3208 & n3214;
  assign n3216 = ~n2571 & n3215;
  assign n3217 = n3213 & ~n3216;
  assign n3218 = n2321 & n3217;
  assign n3219 = n1951 & n2320;
  assign n3220 = ~n2832 & ~n3064;
  assign n3221 = ~n2571 & n3208;
  assign n3222 = ~n3210 & ~n3221;
  assign n3223 = n3220 & ~n3222;
  assign n3224 = n2832 & n3064;
  assign n3225 = ~n3208 & n3224;
  assign n3226 = n3065 & n3222;
  assign n3227 = ~n3225 & ~n3226;
  assign n3228 = ~n3223 & n3227;
  assign n3229 = ~n3208 & n3220;
  assign n3230 = n3229 ^ n3208;
  assign n3231 = n3230 ^ n3229;
  assign n3232 = n3229 ^ n3214;
  assign n3233 = n3232 ^ n3229;
  assign n3234 = n3231 & n3233;
  assign n3235 = n3234 ^ n3229;
  assign n3236 = n2571 & n3235;
  assign n3237 = n3236 ^ n3229;
  assign n3238 = n3228 & ~n3237;
  assign n3239 = n3219 & ~n3238;
  assign n3240 = ~n3218 & ~n3239;
  assign n3241 = ~n1951 & ~n2320;
  assign n3242 = n3208 ^ n2571;
  assign n3243 = n3242 ^ n3064;
  assign n3244 = n3243 ^ n3208;
  assign n3245 = n3064 ^ n2832;
  assign n3246 = n3245 ^ n2832;
  assign n3247 = n3208 ^ n2832;
  assign n3248 = n3247 ^ n2832;
  assign n3249 = n3246 & n3248;
  assign n3250 = n3249 ^ n2832;
  assign n3251 = n3244 & ~n3250;
  assign n3252 = n3251 ^ n3242;
  assign n3253 = n3241 & n3252;
  assign n3254 = ~n1951 & n2320;
  assign n3255 = n2571 & n3220;
  assign n3256 = n3208 & n3224;
  assign n3257 = n3064 & ~n3222;
  assign n3258 = ~n3256 & ~n3257;
  assign n3259 = ~n3255 & n3258;
  assign n3260 = ~n3216 & n3259;
  assign n3261 = n3254 & ~n3260;
  assign n3262 = ~n3253 & ~n3261;
  assign n3263 = n3240 & n3262;
  assign n3264 = n3263 ^ n2908;
  assign n3265 = n3264 ^ x117;
  assign n3266 = n2600 ^ x105;
  assign n3267 = n1812 & ~n1830;
  assign n3268 = n1834 & n2617;
  assign n3269 = ~n3267 & ~n3268;
  assign n3270 = n1825 & ~n2229;
  assign n3271 = n2226 & n2626;
  assign n3272 = ~n1862 & n3271;
  assign n3273 = ~n1848 & n3272;
  assign n3274 = n1742 & ~n3273;
  assign n3275 = ~n1847 & n1873;
  assign n3276 = ~n1837 & n3275;
  assign n3277 = n3276 ^ n1841;
  assign n3278 = n1841 ^ n1741;
  assign n3279 = n3278 ^ n1841;
  assign n3280 = n3277 & n3279;
  assign n3281 = n3280 ^ n1841;
  assign n3282 = n1870 & ~n3281;
  assign n3283 = ~n3274 & ~n3282;
  assign n3284 = ~n3270 & n3283;
  assign n3285 = n3269 & n3284;
  assign n3286 = n1819 & n3285;
  assign n3287 = n2603 & n3286;
  assign n3288 = n3287 ^ x18;
  assign n3289 = n3288 ^ x104;
  assign n3290 = n3266 & n3289;
  assign n3291 = n2865 ^ x122;
  assign n3292 = n1558 & n1670;
  assign n3293 = n1673 & n1689;
  assign n3294 = ~n3292 & ~n3293;
  assign n3295 = n1685 & ~n1711;
  assign n3296 = ~n1699 & ~n1710;
  assign n3297 = n1664 & ~n3296;
  assign n3298 = ~n3295 & ~n3297;
  assign n3299 = n3294 & n3298;
  assign n3300 = n1559 & ~n1692;
  assign n3301 = ~n1667 & ~n1703;
  assign n3302 = n1698 & ~n3301;
  assign n3303 = n1698 & ~n2071;
  assign n3304 = ~n1662 & ~n1676;
  assign n3305 = n1692 & n3304;
  assign n3306 = n1664 & ~n3305;
  assign n3307 = ~n3303 & ~n3306;
  assign n3308 = n1692 & ~n1702;
  assign n3309 = n1685 & ~n3308;
  assign n3310 = ~n1699 & n1711;
  assign n3311 = ~n1673 & n3310;
  assign n3312 = n1559 & ~n3311;
  assign n3313 = ~n3309 & ~n3312;
  assign n3314 = n3307 & n3313;
  assign n3315 = ~n1736 & n3314;
  assign n3316 = ~n3302 & n3315;
  assign n3317 = ~n3300 & n3316;
  assign n3318 = n3299 & n3317;
  assign n3319 = ~n1677 & n3318;
  assign n3320 = ~n2064 & n3319;
  assign n3321 = n1669 & n3320;
  assign n3322 = n3321 ^ x10;
  assign n3323 = n3322 ^ x66;
  assign n3324 = ~n3291 & ~n3323;
  assign n3325 = n2667 ^ x98;
  assign n3326 = n2933 ^ x80;
  assign n3327 = n3325 & n3326;
  assign n3328 = n3324 & n3327;
  assign n3329 = n3291 & ~n3323;
  assign n3330 = ~n3325 & n3326;
  assign n3331 = n3329 & n3330;
  assign n3332 = ~n3328 & ~n3331;
  assign n3333 = n3290 & ~n3332;
  assign n3334 = ~n3266 & ~n3289;
  assign n3335 = ~n3291 & n3334;
  assign n3336 = ~n3266 & n3289;
  assign n3337 = n3329 & n3336;
  assign n3338 = ~n3335 & ~n3337;
  assign n3339 = n3291 & n3323;
  assign n3340 = n3289 & n3339;
  assign n3341 = n3334 & n3339;
  assign n3342 = n3266 & ~n3289;
  assign n3343 = n3329 & n3342;
  assign n3344 = ~n3341 & ~n3343;
  assign n3345 = ~n3340 & n3344;
  assign n3346 = n3338 & n3345;
  assign n3347 = n3327 & ~n3346;
  assign n3348 = ~n3291 & n3342;
  assign n3349 = ~n3291 & n3323;
  assign n3350 = n3336 & n3349;
  assign n3351 = ~n3348 & ~n3350;
  assign n3352 = n3339 ^ n3323;
  assign n3353 = n3266 & ~n3352;
  assign n3354 = n3353 ^ n3323;
  assign n3355 = ~n3289 & ~n3354;
  assign n3356 = n3351 & ~n3355;
  assign n3357 = ~n3337 & n3356;
  assign n3358 = n3330 & ~n3357;
  assign n3359 = ~n3347 & ~n3358;
  assign n3360 = n3266 & n3339;
  assign n3361 = n3291 & n3334;
  assign n3362 = n3349 ^ n3324;
  assign n3363 = n3349 ^ n3336;
  assign n3364 = n3363 ^ n3349;
  assign n3365 = n3362 & ~n3364;
  assign n3366 = n3365 ^ n3349;
  assign n3367 = ~n3361 & ~n3366;
  assign n3368 = ~n3360 & n3367;
  assign n3369 = n3368 ^ n3325;
  assign n3370 = n3369 ^ n3368;
  assign n3371 = n3323 ^ n3289;
  assign n3372 = n3323 ^ n3291;
  assign n3373 = n3372 ^ n3291;
  assign n3374 = n3289 ^ n3266;
  assign n3375 = n3374 ^ n3291;
  assign n3376 = n3375 ^ n3291;
  assign n3377 = n3373 & n3376;
  assign n3378 = n3377 ^ n3291;
  assign n3379 = n3371 & ~n3378;
  assign n3380 = n3379 ^ n3374;
  assign n3381 = n3380 ^ n3368;
  assign n3382 = ~n3370 & ~n3381;
  assign n3383 = n3382 ^ n3368;
  assign n3384 = ~n3326 & n3383;
  assign n3385 = n3359 & ~n3384;
  assign n3386 = ~n3333 & n3385;
  assign n3387 = n3386 ^ n719;
  assign n3388 = n3387 ^ x91;
  assign n3389 = n2319 ^ x118;
  assign n3390 = n3388 & n3389;
  assign n3391 = n3151 & n3178;
  assign n3392 = n3164 & n3184;
  assign n3393 = n3164 & n3178;
  assign n3394 = n3144 & n3167;
  assign n3395 = ~n3393 & ~n3394;
  assign n3396 = n3166 & ~n3183;
  assign n3397 = ~n3153 & n3185;
  assign n3398 = ~n3160 & n3397;
  assign n3399 = ~n3135 & n3398;
  assign n3400 = n3144 & ~n3399;
  assign n3401 = ~n3396 & ~n3400;
  assign n3402 = ~n3149 & n3164;
  assign n3403 = ~n3128 & ~n3174;
  assign n3404 = ~n3148 & n3403;
  assign n3405 = n3151 & ~n3404;
  assign n3406 = ~n3152 & n3182;
  assign n3407 = ~n3157 & n3406;
  assign n3408 = n3070 & ~n3407;
  assign n3409 = ~n3405 & ~n3408;
  assign n3410 = ~n3402 & n3409;
  assign n3411 = n3401 & n3410;
  assign n3412 = n3170 & n3411;
  assign n3413 = n3395 & n3412;
  assign n3414 = n3156 & n3413;
  assign n3415 = n3143 & n3414;
  assign n3416 = ~n3392 & n3415;
  assign n3417 = ~n3391 & n3416;
  assign n3418 = n3417 ^ n1807;
  assign n3419 = n3418 ^ x125;
  assign n3420 = n2908 ^ x86;
  assign n3421 = n1884 ^ x68;
  assign n3422 = ~n3420 & n3421;
  assign n3423 = ~n2056 & ~n2648;
  assign n3424 = ~n3078 & ~n3423;
  assign n3425 = n2040 & n3075;
  assign n3426 = ~n2053 & n3425;
  assign n3427 = n2023 & ~n3426;
  assign n3428 = ~n3424 & ~n3427;
  assign n3429 = ~n1952 & n2001;
  assign n3430 = n1954 & n2000;
  assign n3431 = ~n2016 & ~n3430;
  assign n3432 = ~n2038 & ~n3431;
  assign n3433 = ~n2019 & n3089;
  assign n3434 = n1997 & ~n3433;
  assign n3435 = ~n2018 & n3081;
  assign n3436 = ~n2640 & n3435;
  assign n3437 = n2016 & ~n3436;
  assign n3438 = ~n3434 & ~n3437;
  assign n3439 = ~n3432 & n3438;
  assign n3440 = ~n3429 & n3439;
  assign n3441 = n3428 & n3440;
  assign n3442 = n2647 & n3441;
  assign n3443 = n2642 & n3442;
  assign n3444 = ~n2060 & n3443;
  assign n3445 = n3444 ^ x20;
  assign n3446 = n3445 ^ x75;
  assign n3447 = n2895 ^ x69;
  assign n3448 = ~n3446 & n3447;
  assign n3449 = n680 ^ x125;
  assign n3450 = n2364 & n2478;
  assign n3451 = n2468 & ~n2910;
  assign n3452 = ~n3450 & ~n3451;
  assign n3453 = n2366 & n2422;
  assign n3454 = ~n2460 & ~n2464;
  assign n3455 = n2436 & ~n3454;
  assign n3456 = n2436 & ~n2919;
  assign n3457 = n2434 & ~n2475;
  assign n3458 = ~n3456 & ~n3457;
  assign n3459 = ~n2482 & n3454;
  assign n3460 = ~n2473 & n3459;
  assign n3461 = ~n2438 & n3460;
  assign n3462 = n2427 & ~n3461;
  assign n3463 = n2434 & ~n2693;
  assign n3464 = n2366 & n2473;
  assign n3465 = ~n2469 & ~n2910;
  assign n3466 = ~n3464 & ~n3465;
  assign n3467 = ~n3463 & n3466;
  assign n3468 = ~n2433 & n3467;
  assign n3469 = ~n3462 & n3468;
  assign n3470 = n3458 & n3469;
  assign n3471 = ~n2928 & n3470;
  assign n3472 = ~n2431 & n3471;
  assign n3473 = ~n3455 & n3472;
  assign n3474 = ~n3453 & n3473;
  assign n3475 = n3452 & n3474;
  assign n3476 = n2456 & n3475;
  assign n3477 = n3476 ^ x12;
  assign n3478 = n3477 ^ x92;
  assign n3479 = ~n3449 & n3478;
  assign n3480 = n3448 & n3479;
  assign n3481 = n3422 & n3480;
  assign n3482 = n3446 & ~n3447;
  assign n3483 = n3449 & n3478;
  assign n3484 = n3482 & n3483;
  assign n3485 = ~n3420 & ~n3421;
  assign n3486 = n3484 & n3485;
  assign n3487 = ~n3481 & ~n3486;
  assign n3488 = n3420 & n3421;
  assign n3489 = ~n3485 & ~n3488;
  assign n3490 = ~n3446 & ~n3447;
  assign n3491 = ~n3449 & ~n3478;
  assign n3492 = n3490 & n3491;
  assign n3493 = n3449 & ~n3478;
  assign n3494 = n3482 & n3493;
  assign n3495 = ~n3492 & ~n3494;
  assign n3496 = ~n3489 & ~n3495;
  assign n3497 = n3479 & n3490;
  assign n3498 = n3490 & n3493;
  assign n3499 = ~n3497 & ~n3498;
  assign n3500 = n3488 & ~n3499;
  assign n3501 = n3446 & n3447;
  assign n3502 = n3479 & n3501;
  assign n3503 = n3448 & n3493;
  assign n3504 = ~n3502 & ~n3503;
  assign n3505 = n3483 & n3490;
  assign n3506 = ~n3492 & ~n3505;
  assign n3507 = ~n3497 & n3506;
  assign n3508 = ~n3494 & n3507;
  assign n3509 = n3504 & n3508;
  assign n3510 = n3422 & ~n3509;
  assign n3511 = n3448 & n3483;
  assign n3512 = ~n3502 & ~n3511;
  assign n3513 = n3483 & n3501;
  assign n3514 = n3491 & n3501;
  assign n3515 = ~n3513 & ~n3514;
  assign n3516 = n3512 & n3515;
  assign n3517 = n3488 & ~n3516;
  assign n3518 = ~n3480 & ~n3511;
  assign n3519 = n3504 & n3518;
  assign n3520 = n3485 & ~n3519;
  assign n3521 = ~n3517 & ~n3520;
  assign n3522 = ~n3510 & n3521;
  assign n3534 = n3493 & n3501;
  assign n3523 = n3447 ^ n3446;
  assign n3524 = n3523 ^ n3447;
  assign n3525 = n3524 ^ n3478;
  assign n3526 = n3478 ^ n3449;
  assign n3527 = n3526 ^ n3449;
  assign n3528 = n3449 ^ n3447;
  assign n3529 = n3528 ^ n3449;
  assign n3530 = ~n3527 & n3529;
  assign n3531 = n3530 ^ n3449;
  assign n3532 = n3525 & n3531;
  assign n3533 = n3532 ^ n3523;
  assign n3535 = n3534 ^ n3533;
  assign n3536 = n3535 ^ n3534;
  assign n3537 = n3534 ^ n3421;
  assign n3538 = n3537 ^ n3534;
  assign n3539 = n3536 & ~n3538;
  assign n3540 = n3539 ^ n3534;
  assign n3541 = n3420 & n3540;
  assign n3542 = n3541 ^ n3534;
  assign n3543 = n3522 & ~n3542;
  assign n3544 = ~n3500 & n3543;
  assign n3545 = ~n3496 & n3544;
  assign n3546 = n3487 & n3545;
  assign n3547 = n3546 ^ n1770;
  assign n3548 = n3547 ^ x77;
  assign n3549 = ~n3419 & ~n3548;
  assign n3550 = n3390 & n3549;
  assign n3551 = n2512 & n2529;
  assign n3552 = n2324 & n2554;
  assign n3553 = ~n3551 & ~n3552;
  assign n3554 = n2504 & n2521;
  assign n3555 = n2324 & n2509;
  assign n3556 = ~n3554 & ~n3555;
  assign n3557 = n2504 & ~n2545;
  assign n3558 = n3556 & ~n3557;
  assign n3559 = n2323 & n2507;
  assign n3560 = n2514 & n2536;
  assign n3561 = ~n3559 & ~n3560;
  assign n3562 = n2324 & n2553;
  assign n3563 = ~n2516 & ~n2527;
  assign n3564 = ~n2520 & ~n3563;
  assign n3565 = ~n2553 & ~n2557;
  assign n3566 = ~n2521 & n3565;
  assign n3567 = ~n2509 & n3566;
  assign n3568 = n2529 & ~n3567;
  assign n3569 = n2554 ^ n2323;
  assign n3570 = n2533 ^ n2322;
  assign n3571 = n3570 ^ n2533;
  assign n3572 = n2537 & ~n2557;
  assign n3573 = n3572 ^ n2533;
  assign n3574 = ~n3571 & ~n3573;
  assign n3575 = n3574 ^ n2533;
  assign n3576 = n3575 ^ n2554;
  assign n3577 = ~n3569 & n3576;
  assign n3578 = n3577 ^ n3574;
  assign n3579 = n3578 ^ n2533;
  assign n3580 = n3579 ^ n2323;
  assign n3581 = ~n2554 & ~n3580;
  assign n3582 = n3581 ^ n2554;
  assign n3583 = n3582 ^ n2323;
  assign n3584 = ~n3568 & n3583;
  assign n3585 = ~n3564 & n3584;
  assign n3586 = ~n3562 & n3585;
  assign n3587 = n3561 & n3586;
  assign n3588 = n3558 & n3587;
  assign n3589 = n2547 & n3588;
  assign n3590 = n3553 & n3589;
  assign n3591 = n2521 ^ n2322;
  assign n3592 = n3591 ^ n2521;
  assign n3593 = n2533 ^ n2521;
  assign n3594 = n3592 & n3593;
  assign n3595 = n3594 ^ n2521;
  assign n3596 = ~n2323 & n3595;
  assign n3597 = n3590 & ~n3596;
  assign n3598 = ~n2542 & n3597;
  assign n3599 = n3598 ^ n917;
  assign n3600 = n3599 ^ x94;
  assign n3601 = n3550 & ~n3600;
  assign n3602 = ~n3419 & n3548;
  assign n3603 = n3388 & ~n3389;
  assign n3604 = n3602 & n3603;
  assign n3605 = n3419 & n3548;
  assign n3606 = ~n3388 & ~n3389;
  assign n3607 = n3605 & n3606;
  assign n3608 = ~n3604 & ~n3607;
  assign n3609 = n3603 & n3605;
  assign n3610 = n3419 & ~n3548;
  assign n3611 = n3606 & n3610;
  assign n3612 = ~n3609 & ~n3611;
  assign n3613 = n3608 & n3612;
  assign n3614 = n2831 ^ x108;
  assign n3615 = n3600 & ~n3614;
  assign n3616 = ~n3613 & n3615;
  assign n3617 = ~n3600 & ~n3614;
  assign n3618 = n3419 ^ n3389;
  assign n3619 = n3618 ^ n3388;
  assign n3620 = n3619 ^ n3389;
  assign n3621 = n3620 ^ n3548;
  assign n3622 = n3618 ^ n3389;
  assign n3623 = n3618 ^ n3548;
  assign n3624 = ~n3622 & n3623;
  assign n3625 = n3624 ^ n3618;
  assign n3626 = ~n3621 & ~n3625;
  assign n3627 = n3626 ^ n3618;
  assign n3628 = n3617 & ~n3627;
  assign n3629 = n3390 & n3610;
  assign n3630 = n3600 & n3614;
  assign n3631 = ~n3617 & ~n3630;
  assign n3632 = n3629 & ~n3631;
  assign n3633 = ~n3628 & ~n3632;
  assign n3634 = ~n3388 & n3389;
  assign n3635 = n3605 & n3634;
  assign n3636 = n3602 & n3634;
  assign n3637 = n3390 & n3602;
  assign n3638 = ~n3636 & ~n3637;
  assign n3639 = ~n3635 & n3638;
  assign n3640 = n3614 & ~n3639;
  assign n3641 = n3549 & n3634;
  assign n3642 = ~n3629 & ~n3641;
  assign n3643 = ~n3550 & ~n3617;
  assign n3644 = n3642 & n3643;
  assign n3645 = ~n3635 & n3644;
  assign n3646 = n3615 & ~n3645;
  assign n3647 = ~n3600 & n3614;
  assign n3648 = n3549 & n3603;
  assign n3649 = n3612 & ~n3648;
  assign n3650 = n3602 & n3606;
  assign n3651 = n3630 & n3650;
  assign n3652 = n3603 & n3610;
  assign n3653 = n3647 & n3652;
  assign n3654 = ~n3651 & ~n3653;
  assign n3655 = n3649 & n3654;
  assign n3656 = ~n3647 & n3655;
  assign n3657 = n3549 & n3606;
  assign n3658 = ~n3609 & ~n3650;
  assign n3659 = ~n3657 & n3658;
  assign n3660 = ~n3630 & n3659;
  assign n3661 = n3614 & ~n3660;
  assign n3662 = n3654 & ~n3661;
  assign n3663 = ~n3656 & ~n3662;
  assign n3664 = ~n3646 & ~n3663;
  assign n3665 = ~n3640 & n3664;
  assign n3666 = n3633 & n3665;
  assign n3667 = ~n3616 & n3666;
  assign n3668 = ~n3601 & n3667;
  assign n3669 = n3668 ^ n1884;
  assign n3670 = n3669 ^ x67;
  assign n3671 = ~n3265 & ~n3670;
  assign n3672 = ~n2248 & n2309;
  assign n3673 = n2274 & ~n3672;
  assign n3674 = n2172 ^ n2135;
  assign n3675 = n3674 ^ n2207;
  assign n3676 = n3675 ^ n2172;
  assign n3677 = n3676 ^ n2207;
  assign n3678 = n3677 ^ n2242;
  assign n3679 = n2242 ^ n2172;
  assign n3680 = n2207 ^ n2172;
  assign n3681 = ~n3679 & ~n3680;
  assign n3682 = n3681 ^ n2172;
  assign n3683 = ~n3678 & ~n3682;
  assign n3684 = n3683 ^ n3675;
  assign n3685 = ~n2282 & ~n3684;
  assign n3686 = n2304 & ~n3685;
  assign n3687 = ~n3673 & ~n3686;
  assign n3688 = ~n2263 & n2287;
  assign n3689 = n2097 & ~n3688;
  assign n3690 = ~n2252 & ~n2282;
  assign n3691 = n2274 & ~n3690;
  assign n3692 = ~n2097 & ~n2268;
  assign n3693 = ~n2271 & ~n3692;
  assign n3694 = ~n3691 & ~n3693;
  assign n3695 = ~n2246 & ~n2274;
  assign n3696 = n2259 & ~n3695;
  assign n3697 = ~n2248 & ~n2264;
  assign n3698 = n2279 & n3697;
  assign n3699 = ~n2286 & n3698;
  assign n3700 = n2246 & ~n3699;
  assign n3701 = ~n3696 & ~n3700;
  assign n3702 = n3694 & n3701;
  assign n3703 = ~n3689 & n3702;
  assign n3704 = n3687 & n3703;
  assign n3705 = ~n2257 & n3704;
  assign n3706 = ~n2245 & n3705;
  assign n3707 = n3706 ^ n607;
  assign n3708 = n3707 ^ x123;
  assign n3709 = n1950 ^ x96;
  assign n3710 = ~n3708 & ~n3709;
  assign n3711 = n3326 & ~n3344;
  assign n3712 = n3266 & n3349;
  assign n3713 = n3338 & ~n3712;
  assign n3714 = n3330 & ~n3713;
  assign n3715 = ~n3711 & ~n3714;
  assign n3716 = n3325 & ~n3326;
  assign n3717 = n3339 & n3342;
  assign n3718 = n3349 ^ n3290;
  assign n3719 = n3718 ^ n3349;
  assign n3720 = n3362 & ~n3719;
  assign n3721 = n3720 ^ n3349;
  assign n3722 = ~n3717 & ~n3721;
  assign n3723 = ~n3337 & n3722;
  assign n3724 = n3344 & n3723;
  assign n3725 = n3716 & n3724;
  assign n3726 = ~n3333 & ~n3725;
  assign n3727 = n3336 & ~n3372;
  assign n3728 = n3351 & ~n3727;
  assign n3729 = n3327 & ~n3728;
  assign n3730 = ~n3325 & ~n3326;
  assign n3731 = n3336 & n3339;
  assign n3732 = n3722 & ~n3731;
  assign n3733 = n3338 & n3732;
  assign n3734 = n3730 & ~n3733;
  assign n3735 = ~n3729 & ~n3734;
  assign n3736 = n3726 & n3735;
  assign n3737 = n3715 & n3736;
  assign n3738 = n3737 ^ n527;
  assign n3739 = n3738 ^ x114;
  assign n3740 = n3485 & n3498;
  assign n3741 = ~n3494 & ~n3505;
  assign n3742 = n3488 & ~n3741;
  assign n3743 = ~n3740 & ~n3742;
  assign n3744 = n3420 & ~n3421;
  assign n3745 = n3479 & n3482;
  assign n3746 = ~n3494 & ~n3745;
  assign n3747 = n3506 & n3746;
  assign n3748 = n3744 & ~n3747;
  assign n3749 = ~n3503 & n3515;
  assign n3750 = n3422 & ~n3749;
  assign n3751 = ~n3497 & ~n3745;
  assign n3752 = ~n3489 & ~n3751;
  assign n3753 = n3448 & n3491;
  assign n3754 = ~n3511 & ~n3753;
  assign n3755 = n3504 & n3754;
  assign n3756 = n3485 & ~n3755;
  assign n3757 = n3482 & n3491;
  assign n3758 = ~n3484 & ~n3757;
  assign n3759 = n3495 & n3758;
  assign n3760 = n3422 & ~n3759;
  assign n3761 = ~n3756 & ~n3760;
  assign n3762 = ~n3752 & n3761;
  assign n3763 = ~n3488 & n3518;
  assign n3764 = ~n3534 & ~n3753;
  assign n3765 = ~n3744 & n3764;
  assign n3766 = ~n3763 & ~n3765;
  assign n3767 = n3515 & ~n3766;
  assign n3768 = n3420 & ~n3767;
  assign n3769 = n3762 & ~n3768;
  assign n3770 = ~n3750 & n3769;
  assign n3771 = ~n3748 & n3770;
  assign n3772 = n3743 & n3771;
  assign n3773 = n3487 & n3772;
  assign n3774 = n3773 ^ n456;
  assign n3775 = n3774 ^ x113;
  assign n3776 = ~n3739 & ~n3775;
  assign n3777 = n3710 & n3776;
  assign n3778 = ~n3012 & ~n3025;
  assign n3779 = n3028 & ~n3778;
  assign n3780 = n2991 & n3057;
  assign n3781 = ~n2999 & ~n3012;
  assign n3782 = n2897 & ~n3781;
  assign n3783 = ~n3780 & ~n3782;
  assign n3784 = ~n3779 & n3783;
  assign n3785 = ~n3003 & n3784;
  assign n3786 = n2989 & n3025;
  assign n3787 = n2897 & n3057;
  assign n3788 = ~n3786 & ~n3787;
  assign n3789 = ~n2987 & ~n3024;
  assign n3790 = n2991 & ~n3789;
  assign n3791 = n2989 & ~n3036;
  assign n3792 = ~n3006 & ~n3035;
  assign n3793 = n3030 & n3792;
  assign n3794 = n2991 & ~n3793;
  assign n3796 = n2985 ^ n2934;
  assign n3798 = n3796 ^ n2934;
  assign n3799 = n2909 & ~n3798;
  assign n3795 = n2985 ^ n2956;
  assign n3797 = ~n3795 & n3796;
  assign n3800 = n3799 ^ n3797;
  assign n3801 = n3028 & n3800;
  assign n3802 = ~n3794 & ~n3801;
  assign n3803 = ~n3791 & n3802;
  assign n3804 = n3007 ^ n2897;
  assign n3805 = n3007 ^ n2989;
  assign n3806 = n3805 ^ n2989;
  assign n3807 = ~n3001 & ~n3013;
  assign n3808 = ~n2994 & n3807;
  assign n3809 = n3808 ^ n2989;
  assign n3810 = ~n3806 & n3809;
  assign n3811 = n3810 ^ n2989;
  assign n3812 = n3804 & n3811;
  assign n3813 = n3812 ^ n2897;
  assign n3814 = n3803 & ~n3813;
  assign n3815 = ~n3790 & n3814;
  assign n3816 = n3788 & n3815;
  assign n3817 = n2996 & n3816;
  assign n3818 = n3785 & n3817;
  assign n3819 = ~n3061 & n3818;
  assign n3820 = n3819 ^ n294;
  assign n3821 = n3820 ^ x120;
  assign n3822 = n3207 ^ x81;
  assign n3823 = n3821 & n3822;
  assign n3824 = n3777 & n3823;
  assign n3825 = n3708 & ~n3709;
  assign n3826 = ~n3739 & n3775;
  assign n3827 = n3825 & n3826;
  assign n3828 = n3708 & n3709;
  assign n3829 = n3739 & n3775;
  assign n3830 = n3828 & n3829;
  assign n3831 = ~n3827 & ~n3830;
  assign n3832 = ~n3821 & n3822;
  assign n3833 = ~n3831 & n3832;
  assign n3834 = ~n3824 & ~n3833;
  assign n3835 = ~n3708 & n3709;
  assign n3836 = n3829 & n3835;
  assign n3837 = n3823 & n3836;
  assign n3838 = n3826 & n3835;
  assign n3839 = n3739 & ~n3775;
  assign n3840 = n3710 & n3839;
  assign n3841 = ~n3838 & ~n3840;
  assign n3842 = n3823 & ~n3841;
  assign n3843 = n3821 & ~n3822;
  assign n3844 = n3776 & n3828;
  assign n3845 = n3825 & n3839;
  assign n3846 = ~n3844 & ~n3845;
  assign n3847 = n3831 & n3846;
  assign n3848 = n3843 & ~n3847;
  assign n3849 = n3776 & n3835;
  assign n3850 = n3835 & n3839;
  assign n3851 = ~n3840 & ~n3850;
  assign n3852 = ~n3843 & n3851;
  assign n3853 = n3710 & n3829;
  assign n3854 = n3710 & n3826;
  assign n3855 = ~n3853 & ~n3854;
  assign n3856 = ~n3821 & ~n3822;
  assign n3857 = n3855 & ~n3856;
  assign n3858 = ~n3852 & ~n3857;
  assign n3859 = ~n3849 & ~n3858;
  assign n3860 = ~n3836 & n3859;
  assign n3861 = ~n3822 & ~n3860;
  assign n3862 = ~n3848 & ~n3861;
  assign n3863 = ~n3842 & n3862;
  assign n3864 = n3822 ^ n3821;
  assign n3868 = n3776 & n3825;
  assign n3869 = ~n3853 & ~n3868;
  assign n3870 = ~n3850 & ~n3854;
  assign n3871 = ~n3849 & n3870;
  assign n3872 = ~n3840 & n3871;
  assign n3873 = n3869 & n3872;
  assign n3865 = n3739 ^ n3709;
  assign n3866 = n3865 ^ n3775;
  assign n3867 = n3708 & ~n3866;
  assign n3874 = n3873 ^ n3867;
  assign n3875 = n3874 ^ n3867;
  assign n3876 = n3867 ^ n3822;
  assign n3877 = n3876 ^ n3867;
  assign n3878 = ~n3875 & n3877;
  assign n3879 = n3878 ^ n3867;
  assign n3880 = n3864 & n3879;
  assign n3881 = n3880 ^ n3867;
  assign n3882 = n3863 & ~n3881;
  assign n3883 = ~n3837 & n3882;
  assign n3884 = n3834 & n3883;
  assign n3885 = n3884 ^ n680;
  assign n3886 = n3885 ^ x93;
  assign n3887 = n681 & ~n1071;
  assign n3888 = ~n1072 & ~n3887;
  assign n3889 = n1888 & n1893;
  assign n3890 = ~n1911 & ~n3889;
  assign n3891 = ~n3888 & ~n3890;
  assign n3892 = n1917 & n1940;
  assign n3893 = ~n3891 & ~n3892;
  assign n3894 = n1072 & n1906;
  assign n3895 = ~n1907 & n1923;
  assign n3896 = n3887 & ~n3895;
  assign n3897 = ~n3894 & ~n3896;
  assign n3898 = ~n1899 & n1921;
  assign n3899 = n1905 & ~n3898;
  assign n3900 = n1889 ^ n1071;
  assign n3904 = n1895 & n1909;
  assign n3901 = ~n1894 & ~n1918;
  assign n3902 = ~n1907 & n3901;
  assign n3903 = ~n1908 & n3902;
  assign n3905 = n3904 ^ n3903;
  assign n3906 = n3904 ^ n681;
  assign n3907 = n3906 ^ n3904;
  assign n3908 = n3905 & ~n3907;
  assign n3909 = n3908 ^ n3904;
  assign n3910 = n3909 ^ n1889;
  assign n3911 = ~n3900 & ~n3910;
  assign n3912 = n3911 ^ n3908;
  assign n3913 = n3912 ^ n3904;
  assign n3914 = n3913 ^ n1071;
  assign n3915 = ~n1889 & n3914;
  assign n3916 = n3915 ^ n1889;
  assign n3917 = n3916 ^ n1071;
  assign n3918 = ~n3899 & n3917;
  assign n3919 = n3897 & n3918;
  assign n3920 = n3893 & n3919;
  assign n3921 = n3920 ^ n1577;
  assign n3922 = n3921 ^ x98;
  assign n3923 = ~n2522 & n3565;
  assign n3924 = n2324 & ~n3923;
  assign n3925 = ~n2554 & n3565;
  assign n3926 = n2504 & ~n3925;
  assign n3927 = n2512 & ~n2520;
  assign n3928 = n2323 & n2516;
  assign n3929 = ~n3927 & ~n3928;
  assign n3930 = ~n2540 & n2550;
  assign n3931 = n2534 & n3930;
  assign n3932 = ~n2553 & n3931;
  assign n3933 = n2514 & ~n3932;
  assign n3934 = ~n2540 & n3572;
  assign n3935 = ~n2507 & n3934;
  assign n3936 = ~n2512 & n3935;
  assign n3937 = n2529 & ~n3936;
  assign n3938 = ~n3933 & ~n3937;
  assign n3939 = n3929 & n3938;
  assign n3940 = ~n3926 & n3939;
  assign n3941 = ~n3924 & n3940;
  assign n3942 = ~n2511 & n3941;
  assign n3943 = n3556 & n3942;
  assign n3944 = n2548 & n3943;
  assign n3945 = ~n2503 & n3944;
  assign n3946 = n3945 ^ n1411;
  assign n3947 = n3946 ^ x105;
  assign n3948 = ~n3922 & n3947;
  assign n3949 = n2989 & n3029;
  assign n3950 = ~n2994 & ~n3006;
  assign n3951 = n3017 & n3950;
  assign n3952 = ~n2989 & n3951;
  assign n3953 = ~n2897 & ~n3012;
  assign n3954 = ~n3004 & n3953;
  assign n3955 = n3792 & n3954;
  assign n3956 = ~n3011 & ~n3955;
  assign n3957 = ~n3952 & n3956;
  assign n3960 = ~n2999 & ~n3024;
  assign n3958 = n3008 & ~n3035;
  assign n3959 = ~n3016 & n3958;
  assign n3961 = n3960 ^ n3959;
  assign n3962 = n3960 ^ n3028;
  assign n3963 = n3960 & n3962;
  assign n3964 = n3963 ^ n3960;
  assign n3965 = n3961 & n3964;
  assign n3966 = n3965 ^ n3963;
  assign n3967 = n3966 ^ n3960;
  assign n3968 = n3967 ^ n3028;
  assign n3969 = ~n3957 & n3968;
  assign n3970 = n3969 ^ n3957;
  assign n3971 = ~n3949 & ~n3970;
  assign n3972 = ~n3011 & n3031;
  assign n3973 = n3026 & n3807;
  assign n3974 = ~n3007 & n3973;
  assign n3975 = ~n3035 & n3974;
  assign n3976 = ~n3029 & n3975;
  assign n3977 = n2991 & ~n3976;
  assign n3978 = ~n3972 & ~n3977;
  assign n3979 = n3971 & n3978;
  assign n3980 = n3785 & n3979;
  assign n3981 = ~n2988 & n3980;
  assign n3982 = n3981 ^ n2390;
  assign n3983 = n3982 ^ x112;
  assign n3984 = n3512 & n3764;
  assign n3985 = n3744 & ~n3984;
  assign n3986 = ~n3484 & n3506;
  assign n3987 = ~n3745 & n3986;
  assign n3988 = n3422 & ~n3987;
  assign n3989 = ~n3985 & ~n3988;
  assign n3990 = n3504 & ~n3513;
  assign n3991 = ~n3489 & ~n3990;
  assign n3997 = ~n3485 & ~n3757;
  assign n3998 = n3746 & n3997;
  assign n3999 = ~n3498 & n3998;
  assign n3992 = ~n3480 & ~n3514;
  assign n3993 = n3765 & n3992;
  assign n3994 = ~n3514 & n3986;
  assign n3995 = ~n3422 & n3994;
  assign n3996 = ~n3993 & ~n3995;
  assign n4000 = n3999 ^ n3996;
  assign n4001 = n4000 ^ n3996;
  assign n4002 = n3499 & ~n3514;
  assign n4003 = ~n3494 & n4002;
  assign n4004 = ~n3488 & n4003;
  assign n4005 = n4004 ^ n3996;
  assign n4006 = n4005 ^ n3996;
  assign n4007 = ~n4001 & ~n4006;
  assign n4008 = n4007 ^ n3996;
  assign n4009 = ~n3489 & n4008;
  assign n4010 = n4009 ^ n3996;
  assign n4011 = ~n3991 & ~n4010;
  assign n4012 = n3989 & n4011;
  assign n4013 = n3421 ^ n3420;
  assign n4014 = n3480 ^ n3421;
  assign n4015 = n4014 ^ n3480;
  assign n4016 = n3753 ^ n3480;
  assign n4017 = n4015 & n4016;
  assign n4018 = n4017 ^ n3480;
  assign n4019 = ~n4013 & n4018;
  assign n4020 = n4012 & ~n4019;
  assign n4021 = n4020 ^ n1309;
  assign n4022 = n4021 ^ x72;
  assign n4023 = ~n3983 & n4022;
  assign n4024 = n3324 & n3716;
  assign n4025 = n3329 & n3730;
  assign n4026 = ~n4024 & ~n4025;
  assign n4027 = n3290 & ~n4026;
  assign n4028 = n3330 & n3733;
  assign n4029 = ~n3713 & n3730;
  assign n4030 = ~n4028 & ~n4029;
  assign n4031 = n3716 & ~n3728;
  assign n4032 = n3327 & ~n3723;
  assign n4033 = ~n4031 & ~n4032;
  assign n4034 = n4030 & n4033;
  assign n4035 = ~n4027 & n4034;
  assign n4036 = n3344 & n4035;
  assign n4037 = n4036 ^ n1518;
  assign n4038 = n4037 ^ x74;
  assign n4039 = n3070 & n3184;
  assign n4040 = n3138 & ~n3153;
  assign n4041 = n3151 & ~n4040;
  assign n4042 = ~n4039 & ~n4041;
  assign n4043 = n3144 & n3178;
  assign n4044 = ~n3160 & ~n3171;
  assign n4045 = n3164 & ~n4044;
  assign n4046 = ~n4043 & ~n4045;
  assign n4047 = ~n3166 & n3403;
  assign n4048 = n3070 & ~n4047;
  assign n4060 = ~n3166 & ~n3184;
  assign n4061 = ~n3144 & n4060;
  assign n4062 = ~n3135 & n3154;
  assign n4063 = ~n3151 & n4062;
  assign n4064 = ~n4061 & ~n4063;
  assign n4065 = ~n3174 & ~n4064;
  assign n4049 = n3157 ^ n3149;
  assign n4050 = n3164 ^ n3149;
  assign n4051 = n4050 ^ n3164;
  assign n4052 = ~n3070 & ~n3148;
  assign n4053 = n4052 ^ n3164;
  assign n4054 = ~n4051 & n4053;
  assign n4055 = n4054 ^ n3164;
  assign n4056 = ~n4049 & ~n4055;
  assign n4057 = n4056 ^ n3157;
  assign n4058 = ~n3152 & ~n4057;
  assign n4059 = ~n3137 & n4058;
  assign n4066 = n4065 ^ n4059;
  assign n4067 = ~n3183 & n4066;
  assign n4068 = n4067 ^ n4065;
  assign n4069 = ~n3391 & n4068;
  assign n4070 = ~n4048 & n4069;
  assign n4071 = n4046 & n4070;
  assign n4072 = n3395 & n4071;
  assign n4073 = n4042 & n4072;
  assign n4074 = n3163 & n4073;
  assign n4075 = ~n3392 & n4074;
  assign n4076 = n4075 ^ n2419;
  assign n4077 = n4076 ^ x122;
  assign n4078 = n4038 & n4077;
  assign n4079 = n4023 & n4078;
  assign n4080 = n3948 & n4079;
  assign n4081 = ~n3922 & ~n3947;
  assign n4082 = ~n3983 & ~n4022;
  assign n4083 = n4078 & n4082;
  assign n4084 = n3983 & n4022;
  assign n4085 = ~n4038 & ~n4077;
  assign n4086 = n4084 & n4085;
  assign n4087 = ~n4083 & ~n4086;
  assign n4088 = n4081 & ~n4087;
  assign n4089 = ~n4080 & ~n4088;
  assign n4090 = n3922 & ~n3947;
  assign n4091 = n4023 & n4085;
  assign n4092 = n4090 & n4091;
  assign n4093 = n3922 & n3947;
  assign n4094 = n3983 & ~n4022;
  assign n4095 = ~n4038 & n4077;
  assign n4096 = n4094 & n4095;
  assign n4097 = n4093 & n4096;
  assign n4098 = n4038 & ~n4077;
  assign n4099 = n4082 & n4098;
  assign n4100 = n4093 & n4099;
  assign n4101 = ~n4097 & ~n4100;
  assign n4102 = n4078 & n4094;
  assign n4103 = n4081 & n4102;
  assign n4104 = n4023 & n4095;
  assign n4105 = n4085 & n4094;
  assign n4106 = ~n4104 & ~n4105;
  assign n4107 = n4093 & ~n4106;
  assign n4108 = ~n4103 & ~n4107;
  assign n4109 = n4078 & n4084;
  assign n4110 = ~n4079 & ~n4109;
  assign n4111 = ~n4091 & n4110;
  assign n4112 = n4093 & ~n4111;
  assign n4113 = n4084 & n4095;
  assign n4114 = ~n4079 & ~n4113;
  assign n4115 = n4084 & n4098;
  assign n4116 = ~n4091 & ~n4105;
  assign n4117 = ~n4115 & n4116;
  assign n4118 = n4114 & n4117;
  assign n4119 = n4081 & ~n4118;
  assign n4120 = ~n4112 & ~n4119;
  assign n4121 = n4082 & n4095;
  assign n4122 = n3922 & n4121;
  assign n4123 = n4094 & n4098;
  assign n4124 = ~n4109 & ~n4123;
  assign n4125 = ~n4083 & n4124;
  assign n4126 = n3948 & ~n4125;
  assign n4127 = n3947 ^ n3922;
  assign n4128 = n4082 & n4085;
  assign n4129 = ~n4086 & ~n4128;
  assign n4130 = n4127 & ~n4129;
  assign n4131 = ~n4096 & ~n4113;
  assign n4132 = n3948 & ~n4131;
  assign n4133 = n4023 & n4098;
  assign n4134 = n4124 & ~n4133;
  assign n4135 = ~n4102 & n4134;
  assign n4136 = n4090 & ~n4135;
  assign n4137 = ~n4132 & ~n4136;
  assign n4138 = ~n4130 & n4137;
  assign n4139 = ~n4126 & n4138;
  assign n4140 = ~n4122 & n4139;
  assign n4141 = n4120 & n4140;
  assign n4142 = n4108 & n4141;
  assign n4143 = n4101 & n4142;
  assign n4144 = ~n4092 & n4143;
  assign n4145 = n4089 & n4144;
  assign n4146 = n4145 ^ n3477;
  assign n4147 = n4146 ^ x91;
  assign n4148 = n3886 & n4147;
  assign n4149 = n4037 ^ x117;
  assign n4150 = n3149 & ~n3167;
  assign n4151 = n3151 & ~n4150;
  assign n4152 = ~n3166 & n3406;
  assign n4153 = n3164 & ~n4152;
  assign n4154 = ~n4151 & ~n4153;
  assign n4155 = ~n3146 & n3182;
  assign n4156 = n3154 & n4155;
  assign n4157 = n3144 & ~n4156;
  assign n4158 = ~n3157 & ~n3174;
  assign n4159 = n4158 ^ n3070;
  assign n4160 = n4158 ^ n3164;
  assign n4161 = n4160 ^ n3164;
  assign n4162 = n3168 & ~n3178;
  assign n4163 = n4162 ^ n3164;
  assign n4164 = n4161 & n4163;
  assign n4165 = n4164 ^ n3164;
  assign n4166 = ~n4159 & n4165;
  assign n4167 = n4166 ^ n3070;
  assign n4168 = ~n4157 & ~n4167;
  assign n4169 = n4154 & n4168;
  assign n4170 = ~n3202 & n4169;
  assign n4171 = ~n3162 & n4170;
  assign n4172 = n4042 & n4171;
  assign n4173 = ~n3142 & n4172;
  assign n4174 = ~n3392 & n4173;
  assign n4175 = ~n3391 & n4174;
  assign n4176 = n4175 ^ n1557;
  assign n4177 = n4176 ^ x68;
  assign n4178 = ~n4149 & n4177;
  assign n4179 = n2271 & ~n2308;
  assign n4180 = n2097 & ~n4179;
  assign n4181 = ~n2244 & ~n2277;
  assign n4182 = n2261 & n2270;
  assign n4183 = n4181 & n4182;
  assign n4184 = n2246 & ~n4183;
  assign n4185 = ~n4180 & ~n4184;
  assign n4186 = ~n2248 & ~n2282;
  assign n4187 = n2063 & ~n4186;
  assign n4188 = ~n2256 & ~n2282;
  assign n4189 = n2266 & n4188;
  assign n4190 = n2278 & n4189;
  assign n4191 = n2304 & ~n4190;
  assign n4192 = ~n4187 & ~n4191;
  assign n4193 = n4185 & n4192;
  assign n4194 = n2274 ^ n2263;
  assign n4195 = n2263 ^ n2246;
  assign n4196 = n4195 ^ n2246;
  assign n4197 = ~n2252 & ~n2256;
  assign n4198 = ~n2275 & n4197;
  assign n4199 = n2287 & n4198;
  assign n4200 = n4199 ^ n2246;
  assign n4201 = ~n4196 & n4200;
  assign n4202 = n4201 ^ n2246;
  assign n4203 = n4194 & n4202;
  assign n4204 = n4203 ^ n2274;
  assign n4205 = n4193 & ~n4204;
  assign n4206 = n2254 & n4205;
  assign n4207 = ~n2245 & n4206;
  assign n4208 = n4207 ^ n1659;
  assign n4209 = n4208 ^ x85;
  assign n4210 = n3921 ^ x78;
  assign n4211 = ~n4209 & n4210;
  assign n4212 = n2780 & n2808;
  assign n4213 = n2760 & ~n2797;
  assign n4214 = ~n4212 & ~n4213;
  assign n4215 = ~n2784 & n2787;
  assign n4216 = n2639 & ~n2796;
  assign n4217 = ~n4215 & ~n4216;
  assign n4218 = n2765 & ~n2786;
  assign n4219 = n2780 & ~n4218;
  assign n4220 = ~n2803 & n4218;
  assign n4221 = ~n2790 & n4220;
  assign n4222 = n2639 & ~n4221;
  assign n4223 = ~n4219 & ~n4222;
  assign n4224 = ~n2771 & ~n2790;
  assign n4225 = ~n2786 & n4224;
  assign n4226 = ~n2805 & n4225;
  assign n4227 = n2767 & ~n4226;
  assign n4228 = ~n2794 & ~n2805;
  assign n4229 = ~n2767 & n4228;
  assign n4230 = ~n2758 & n2804;
  assign n4231 = ~n2780 & n4230;
  assign n4232 = ~n4229 & ~n4231;
  assign n4233 = ~n2803 & ~n2808;
  assign n4234 = ~n2777 & n4233;
  assign n4235 = ~n2764 & n4234;
  assign n4236 = n2760 & ~n4235;
  assign n4237 = ~n4232 & ~n4236;
  assign n4238 = ~n2795 & n4237;
  assign n4239 = ~n4227 & n4238;
  assign n4240 = n4223 & n4239;
  assign n4241 = n4217 & n4240;
  assign n4242 = n4214 & n4241;
  assign n4243 = ~n2759 & n4242;
  assign n4244 = n4243 ^ n1597;
  assign n4245 = n4244 ^ x67;
  assign n4246 = ~n3505 & n3512;
  assign n4247 = n3485 & ~n4246;
  assign n4248 = ~n3534 & n3758;
  assign n4249 = ~n3497 & n4248;
  assign n4250 = n3422 & ~n4249;
  assign n4251 = ~n4247 & ~n4250;
  assign n4252 = ~n3489 & n3514;
  assign n4253 = ~n3480 & n3504;
  assign n4254 = n3488 & ~n4253;
  assign n4255 = n3422 & n3448;
  assign n4256 = n3488 & ~n3747;
  assign n4257 = ~n4255 & ~n4256;
  assign n4258 = ~n3513 & n3764;
  assign n4259 = ~n3480 & n4258;
  assign n4260 = n3744 & ~n4259;
  assign n4261 = n3506 & n3997;
  assign n4262 = ~n3492 & n3746;
  assign n4263 = ~n3744 & n4262;
  assign n4264 = ~n4261 & ~n4263;
  assign n4265 = ~n3498 & ~n4264;
  assign n4266 = ~n3421 & ~n4265;
  assign n4267 = ~n4260 & ~n4266;
  assign n4268 = n4257 & n4267;
  assign n4269 = ~n4254 & n4268;
  assign n4270 = ~n4252 & n4269;
  assign n4271 = n4251 & n4270;
  assign n4272 = n4271 ^ n1624;
  assign n4273 = n4272 ^ x100;
  assign n4274 = ~n4245 & n4273;
  assign n4275 = n4211 & n4274;
  assign n4276 = n4178 & n4275;
  assign n4277 = ~n4149 & ~n4177;
  assign n4278 = ~n4245 & ~n4273;
  assign n4279 = n4211 & n4278;
  assign n4280 = ~n4209 & ~n4210;
  assign n4281 = n4245 & ~n4273;
  assign n4282 = n4280 & n4281;
  assign n4283 = ~n4279 & ~n4282;
  assign n4284 = n4277 & ~n4283;
  assign n4285 = ~n4276 & ~n4284;
  assign n4286 = n4149 & ~n4177;
  assign n4287 = n4245 & n4273;
  assign n4288 = n4280 & n4287;
  assign n4289 = n4209 & n4210;
  assign n4290 = n4273 & n4289;
  assign n4291 = n4245 & n4290;
  assign n4292 = ~n4288 & ~n4291;
  assign n4293 = n4286 & ~n4292;
  assign n4294 = n4274 & n4280;
  assign n4295 = n4209 & ~n4210;
  assign n4296 = n4274 & n4295;
  assign n4297 = ~n4291 & ~n4296;
  assign n4298 = ~n4294 & n4297;
  assign n4299 = n4178 & ~n4298;
  assign n4300 = n4211 & n4287;
  assign n4301 = n4286 & n4300;
  assign n4302 = n4281 & n4289;
  assign n4303 = n4302 ^ n4149;
  assign n4304 = n4303 ^ n4302;
  assign n4305 = n4211 & n4281;
  assign n4306 = n4278 & n4280;
  assign n4307 = n4278 & n4295;
  assign n4308 = ~n4306 & ~n4307;
  assign n4309 = ~n4305 & n4308;
  assign n4310 = n4309 ^ n4302;
  assign n4311 = n4304 & ~n4310;
  assign n4312 = n4311 ^ n4302;
  assign n4313 = n4177 & n4312;
  assign n4314 = ~n4301 & ~n4313;
  assign n4315 = ~n4149 & n4307;
  assign n4316 = n4278 & n4289;
  assign n4317 = n4277 & n4316;
  assign n4318 = ~n4315 & ~n4317;
  assign n4319 = n4286 & n4296;
  assign n4320 = n4149 & n4177;
  assign n4321 = ~n4245 & n4290;
  assign n4322 = n4287 & n4295;
  assign n4323 = ~n4321 & ~n4322;
  assign n4324 = ~n4282 & n4323;
  assign n4325 = n4281 & n4295;
  assign n4326 = ~n4275 & ~n4325;
  assign n4327 = n4324 & n4326;
  assign n4328 = n4320 & ~n4327;
  assign n4329 = ~n4305 & ~n4325;
  assign n4330 = n4178 & ~n4329;
  assign n4331 = n4294 ^ n4177;
  assign n4334 = ~n4300 & n4323;
  assign n4332 = ~n4302 & ~n4316;
  assign n4333 = ~n4282 & n4332;
  assign n4335 = n4334 ^ n4333;
  assign n4336 = n4334 ^ n4149;
  assign n4337 = n4336 ^ n4334;
  assign n4338 = n4335 & n4337;
  assign n4339 = n4338 ^ n4334;
  assign n4340 = n4339 ^ n4294;
  assign n4341 = n4331 & ~n4340;
  assign n4342 = n4341 ^ n4338;
  assign n4343 = n4342 ^ n4334;
  assign n4344 = n4343 ^ n4177;
  assign n4345 = ~n4294 & ~n4344;
  assign n4346 = n4345 ^ n4294;
  assign n4347 = n4346 ^ n4177;
  assign n4348 = ~n4330 & ~n4347;
  assign n4349 = ~n4328 & n4348;
  assign n4350 = ~n4319 & n4349;
  assign n4351 = n4318 & n4350;
  assign n4352 = n4314 & n4351;
  assign n4353 = ~n4299 & n4352;
  assign n4354 = ~n4293 & n4353;
  assign n4355 = n4285 & n4354;
  assign n4356 = n4355 ^ n2895;
  assign n4357 = n4356 ^ x100;
  assign n4358 = n2767 & n2786;
  assign n4359 = n2639 & ~n2765;
  assign n4360 = ~n4358 & ~n4359;
  assign n4361 = ~n2828 & n4360;
  assign n4362 = ~n2777 & n2809;
  assign n4363 = n2639 & ~n4362;
  assign n4364 = ~n2794 & n2806;
  assign n4365 = ~n2795 & n4364;
  assign n4366 = ~n2762 & n4365;
  assign n4367 = n2767 & ~n4366;
  assign n4368 = ~n4363 & ~n4367;
  assign n4369 = n2772 & ~n2808;
  assign n4370 = ~n2802 & n4228;
  assign n4371 = ~n2775 & n4370;
  assign n4372 = ~n2760 & n4371;
  assign n4373 = ~n2805 & n4231;
  assign n4374 = ~n4372 & ~n4373;
  assign n4375 = n4369 & ~n4374;
  assign n4376 = ~n2784 & n4375;
  assign n4377 = n4376 ^ n2784;
  assign n4378 = n4368 & n4377;
  assign n4379 = n4217 & n4378;
  assign n4380 = n4361 & n4379;
  assign n4381 = n4380 ^ n836;
  assign n4382 = n4381 ^ x84;
  assign n4383 = n4272 ^ x110;
  assign n4384 = ~n4382 & n4383;
  assign n4385 = ~n3356 & n3730;
  assign n4386 = ~n3326 & n3337;
  assign n4387 = ~n3335 & n3345;
  assign n4388 = n3716 & ~n4387;
  assign n4389 = ~n4386 & ~n4388;
  assign n4390 = ~n4385 & n4389;
  assign n4391 = n3326 & ~n3383;
  assign n4392 = n4390 & ~n4391;
  assign n4393 = ~n4027 & n4392;
  assign n4394 = n4393 ^ n1965;
  assign n4395 = n4394 ^ x124;
  assign n4396 = n4176 ^ x101;
  assign n4397 = n4395 & ~n4396;
  assign n4398 = n2897 & ~n3017;
  assign n4399 = ~n3013 & n3038;
  assign n4400 = ~n3016 & n4399;
  assign n4401 = n3028 & ~n4400;
  assign n4402 = ~n4398 & ~n4401;
  assign n4403 = n2991 & ~n3778;
  assign n4404 = ~n3006 & ~n3016;
  assign n4405 = n2989 & ~n4404;
  assign n4406 = ~n2987 & n3030;
  assign n4407 = ~n3012 & n4406;
  assign n4408 = n3028 & ~n4407;
  assign n4409 = n3017 & n3792;
  assign n4410 = n2991 & ~n4409;
  assign n4411 = ~n4408 & ~n4410;
  assign n4412 = n3032 & n3953;
  assign n4413 = ~n2989 & n3030;
  assign n4414 = ~n4412 & ~n4413;
  assign n4415 = ~n3024 & ~n4414;
  assign n4416 = ~n3011 & ~n4415;
  assign n4417 = n4411 & ~n4416;
  assign n4418 = ~n2988 & n4417;
  assign n4419 = ~n4405 & n4418;
  assign n4420 = ~n4403 & n4419;
  assign n4421 = n4402 & n4420;
  assign n4422 = ~n3790 & n4421;
  assign n4423 = n3788 & n4422;
  assign n4424 = ~n3061 & n4423;
  assign n4425 = n4424 ^ n750;
  assign n4426 = n4425 ^ x75;
  assign n4427 = n2504 & n2509;
  assign n4428 = ~n2527 & n2545;
  assign n4429 = ~n2512 & n4428;
  assign n4430 = n2514 & ~n4429;
  assign n4431 = ~n4427 & ~n4430;
  assign n4432 = ~n2520 & ~n2558;
  assign n4433 = ~n2507 & ~n2557;
  assign n4434 = n2324 & ~n4433;
  assign n4435 = n2534 & n3565;
  assign n4436 = n2504 & ~n4435;
  assign n4438 = n2500 ^ n2326;
  assign n4437 = n2363 ^ n2325;
  assign n4439 = n4438 ^ n4437;
  assign n4440 = n4439 ^ n2500;
  assign n4441 = n4438 ^ n2363;
  assign n4442 = n2500 ^ n2363;
  assign n4443 = n4442 ^ n2363;
  assign n4444 = ~n4441 & n4443;
  assign n4445 = n4444 ^ n2363;
  assign n4446 = n4440 & ~n4445;
  assign n4447 = n4446 ^ n4438;
  assign n4448 = n2529 & n4447;
  assign n4449 = ~n4436 & ~n4448;
  assign n4450 = ~n4434 & n4449;
  assign n4451 = ~n4432 & n4450;
  assign n4452 = n4431 & n4451;
  assign n4453 = n3553 & n4452;
  assign n4454 = ~n3596 & n4453;
  assign n4455 = n3558 & n4454;
  assign n4456 = ~n2503 & n4455;
  assign n4457 = ~n2542 & n4456;
  assign n4458 = n4457 ^ n1988;
  assign n4459 = n4458 ^ x86;
  assign n4460 = n4426 & ~n4459;
  assign n4461 = n4397 & n4460;
  assign n4462 = ~n4395 & n4396;
  assign n4463 = n4460 & n4462;
  assign n4464 = ~n4461 & ~n4463;
  assign n4465 = n4384 & ~n4464;
  assign n4466 = n4382 & n4383;
  assign n4467 = n4426 & n4459;
  assign n4468 = n4397 & n4467;
  assign n4469 = n4395 & n4396;
  assign n4470 = n4460 & n4469;
  assign n4471 = ~n4468 & ~n4470;
  assign n4472 = n4466 & ~n4471;
  assign n4473 = ~n4465 & ~n4472;
  assign n4474 = n4462 & n4467;
  assign n4475 = n4466 & n4474;
  assign n4476 = ~n4382 & ~n4383;
  assign n4477 = ~n4426 & ~n4459;
  assign n4478 = n4397 & n4477;
  assign n4479 = n4462 & n4477;
  assign n4480 = ~n4478 & ~n4479;
  assign n4481 = n4476 & ~n4480;
  assign n4482 = ~n4475 & ~n4481;
  assign n4483 = n4461 & n4466;
  assign n4484 = ~n4426 & n4459;
  assign n4485 = n4462 & n4484;
  assign n4486 = ~n4395 & ~n4396;
  assign n4487 = n4484 & n4486;
  assign n4488 = ~n4485 & ~n4487;
  assign n4489 = n4476 & ~n4488;
  assign n4490 = ~n4483 & ~n4489;
  assign n4491 = n4382 & ~n4383;
  assign n4492 = n4460 & n4486;
  assign n4493 = n4467 & n4469;
  assign n4494 = n4467 & n4486;
  assign n4495 = ~n4493 & ~n4494;
  assign n4496 = ~n4492 & n4495;
  assign n4497 = ~n4463 & n4496;
  assign n4498 = n4491 & ~n4497;
  assign n4499 = n4469 & n4484;
  assign n4500 = n4477 & n4486;
  assign n4501 = ~n4499 & ~n4500;
  assign n4502 = n4466 & ~n4501;
  assign n4503 = n4474 & n4476;
  assign n4504 = ~n4470 & ~n4493;
  assign n4505 = n4384 & ~n4504;
  assign n4506 = n4397 & n4484;
  assign n4507 = n4469 & n4477;
  assign n4508 = ~n4487 & ~n4499;
  assign n4509 = ~n4507 & n4508;
  assign n4510 = ~n4506 & n4509;
  assign n4511 = n4491 & ~n4510;
  assign n4512 = ~n4505 & ~n4511;
  assign n4513 = ~n4479 & ~n4506;
  assign n4514 = n4466 & ~n4513;
  assign n4515 = n4492 ^ n4382;
  assign n4516 = n4488 & ~n4499;
  assign n4517 = n4516 ^ n4471;
  assign n4518 = n4516 ^ n4383;
  assign n4519 = n4518 ^ n4516;
  assign n4520 = n4517 & ~n4519;
  assign n4521 = n4520 ^ n4516;
  assign n4522 = n4521 ^ n4492;
  assign n4523 = n4515 & ~n4522;
  assign n4524 = n4523 ^ n4520;
  assign n4525 = n4524 ^ n4516;
  assign n4526 = n4525 ^ n4382;
  assign n4527 = ~n4492 & ~n4526;
  assign n4528 = n4527 ^ n4492;
  assign n4529 = n4528 ^ n4382;
  assign n4530 = ~n4514 & ~n4529;
  assign n4531 = n4512 & n4530;
  assign n4532 = ~n4503 & n4531;
  assign n4533 = ~n4502 & n4532;
  assign n4534 = ~n4498 & n4533;
  assign n4535 = n4490 & n4534;
  assign n4536 = n4482 & n4535;
  assign n4537 = n4473 & n4536;
  assign n4538 = n4537 ^ n3445;
  assign n4539 = n4538 ^ x110;
  assign n4540 = n4357 & n4539;
  assign n4541 = n4148 & n4540;
  assign n4542 = ~n3886 & n4147;
  assign n4543 = n4357 & ~n4539;
  assign n4544 = n4542 & n4543;
  assign n4545 = ~n4541 & ~n4544;
  assign n4546 = n3671 & ~n4545;
  assign n4547 = ~n3265 & n3670;
  assign n4548 = ~n4357 & n4539;
  assign n4549 = n4542 & n4548;
  assign n4550 = n4547 & n4549;
  assign n4551 = n3265 & ~n3670;
  assign n4552 = ~n3886 & ~n4147;
  assign n4553 = ~n4357 & ~n4539;
  assign n4554 = n4552 & n4553;
  assign n4555 = n4551 & n4554;
  assign n4556 = n3265 & n3670;
  assign n4557 = ~n3671 & ~n4556;
  assign n4558 = n4548 & n4552;
  assign n4559 = n3886 & ~n4147;
  assign n4560 = n4553 & n4559;
  assign n4561 = ~n4558 & ~n4560;
  assign n4562 = ~n4557 & ~n4561;
  assign n4563 = ~n4555 & ~n4562;
  assign n4564 = ~n4550 & n4563;
  assign n4565 = n4544 & n4556;
  assign n4566 = n4543 & n4559;
  assign n4567 = n4547 & n4566;
  assign n4568 = ~n4565 & ~n4567;
  assign n4569 = n4548 & n4559;
  assign n4570 = n3671 & n4569;
  assign n4571 = n4551 & n4558;
  assign n4572 = ~n4570 & ~n4571;
  assign n4573 = n4148 & n4548;
  assign n4574 = n4551 & n4573;
  assign n4575 = n4547 & n4554;
  assign n4576 = ~n4574 & ~n4575;
  assign n4577 = n4572 & n4576;
  assign n4578 = n4540 & n4552;
  assign n4579 = ~n4569 & ~n4578;
  assign n4580 = n4551 & ~n4579;
  assign n4581 = n4540 & n4542;
  assign n4582 = n4540 & n4559;
  assign n4583 = ~n4581 & ~n4582;
  assign n4584 = n4148 & n4553;
  assign n4585 = ~n4541 & ~n4584;
  assign n4586 = ~n4578 & n4585;
  assign n4587 = n4583 & n4586;
  assign n4588 = n4547 & ~n4587;
  assign n4589 = ~n4580 & ~n4588;
  assign n4590 = n4543 & n4552;
  assign n4591 = ~n4573 & ~n4590;
  assign n4592 = n3671 & ~n4591;
  assign n4596 = n4583 & ~n4590;
  assign n4593 = n4148 & n4543;
  assign n4594 = ~n4581 & ~n4593;
  assign n4595 = ~n4566 & n4594;
  assign n4597 = n4596 ^ n4595;
  assign n4598 = n4596 ^ n3670;
  assign n4599 = n4598 ^ n4596;
  assign n4600 = n4597 & ~n4599;
  assign n4601 = n4600 ^ n4596;
  assign n4602 = n3265 & ~n4601;
  assign n4603 = ~n4592 & ~n4602;
  assign n4604 = n4589 & n4603;
  assign n4605 = n4577 & n4604;
  assign n4606 = n4542 & n4553;
  assign n4607 = n4606 ^ n4556;
  assign n4608 = n4606 ^ n3671;
  assign n4609 = n4608 ^ n3671;
  assign n4610 = n4573 ^ n3671;
  assign n4611 = ~n4609 & ~n4610;
  assign n4612 = n4611 ^ n3671;
  assign n4613 = n4607 & n4612;
  assign n4614 = n4613 ^ n4556;
  assign n4615 = n4605 & ~n4614;
  assign n4616 = n4568 & n4615;
  assign n4617 = n4564 & n4616;
  assign n4618 = ~n4546 & n4617;
  assign n4619 = n4618 ^ n4272;
  assign n4620 = n4619 ^ x78;
  assign n4621 = n4466 & n4492;
  assign n4622 = n4466 & n4478;
  assign n4623 = n4384 & ~n4513;
  assign n4624 = ~n4622 & ~n4623;
  assign n4625 = ~n4468 & n4509;
  assign n4626 = n4384 & ~n4625;
  assign n4627 = ~n4485 & ~n4494;
  assign n4628 = n4513 & n4627;
  assign n4629 = n4466 & ~n4628;
  assign n4630 = ~n4626 & ~n4629;
  assign n4631 = ~n4463 & ~n4494;
  assign n4632 = ~n4478 & ~n4485;
  assign n4633 = ~n4470 & n4513;
  assign n4634 = n4632 & n4633;
  assign n4635 = n4631 & n4634;
  assign n4636 = ~n4499 & n4635;
  assign n4637 = n4491 & n4636;
  assign n4638 = n4396 ^ n4395;
  assign n4639 = n4638 ^ n4396;
  assign n4640 = n4639 ^ n4459;
  assign n4641 = ~n4426 & ~n4640;
  assign n4642 = n4641 ^ n4638;
  assign n4643 = n4476 & ~n4642;
  assign n4644 = ~n4637 & ~n4643;
  assign n4645 = n4630 & n4644;
  assign n4646 = n4624 & n4645;
  assign n4647 = ~n4621 & n4646;
  assign n4648 = n4473 & n4647;
  assign n4649 = n4648 ^ n2667;
  assign n4650 = n4649 ^ x80;
  assign n4651 = n4081 & n4099;
  assign n4652 = n4090 & n4096;
  assign n4653 = ~n4092 & ~n4652;
  assign n4654 = ~n4086 & n4114;
  assign n4655 = ~n4121 & n4654;
  assign n4656 = ~n4123 & n4655;
  assign n4657 = n4093 & ~n4656;
  assign n4658 = ~n4083 & ~n4115;
  assign n4659 = ~n4104 & ~n4128;
  assign n4660 = ~n4109 & n4659;
  assign n4661 = n4658 & n4660;
  assign n4662 = n4090 & ~n4661;
  assign n4663 = ~n4657 & ~n4662;
  assign n4664 = n4038 ^ n3983;
  assign n4665 = n4022 ^ n3983;
  assign n4666 = n4665 ^ n4077;
  assign n4667 = ~n4664 & n4666;
  assign n4668 = n4081 & n4667;
  assign n4669 = n4106 & n4129;
  assign n4670 = ~n4133 & n4669;
  assign n4671 = ~n4113 & n4670;
  assign n4672 = n3948 & ~n4671;
  assign n4673 = ~n4668 & ~n4672;
  assign n4674 = n4663 & n4673;
  assign n4675 = n4653 & n4674;
  assign n4676 = n4101 & n4675;
  assign n4677 = ~n4651 & n4676;
  assign n4678 = n4089 & n4677;
  assign n4679 = ~n4102 & n4678;
  assign n4680 = n4679 ^ n2716;
  assign n4681 = n4680 ^ x107;
  assign n4682 = n4650 & ~n4681;
  assign n4683 = n3221 & ~n3224;
  assign n4684 = ~n3220 & n4683;
  assign n4685 = n3210 ^ n2571;
  assign n4686 = n4685 ^ n3210;
  assign n4687 = n3210 ^ n2832;
  assign n4688 = n4687 ^ n3210;
  assign n4689 = n4686 & n4688;
  assign n4690 = n4689 ^ n3210;
  assign n4691 = n3064 & n4690;
  assign n4692 = n4691 ^ n3210;
  assign n4693 = ~n4684 & ~n4692;
  assign n4694 = ~n3226 & n4693;
  assign n4695 = n2321 & n4694;
  assign n4696 = n2832 & n3210;
  assign n4697 = ~n3221 & n3224;
  assign n4698 = ~n3229 & ~n4697;
  assign n4699 = ~n4696 & n4698;
  assign n4700 = ~n4684 & n4699;
  assign n4701 = n3241 & ~n4700;
  assign n4702 = ~n4695 & ~n4701;
  assign n4703 = n3224 ^ n3214;
  assign n4704 = ~n3208 & n4703;
  assign n4705 = n4704 ^ n3224;
  assign n4706 = ~n3237 & ~n4705;
  assign n4707 = ~n3226 & n4706;
  assign n4708 = n3219 & ~n4707;
  assign n4709 = n2832 & n3221;
  assign n4710 = ~n3255 & ~n4709;
  assign n4711 = n3227 & n4710;
  assign n4712 = n3254 & ~n4711;
  assign n4713 = ~n4708 & ~n4712;
  assign n4714 = n4702 & n4713;
  assign n4715 = n4714 ^ n2681;
  assign n4716 = n4715 ^ x98;
  assign n4717 = n3387 ^ x70;
  assign n4718 = n4425 ^ x83;
  assign n4719 = ~n4717 & n4718;
  assign n4720 = n2304 & ~n4182;
  assign n4721 = ~n2259 & n4188;
  assign n4722 = ~n2263 & n4721;
  assign n4723 = n2274 & ~n4722;
  assign n4724 = ~n4720 & ~n4723;
  assign n4725 = n2265 & ~n2286;
  assign n4726 = n2246 & ~n4725;
  assign n4727 = ~n2268 & ~n2275;
  assign n4728 = n2097 & ~n4727;
  assign n4729 = n3697 & n4181;
  assign n4730 = n2304 & ~n4729;
  assign n4731 = ~n4728 & ~n4730;
  assign n4732 = n2261 & n4197;
  assign n4733 = n2246 & ~n4732;
  assign n4736 = ~n2264 & ~n2308;
  assign n4737 = ~n2286 & n4736;
  assign n4734 = ~n2244 & ~n2308;
  assign n4735 = n2278 & n4734;
  assign n4738 = n4737 ^ n4735;
  assign n4739 = n4737 ^ n2096;
  assign n4740 = n4739 ^ n4737;
  assign n4741 = n4738 & n4740;
  assign n4742 = n4741 ^ n4737;
  assign n4743 = n2063 & ~n4742;
  assign n4744 = ~n4733 & ~n4743;
  assign n4745 = n4731 & n4744;
  assign n4746 = ~n2245 & n4745;
  assign n4747 = ~n4726 & n4746;
  assign n4748 = n4724 & n4747;
  assign n4749 = ~n2257 & n4748;
  assign n4750 = n2254 & n4749;
  assign n4751 = n4750 ^ n953;
  assign n4752 = n4751 ^ x76;
  assign n4753 = n1886 & n1897;
  assign n4754 = ~n1887 & ~n4753;
  assign n4755 = n1072 & ~n4754;
  assign n4756 = ~n1889 & ~n1920;
  assign n4757 = n1917 & ~n4756;
  assign n4758 = ~n4755 & ~n4757;
  assign n4759 = ~n1894 & ~n1896;
  assign n4760 = n3887 & ~n4759;
  assign n4761 = ~n1899 & ~n1912;
  assign n4762 = n1917 & ~n4761;
  assign n4763 = ~n4760 & ~n4762;
  assign n4764 = ~n1072 & ~n1917;
  assign n4765 = ~n1908 & ~n1918;
  assign n4766 = n4764 & ~n4765;
  assign n4767 = ~n1892 & ~n1907;
  assign n4768 = n1071 & ~n4767;
  assign n4769 = n1913 & ~n1919;
  assign n4770 = n3887 & ~n4769;
  assign n4771 = n1917 & n4753;
  assign n4772 = ~n1912 & ~n4771;
  assign n4773 = ~n1906 & n4772;
  assign n4774 = n1900 & n4773;
  assign n4775 = ~n1917 & n4774;
  assign n4776 = ~n1887 & ~n1892;
  assign n4777 = ~n1896 & n4776;
  assign n4778 = n1917 & ~n4777;
  assign n4779 = ~n4771 & ~n4778;
  assign n4780 = ~n1905 & n4779;
  assign n4781 = ~n4775 & ~n4780;
  assign n4782 = ~n4770 & ~n4781;
  assign n4783 = n1906 ^ n1072;
  assign n4784 = n3887 ^ n1906;
  assign n4785 = n4784 ^ n3887;
  assign n4786 = n1921 & ~n3889;
  assign n4787 = n4786 ^ n3887;
  assign n4788 = ~n4785 & n4787;
  assign n4789 = n4788 ^ n3887;
  assign n4790 = n4783 & n4789;
  assign n4791 = n4790 ^ n1072;
  assign n4792 = n4782 & ~n4791;
  assign n4793 = ~n4768 & n4792;
  assign n4794 = ~n4766 & n4793;
  assign n4795 = n4763 & n4794;
  assign n4796 = n4758 & n4795;
  assign n4797 = n4796 ^ n991;
  assign n4798 = n4797 ^ x126;
  assign n4799 = n4752 & n4798;
  assign n4800 = n4381 ^ x109;
  assign n4801 = n3599 ^ x116;
  assign n4802 = ~n4800 & n4801;
  assign n4803 = n4799 & n4802;
  assign n4804 = n4719 & n4803;
  assign n4805 = n4717 & n4718;
  assign n4806 = ~n4752 & ~n4798;
  assign n4807 = n4800 & ~n4801;
  assign n4808 = n4806 & n4807;
  assign n4809 = n4752 & ~n4798;
  assign n4810 = ~n4800 & ~n4801;
  assign n4811 = n4809 & n4810;
  assign n4812 = ~n4808 & ~n4811;
  assign n4813 = n4805 & ~n4812;
  assign n4814 = ~n4804 & ~n4813;
  assign n4815 = n4806 & n4810;
  assign n4816 = n4807 & n4809;
  assign n4817 = ~n4815 & ~n4816;
  assign n4818 = n4719 & ~n4817;
  assign n4819 = ~n4717 & ~n4718;
  assign n4820 = ~n4752 & n4798;
  assign n4821 = n4801 & n4820;
  assign n4822 = ~n4811 & ~n4816;
  assign n4823 = n4802 & n4809;
  assign n4824 = n4799 & n4810;
  assign n4825 = n4807 & n4820;
  assign n4826 = ~n4824 & ~n4825;
  assign n4827 = ~n4823 & n4826;
  assign n4828 = n4822 & n4827;
  assign n4829 = ~n4821 & n4828;
  assign n4830 = n4819 & ~n4829;
  assign n4831 = n4717 & ~n4718;
  assign n4832 = n4810 & n4820;
  assign n4833 = n4799 & n4807;
  assign n4834 = ~n4832 & ~n4833;
  assign n4835 = n4812 & n4834;
  assign n4836 = n4831 & ~n4835;
  assign n4837 = n4800 & n4801;
  assign n4838 = n4799 & n4837;
  assign n4839 = n4831 & n4838;
  assign n4840 = ~n4805 & ~n4819;
  assign n4841 = n4809 & n4837;
  assign n4842 = n4802 & n4806;
  assign n4843 = ~n4841 & ~n4842;
  assign n4844 = n4840 & ~n4843;
  assign n4845 = ~n4839 & ~n4844;
  assign n4846 = n4820 & n4837;
  assign n4847 = n4719 & n4846;
  assign n4848 = n4806 & n4837;
  assign n4849 = n4802 & n4820;
  assign n4850 = ~n4848 & ~n4849;
  assign n4851 = ~n4824 & ~n4833;
  assign n4852 = n4850 & n4851;
  assign n4853 = n4805 & ~n4852;
  assign n4854 = ~n4847 & ~n4853;
  assign n4855 = n4845 & n4854;
  assign n4856 = ~n4836 & n4855;
  assign n4857 = ~n4830 & n4856;
  assign n4858 = ~n4818 & n4857;
  assign n4859 = n4814 & n4858;
  assign n4860 = n4843 ^ n4717;
  assign n4861 = n4860 ^ n4843;
  assign n4862 = ~n4808 & ~n4832;
  assign n4863 = n4862 ^ n4843;
  assign n4864 = ~n4861 & n4863;
  assign n4865 = n4864 ^ n4843;
  assign n4866 = n4718 & ~n4865;
  assign n4867 = n4859 & ~n4866;
  assign n4868 = n4803 ^ n4717;
  assign n4869 = n4868 ^ n4803;
  assign n4870 = n4838 ^ n4803;
  assign n4871 = ~n4869 & n4870;
  assign n4872 = n4871 ^ n4803;
  assign n4873 = ~n4718 & n4872;
  assign n4874 = n4867 & ~n4873;
  assign n4875 = n4874 ^ n2755;
  assign n4876 = n4875 ^ x97;
  assign n4877 = n4716 & n4876;
  assign n4878 = n4682 & n4877;
  assign n5011 = n3630 & n3657;
  assign n5012 = ~n3648 & ~n3652;
  assign n5013 = ~n3631 & ~n5012;
  assign n5014 = ~n5011 & ~n5013;
  assign n5015 = ~n3607 & ~n3641;
  assign n5016 = n3617 & ~n5015;
  assign n5017 = ~n3604 & n3612;
  assign n5018 = n3647 & ~n5017;
  assign n5019 = n3390 & n3605;
  assign n5020 = ~n3636 & ~n5019;
  assign n5021 = ~n3641 & n5020;
  assign n5022 = ~n3550 & n5021;
  assign n5023 = n3647 & ~n5022;
  assign n5024 = ~n3629 & n3639;
  assign n5025 = ~n3648 & n5024;
  assign n5026 = n3608 & n5025;
  assign n5027 = ~n3657 & n5026;
  assign n5028 = n3615 & ~n5027;
  assign n5029 = ~n5023 & ~n5028;
  assign n5030 = n3610 & n3634;
  assign n5031 = ~n3637 & ~n5030;
  assign n5032 = n3550 & n3630;
  assign n5033 = ~n3635 & ~n5019;
  assign n5034 = n5033 ^ n3609;
  assign n5035 = n5033 ^ n3630;
  assign n5036 = n5035 ^ n3630;
  assign n5037 = n3643 ^ n3630;
  assign n5038 = ~n5036 & n5037;
  assign n5039 = n5038 ^ n3630;
  assign n5040 = ~n5034 & ~n5039;
  assign n5041 = n5040 ^ n3609;
  assign n5042 = ~n5032 & ~n5041;
  assign n5043 = n5031 & n5042;
  assign n5044 = ~n3631 & ~n5043;
  assign n5045 = n5029 & ~n5044;
  assign n5046 = ~n5018 & n5045;
  assign n5047 = ~n5016 & n5046;
  assign n5048 = n5014 & n5047;
  assign n5049 = n3654 & n5048;
  assign n5050 = n5049 ^ n2637;
  assign n5051 = n5050 ^ x104;
  assign n4879 = n3707 ^ x65;
  assign n4880 = n4021 ^ x121;
  assign n4881 = n4879 & ~n4880;
  assign n4882 = n1071 & n1908;
  assign n4883 = ~n1895 & n1905;
  assign n4884 = ~n4882 & ~n4883;
  assign n4885 = ~n1892 & n1909;
  assign n4886 = n3887 & ~n4885;
  assign n4887 = ~n1906 & n3902;
  assign n4888 = n1917 & ~n4887;
  assign n4889 = ~n4886 & ~n4888;
  assign n4890 = ~n1072 & ~n4771;
  assign n4891 = n4756 & n4773;
  assign n4892 = ~n4890 & ~n4891;
  assign n4893 = n1913 & ~n3889;
  assign n4894 = ~n1899 & n4893;
  assign n4895 = n4764 & ~n4894;
  assign n4896 = ~n4892 & ~n4895;
  assign n4897 = n4889 & n4896;
  assign n4898 = n4764 ^ n1896;
  assign n4899 = n4898 ^ n1896;
  assign n4900 = n1919 ^ n1896;
  assign n4901 = n4899 & n4900;
  assign n4902 = n4901 ^ n1896;
  assign n4903 = n4897 & ~n4902;
  assign n4904 = n4884 & n4903;
  assign n4905 = n4758 & n4904;
  assign n4906 = n4905 ^ n1375;
  assign n4907 = n4906 ^ x97;
  assign n4908 = n3820 ^ x107;
  assign n4909 = n4907 & n4908;
  assign n4910 = ~n2784 & ~n4225;
  assign n4911 = ~n2787 & ~n2805;
  assign n4912 = n2760 & ~n4911;
  assign n4913 = n2796 & n2806;
  assign n4914 = n2780 & ~n4913;
  assign n4915 = ~n4912 & ~n4914;
  assign n4916 = ~n4910 & n4915;
  assign n4917 = ~n2769 & n2804;
  assign n4918 = ~n2787 & n4917;
  assign n4919 = n2639 & ~n4918;
  assign n4920 = ~n2775 & n4234;
  assign n4921 = ~n2758 & n4920;
  assign n4922 = n2767 & ~n4921;
  assign n4923 = ~n4919 & ~n4922;
  assign n4924 = n4916 & n4923;
  assign n4925 = n4214 & n4924;
  assign n4926 = n4361 & n4925;
  assign n4927 = ~n2759 & n4926;
  assign n4928 = n4927 ^ n1339;
  assign n4929 = n4928 ^ x90;
  assign n4930 = n3946 ^ x80;
  assign n4931 = n4929 & n4930;
  assign n4932 = n4909 & n4931;
  assign n4933 = n4907 & ~n4908;
  assign n4934 = ~n4929 & n4930;
  assign n4935 = n4933 & n4934;
  assign n4936 = ~n4932 & ~n4935;
  assign n4937 = n4881 & ~n4936;
  assign n4938 = ~n4879 & n4880;
  assign n4939 = n4909 & ~n4930;
  assign n4940 = n4929 & n4939;
  assign n4941 = ~n4907 & ~n4930;
  assign n4942 = ~n4908 & n4941;
  assign n4943 = ~n4929 & n4942;
  assign n4944 = ~n4940 & ~n4943;
  assign n4945 = n4938 & ~n4944;
  assign n4946 = ~n4937 & ~n4945;
  assign n4947 = n4881 & n4943;
  assign n4948 = n4931 & n4933;
  assign n4949 = ~n4907 & n4931;
  assign n4950 = n4908 & n4949;
  assign n4951 = ~n4948 & ~n4950;
  assign n4952 = n4938 & ~n4951;
  assign n4953 = ~n4947 & ~n4952;
  assign n4954 = n4879 & n4880;
  assign n4955 = ~n4908 & n4949;
  assign n4956 = n4954 & n4955;
  assign n4957 = n4950 & n4954;
  assign n4958 = ~n4956 & ~n4957;
  assign n4959 = ~n4929 & n4939;
  assign n4960 = n4881 & n4959;
  assign n4961 = ~n4879 & ~n4880;
  assign n4962 = ~n4951 & n4961;
  assign n4963 = ~n4960 & ~n4962;
  assign n4964 = ~n4881 & ~n4938;
  assign n4965 = ~n4907 & n4934;
  assign n4966 = n4908 & n4965;
  assign n4967 = ~n4935 & ~n4966;
  assign n4968 = ~n4930 & n4933;
  assign n4969 = n4929 & n4968;
  assign n4970 = n4929 & n4942;
  assign n4971 = ~n4959 & ~n4970;
  assign n4972 = ~n4969 & n4971;
  assign n4973 = ~n4940 & n4972;
  assign n4974 = ~n4961 & n4973;
  assign n4975 = n4908 & n4941;
  assign n4976 = ~n4929 & n4975;
  assign n4977 = ~n4969 & ~n4976;
  assign n4978 = ~n4940 & n4977;
  assign n4979 = ~n4954 & ~n4970;
  assign n4980 = ~n4972 & ~n4979;
  assign n4981 = n4978 & ~n4980;
  assign n4982 = ~n4974 & ~n4981;
  assign n4983 = n4967 & ~n4982;
  assign n4984 = n4964 & n4983;
  assign n4985 = n4984 ^ n4964;
  assign n4986 = n4963 & ~n4985;
  assign n4987 = ~n4929 & n4968;
  assign n4988 = n4929 & n4975;
  assign n4989 = ~n4987 & ~n4988;
  assign n4990 = n4989 ^ n4938;
  assign n4991 = n4989 ^ n4881;
  assign n4992 = n4991 ^ n4881;
  assign n4993 = n4909 & n4934;
  assign n4994 = ~n4908 & n4965;
  assign n4995 = ~n4993 & ~n4994;
  assign n4996 = n4995 ^ n4881;
  assign n4997 = n4992 & n4996;
  assign n4998 = n4997 ^ n4881;
  assign n4999 = ~n4990 & n4998;
  assign n5000 = n4999 ^ n4938;
  assign n5001 = n4986 & ~n5000;
  assign n5002 = n4958 & n5001;
  assign n5003 = n4953 & n5002;
  assign n5004 = ~n4955 & ~n4966;
  assign n5005 = n4881 & n5004;
  assign n5006 = n5005 ^ n4881;
  assign n5007 = n5003 & ~n5006;
  assign n5008 = n4946 & n5007;
  assign n5009 = n5008 ^ n2600;
  assign n5010 = n5009 ^ x65;
  assign n5052 = n5051 ^ n5010;
  assign n5053 = n4878 & ~n5052;
  assign n5054 = n4682 & ~n4716;
  assign n5055 = ~n4876 & n5054;
  assign n5056 = n5010 & ~n5051;
  assign n5057 = n5055 & n5056;
  assign n5058 = n5010 & n5051;
  assign n5059 = n4681 & n4716;
  assign n5060 = ~n4876 & n5059;
  assign n5061 = n4650 & n5060;
  assign n5062 = n5058 & n5061;
  assign n5063 = ~n5010 & n5051;
  assign n5064 = n4878 & n5063;
  assign n5065 = ~n5062 & ~n5064;
  assign n5066 = ~n4681 & ~n4716;
  assign n5067 = ~n4650 & ~n4876;
  assign n5068 = n5066 & n5067;
  assign n5069 = n5058 & n5068;
  assign n5070 = n4681 & ~n4716;
  assign n5071 = n4876 & n5070;
  assign n5072 = ~n4650 & n5071;
  assign n5073 = n4681 & n4877;
  assign n5074 = n4650 & n5073;
  assign n5075 = ~n5072 & ~n5074;
  assign n5076 = n5056 & ~n5075;
  assign n5077 = ~n5069 & ~n5076;
  assign n5078 = n4876 & n5066;
  assign n5079 = ~n4650 & n5078;
  assign n5080 = ~n4681 & n4877;
  assign n5081 = ~n4650 & n5080;
  assign n5082 = ~n5079 & ~n5081;
  assign n5083 = n5063 & ~n5082;
  assign n5084 = n4876 & n5054;
  assign n5085 = n4716 & n5067;
  assign n5086 = ~n4681 & n5085;
  assign n5087 = ~n5084 & ~n5086;
  assign n5088 = n5058 & ~n5087;
  assign n5089 = ~n5083 & ~n5088;
  assign n5090 = ~n5010 & ~n5051;
  assign n5091 = n4682 & n4716;
  assign n5092 = ~n4876 & n5091;
  assign n5093 = ~n5086 & ~n5092;
  assign n5094 = n5090 & ~n5093;
  assign n5095 = ~n5079 & ~n5092;
  assign n5096 = n5056 & ~n5095;
  assign n5097 = n5059 & n5067;
  assign n5098 = ~n4876 & n5070;
  assign n5099 = n4650 & n5098;
  assign n5100 = ~n5097 & ~n5099;
  assign n5101 = n5063 & ~n5100;
  assign n5102 = ~n5096 & ~n5101;
  assign n5103 = n5061 & n5090;
  assign n5104 = n5063 & ~n5075;
  assign n5105 = n5056 & n5086;
  assign n5106 = n4650 & n5071;
  assign n5107 = ~n4650 & n5073;
  assign n5108 = n5067 & n5070;
  assign n5109 = ~n5107 & ~n5108;
  assign n5110 = ~n5106 & n5109;
  assign n5111 = ~n5052 & ~n5110;
  assign n5112 = ~n5105 & ~n5111;
  assign n5113 = ~n5104 & n5112;
  assign n5114 = ~n5103 & n5113;
  assign n5115 = n5102 & n5114;
  assign n5116 = ~n5094 & n5115;
  assign n5117 = n5089 & n5116;
  assign n5118 = ~n5081 & ~n5108;
  assign n5119 = n5118 ^ n5055;
  assign n5120 = n5119 ^ n5055;
  assign n5121 = n5055 ^ n5051;
  assign n5122 = n5121 ^ n5055;
  assign n5123 = ~n5120 & ~n5122;
  assign n5124 = n5123 ^ n5055;
  assign n5125 = n5010 & n5124;
  assign n5126 = n5125 ^ n5055;
  assign n5127 = n5117 & ~n5126;
  assign n5128 = n5077 & n5127;
  assign n5129 = n5065 & n5128;
  assign n5130 = ~n5057 & n5129;
  assign n5131 = ~n5053 & n5130;
  assign n5132 = n5131 ^ n4381;
  assign n5133 = n5132 ^ x83;
  assign n5134 = ~n4620 & n5133;
  assign n5135 = n3836 & n3856;
  assign n5136 = n3777 & n3843;
  assign n5137 = ~n5135 & ~n5136;
  assign n5138 = ~n3838 & ~n3853;
  assign n5139 = n3856 & ~n5138;
  assign n5140 = n3840 & ~n3864;
  assign n5141 = ~n5139 & ~n5140;
  assign n5142 = n3843 & ~n3871;
  assign n5143 = ~n3854 & ~n3868;
  assign n5144 = n3823 & ~n5143;
  assign n5145 = n3825 & n3829;
  assign n5146 = n3826 & n3828;
  assign n5147 = ~n3845 & ~n5146;
  assign n5148 = ~n5145 & n5147;
  assign n5149 = ~n3827 & n5148;
  assign n5150 = n3832 & ~n5149;
  assign n5151 = n3830 & n3843;
  assign n5152 = ~n3777 & ~n3849;
  assign n5153 = n3832 & ~n5152;
  assign n5154 = ~n5151 & ~n5153;
  assign n5155 = ~n3850 & ~n3853;
  assign n5156 = n3832 & ~n5155;
  assign n5157 = n3843 & ~n5148;
  assign n5158 = ~n5156 & ~n5157;
  assign n5159 = n5154 & n5158;
  assign n5160 = ~n5150 & n5159;
  assign n5161 = n3828 & n3839;
  assign n5162 = ~n3844 & ~n5161;
  assign n5163 = n3831 & n5162;
  assign n5164 = n5163 ^ n3822;
  assign n5165 = n5164 ^ n5163;
  assign n5166 = n3708 & n3826;
  assign n5167 = n5162 & ~n5166;
  assign n5168 = n5167 ^ n5163;
  assign n5169 = ~n5165 & n5168;
  assign n5170 = n5169 ^ n5163;
  assign n5171 = ~n3864 & ~n5170;
  assign n5172 = n5160 & ~n5171;
  assign n5173 = ~n5144 & n5172;
  assign n5174 = ~n5142 & n5173;
  assign n5175 = n5141 & n5174;
  assign n5176 = n5137 & n5175;
  assign n5177 = ~n3837 & n5176;
  assign n5178 = n5177 ^ n2865;
  assign n5179 = n5178 ^ x92;
  assign n5180 = n4356 ^ x78;
  assign n5181 = n5179 & ~n5180;
  assign n5182 = n3264 ^ x75;
  assign n5183 = ~n4840 & ~n4862;
  assign n5184 = n4719 & ~n4851;
  assign n5185 = ~n5183 & ~n5184;
  assign n5186 = ~n4821 & ~n4842;
  assign n5187 = n4831 & ~n5186;
  assign n5188 = ~n4803 & ~n4846;
  assign n5189 = ~n4823 & n5188;
  assign n5190 = ~n4848 & n5189;
  assign n5191 = ~n4816 & n5190;
  assign n5192 = n4819 & ~n5191;
  assign n5193 = ~n5187 & ~n5192;
  assign n5194 = n4827 & ~n4838;
  assign n5195 = n4805 & ~n5194;
  assign n5196 = n4719 & ~n5190;
  assign n5197 = ~n4815 & n4822;
  assign n5198 = ~n4833 & n5197;
  assign n5199 = n4831 & ~n5198;
  assign n5200 = ~n5196 & ~n5199;
  assign n5201 = ~n5195 & n5200;
  assign n5202 = n5193 & n5201;
  assign n5203 = n5185 & n5202;
  assign n5204 = ~n4866 & n5203;
  assign n5205 = ~n4873 & n5204;
  assign n5206 = n5205 ^ n2984;
  assign n5207 = n5206 ^ x124;
  assign n5208 = n5182 & ~n5207;
  assign n5209 = n4949 & n4961;
  assign n5210 = n4935 & n4938;
  assign n5211 = ~n5209 & ~n5210;
  assign n5212 = ~n4936 & n4961;
  assign n5213 = ~n4948 & ~n4993;
  assign n5214 = ~n4966 & n5213;
  assign n5215 = n4880 & ~n5214;
  assign n5216 = n4978 & ~n4987;
  assign n5217 = n4954 & ~n5216;
  assign n5218 = n4971 & ~n4987;
  assign n5219 = ~n4940 & n5218;
  assign n5220 = n4961 & ~n5219;
  assign n5221 = ~n5217 & ~n5220;
  assign n5222 = n4938 & n4941;
  assign n5223 = n4930 ^ n4929;
  assign n5224 = n5223 ^ n4907;
  assign n5225 = n5224 ^ n4908;
  assign n5226 = n5225 ^ n4930;
  assign n5227 = n4930 ^ n4908;
  assign n5228 = n5227 ^ n4908;
  assign n5229 = n4908 ^ n4907;
  assign n5230 = n5229 ^ n4908;
  assign n5231 = n5228 & ~n5230;
  assign n5232 = n5231 ^ n4908;
  assign n5233 = n5226 & ~n5232;
  assign n5234 = n5233 ^ n5223;
  assign n5235 = n4881 & n5234;
  assign n5236 = ~n5222 & ~n5235;
  assign n5237 = n5221 & n5236;
  assign n5238 = ~n5006 & n5237;
  assign n5239 = ~n5215 & n5238;
  assign n5240 = ~n5212 & n5239;
  assign n5241 = n5211 & n5240;
  assign n5242 = ~n4956 & n5241;
  assign n5243 = n5242 ^ n2955;
  assign n5244 = n5243 ^ x109;
  assign n5245 = n4081 & n4096;
  assign n5246 = n4113 & n4127;
  assign n5247 = n4090 & n4123;
  assign n5248 = ~n5246 & ~n5247;
  assign n5249 = ~n5245 & n5248;
  assign n5250 = ~n4102 & n4658;
  assign n5251 = n4660 & n5250;
  assign n5252 = ~n4099 & n5251;
  assign n5253 = n5252 ^ n4086;
  assign n5254 = n5253 ^ n4086;
  assign n5255 = n4086 ^ n3947;
  assign n5256 = n5255 ^ n4086;
  assign n5257 = ~n5254 & n5256;
  assign n5258 = n5257 ^ n4086;
  assign n5259 = ~n3922 & n5258;
  assign n5260 = n5259 ^ n4086;
  assign n5261 = ~n4123 & ~n4133;
  assign n5262 = ~n4079 & n5261;
  assign n5263 = n5262 ^ n4110;
  assign n5264 = n4127 ^ n3947;
  assign n5265 = n5262 ^ n3947;
  assign n5266 = ~n5264 & n5265;
  assign n5267 = n5266 ^ n3947;
  assign n5268 = n5263 & n5267;
  assign n5269 = n5268 ^ n4110;
  assign n5270 = ~n4083 & n5269;
  assign n5271 = n5270 ^ n3947;
  assign n5272 = n5271 ^ n5270;
  assign n5273 = ~n4133 & n4655;
  assign n5274 = n5273 ^ n5270;
  assign n5275 = n5274 ^ n5270;
  assign n5276 = ~n5272 & ~n5275;
  assign n5277 = n5276 ^ n5270;
  assign n5278 = ~n3922 & ~n5277;
  assign n5279 = n5278 ^ n5270;
  assign n5280 = ~n5260 & n5279;
  assign n5281 = n4108 & n5280;
  assign n5282 = n4653 & n5281;
  assign n5283 = n5249 & n5282;
  assign n5284 = ~n4651 & n5283;
  assign n5285 = ~n4097 & n5284;
  assign n5286 = n5285 ^ n2933;
  assign n5287 = n5286 ^ x102;
  assign n5288 = n5244 & ~n5287;
  assign n5289 = n5208 & n5288;
  assign n5290 = n5181 & n5289;
  assign n5291 = n5179 & n5180;
  assign n5292 = ~n5182 & n5207;
  assign n5293 = ~n5244 & ~n5287;
  assign n5294 = n5292 & n5293;
  assign n5295 = n5182 & n5207;
  assign n5296 = n5288 & n5295;
  assign n5297 = ~n5294 & ~n5296;
  assign n5298 = n5291 & ~n5297;
  assign n5299 = ~n5290 & ~n5298;
  assign n5300 = ~n5179 & ~n5180;
  assign n5301 = n5244 & n5287;
  assign n5302 = n5295 & n5301;
  assign n5303 = ~n5182 & ~n5207;
  assign n5304 = n5301 & n5303;
  assign n5305 = ~n5302 & ~n5304;
  assign n5306 = n5300 & ~n5305;
  assign n5307 = ~n5244 & n5287;
  assign n5308 = n5295 & n5307;
  assign n5309 = n5292 & n5307;
  assign n5310 = ~n5308 & ~n5309;
  assign n5311 = n5181 & ~n5310;
  assign n5312 = ~n5179 & n5180;
  assign n5313 = n5293 & n5295;
  assign n5314 = n5288 & n5303;
  assign n5315 = ~n5313 & ~n5314;
  assign n5316 = n5312 & ~n5315;
  assign n5317 = ~n5311 & ~n5316;
  assign n5318 = n5208 & n5307;
  assign n5319 = n5300 & n5318;
  assign n5320 = n5296 & n5312;
  assign n5321 = ~n5319 & ~n5320;
  assign n5322 = n5303 & n5307;
  assign n5323 = n5300 & n5322;
  assign n5324 = n5208 & n5293;
  assign n5325 = ~n5181 & ~n5312;
  assign n5326 = n5324 & n5325;
  assign n5327 = ~n5323 & ~n5326;
  assign n5328 = n5292 & n5301;
  assign n5329 = n5208 & n5301;
  assign n5330 = ~n5328 & ~n5329;
  assign n5331 = n5310 & n5330;
  assign n5332 = ~n5314 & n5331;
  assign n5333 = n5291 & ~n5332;
  assign n5334 = n5293 & n5303;
  assign n5335 = n5297 & ~n5334;
  assign n5336 = ~n5328 & n5335;
  assign n5337 = n5181 & ~n5336;
  assign n5338 = ~n5333 & ~n5337;
  assign n5339 = n5318 & ~n5325;
  assign n5340 = ~n5294 & ~n5313;
  assign n5341 = ~n5329 & n5340;
  assign n5342 = n5300 & ~n5341;
  assign n5343 = n5288 & n5292;
  assign n5344 = ~n5322 & ~n5343;
  assign n5345 = n5330 & n5344;
  assign n5346 = n5312 & ~n5345;
  assign n5347 = ~n5342 & ~n5346;
  assign n5348 = ~n5339 & n5347;
  assign n5349 = n5338 & n5348;
  assign n5350 = n5327 & n5349;
  assign n5351 = n5321 & n5350;
  assign n5352 = n5317 & n5351;
  assign n5353 = ~n5306 & n5352;
  assign n5354 = n5299 & n5353;
  assign n5355 = n5354 ^ n4425;
  assign n5356 = n5355 ^ x110;
  assign n5357 = n4680 ^ x114;
  assign n5358 = ~n4840 & n4841;
  assign n5359 = n4719 & ~n4822;
  assign n5360 = ~n5358 & ~n5359;
  assign n5361 = n4800 ^ n4798;
  assign n5362 = n5361 ^ n4752;
  assign n5363 = n4801 & n5362;
  assign n5364 = n4831 & n5363;
  assign n5365 = ~n4815 & ~n4825;
  assign n5366 = ~n4819 & n5365;
  assign n5367 = ~n4840 & ~n5366;
  assign n5368 = n5367 ^ n4805;
  assign n5369 = n5367 ^ n4812;
  assign n5370 = n5369 ^ n4812;
  assign n5371 = ~n4808 & n4826;
  assign n5372 = ~n4842 & n5371;
  assign n5373 = n5372 ^ n4812;
  assign n5374 = n5370 & ~n5373;
  assign n5375 = n5374 ^ n4812;
  assign n5376 = n5368 & n5375;
  assign n5377 = n5376 ^ n4805;
  assign n5378 = ~n5364 & ~n5377;
  assign n5379 = n5360 & n5378;
  assign n5380 = n4819 & ~n5189;
  assign n5386 = ~n4821 & ~n4823;
  assign n5381 = ~n4803 & n4850;
  assign n5382 = n4719 & ~n5381;
  assign n5383 = n4834 & ~n5382;
  assign n5384 = ~n4816 & n5383;
  assign n5385 = ~n4842 & n5384;
  assign n5387 = n5386 ^ n5385;
  assign n5388 = n5387 ^ n5386;
  assign n5389 = n5386 ^ n4819;
  assign n5390 = n5389 ^ n5386;
  assign n5391 = ~n5388 & ~n5390;
  assign n5392 = n5391 ^ n5386;
  assign n5393 = ~n4805 & ~n5392;
  assign n5394 = n5393 ^ n5386;
  assign n5395 = ~n5380 & n5394;
  assign n5396 = n5379 & n5395;
  assign n5397 = n5396 ^ n2171;
  assign n5398 = n5397 ^ x105;
  assign n5399 = ~n5357 & n5398;
  assign n5400 = ~n3844 & n5147;
  assign n5401 = ~n3836 & n5400;
  assign n5402 = n3856 & ~n5401;
  assign n5403 = ~n3822 & ~n3869;
  assign n5404 = ~n3864 & ~n3870;
  assign n5405 = n5147 & n5162;
  assign n5406 = n3823 & ~n5405;
  assign n5407 = ~n5404 & ~n5406;
  assign n5408 = ~n5145 & ~n5161;
  assign n5409 = n3841 & n5408;
  assign n5410 = n3832 & ~n5409;
  assign n5411 = ~n3838 & n3846;
  assign n5412 = ~n3777 & n5411;
  assign n5413 = ~n3850 & n5412;
  assign n5414 = n3843 & ~n5413;
  assign n5415 = ~n5410 & ~n5414;
  assign n5416 = n5407 & n5415;
  assign n5417 = n5154 & n5416;
  assign n5418 = ~n5403 & n5417;
  assign n5419 = ~n5402 & n5418;
  assign n5420 = n3834 & n5419;
  assign n5421 = ~n3837 & n5420;
  assign n5422 = n5421 ^ n3124;
  assign n5423 = n5422 ^ x74;
  assign n5424 = n4286 & n4305;
  assign n5425 = ~n4149 & n4300;
  assign n5426 = n4286 & n4306;
  assign n5427 = ~n5425 & ~n5426;
  assign n5428 = ~n4149 & ~n4332;
  assign n5429 = ~n4294 & ~n4322;
  assign n5430 = n4308 & n5429;
  assign n5431 = n4178 & ~n5430;
  assign n5432 = ~n5428 & ~n5431;
  assign n5433 = ~n4302 & n4326;
  assign n5434 = ~n4296 & n5433;
  assign n5435 = n4286 & ~n5434;
  assign n5436 = ~n4288 & n4297;
  assign n5437 = n4277 & ~n5436;
  assign n5438 = ~n4316 & n4324;
  assign n5439 = ~n4288 & ~n4306;
  assign n5440 = ~n4300 & n5439;
  assign n5441 = ~n4279 & n5440;
  assign n5442 = n5438 & n5441;
  assign n5443 = n4320 & ~n5442;
  assign n5444 = ~n5437 & ~n5443;
  assign n5445 = ~n5435 & n5444;
  assign n5446 = n5432 & n5445;
  assign n5447 = n5427 & n5446;
  assign n5448 = ~n4293 & n5447;
  assign n5449 = ~n5424 & n5448;
  assign n5450 = n4285 & n5449;
  assign n5451 = n5450 ^ n2095;
  assign n5452 = n5451 ^ x64;
  assign n5453 = ~n5423 & n5452;
  assign n5454 = ~n4461 & n4495;
  assign n5455 = n4476 & ~n5454;
  assign n5456 = ~n4384 & ~n4491;
  assign n5457 = ~n4500 & ~n4507;
  assign n5458 = n4488 & n5457;
  assign n5459 = ~n5456 & ~n5458;
  assign n5460 = ~n5455 & ~n5459;
  assign n5461 = n4480 & n4508;
  assign n5462 = n4466 & ~n5461;
  assign n5463 = ~n4470 & n4631;
  assign n5464 = ~n4506 & n5463;
  assign n5465 = n4384 & ~n5464;
  assign n5466 = ~n4492 & ~n4499;
  assign n5467 = n4476 & ~n5466;
  assign n5468 = n4471 & ~n4621;
  assign n5469 = ~n4506 & n5468;
  assign n5470 = ~n4463 & n5469;
  assign n5471 = ~n4468 & ~n4492;
  assign n5472 = ~n4463 & n5471;
  assign n5473 = n4466 & ~n5472;
  assign n5474 = ~n4491 & ~n5473;
  assign n5475 = ~n5470 & ~n5474;
  assign n5476 = ~n5467 & ~n5475;
  assign n5477 = ~n5465 & n5476;
  assign n5478 = n4482 & n5477;
  assign n5479 = ~n5462 & n5478;
  assign n5480 = n5460 & n5479;
  assign n5481 = ~n4503 & n5480;
  assign n5482 = n5481 ^ n3100;
  assign n5483 = n5482 ^ x81;
  assign n5484 = n5050 ^ x120;
  assign n5485 = ~n5483 & n5484;
  assign n5486 = n5453 & n5485;
  assign n5487 = n5399 & n5486;
  assign n5488 = n5357 & ~n5398;
  assign n5489 = n5423 & ~n5452;
  assign n5490 = n5485 & n5489;
  assign n5491 = n5488 & n5490;
  assign n5492 = ~n5357 & ~n5398;
  assign n5493 = n5423 & n5452;
  assign n5494 = n5483 & n5484;
  assign n5495 = n5493 & n5494;
  assign n5496 = n5485 & n5493;
  assign n5497 = n5483 & ~n5484;
  assign n5498 = n5453 & n5497;
  assign n5499 = ~n5496 & ~n5498;
  assign n5500 = ~n5495 & n5499;
  assign n5501 = n5492 & ~n5500;
  assign n5502 = ~n5491 & ~n5501;
  assign n5503 = n5489 & n5497;
  assign n5504 = n5492 & n5503;
  assign n5505 = n5357 & n5398;
  assign n5506 = ~n5483 & ~n5484;
  assign n5507 = n5493 & n5506;
  assign n5508 = n5505 & n5507;
  assign n5509 = n5489 & n5494;
  assign n5510 = ~n5423 & ~n5452;
  assign n5511 = n5506 & n5510;
  assign n5512 = ~n5509 & ~n5511;
  assign n5513 = n5399 & ~n5512;
  assign n5514 = ~n5508 & ~n5513;
  assign n5515 = ~n5504 & n5514;
  assign n5516 = n5494 & n5510;
  assign n5517 = n5489 & n5506;
  assign n5518 = ~n5516 & ~n5517;
  assign n5519 = n5505 & ~n5518;
  assign n5520 = n5493 & n5497;
  assign n5521 = ~n5496 & ~n5520;
  assign n5522 = n5399 & ~n5521;
  assign n5523 = ~n5519 & ~n5522;
  assign n5524 = n5495 & n5505;
  assign n5525 = n5488 & n5503;
  assign n5526 = ~n5524 & ~n5525;
  assign n5527 = ~n5507 & n5518;
  assign n5528 = n5399 & ~n5527;
  assign n5529 = n5453 & n5494;
  assign n5530 = ~n5520 & ~n5529;
  assign n5531 = n5499 & n5530;
  assign n5532 = ~n5511 & n5531;
  assign n5533 = n5488 & ~n5532;
  assign n5534 = ~n5528 & ~n5533;
  assign n5535 = n5497 & n5510;
  assign n5536 = n5485 & n5510;
  assign n5537 = n5453 & n5506;
  assign n5538 = ~n5536 & ~n5537;
  assign n5539 = ~n5535 & n5538;
  assign n5540 = n5539 ^ n5492;
  assign n5541 = n5539 ^ n5505;
  assign n5542 = n5541 ^ n5505;
  assign n5543 = n5505 ^ n5490;
  assign n5544 = n5542 & ~n5543;
  assign n5545 = n5544 ^ n5505;
  assign n5546 = ~n5540 & n5545;
  assign n5547 = n5546 ^ n5492;
  assign n5548 = n5534 & ~n5547;
  assign n5549 = n5526 & n5548;
  assign n5550 = n5523 & n5549;
  assign n5551 = n5515 & n5550;
  assign n5552 = n5502 & n5551;
  assign n5553 = ~n5487 & n5552;
  assign n5554 = n5486 ^ n5398;
  assign n5555 = n5554 ^ n5486;
  assign n5556 = n5509 ^ n5486;
  assign n5557 = n5555 & n5556;
  assign n5558 = n5557 ^ n5486;
  assign n5559 = n5357 & n5558;
  assign n5560 = n5553 & ~n5559;
  assign n5561 = n5560 ^ n4176;
  assign n5562 = n5561 ^ x69;
  assign n5563 = ~n5356 & ~n5562;
  assign n5564 = n4649 ^ x66;
  assign n5565 = n5286 ^ x113;
  assign n5566 = ~n5564 & n5565;
  assign n5567 = ~n4149 & n4325;
  assign n5568 = ~n4290 & n4298;
  assign n5569 = ~n4305 & n5568;
  assign n5570 = n4277 & ~n5569;
  assign n5571 = ~n5567 & ~n5570;
  assign n5572 = ~n4296 & n5441;
  assign n5573 = n4178 & ~n5572;
  assign n5574 = n4292 & n5429;
  assign n5575 = ~n4316 & n5574;
  assign n5576 = n4320 & ~n5575;
  assign n5577 = n4297 & ~n4325;
  assign n5578 = ~n4290 & n5577;
  assign n5579 = ~n4279 & n5578;
  assign n5580 = ~n4282 & n5579;
  assign n5581 = n4286 & ~n5580;
  assign n5582 = ~n5576 & ~n5581;
  assign n5583 = ~n5573 & n5582;
  assign n5584 = n5571 & n5583;
  assign n5585 = n4314 & n5584;
  assign n5586 = ~n5424 & n5585;
  assign n5587 = n4285 & n5586;
  assign n5588 = n5587 ^ n3322;
  assign n5589 = n5588 ^ x99;
  assign n5590 = n5178 ^ x90;
  assign n5591 = n5589 & n5590;
  assign n5592 = n5009 ^ x73;
  assign n5593 = n5591 & ~n5592;
  assign n5594 = ~n3600 & ~n5031;
  assign n5595 = ~n3550 & ~n3635;
  assign n5596 = ~n3631 & ~n5595;
  assign n5597 = ~n3609 & n3642;
  assign n5598 = n3630 & ~n5597;
  assign n5599 = n5015 & n5020;
  assign n5600 = ~n3657 & n5599;
  assign n5601 = n3647 & ~n5600;
  assign n5602 = ~n5598 & ~n5601;
  assign n5603 = ~n3604 & ~n3652;
  assign n5604 = ~n3615 & ~n3630;
  assign n5605 = ~n5603 & ~n5604;
  assign n5606 = ~n3617 & n3654;
  assign n5607 = ~n3650 & n3655;
  assign n5608 = ~n5606 & ~n5607;
  assign n5609 = ~n3611 & ~n3657;
  assign n5610 = n5609 ^ n5599;
  assign n5611 = n5599 ^ n3615;
  assign n5612 = n5599 & n5611;
  assign n5613 = n5612 ^ n5599;
  assign n5614 = n5610 & n5613;
  assign n5615 = n5614 ^ n5612;
  assign n5616 = n5615 ^ n5599;
  assign n5617 = n5616 ^ n3615;
  assign n5618 = ~n5608 & n5617;
  assign n5619 = n5618 ^ n5608;
  assign n5620 = ~n5605 & ~n5619;
  assign n5621 = n5602 & n5620;
  assign n5622 = ~n5596 & n5621;
  assign n5623 = ~n5594 & n5622;
  assign n5624 = n5623 ^ n3288;
  assign n5625 = n5624 ^ x72;
  assign n5626 = n5590 & n5625;
  assign n5627 = ~n5589 & n5592;
  assign n5628 = ~n5626 & n5627;
  assign n5629 = n5625 ^ n5592;
  assign n5630 = ~n5590 & n5629;
  assign n5631 = ~n5628 & ~n5630;
  assign n5632 = ~n5593 & n5631;
  assign n5633 = n5566 & n5632;
  assign n5634 = n5564 & n5565;
  assign n5635 = n5591 & n5592;
  assign n5636 = ~n5589 & n5630;
  assign n5637 = ~n5635 & ~n5636;
  assign n5638 = ~n5589 & ~n5592;
  assign n5639 = n5590 & n5638;
  assign n5640 = ~n5625 & n5639;
  assign n5641 = ~n5590 & n5625;
  assign n5642 = n5627 & n5641;
  assign n5643 = ~n5592 & n5625;
  assign n5644 = ~n5626 & ~n5643;
  assign n5645 = n5589 & ~n5644;
  assign n5646 = ~n5642 & ~n5645;
  assign n5647 = ~n5640 & n5646;
  assign n5648 = n5637 & n5647;
  assign n5649 = n5634 & ~n5648;
  assign n5650 = ~n5633 & ~n5649;
  assign n5651 = n5564 & ~n5565;
  assign n5652 = n5629 ^ n5592;
  assign n5653 = n5625 ^ n5590;
  assign n5654 = n5653 ^ n5592;
  assign n5655 = n5654 ^ n5592;
  assign n5656 = n5655 ^ n5592;
  assign n5657 = n5652 & n5656;
  assign n5658 = n5657 ^ n5592;
  assign n5659 = ~n5589 & n5658;
  assign n5660 = n5659 ^ n5654;
  assign n5661 = n5651 & ~n5660;
  assign n5662 = ~n5564 & ~n5565;
  assign n5663 = ~n5590 & ~n5625;
  assign n5664 = n5589 & n5663;
  assign n5665 = n5626 & n5627;
  assign n5666 = ~n5664 & ~n5665;
  assign n5667 = n5647 & n5666;
  assign n5668 = n5662 & ~n5667;
  assign n5669 = ~n5661 & ~n5668;
  assign n5670 = n5650 & n5669;
  assign n5671 = n5670 ^ n4394;
  assign n5672 = n5671 ^ x92;
  assign n5673 = ~n3225 & n4710;
  assign n5674 = n5673 ^ n2320;
  assign n5675 = n5674 ^ n5673;
  assign n5676 = n5673 ^ n4700;
  assign n5677 = n5675 & ~n5676;
  assign n5678 = n5677 ^ n5673;
  assign n5679 = ~n1951 & ~n5678;
  assign n5680 = n4706 ^ n2320;
  assign n5681 = n5680 ^ n4706;
  assign n5682 = n4706 ^ n4694;
  assign n5683 = n5681 & n5682;
  assign n5684 = n5683 ^ n4706;
  assign n5685 = n1951 & ~n5684;
  assign n5686 = ~n5679 & ~n5685;
  assign n5687 = ~n3226 & n5686;
  assign n5688 = n5687 ^ n2134;
  assign n5689 = n5688 ^ x101;
  assign n5690 = n4881 & n4966;
  assign n5691 = n4938 & ~n5004;
  assign n5692 = n4950 & n4961;
  assign n5693 = ~n4969 & ~n4988;
  assign n5694 = n4951 & n5693;
  assign n5695 = ~n4993 & n5694;
  assign n5696 = n4881 & ~n5695;
  assign n5697 = ~n5692 & ~n5696;
  assign n5698 = ~n4932 & ~n4994;
  assign n5699 = n4964 & ~n5698;
  assign n5700 = n4977 & n4989;
  assign n5701 = ~n4880 & n5700;
  assign n5702 = ~n4976 & ~n4987;
  assign n5703 = ~n4961 & n5702;
  assign n5704 = ~n5700 & ~n5703;
  assign n5705 = n4964 & n5704;
  assign n5706 = n4971 & ~n5705;
  assign n5707 = ~n5701 & ~n5706;
  assign n5708 = ~n5699 & ~n5707;
  assign n5709 = n5697 & n5708;
  assign n5710 = n4940 ^ n4935;
  assign n5711 = n5710 ^ n4935;
  assign n5712 = n4935 ^ n4879;
  assign n5713 = n5712 ^ n4935;
  assign n5714 = n5711 & n5713;
  assign n5715 = n5714 ^ n4935;
  assign n5716 = n4880 & n5715;
  assign n5717 = n5716 ^ n4935;
  assign n5718 = n5709 & ~n5717;
  assign n5719 = ~n4945 & n5718;
  assign n5720 = ~n5691 & n5719;
  assign n5721 = n4953 & n5720;
  assign n5722 = ~n4956 & n5721;
  assign n5723 = ~n5690 & n5722;
  assign n5724 = n5723 ^ n1499;
  assign n5725 = n5724 ^ x83;
  assign n5726 = n5689 & ~n5725;
  assign n5727 = ~n3838 & ~n3850;
  assign n5728 = n3823 & ~n5727;
  assign n5729 = n3870 & n5412;
  assign n5730 = n3832 & ~n5729;
  assign n5731 = ~n5728 & ~n5730;
  assign n5732 = ~n3849 & ~n3868;
  assign n5733 = n3856 & ~n5732;
  assign n5734 = n3841 & n5401;
  assign n5735 = n3843 & ~n5734;
  assign n5736 = ~n3839 & n3869;
  assign n5737 = ~n3829 & n5736;
  assign n5738 = ~n3856 & n5737;
  assign n5739 = n3823 & ~n3869;
  assign n5740 = n5163 & ~n5739;
  assign n5741 = ~n5738 & ~n5740;
  assign n5742 = ~n3864 & n5741;
  assign n5743 = ~n5735 & ~n5742;
  assign n5744 = ~n5733 & n5743;
  assign n5745 = n5731 & n5744;
  assign n5746 = n5137 & n5745;
  assign n5747 = n3834 & n5746;
  assign n5748 = ~n3854 & n5747;
  assign n5749 = n5748 ^ n2362;
  assign n5750 = n5749 ^ x118;
  assign n5751 = n4476 & n4636;
  assign n5752 = ~n4507 & n4631;
  assign n5753 = n5752 ^ n4383;
  assign n5754 = n5753 ^ n5752;
  assign n5755 = n4633 & n5457;
  assign n5756 = ~n4461 & n5755;
  assign n5757 = n5756 ^ n5752;
  assign n5758 = ~n5754 & n5757;
  assign n5759 = n5758 ^ n5752;
  assign n5760 = n4382 & ~n5759;
  assign n5761 = ~n5751 & ~n5760;
  assign n5762 = n4495 ^ n4384;
  assign n5763 = n4495 ^ n4491;
  assign n5764 = n5763 ^ n4491;
  assign n5765 = n4632 ^ n4491;
  assign n5766 = n5764 & n5765;
  assign n5767 = n5766 ^ n4491;
  assign n5768 = ~n5762 & n5767;
  assign n5769 = n5768 ^ n4384;
  assign n5770 = n5761 & ~n5769;
  assign n5771 = n4624 & n5770;
  assign n5772 = ~n4502 & n5771;
  assign n5773 = n4473 & n5772;
  assign n5774 = n5773 ^ n2062;
  assign n5775 = n5774 ^ x125;
  assign n5776 = n5750 & n5775;
  assign n5777 = n3922 & n4099;
  assign n5778 = n4127 & ~n5250;
  assign n5779 = ~n5777 & ~n5778;
  assign n5780 = n4106 & n4110;
  assign n5781 = n4081 & ~n5780;
  assign n5782 = ~n4096 & n4116;
  assign n5783 = n3948 & ~n5782;
  assign n5784 = ~n5781 & ~n5783;
  assign n5785 = n4090 & n4121;
  assign n5786 = n4134 & n4659;
  assign n5787 = ~n4113 & n5786;
  assign n5788 = n4093 & ~n5787;
  assign n5789 = ~n5785 & ~n5788;
  assign n5790 = n5784 & n5789;
  assign n5791 = n5779 & n5790;
  assign n5792 = n5249 & n5791;
  assign n5793 = ~n4651 & n5792;
  assign n5794 = ~n4092 & n5793;
  assign n5795 = ~n4097 & n5794;
  assign n5796 = n4089 & n5795;
  assign n5797 = n5796 ^ n2499;
  assign n5798 = n5797 ^ x69;
  assign n5799 = n4717 & ~n4834;
  assign n5800 = ~n4811 & ~n4825;
  assign n5801 = n4862 & n5800;
  assign n5802 = n4819 & ~n5801;
  assign n5803 = ~n4824 & ~n4848;
  assign n5804 = ~n4821 & n5803;
  assign n5805 = ~n4838 & n5804;
  assign n5806 = n4719 & ~n5805;
  assign n5807 = ~n4841 & n5365;
  assign n5808 = n4850 & n5807;
  assign n5809 = n4831 & ~n5808;
  assign n5810 = n4805 & ~n5189;
  assign n5811 = ~n4833 & ~n5810;
  assign n5812 = ~n4823 & n5811;
  assign n5813 = ~n4842 & n5812;
  assign n5814 = ~n4840 & ~n5813;
  assign n5815 = ~n5809 & ~n5814;
  assign n5816 = ~n5806 & n5815;
  assign n5817 = ~n4818 & n5816;
  assign n5818 = ~n4873 & n5817;
  assign n5819 = ~n5802 & n5818;
  assign n5820 = ~n5799 & n5819;
  assign n5821 = n4814 & n5820;
  assign n5822 = n5821 ^ n1070;
  assign n5823 = n5822 ^ x84;
  assign n5824 = n5798 & n5823;
  assign n5825 = n5776 & n5824;
  assign n5826 = n5750 & ~n5775;
  assign n5827 = ~n5798 & n5823;
  assign n5828 = n5826 & n5827;
  assign n5829 = ~n5825 & ~n5828;
  assign n5830 = n5726 & ~n5829;
  assign n5831 = n5689 & n5725;
  assign n5832 = ~n5750 & ~n5775;
  assign n5833 = ~n5798 & ~n5823;
  assign n5834 = n5832 & n5833;
  assign n5835 = n5776 & n5833;
  assign n5836 = ~n5834 & ~n5835;
  assign n5837 = n5831 & ~n5836;
  assign n5838 = n5726 & n5835;
  assign n5839 = ~n5689 & n5725;
  assign n5840 = n5825 & n5839;
  assign n5841 = ~n5750 & n5775;
  assign n5842 = n5798 & ~n5823;
  assign n5843 = n5841 & n5842;
  assign n5844 = n5726 & n5843;
  assign n5845 = ~n5840 & ~n5844;
  assign n5846 = n5776 & n5842;
  assign n5847 = ~n5689 & n5846;
  assign n5848 = n5776 & n5827;
  assign n5849 = n5827 & n5832;
  assign n5850 = ~n5848 & ~n5849;
  assign n5851 = n5839 & ~n5850;
  assign n5852 = ~n5847 & ~n5851;
  assign n5853 = n5826 & n5833;
  assign n5854 = ~n5726 & ~n5839;
  assign n5855 = n5853 & ~n5854;
  assign n5856 = n5824 & n5826;
  assign n5857 = n5824 & n5841;
  assign n5858 = ~n5856 & ~n5857;
  assign n5859 = ~n5834 & n5858;
  assign n5860 = n5726 & ~n5859;
  assign n5861 = ~n5855 & ~n5860;
  assign n5862 = n5824 & n5832;
  assign n5863 = ~n5857 & ~n5862;
  assign n5864 = n5829 & n5863;
  assign n5865 = n5831 & ~n5864;
  assign n5866 = n5833 & n5841;
  assign n5867 = n5826 & n5842;
  assign n5868 = ~n5866 & ~n5867;
  assign n5869 = n5854 & ~n5868;
  assign n5870 = ~n5865 & ~n5869;
  assign n5871 = ~n5689 & ~n5725;
  assign n5872 = n5832 & n5842;
  assign n5873 = n5827 & n5841;
  assign n5874 = ~n5862 & ~n5873;
  assign n5875 = n5850 & n5874;
  assign n5876 = ~n5872 & n5875;
  assign n5877 = n5871 & ~n5876;
  assign n5878 = ~n5843 & ~n5866;
  assign n5879 = ~n5862 & n5878;
  assign n5880 = n5839 & ~n5879;
  assign n5881 = ~n5877 & ~n5880;
  assign n5882 = n5870 & n5881;
  assign n5883 = n5861 & n5882;
  assign n5884 = n5852 & n5883;
  assign n5885 = n5845 & n5884;
  assign n5886 = ~n5838 & n5885;
  assign n5887 = ~n5837 & n5886;
  assign n5888 = ~n5830 & n5887;
  assign n5889 = n5888 ^ n4458;
  assign n5890 = n5889 ^ x117;
  assign n5891 = ~n5672 & n5890;
  assign n5892 = n5563 & n5891;
  assign n5893 = n5134 & n5892;
  assign n5894 = n4620 & n5133;
  assign n5895 = n5356 & ~n5562;
  assign n5896 = n5672 & n5890;
  assign n5897 = n5895 & n5896;
  assign n5898 = n5894 & n5897;
  assign n5899 = n5891 & n5895;
  assign n5900 = n5356 & n5562;
  assign n5901 = ~n5672 & ~n5890;
  assign n5902 = n5900 & n5901;
  assign n5903 = ~n5899 & ~n5902;
  assign n5904 = n5894 & ~n5903;
  assign n5905 = n4620 & ~n5133;
  assign n5906 = n5672 & ~n5890;
  assign n5907 = n5900 & n5906;
  assign n5908 = n5895 & n5901;
  assign n5909 = ~n5907 & ~n5908;
  assign n5910 = n5905 & ~n5909;
  assign n5911 = ~n5904 & ~n5910;
  assign n5912 = ~n5898 & n5911;
  assign n5913 = n5563 & n5901;
  assign n5914 = n5894 & n5913;
  assign n5915 = n5133 ^ n4620;
  assign n5916 = n5891 & n5900;
  assign n5917 = ~n5897 & ~n5916;
  assign n5918 = n5915 & ~n5917;
  assign n5919 = ~n5356 & n5562;
  assign n5920 = n5906 & n5919;
  assign n5921 = ~n5908 & ~n5920;
  assign n5922 = ~n5902 & n5921;
  assign n5923 = n5134 & ~n5922;
  assign n5924 = ~n5918 & ~n5923;
  assign n5925 = n5891 & n5919;
  assign n5926 = ~n5907 & ~n5925;
  assign n5927 = n5894 & ~n5926;
  assign n5928 = n5896 & n5919;
  assign n5929 = ~n5913 & ~n5920;
  assign n5930 = ~n5928 & n5929;
  assign n5931 = ~n5892 & n5930;
  assign n5932 = n5905 & ~n5931;
  assign n5933 = ~n5927 & ~n5932;
  assign n5934 = n5924 & n5933;
  assign n5945 = n5563 & n5906;
  assign n5946 = n5901 & n5919;
  assign n5947 = ~n5945 & ~n5946;
  assign n5935 = n5890 ^ n5562;
  assign n5936 = n5890 ^ n5356;
  assign n5937 = n5936 ^ n5356;
  assign n5938 = n5672 ^ n5356;
  assign n5939 = n5938 ^ n5356;
  assign n5940 = n5937 & ~n5939;
  assign n5941 = n5940 ^ n5356;
  assign n5942 = n5935 & n5941;
  assign n5943 = n5930 & ~n5942;
  assign n5944 = ~n5925 & n5943;
  assign n5948 = n5947 ^ n5944;
  assign n5949 = n5948 ^ n5947;
  assign n5950 = n5947 ^ n4620;
  assign n5951 = n5950 ^ n5947;
  assign n5952 = n5949 & ~n5951;
  assign n5953 = n5952 ^ n5947;
  assign n5954 = ~n5133 & ~n5953;
  assign n5955 = n5954 ^ n5947;
  assign n5956 = n5934 & n5955;
  assign n5957 = ~n5914 & n5956;
  assign n5958 = n5912 & n5957;
  assign n5959 = ~n5893 & n5958;
  assign n5960 = n5959 ^ n5774;
  assign n5961 = n5960 ^ x115;
  assign n5962 = n5063 & n5074;
  assign n5963 = ~n5062 & ~n5962;
  assign n5964 = n5056 & n5068;
  assign n5965 = ~n5103 & ~n5964;
  assign n5966 = ~n5052 & n5099;
  assign n5967 = n5058 & ~n5075;
  assign n5968 = ~n5966 & ~n5967;
  assign n5969 = n5010 ^ n4650;
  assign n5970 = n5969 ^ n5010;
  assign n5971 = n5090 ^ n5010;
  assign n5972 = ~n5970 & ~n5971;
  assign n5973 = n5972 ^ n5010;
  assign n5974 = n5071 & ~n5973;
  assign n5975 = n5968 & ~n5974;
  assign n5976 = ~n5097 & ~n5107;
  assign n5977 = n5063 & ~n5976;
  assign n5978 = ~n5081 & ~n5092;
  assign n5979 = n5056 & ~n5978;
  assign n5980 = n5058 & n5079;
  assign n5981 = n5063 & n5068;
  assign n5982 = ~n5980 & ~n5981;
  assign n5983 = ~n5055 & n5095;
  assign n5984 = n5063 & ~n5983;
  assign n5985 = ~n5072 & n5976;
  assign n5986 = ~n5106 & n5985;
  assign n5987 = n5056 & ~n5986;
  assign n5988 = ~n5984 & ~n5987;
  assign n5989 = ~n5086 & ~n5108;
  assign n5990 = n5058 & ~n5989;
  assign n5991 = ~n5081 & n5087;
  assign n5992 = n5090 & ~n5991;
  assign n5993 = ~n5990 & ~n5992;
  assign n5994 = n5988 & n5993;
  assign n5995 = n5982 & n5994;
  assign n5996 = ~n5053 & n5995;
  assign n5997 = ~n5979 & n5996;
  assign n5998 = ~n5977 & n5997;
  assign n5999 = n5975 & n5998;
  assign n6000 = n5965 & n5999;
  assign n6001 = n5963 & n6000;
  assign n6002 = ~n5057 & n6001;
  assign n6003 = n6002 ^ n2831;
  assign n6004 = n6003 ^ x74;
  assign n6005 = n5399 & n5537;
  assign n6006 = n5503 & n5505;
  assign n6007 = ~n6005 & ~n6006;
  assign n6008 = n5399 & n5490;
  assign n6009 = n5492 & n5509;
  assign n6010 = ~n6008 & ~n6009;
  assign n6011 = n5488 & n5535;
  assign n6012 = n5492 & n5520;
  assign n6013 = ~n6011 & ~n6012;
  assign n6014 = ~n5517 & ~n5536;
  assign n6015 = n5492 & ~n6014;
  assign n6016 = ~n5529 & ~n5535;
  assign n6017 = n5399 & ~n6016;
  assign n6018 = ~n6015 & ~n6017;
  assign n6019 = ~n5492 & ~n5505;
  assign n6020 = ~n5486 & n5499;
  assign n6021 = ~n6019 & ~n6020;
  assign n6022 = ~n5511 & ~n5516;
  assign n6023 = ~n5490 & ~n5498;
  assign n6024 = ~n5507 & n6023;
  assign n6025 = n6022 & n6024;
  assign n6026 = ~n5495 & n6025;
  assign n6027 = n5488 & ~n6026;
  assign n6028 = ~n6021 & ~n6027;
  assign n6029 = n6018 & n6028;
  assign n6030 = n6013 & n6029;
  assign n6031 = n5523 & n6030;
  assign n6032 = n6010 & n6031;
  assign n6033 = n5515 & n6032;
  assign n6034 = n6007 & n6033;
  assign n6035 = ~n5559 & n6034;
  assign n6036 = n6035 ^ n3207;
  assign n6037 = n6036 ^ x122;
  assign n6038 = n6004 & ~n6037;
  assign n6039 = n5291 & n5318;
  assign n6040 = n5289 & n5312;
  assign n6041 = ~n6039 & ~n6040;
  assign n6042 = n5181 & n5304;
  assign n6043 = n5244 ^ n5182;
  assign n6044 = n6043 ^ n5207;
  assign n6045 = n5207 & n5287;
  assign n6046 = n6044 & n6045;
  assign n6047 = n6046 ^ n6044;
  assign n6048 = ~n5308 & ~n6047;
  assign n6049 = n5300 & ~n6048;
  assign n6050 = ~n5313 & n5330;
  assign n6051 = ~n5322 & n6050;
  assign n6052 = ~n5289 & n6051;
  assign n6053 = n5291 & ~n6052;
  assign n6054 = ~n5302 & n5344;
  assign n6055 = ~n5309 & n6054;
  assign n6056 = ~n5334 & n6055;
  assign n6057 = ~n5325 & ~n6056;
  assign n6058 = ~n6053 & ~n6057;
  assign n6059 = ~n6049 & n6058;
  assign n6060 = ~n6042 & n6059;
  assign n6061 = n5328 ^ n5180;
  assign n6062 = n6061 ^ n5328;
  assign n6063 = n5334 ^ n5328;
  assign n6064 = n6062 & n6063;
  assign n6065 = n6064 ^ n5328;
  assign n6066 = ~n5179 & n6065;
  assign n6067 = n6060 & ~n6066;
  assign n6068 = n6041 & n6067;
  assign n6069 = n5317 & n6068;
  assign n6070 = n5299 & n6069;
  assign n6071 = n6070 ^ n3063;
  assign n6072 = n6071 ^ x121;
  assign n6073 = n5726 & n5853;
  assign n6074 = n5839 & ~n5874;
  assign n6075 = ~n6073 & ~n6074;
  assign n6076 = ~n5863 & n5871;
  assign n6077 = n5726 & ~n5868;
  assign n6078 = ~n6076 & ~n6077;
  assign n6079 = n5831 & n5856;
  assign n6080 = n5826 & n5831;
  assign n6081 = n5750 & n5839;
  assign n6082 = ~n6080 & ~n6081;
  assign n6083 = n5827 & ~n6082;
  assign n6084 = ~n6079 & ~n6083;
  assign n6085 = ~n5825 & ~n5849;
  assign n6086 = n5854 & ~n6085;
  assign n6087 = n5839 & n5846;
  assign n6088 = ~n5848 & ~n5862;
  assign n6089 = n5726 & ~n6088;
  assign n6090 = ~n6087 & ~n6089;
  assign n6091 = ~n5835 & ~n5853;
  assign n6092 = n5868 & n6091;
  assign n6093 = n5871 & ~n6092;
  assign n6094 = ~n5834 & n5868;
  assign n6095 = n5839 & ~n6094;
  assign n6096 = ~n6093 & ~n6095;
  assign n6097 = ~n5825 & ~n5857;
  assign n6098 = n6097 ^ n5725;
  assign n6099 = n6098 ^ n6097;
  assign n6100 = ~n5843 & ~n5872;
  assign n6101 = n6100 ^ n6097;
  assign n6102 = n6099 & n6101;
  assign n6103 = n6102 ^ n6097;
  assign n6104 = n5689 & ~n6103;
  assign n6105 = n6096 & ~n6104;
  assign n6106 = n6090 & n6105;
  assign n6107 = ~n5837 & n6106;
  assign n6108 = ~n6086 & n6107;
  assign n6109 = n6084 & n6108;
  assign n6110 = n6078 & n6109;
  assign n6111 = n6075 & n6110;
  assign n6112 = ~n5838 & n6111;
  assign n6113 = n6112 ^ n2570;
  assign n6114 = n6113 ^ x112;
  assign n6115 = ~n6072 & n6114;
  assign n6116 = n6038 & n6115;
  assign n6117 = n6004 & n6037;
  assign n6118 = ~n6114 & n6117;
  assign n6119 = ~n6072 & n6118;
  assign n6120 = ~n6116 & ~n6119;
  assign n6121 = n5451 ^ x89;
  assign n6122 = n5774 ^ x82;
  assign n6123 = ~n6121 & ~n6122;
  assign n6124 = n4932 & n4954;
  assign n6125 = n4938 & ~n5693;
  assign n6126 = ~n6124 & ~n6125;
  assign n6127 = n4948 & n4961;
  assign n6128 = ~n4950 & n4977;
  assign n6129 = ~n4987 & n6128;
  assign n6130 = n4881 & ~n6129;
  assign n6131 = ~n6127 & ~n6130;
  assign n6132 = n6126 & n6131;
  assign n6133 = ~n4943 & ~n4959;
  assign n6134 = n4977 & n6133;
  assign n6135 = ~n4961 & n6134;
  assign n6136 = ~n4994 & n5702;
  assign n6137 = ~n4954 & n6136;
  assign n6138 = ~n4940 & n6137;
  assign n6139 = ~n6135 & ~n6138;
  assign n6140 = n6139 ^ n4994;
  assign n6141 = n6140 ^ n4994;
  assign n6142 = n4994 ^ n4993;
  assign n6143 = n6142 ^ n4994;
  assign n6144 = ~n6141 & ~n6143;
  assign n6145 = n6144 ^ n4994;
  assign n6146 = n4964 & ~n6145;
  assign n6147 = n6146 ^ n4994;
  assign n6148 = n6132 & ~n6147;
  assign n6149 = ~n5691 & n6148;
  assign n6150 = n4958 & n6149;
  assign n6151 = n5211 & n6150;
  assign n6152 = n4946 & n6151;
  assign n6153 = ~n5690 & n6152;
  assign n6154 = n6153 ^ n2206;
  assign n6155 = n6154 ^ x106;
  assign n6156 = n5688 ^ x123;
  assign n6157 = ~n3642 & n3647;
  assign n6158 = ~n3607 & n5012;
  assign n6159 = ~n3609 & n6158;
  assign n6160 = n3615 & ~n6159;
  assign n6161 = ~n6157 & ~n6160;
  assign n6162 = ~n3631 & n5019;
  assign n6163 = ~n3636 & n5031;
  assign n6164 = n3617 & ~n6163;
  assign n6165 = n3630 & n3635;
  assign n6166 = n3608 & ~n3652;
  assign n6167 = ~n3650 & n6166;
  assign n6168 = n3647 & ~n6167;
  assign n6169 = ~n6165 & ~n6168;
  assign n6172 = ~n3550 & ~n3637;
  assign n6170 = n3642 & ~n5030;
  assign n6171 = ~n3636 & n6170;
  assign n6173 = n6172 ^ n6171;
  assign n6174 = n6173 ^ n6172;
  assign n6175 = n6172 ^ n3600;
  assign n6176 = n6175 ^ n6172;
  assign n6177 = ~n6174 & n6176;
  assign n6178 = n6177 ^ n6172;
  assign n6179 = ~n3614 & ~n6178;
  assign n6180 = n6179 ^ n6172;
  assign n6181 = n3614 ^ n3600;
  assign n6183 = n3608 & ~n3611;
  assign n6184 = ~n3550 & n6183;
  assign n6182 = ~n3657 & n5017;
  assign n6185 = n6184 ^ n6182;
  assign n6186 = n6184 ^ n3600;
  assign n6187 = n6186 ^ n6184;
  assign n6188 = n6185 & n6187;
  assign n6189 = n6188 ^ n6184;
  assign n6190 = ~n6181 & ~n6189;
  assign n6191 = n6180 & ~n6190;
  assign n6192 = n6169 & n6191;
  assign n6193 = ~n6164 & n6192;
  assign n6194 = ~n6162 & n6193;
  assign n6195 = n6161 & n6194;
  assign n6196 = n6195 ^ n2241;
  assign n6197 = n6196 ^ x96;
  assign n6198 = n6156 & ~n6197;
  assign n6199 = n5397 ^ x121;
  assign n6200 = n6198 & ~n6199;
  assign n6201 = ~n6155 & n6200;
  assign n6202 = n6123 & n6201;
  assign n6203 = n6121 & ~n6122;
  assign n6204 = n6155 & n6199;
  assign n6205 = ~n6156 & n6204;
  assign n6206 = n6197 & n6205;
  assign n6207 = n6203 & n6206;
  assign n6208 = ~n6202 & ~n6207;
  assign n6209 = n6121 & n6122;
  assign n6210 = ~n6156 & ~n6199;
  assign n6211 = n6197 & n6210;
  assign n6212 = n6155 & n6211;
  assign n6213 = n6209 & n6212;
  assign n6214 = n6156 & n6197;
  assign n6215 = ~n6199 & n6214;
  assign n6216 = n6155 & n6215;
  assign n6217 = ~n6155 & n6199;
  assign n6218 = n6214 & n6217;
  assign n6219 = ~n6216 & ~n6218;
  assign n6220 = n6203 & ~n6219;
  assign n6221 = ~n6213 & ~n6220;
  assign n6222 = ~n6155 & n6215;
  assign n6223 = ~n6197 & n6204;
  assign n6224 = n6156 & n6223;
  assign n6225 = ~n6222 & ~n6224;
  assign n6226 = n6209 & ~n6225;
  assign n6227 = n6155 & n6200;
  assign n6228 = n6203 & n6227;
  assign n6229 = ~n6155 & n6211;
  assign n6230 = ~n6223 & ~n6229;
  assign n6231 = n6209 & ~n6230;
  assign n6232 = ~n6228 & ~n6231;
  assign n6233 = ~n6156 & n6217;
  assign n6234 = n6197 & n6233;
  assign n6235 = ~n6227 & ~n6234;
  assign n6236 = n6209 & ~n6235;
  assign n6237 = ~n6197 & n6210;
  assign n6238 = n6155 & n6237;
  assign n6239 = ~n6224 & ~n6238;
  assign n6240 = ~n6216 & n6239;
  assign n6241 = n6123 & ~n6240;
  assign n6242 = ~n6121 & n6122;
  assign n6243 = n6204 & n6214;
  assign n6244 = ~n6222 & ~n6243;
  assign n6245 = ~n6224 & ~n6227;
  assign n6246 = n6244 & n6245;
  assign n6247 = n6242 & ~n6246;
  assign n6248 = ~n6241 & ~n6247;
  assign n6249 = ~n6236 & n6248;
  assign n6250 = ~n6212 & ~n6234;
  assign n6251 = ~n6206 & n6250;
  assign n6252 = n6251 ^ n6122;
  assign n6253 = n6252 ^ n6251;
  assign n6254 = ~n6156 & n6223;
  assign n6255 = ~n6155 & n6237;
  assign n6256 = ~n6254 & ~n6255;
  assign n6257 = ~n6243 & n6256;
  assign n6258 = ~n6201 & n6257;
  assign n6259 = n6258 ^ n6251;
  assign n6260 = n6259 ^ n6251;
  assign n6261 = ~n6253 & ~n6260;
  assign n6262 = n6261 ^ n6251;
  assign n6263 = n6121 & ~n6262;
  assign n6264 = n6263 ^ n6251;
  assign n6265 = n6249 & n6264;
  assign n6266 = n6122 ^ n6121;
  assign n6268 = n6198 & n6217;
  assign n6267 = ~n6197 & n6233;
  assign n6269 = n6268 ^ n6267;
  assign n6270 = n6269 ^ n6268;
  assign n6271 = n6268 ^ n6122;
  assign n6272 = n6271 ^ n6268;
  assign n6273 = n6270 & n6272;
  assign n6274 = n6273 ^ n6268;
  assign n6275 = n6266 & n6274;
  assign n6276 = n6275 ^ n6268;
  assign n6277 = n6265 & ~n6276;
  assign n6278 = n6232 & n6277;
  assign n6279 = ~n6226 & n6278;
  assign n6280 = n6221 & n6279;
  assign n6281 = n6208 & n6280;
  assign n6282 = n6281 ^ n2319;
  assign n6283 = n6282 ^ x97;
  assign n6284 = ~n3252 & n3254;
  assign n6285 = ~n3217 & n3219;
  assign n6286 = ~n6284 & ~n6285;
  assign n6287 = n2321 & ~n3238;
  assign n6288 = n3241 & ~n3260;
  assign n6289 = ~n6287 & ~n6288;
  assign n6290 = n6286 & n6289;
  assign n6291 = n6290 ^ n1276;
  assign n6292 = n6291 ^ x108;
  assign n6293 = n3669 ^ x126;
  assign n6294 = ~n6292 & ~n6293;
  assign n6295 = ~n4279 & n4333;
  assign n6296 = n4178 & ~n6295;
  assign n6298 = n4273 ^ n4209;
  assign n6297 = ~n4210 & n4245;
  assign n6299 = n6298 ^ n6297;
  assign n6300 = n4320 & ~n6299;
  assign n6301 = ~n6296 & ~n6300;
  assign n6302 = n4286 & ~n5438;
  assign n6303 = ~n4307 & n5434;
  assign n6304 = ~n4294 & n6303;
  assign n6305 = ~n4279 & n6304;
  assign n6306 = n4277 & ~n6305;
  assign n6307 = ~n6302 & ~n6306;
  assign n6308 = n6301 & n6307;
  assign n6309 = n5427 & n6308;
  assign n6310 = ~n4299 & n6309;
  assign n6311 = ~n4293 & n6310;
  assign n6312 = ~n5424 & n6311;
  assign n6313 = n6312 ^ n1738;
  assign n6314 = n6313 ^ x70;
  assign n6315 = n5724 ^ x85;
  assign n6316 = ~n6314 & n6315;
  assign n6317 = n6294 & n6316;
  assign n6318 = n3885 ^ x68;
  assign n6319 = n5822 ^ x94;
  assign n6320 = n6318 & n6319;
  assign n6321 = n6317 & n6320;
  assign n6322 = n6314 & ~n6315;
  assign n6323 = n6294 & n6322;
  assign n6324 = ~n6318 & ~n6319;
  assign n6325 = n6323 & n6324;
  assign n6326 = ~n6321 & ~n6325;
  assign n6327 = n6292 & ~n6293;
  assign n6328 = n6322 & n6327;
  assign n6329 = n6320 & n6328;
  assign n6330 = ~n6318 & n6319;
  assign n6331 = ~n6292 & n6293;
  assign n6332 = n6316 & n6331;
  assign n6333 = n6292 & n6293;
  assign n6334 = ~n6314 & ~n6315;
  assign n6335 = n6333 & n6334;
  assign n6336 = ~n6332 & ~n6335;
  assign n6337 = n6330 & ~n6336;
  assign n6338 = n6316 & n6333;
  assign n6339 = n6322 & n6333;
  assign n6340 = ~n6338 & ~n6339;
  assign n6341 = n6320 & ~n6340;
  assign n6342 = ~n6337 & ~n6341;
  assign n6343 = ~n6329 & n6342;
  assign n6344 = n6331 & n6334;
  assign n6345 = n6324 & n6344;
  assign n6346 = n6327 & n6334;
  assign n6347 = n6320 & n6346;
  assign n6348 = ~n6345 & ~n6347;
  assign n6349 = n6314 & n6315;
  assign n6350 = n6327 & n6349;
  assign n6351 = ~n6323 & ~n6350;
  assign n6352 = ~n6339 & n6351;
  assign n6353 = ~n6317 & n6352;
  assign n6354 = n6330 & ~n6353;
  assign n6355 = n6333 & n6349;
  assign n6356 = n6322 & n6331;
  assign n6357 = ~n6355 & ~n6356;
  assign n6358 = ~n6317 & n6357;
  assign n6359 = ~n6338 & n6358;
  assign n6360 = n6324 & ~n6359;
  assign n6361 = ~n6354 & ~n6360;
  assign n6362 = n6316 & n6327;
  assign n6363 = ~n6328 & ~n6362;
  assign n6364 = ~n6318 & ~n6363;
  assign n6365 = n6294 & n6349;
  assign n6366 = ~n6344 & ~n6365;
  assign n6367 = ~n6356 & n6366;
  assign n6368 = n6320 & ~n6367;
  assign n6369 = n6318 & ~n6319;
  assign n6370 = ~n6332 & ~n6356;
  assign n6371 = ~n6317 & ~n6346;
  assign n6372 = ~n6328 & n6371;
  assign n6373 = ~n6365 & n6372;
  assign n6374 = n6370 & n6373;
  assign n6375 = ~n6350 & n6374;
  assign n6376 = ~n6338 & n6375;
  assign n6377 = n6369 & n6376;
  assign n6378 = ~n6368 & ~n6377;
  assign n6379 = ~n6364 & n6378;
  assign n6380 = n6361 & n6379;
  assign n6381 = n6348 & n6380;
  assign n6382 = n6343 & n6381;
  assign n6383 = n6326 & n6382;
  assign n6384 = n6383 ^ n1950;
  assign n6385 = n6384 ^ x115;
  assign n6386 = n6283 & ~n6385;
  assign n6387 = ~n6004 & n6037;
  assign n6388 = n6387 ^ n6038;
  assign n6389 = n6072 & n6388;
  assign n6390 = n6389 ^ n6387;
  assign n6391 = ~n6114 & n6390;
  assign n6392 = n6072 & n6114;
  assign n6393 = n6387 & n6392;
  assign n6394 = n6115 & n6117;
  assign n6395 = n6038 & n6392;
  assign n6396 = ~n6004 & ~n6037;
  assign n6397 = ~n6392 & n6396;
  assign n6398 = ~n6395 & ~n6397;
  assign n6399 = ~n6394 & n6398;
  assign n6400 = ~n6393 & n6399;
  assign n6401 = ~n6391 & n6400;
  assign n6402 = n6386 & n6401;
  assign n6403 = ~n6283 & ~n6385;
  assign n6404 = n6115 & n6387;
  assign n6405 = n6072 & ~n6114;
  assign n6406 = n6117 & n6405;
  assign n6407 = ~n6404 & ~n6406;
  assign n6408 = ~n6072 & n6396;
  assign n6409 = n6038 & n6405;
  assign n6410 = ~n6408 & ~n6409;
  assign n6411 = n6407 & n6410;
  assign n6412 = ~n6393 & n6411;
  assign n6413 = n6403 & ~n6412;
  assign n6414 = ~n6402 & ~n6413;
  assign n6415 = ~n6283 & n6385;
  assign n6416 = n6072 & n6396;
  assign n6417 = n6392 ^ n6038;
  assign n6418 = n6417 ^ n6038;
  assign n6419 = n6388 & ~n6418;
  assign n6420 = n6419 ^ n6038;
  assign n6421 = ~n6416 & ~n6420;
  assign n6422 = n6415 & ~n6421;
  assign n6423 = n6283 & n6385;
  assign n6424 = ~n6114 & n6396;
  assign n6425 = ~n6393 & ~n6424;
  assign n6426 = ~n6394 & n6425;
  assign n6427 = ~n6391 & n6426;
  assign n6428 = n6120 & n6427;
  assign n6429 = n6423 & ~n6428;
  assign n6430 = ~n6422 & ~n6429;
  assign n6431 = n6414 & n6430;
  assign n6432 = n6120 & n6431;
  assign n6433 = n6432 ^ n5688;
  assign n6434 = n6433 ^ x120;
  assign n6435 = n6282 ^ x86;
  assign n6436 = n4551 & n4590;
  assign n6437 = n3671 & ~n4583;
  assign n6438 = ~n6436 & ~n6437;
  assign n6439 = n4551 & n4606;
  assign n6440 = n3671 & n4584;
  assign n6441 = n4561 & n4583;
  assign n6442 = n4547 & ~n6441;
  assign n6443 = ~n6440 & ~n6442;
  assign n6444 = ~n6439 & n6443;
  assign n6445 = ~n4573 & ~n4584;
  assign n6446 = n4551 & ~n6445;
  assign n6447 = n4551 & n4578;
  assign n6448 = n4547 & n4573;
  assign n6449 = ~n6447 & ~n6448;
  assign n6450 = n4544 & n4547;
  assign n6451 = n4551 & ~n4583;
  assign n6452 = ~n6450 & ~n6451;
  assign n6453 = n3671 & n4566;
  assign n6454 = ~n4590 & ~n4593;
  assign n6455 = ~n4569 & n6454;
  assign n6456 = ~n4541 & n6455;
  assign n6457 = ~n4549 & n6456;
  assign n6458 = n4556 & ~n6457;
  assign n6459 = ~n6453 & ~n6458;
  assign n6460 = n6452 & n6459;
  assign n6461 = n6449 & n6460;
  assign n6462 = ~n6446 & n6461;
  assign n6463 = n4568 & n6462;
  assign n6464 = n6444 & n6463;
  assign n6465 = n4564 & n6464;
  assign n6466 = n6438 & n6465;
  assign n6467 = ~n4546 & n6466;
  assign n6468 = n6467 ^ n3547;
  assign n6469 = n6468 ^ x108;
  assign n6470 = ~n6435 & n6469;
  assign n6471 = ~n5632 & n5662;
  assign n6472 = n5648 & n5651;
  assign n6473 = ~n6471 & ~n6472;
  assign n6474 = n5634 & ~n5660;
  assign n6475 = n5566 & ~n5667;
  assign n6476 = ~n6474 & ~n6475;
  assign n6477 = n6473 & n6476;
  assign n6478 = n6477 ^ n3387;
  assign n6479 = n6478 ^ x126;
  assign n6480 = ~n5452 & n5506;
  assign n6481 = n5399 & n6480;
  assign n6482 = n5535 & ~n6019;
  assign n6483 = ~n6481 & ~n6482;
  assign n6484 = ~n5529 & ~n5537;
  assign n6485 = ~n5507 & n6484;
  assign n6486 = n5488 & ~n6485;
  assign n6487 = ~n5498 & n5530;
  assign n6488 = n5399 & ~n6487;
  assign n6489 = ~n5486 & n5530;
  assign n6490 = n5505 & ~n6489;
  assign n6491 = ~n6488 & ~n6490;
  assign n6492 = n5507 & ~n6019;
  assign n6493 = ~n5509 & ~n5535;
  assign n6494 = ~n5503 & n6493;
  assign n6495 = n5488 & ~n6494;
  assign n6496 = ~n6492 & ~n6495;
  assign n6497 = n6491 & n6496;
  assign n6498 = n5502 & n6497;
  assign n6499 = ~n5487 & n6498;
  assign n6500 = ~n6486 & n6499;
  assign n6501 = n5536 ^ n5518;
  assign n6502 = n6501 ^ n5536;
  assign n6503 = n5536 ^ n5357;
  assign n6504 = n6503 ^ n5536;
  assign n6505 = ~n6502 & ~n6504;
  assign n6506 = n6505 ^ n5536;
  assign n6507 = ~n5398 & n6506;
  assign n6508 = n6507 ^ n5536;
  assign n6509 = n6500 & ~n6508;
  assign n6510 = n6483 & n6509;
  assign n6511 = ~n6006 & n6510;
  assign n6512 = n6010 & n6511;
  assign n6513 = ~n5559 & n6512;
  assign n6514 = n6513 ^ n3418;
  assign n6515 = n6514 ^ x93;
  assign n6516 = n6479 & ~n6515;
  assign n6517 = n6470 & n6516;
  assign n6518 = n6003 ^ x76;
  assign n6519 = n5839 & n5872;
  assign n6520 = n5853 ^ n5846;
  assign n6521 = n6520 ^ n5846;
  assign n6522 = n5846 ^ n5839;
  assign n6523 = n6522 ^ n5846;
  assign n6524 = n6521 & ~n6523;
  assign n6525 = n6524 ^ n5846;
  assign n6526 = ~n5726 & n6525;
  assign n6527 = n6526 ^ n5846;
  assign n6528 = ~n6519 & ~n6527;
  assign n6529 = n5878 ^ n5725;
  assign n6530 = n6529 ^ n5878;
  assign n6531 = ~n5835 & ~n5867;
  assign n6532 = n6531 ^ n5878;
  assign n6533 = n6530 & n6532;
  assign n6534 = n6533 ^ n5878;
  assign n6535 = ~n5689 & ~n6534;
  assign n6536 = ~n5867 & ~n5873;
  assign n6537 = n6536 ^ n5850;
  assign n6538 = n6536 ^ n5871;
  assign n6539 = n6538 ^ n5871;
  assign n6540 = n5871 ^ n5831;
  assign n6541 = ~n6539 & ~n6540;
  assign n6542 = n6541 ^ n5871;
  assign n6543 = n6537 & ~n6542;
  assign n6544 = n6543 ^ n5850;
  assign n6545 = n5858 & n6544;
  assign n6546 = n5854 & ~n6545;
  assign n6547 = n6075 & ~n6546;
  assign n6548 = n5872 ^ n5854;
  assign n6549 = n6548 ^ n5872;
  assign n6550 = n5872 ^ n5849;
  assign n6551 = ~n6549 & n6550;
  assign n6552 = n6551 ^ n5872;
  assign n6553 = n6547 & ~n6552;
  assign n6554 = ~n6535 & n6553;
  assign n6555 = n5845 & n6554;
  assign n6556 = n6528 & n6555;
  assign n6557 = n6090 & n6556;
  assign n6558 = ~n5837 & n6557;
  assign n6559 = ~n5830 & n6558;
  assign n6560 = n6559 ^ n3599;
  assign n6561 = n6560 ^ x125;
  assign n6562 = n6518 & n6561;
  assign n6563 = n6517 & n6562;
  assign n6564 = ~n6479 & n6515;
  assign n6565 = n6435 & n6469;
  assign n6566 = n6564 & n6565;
  assign n6567 = n6479 & n6515;
  assign n6568 = n6435 & ~n6469;
  assign n6569 = n6567 & n6568;
  assign n6570 = ~n6566 & ~n6569;
  assign n6571 = n6518 & ~n6561;
  assign n6572 = ~n6570 & n6571;
  assign n6573 = ~n6563 & ~n6572;
  assign n6574 = n6516 & n6565;
  assign n6575 = n6564 & n6568;
  assign n6576 = ~n6574 & ~n6575;
  assign n6577 = ~n6569 & n6576;
  assign n6578 = ~n6518 & n6561;
  assign n6579 = ~n6577 & n6578;
  assign n6580 = ~n6479 & ~n6515;
  assign n6581 = n6568 & n6580;
  assign n6582 = n6571 & n6581;
  assign n6583 = ~n6579 & ~n6582;
  assign n6584 = n6516 & n6568;
  assign n6585 = ~n6518 & ~n6561;
  assign n6586 = ~n6562 & ~n6585;
  assign n6587 = n6584 & n6586;
  assign n6588 = ~n6435 & ~n6469;
  assign n6589 = n6567 & n6588;
  assign n6590 = n6470 & n6567;
  assign n6591 = n6564 & n6588;
  assign n6592 = ~n6590 & ~n6591;
  assign n6593 = ~n6589 & n6592;
  assign n6594 = n6562 & ~n6593;
  assign n6595 = n6571 & n6574;
  assign n6596 = n6580 & n6588;
  assign n6597 = n6516 & n6588;
  assign n6598 = ~n6596 & ~n6597;
  assign n6599 = ~n6574 & ~n6584;
  assign n6600 = n6592 & n6599;
  assign n6601 = n6598 & n6600;
  assign n6602 = n6585 & ~n6601;
  assign n6603 = n6565 & n6567;
  assign n6604 = n6565 & n6580;
  assign n6605 = ~n6603 & ~n6604;
  assign n6606 = ~n6586 & ~n6605;
  assign n6607 = ~n6602 & ~n6606;
  assign n6608 = ~n6566 & ~n6581;
  assign n6609 = n6562 & ~n6608;
  assign n6610 = n6470 & n6564;
  assign n6611 = ~n6597 & ~n6610;
  assign n6612 = ~n6591 & n6611;
  assign n6613 = ~n6578 & n6612;
  assign n6614 = n6470 & n6580;
  assign n6615 = ~n6589 & ~n6610;
  assign n6616 = ~n6597 & n6615;
  assign n6617 = ~n6614 & n6616;
  assign n6618 = ~n6571 & n6617;
  assign n6619 = ~n6613 & ~n6618;
  assign n6620 = n6586 & n6619;
  assign n6621 = ~n6609 & ~n6620;
  assign n6622 = n6607 & n6621;
  assign n6623 = ~n6595 & n6622;
  assign n6624 = ~n6594 & n6623;
  assign n6625 = ~n6587 & n6624;
  assign n6626 = n6583 & n6625;
  assign n6627 = n6573 & n6626;
  assign n6628 = n6627 ^ n6196;
  assign n6629 = n6628 ^ x64;
  assign n6630 = n6434 & ~n6629;
  assign n6631 = n6201 & n6209;
  assign n6632 = n6206 & n6209;
  assign n6633 = n6203 & n6224;
  assign n6634 = ~n6632 & ~n6633;
  assign n6635 = n6203 & n6268;
  assign n6636 = ~n6227 & ~n6267;
  assign n6637 = ~n6121 & ~n6636;
  assign n6638 = ~n6234 & ~n6238;
  assign n6639 = ~n6266 & ~n6638;
  assign n6640 = n6230 & ~n6255;
  assign n6641 = ~n6234 & n6640;
  assign n6642 = n6203 & ~n6641;
  assign n6643 = ~n6639 & ~n6642;
  assign n6644 = n6123 & ~n6244;
  assign n6645 = ~n6218 & n6257;
  assign n6646 = ~n6212 & n6645;
  assign n6647 = n6242 & ~n6646;
  assign n6648 = ~n6644 & ~n6647;
  assign n6649 = n6643 & n6648;
  assign n6650 = ~n6637 & n6649;
  assign n6651 = ~n6635 & n6650;
  assign n6652 = n6634 & n6651;
  assign n6653 = ~n6226 & n6652;
  assign n6654 = ~n6631 & n6653;
  assign n6655 = ~n6213 & n6654;
  assign n6656 = n6208 & n6655;
  assign n6657 = ~n6216 & n6656;
  assign n6658 = n6657 ^ n3707;
  assign n6659 = n6658 ^ x98;
  assign n6660 = n4541 & n4551;
  assign n6661 = n4547 & n4584;
  assign n6662 = ~n6660 & ~n6661;
  assign n6663 = ~n4544 & ~n4566;
  assign n6664 = n4551 & ~n6663;
  assign n6665 = n4147 ^ n3886;
  assign n6666 = n6665 ^ n4357;
  assign n6667 = n6666 ^ n4539;
  assign n6668 = n4539 ^ n4147;
  assign n6669 = n6668 ^ n4539;
  assign n6670 = n4539 ^ n4357;
  assign n6671 = n6670 ^ n4539;
  assign n6672 = n6669 & ~n6671;
  assign n6673 = n6672 ^ n4539;
  assign n6674 = ~n6667 & ~n6673;
  assign n6675 = n6674 ^ n3886;
  assign n6676 = n4547 & ~n6675;
  assign n6677 = ~n6664 & ~n6676;
  assign n6678 = ~n4578 & ~n4582;
  assign n6679 = n4556 & ~n6678;
  assign n6680 = ~n4544 & ~n4593;
  assign n6681 = ~n4549 & ~n4590;
  assign n6682 = ~n4556 & n6681;
  assign n6683 = ~n4554 & ~n4606;
  assign n6684 = ~n4569 & n6683;
  assign n6685 = ~n3671 & n6684;
  assign n6686 = ~n6682 & ~n6685;
  assign n6687 = ~n4560 & ~n6686;
  assign n6688 = n6680 & n6687;
  assign n6689 = ~n4557 & n6688;
  assign n6690 = n6689 ^ n4557;
  assign n6691 = ~n6679 & n6690;
  assign n6692 = n6677 & n6691;
  assign n6693 = n6449 & n6692;
  assign n6694 = ~n6446 & n6693;
  assign n6695 = n6662 & n6694;
  assign n6696 = n4572 & n6695;
  assign n6697 = n6438 & n6696;
  assign n6698 = n6697 ^ n4021;
  assign n6699 = n6698 ^ x89;
  assign n6700 = ~n6659 & n6699;
  assign n6701 = n5834 & ~n5854;
  assign n6702 = ~n5856 & ~n5873;
  assign n6703 = ~n5843 & n6702;
  assign n6704 = n5839 & ~n6703;
  assign n6705 = ~n6701 & ~n6704;
  assign n6706 = n5829 & n6088;
  assign n6707 = n5871 & ~n6706;
  assign n6708 = ~n5867 & n5874;
  assign n6709 = n5726 & ~n6708;
  assign n6710 = ~n6707 & ~n6709;
  assign n6711 = n5854 & ~n5878;
  assign n6712 = n5750 & n5827;
  assign n6713 = n5859 & ~n6712;
  assign n6714 = n5831 & ~n6713;
  assign n6715 = ~n6711 & ~n6714;
  assign n6716 = n6710 & n6715;
  assign n6717 = n6705 & n6716;
  assign n6718 = n5852 & n6717;
  assign n6719 = n6528 & n6718;
  assign n6720 = ~n5838 & n6719;
  assign n6721 = ~n5830 & n6720;
  assign n6722 = n6721 ^ n3946;
  assign n6723 = n6722 ^ x113;
  assign n6724 = n5090 & n5108;
  assign n6725 = n5982 & ~n6724;
  assign n6726 = n5058 & n5092;
  assign n6727 = n5077 & ~n6726;
  assign n6728 = ~n5052 & n5106;
  assign n6729 = n5079 & n5090;
  assign n6730 = ~n6728 & ~n6729;
  assign n6731 = n5058 & ~n5100;
  assign n6732 = ~n5084 & ~n5108;
  assign n6733 = n5063 & ~n6732;
  assign n6734 = n5100 & n5978;
  assign n6735 = ~n5010 & ~n6734;
  assign n6736 = n5087 & ~n5107;
  assign n6737 = ~n5061 & n6736;
  assign n6738 = n5056 & ~n6737;
  assign n6739 = ~n6735 & ~n6738;
  assign n6740 = ~n6733 & n6739;
  assign n6741 = ~n6731 & n6740;
  assign n6742 = n6730 & n6741;
  assign n6743 = ~n5964 & n6742;
  assign n6744 = n6727 & n6743;
  assign n6745 = n6725 & n6744;
  assign n6746 = n5963 & n6745;
  assign n6747 = ~n5057 & n6746;
  assign n6748 = ~n5053 & n6747;
  assign n6749 = n6748 ^ n4928;
  assign n6750 = n6749 ^ x123;
  assign n6751 = n6723 & n6750;
  assign n6752 = n6324 & ~n6371;
  assign n6753 = n6319 ^ n6318;
  assign n6754 = n6332 ^ n6319;
  assign n6755 = n6754 ^ n6332;
  assign n6756 = n6338 ^ n6332;
  assign n6757 = n6755 & n6756;
  assign n6758 = n6757 ^ n6332;
  assign n6759 = n6753 & n6758;
  assign n6760 = ~n6752 & ~n6759;
  assign n6761 = n6328 & n6753;
  assign n6762 = n6330 & ~n6370;
  assign n6763 = ~n6761 & ~n6762;
  assign n6764 = ~n6340 & n6369;
  assign n6765 = n6331 & n6349;
  assign n6766 = ~n6335 & ~n6765;
  assign n6767 = n6357 & n6766;
  assign n6768 = ~n6350 & n6767;
  assign n6769 = n6324 & ~n6768;
  assign n6770 = n6315 ^ n6292;
  assign n6771 = n6770 ^ n6292;
  assign n6772 = n6314 ^ n6292;
  assign n6773 = n6772 ^ n6292;
  assign n6774 = n6771 & ~n6773;
  assign n6775 = n6774 ^ n6292;
  assign n6776 = ~n6293 & ~n6775;
  assign n6777 = n6753 & n6776;
  assign n6778 = ~n6344 & ~n6765;
  assign n6779 = n6353 & n6778;
  assign n6780 = ~n6332 & n6779;
  assign n6781 = n6320 & ~n6780;
  assign n6782 = ~n6777 & ~n6781;
  assign n6783 = ~n6769 & n6782;
  assign n6784 = ~n6764 & n6783;
  assign n6785 = n6763 & n6784;
  assign n6786 = n6348 & n6785;
  assign n6787 = n6760 & n6786;
  assign n6788 = n6787 ^ n4906;
  assign n6789 = n6788 ^ x65;
  assign n6790 = ~n5308 & ~n5343;
  assign n6791 = n5300 & ~n6790;
  assign n6792 = n5291 & n5308;
  assign n6793 = n5181 & n5318;
  assign n6794 = ~n6792 & ~n6793;
  assign n6795 = n5291 & n5334;
  assign n6796 = n5181 & n5322;
  assign n6797 = ~n5324 & ~n5343;
  assign n6798 = n5312 & ~n6797;
  assign n6799 = ~n6796 & ~n6798;
  assign n6800 = ~n6795 & n6799;
  assign n6801 = n5289 & n5325;
  assign n6802 = ~n5304 & ~n5318;
  assign n6803 = n5291 & ~n6802;
  assign n6804 = ~n6801 & ~n6803;
  assign n6805 = ~n5313 & n5331;
  assign n6806 = n5312 & ~n6805;
  assign n6807 = ~n5296 & n5315;
  assign n6808 = ~n5302 & n6807;
  assign n6809 = ~n5309 & n6808;
  assign n6810 = n5181 & ~n6809;
  assign n6811 = ~n6806 & ~n6810;
  assign n6812 = n6804 & n6811;
  assign n6813 = ~n6066 & n6812;
  assign n6814 = n5327 & n6813;
  assign n6815 = n6800 & n6814;
  assign n6816 = n6794 & n6815;
  assign n6817 = ~n6791 & n6816;
  assign n6818 = ~n5306 & n6817;
  assign n6819 = n5299 & n6818;
  assign n6820 = n6819 ^ n3820;
  assign n6821 = n6820 ^ x104;
  assign n6822 = n6789 & ~n6821;
  assign n6823 = n6751 & n6822;
  assign n6824 = n6700 & n6823;
  assign n6825 = ~n6789 & n6821;
  assign n6826 = ~n6723 & ~n6750;
  assign n6827 = n6825 & n6826;
  assign n6828 = n6659 & ~n6699;
  assign n6829 = n6827 & n6828;
  assign n6830 = ~n6824 & ~n6829;
  assign n6831 = n6789 & n6821;
  assign n6832 = n6751 & n6831;
  assign n6833 = n6700 & n6832;
  assign n6834 = n6823 & n6828;
  assign n6835 = ~n6723 & n6750;
  assign n6836 = n6831 & n6835;
  assign n6837 = n6822 & n6826;
  assign n6838 = ~n6836 & ~n6837;
  assign n6839 = n6700 & ~n6838;
  assign n6840 = ~n6834 & ~n6839;
  assign n6841 = ~n6833 & n6840;
  assign n6842 = n6723 & ~n6750;
  assign n6843 = n6825 & n6842;
  assign n6844 = ~n6659 & ~n6699;
  assign n6845 = n6843 & n6844;
  assign n6846 = n6659 & n6699;
  assign n6847 = ~n6789 & ~n6821;
  assign n6848 = n6842 & n6847;
  assign n6849 = n6846 & n6848;
  assign n6850 = n6825 & n6835;
  assign n6851 = n6822 & n6835;
  assign n6852 = n6822 & n6842;
  assign n6853 = n6751 & n6825;
  assign n6854 = ~n6852 & ~n6853;
  assign n6855 = ~n6848 & n6854;
  assign n6856 = ~n6832 & n6855;
  assign n6857 = ~n6851 & n6856;
  assign n6858 = ~n6850 & n6857;
  assign n6859 = n6828 & ~n6858;
  assign n6860 = ~n6849 & ~n6859;
  assign n6861 = n6831 & n6842;
  assign n6862 = n6826 & n6847;
  assign n6863 = ~n6827 & ~n6862;
  assign n6864 = ~n6853 & n6863;
  assign n6865 = ~n6861 & n6864;
  assign n6866 = n6700 & ~n6865;
  assign n6867 = ~n6844 & ~n6846;
  assign n6868 = n6751 & n6847;
  assign n6869 = ~n6861 & ~n6868;
  assign n6872 = n6835 & n6847;
  assign n6873 = ~n6836 & ~n6872;
  assign n6874 = ~n6827 & n6873;
  assign n6870 = ~n6850 & ~n6862;
  assign n6871 = ~n6832 & n6870;
  assign n6875 = n6874 ^ n6871;
  assign n6876 = n6699 ^ n6659;
  assign n6877 = n6871 ^ n6699;
  assign n6878 = n6876 & ~n6877;
  assign n6879 = n6878 ^ n6699;
  assign n6880 = n6875 & ~n6879;
  assign n6881 = n6880 ^ n6874;
  assign n6882 = n6869 & n6881;
  assign n6883 = ~n6852 & n6882;
  assign n6884 = ~n6851 & n6883;
  assign n6885 = ~n6867 & ~n6884;
  assign n6886 = ~n6866 & ~n6885;
  assign n6887 = n6860 & n6886;
  assign n6888 = ~n6845 & n6887;
  assign n6889 = n6841 & n6888;
  assign n6890 = n6830 & n6889;
  assign n6891 = n6890 ^ n6154;
  assign n6892 = n6891 ^ x74;
  assign n6893 = n6478 ^ x101;
  assign n6894 = n5355 ^ x118;
  assign n6895 = ~n6893 & n6894;
  assign n6896 = ~n6238 & ~n6267;
  assign n6897 = n6242 & ~n6896;
  assign n6898 = n6123 & ~n6245;
  assign n6899 = ~n6224 & n6244;
  assign n6900 = ~n6206 & n6899;
  assign n6901 = n6203 & ~n6900;
  assign n6902 = ~n6898 & ~n6901;
  assign n6903 = n6197 ^ n6121;
  assign n6904 = n6903 ^ n6121;
  assign n6905 = n6266 ^ n6121;
  assign n6906 = ~n6904 & n6905;
  assign n6907 = n6906 ^ n6121;
  assign n6908 = n6233 & ~n6907;
  assign n6909 = n6902 & ~n6908;
  assign n6910 = n6242 & n6255;
  assign n6911 = n6244 & ~n6268;
  assign n6912 = ~n6216 & n6911;
  assign n6913 = n6242 & ~n6912;
  assign n6914 = n6250 & ~n6255;
  assign n6915 = n6203 & ~n6914;
  assign n6916 = ~n6913 & ~n6915;
  assign n6917 = n6239 & ~n6243;
  assign n6918 = n6917 ^ n6122;
  assign n6919 = n6918 ^ n6917;
  assign n6920 = ~n6206 & n6219;
  assign n6921 = ~n6229 & n6920;
  assign n6922 = n6921 ^ n6917;
  assign n6923 = ~n6919 & n6922;
  assign n6924 = n6923 ^ n6917;
  assign n6925 = ~n6266 & ~n6924;
  assign n6926 = n6916 & ~n6925;
  assign n6927 = ~n6910 & n6926;
  assign n6928 = n6909 & n6927;
  assign n6929 = n6232 & n6928;
  assign n6930 = ~n6897 & n6929;
  assign n6931 = ~n6631 & n6930;
  assign n6932 = ~n6213 & n6931;
  assign n6933 = n6932 ^ n4751;
  assign n6934 = n6933 ^ x75;
  assign n6935 = n6330 & n6355;
  assign n6936 = ~n6363 & n6369;
  assign n6937 = ~n6935 & ~n6936;
  assign n6938 = n6294 & n6334;
  assign n6939 = ~n6350 & ~n6938;
  assign n6940 = n6320 & ~n6939;
  assign n6941 = ~n6357 & n6369;
  assign n6942 = ~n6344 & n6351;
  assign n6943 = n6942 ^ n6319;
  assign n6944 = n6943 ^ n6942;
  assign n6945 = n6340 & n6778;
  assign n6946 = n6945 ^ n6942;
  assign n6947 = n6946 ^ n6942;
  assign n6948 = ~n6944 & ~n6947;
  assign n6949 = n6948 ^ n6942;
  assign n6950 = ~n6753 & ~n6949;
  assign n6951 = n6950 ^ n6942;
  assign n6952 = ~n6941 & n6951;
  assign n6953 = n6766 ^ n6365;
  assign n6954 = n6953 ^ n6365;
  assign n6955 = n6365 ^ n6319;
  assign n6956 = n6955 ^ n6365;
  assign n6957 = ~n6954 & n6956;
  assign n6958 = n6957 ^ n6365;
  assign n6959 = n6318 & n6958;
  assign n6960 = n6959 ^ n6365;
  assign n6961 = n6952 & ~n6960;
  assign n6962 = n6760 & n6961;
  assign n6963 = n6343 & n6962;
  assign n6964 = n6326 & n6963;
  assign n6965 = ~n6940 & n6964;
  assign n6966 = n6937 & n6965;
  assign n6967 = n6966 ^ n4797;
  assign n6968 = n6967 ^ x94;
  assign n6969 = ~n6934 & ~n6968;
  assign n6970 = n5132 ^ x77;
  assign n6971 = n6560 ^ x84;
  assign n6972 = ~n6970 & ~n6971;
  assign n6973 = n6969 & n6972;
  assign n6974 = n6895 & n6973;
  assign n6975 = ~n6893 & ~n6894;
  assign n6976 = n6934 & ~n6968;
  assign n6977 = ~n6970 & n6971;
  assign n6978 = n6976 & n6977;
  assign n6979 = n6970 & n6971;
  assign n6980 = n6969 & n6979;
  assign n6981 = ~n6978 & ~n6980;
  assign n6982 = n6975 & ~n6981;
  assign n6983 = ~n6974 & ~n6982;
  assign n6984 = n6893 & n6894;
  assign n6985 = n6934 & n6968;
  assign n6986 = n6977 & n6985;
  assign n6987 = ~n6980 & ~n6986;
  assign n6988 = n6984 & ~n6987;
  assign n6989 = n6970 & ~n6971;
  assign n6990 = n6969 & n6989;
  assign n6991 = n6975 & n6990;
  assign n6992 = ~n6934 & n6968;
  assign n6993 = n6989 & n6992;
  assign n6994 = n6972 & n6985;
  assign n6995 = ~n6993 & ~n6994;
  assign n6996 = n6984 & ~n6995;
  assign n6997 = ~n6991 & ~n6996;
  assign n6998 = n6893 & ~n6894;
  assign n6999 = ~n6895 & ~n6998;
  assign n7000 = n6979 & n6985;
  assign n7001 = n6999 & n7000;
  assign n7002 = n6969 & n6977;
  assign n7003 = n6893 & n7002;
  assign n7004 = ~n7001 & ~n7003;
  assign n7005 = n6979 & n6992;
  assign n7006 = n6976 & n6979;
  assign n7007 = ~n6986 & ~n7006;
  assign n7008 = ~n7005 & n7007;
  assign n7009 = n6998 & ~n7008;
  assign n7010 = n6977 & n6992;
  assign n7011 = n6972 & n6976;
  assign n7012 = ~n6986 & ~n7011;
  assign n7013 = ~n6993 & n7012;
  assign n7014 = ~n7010 & n7013;
  assign n7015 = n6975 & ~n7014;
  assign n7016 = ~n7009 & ~n7015;
  assign n7017 = n7004 & n7016;
  assign n7018 = n6972 & n6992;
  assign n7019 = ~n6990 & ~n7018;
  assign n7020 = n6984 & ~n7019;
  assign n7021 = n6985 & n6989;
  assign n7022 = n6976 & n6989;
  assign n7023 = ~n6994 & ~n7022;
  assign n7024 = ~n7021 & n7023;
  assign n7025 = n6895 & ~n7024;
  assign n7026 = ~n7002 & ~n7005;
  assign n7027 = ~n7010 & n7026;
  assign n7028 = ~n6998 & n7027;
  assign n7029 = ~n6978 & n7028;
  assign n7030 = n6970 ^ n6934;
  assign n7031 = n6971 ^ n6970;
  assign n7032 = n7031 ^ n6971;
  assign n7033 = n6971 ^ n6968;
  assign n7034 = n7033 ^ n6971;
  assign n7035 = ~n7032 & n7034;
  assign n7036 = n7035 ^ n6971;
  assign n7037 = ~n7030 & ~n7036;
  assign n7038 = ~n6895 & ~n7037;
  assign n7039 = ~n7029 & ~n7038;
  assign n7040 = ~n6999 & n7039;
  assign n7041 = ~n7025 & ~n7040;
  assign n7042 = ~n7020 & n7041;
  assign n7043 = n7017 & n7042;
  assign n7044 = n6997 & n7043;
  assign n7045 = ~n6988 & n7044;
  assign n7046 = n6983 & n7045;
  assign n7047 = n7046 ^ n5397;
  assign n7048 = n7047 ^ x89;
  assign n7049 = ~n6892 & ~n7048;
  assign n7050 = n6630 & n7049;
  assign n7051 = n5961 & n7050;
  assign n7052 = n5592 ^ n5589;
  assign n7053 = n5641 & ~n7052;
  assign n7054 = ~n5626 & ~n5663;
  assign n7055 = ~n5592 & ~n7054;
  assign n7056 = n5589 & n5626;
  assign n7057 = n5627 & n7054;
  assign n7058 = ~n7056 & ~n7057;
  assign n7059 = ~n7055 & n7058;
  assign n7060 = ~n5593 & n7059;
  assign n7061 = n5566 & n7060;
  assign n7062 = n5590 & n5627;
  assign n7063 = ~n5625 & n7062;
  assign n7064 = ~n5592 & n5626;
  assign n7065 = n5666 & ~n7064;
  assign n7066 = ~n7063 & n7065;
  assign n7067 = n5662 & ~n7066;
  assign n7068 = ~n7061 & ~n7067;
  assign n7069 = n5592 ^ n5590;
  assign n7070 = n5629 ^ n5625;
  assign n7071 = n5590 ^ n5589;
  assign n7072 = n7071 ^ n5625;
  assign n7073 = n7072 ^ n5625;
  assign n7074 = n7073 ^ n5625;
  assign n7075 = n7070 & ~n7074;
  assign n7076 = n7075 ^ n5625;
  assign n7077 = n7069 & ~n7076;
  assign n7078 = n7077 ^ n7072;
  assign n7079 = n5634 & n7078;
  assign n7080 = n5592 & n5626;
  assign n7081 = ~n5591 & ~n5638;
  assign n7082 = ~n5625 & ~n7081;
  assign n7083 = ~n7080 & ~n7082;
  assign n7084 = n5651 & ~n7083;
  assign n7085 = ~n7079 & ~n7084;
  assign n7086 = n7068 & n7085;
  assign n7087 = ~n7053 & n7086;
  assign n7088 = n7087 ^ n4037;
  assign n7089 = n7088 ^ x85;
  assign n7090 = n5561 ^ x67;
  assign n7091 = ~n7089 & n7090;
  assign n7092 = n5056 & ~n5100;
  assign n7093 = ~n4878 & ~n5055;
  assign n7094 = n5090 & ~n7093;
  assign n7095 = n5056 & n5084;
  assign n7096 = n5063 & n5106;
  assign n7097 = ~n7095 & ~n7096;
  assign n7098 = ~n5074 & n5118;
  assign n7099 = n7098 ^ n5010;
  assign n7100 = n7099 ^ n7098;
  assign n7101 = n5075 & ~n5099;
  assign n7102 = n7101 ^ n7098;
  assign n7103 = ~n7100 & n7102;
  assign n7104 = n7103 ^ n7098;
  assign n7105 = ~n5052 & ~n7104;
  assign n7106 = n7097 & ~n7105;
  assign n7107 = n5102 & n7106;
  assign n7108 = n5965 & n7107;
  assign n7109 = n5065 & n7108;
  assign n7110 = ~n7094 & n7109;
  assign n7111 = ~n7092 & n7110;
  assign n7112 = n5084 ^ n5063;
  assign n7113 = n5086 ^ n5058;
  assign n7114 = n5063 ^ n5058;
  assign n7115 = n7114 ^ n5058;
  assign n7116 = ~n7113 & n7115;
  assign n7117 = n7116 ^ n5058;
  assign n7118 = n7112 & ~n7117;
  assign n7119 = n7118 ^ n5084;
  assign n7120 = n7111 & ~n7119;
  assign n7121 = n6727 & n7120;
  assign n7122 = n6725 & n7121;
  assign n7123 = ~n5079 & n7122;
  assign n7124 = n7123 ^ n4244;
  assign n7125 = n7124 ^ x102;
  assign n7126 = ~n6362 & n6370;
  assign n7127 = n6320 & ~n7126;
  assign n7128 = ~n6356 & n6373;
  assign n7129 = n6330 & ~n7128;
  assign n7130 = ~n7127 & ~n7129;
  assign n7131 = n6324 & n6376;
  assign n7132 = n6359 & ~n6938;
  assign n7133 = ~n6335 & n7132;
  assign n7134 = n6369 & ~n7133;
  assign n7135 = ~n7131 & ~n7134;
  assign n7136 = n7130 & n7135;
  assign n7137 = ~n6347 & n7136;
  assign n7138 = n6342 & n7137;
  assign n7139 = ~n6940 & n7138;
  assign n7140 = n6937 & n7139;
  assign n7141 = n7140 ^ n3921;
  assign n7142 = n7141 ^ x109;
  assign n7143 = n7125 & n7142;
  assign n7144 = n4619 ^ x68;
  assign n7145 = ~n6229 & n6636;
  assign n7146 = ~n6212 & n7145;
  assign n7147 = n6203 & ~n7146;
  assign n7148 = ~n6209 & ~n6243;
  assign n7149 = ~n6911 & ~n7148;
  assign n7150 = ~n6266 & n7149;
  assign n7151 = n6245 & n6250;
  assign n7152 = n6230 & n7151;
  assign n7153 = n6123 & ~n7152;
  assign n7154 = ~n7150 & ~n7153;
  assign n7155 = ~n7147 & n7154;
  assign n7156 = n6209 & ~n6256;
  assign n7157 = n6156 ^ n6155;
  assign n7158 = n6197 ^ n6156;
  assign n7159 = n7158 ^ n6156;
  assign n7160 = n7157 & n7159;
  assign n7161 = n7160 ^ n6156;
  assign n7162 = n6199 & n7161;
  assign n7163 = n7162 ^ n6156;
  assign n7164 = n6242 & n7163;
  assign n7165 = ~n7156 & ~n7164;
  assign n7166 = n7155 & n7165;
  assign n7167 = ~n6897 & n7166;
  assign n7168 = n6634 & n7167;
  assign n7169 = n6221 & n7168;
  assign n7170 = ~n6631 & n7169;
  assign n7171 = n6208 & n7170;
  assign n7172 = n7171 ^ n4208;
  assign n7173 = n7172 ^ x116;
  assign n7174 = ~n7144 & ~n7173;
  assign n7175 = n7143 & n7174;
  assign n7176 = n7091 & n7175;
  assign n7177 = ~n7144 & n7173;
  assign n7178 = ~n7125 & ~n7142;
  assign n7179 = n7177 & n7178;
  assign n7180 = n7090 & n7179;
  assign n7181 = ~n7176 & ~n7180;
  assign n7182 = ~n7125 & n7142;
  assign n7183 = n7174 & n7182;
  assign n7184 = n7174 & n7178;
  assign n7185 = ~n7183 & ~n7184;
  assign n7186 = n7091 & ~n7185;
  assign n7187 = n7089 & n7090;
  assign n7188 = ~n7089 & ~n7090;
  assign n7189 = ~n7187 & ~n7188;
  assign n7190 = n7142 ^ n7125;
  assign n7191 = n7177 & n7190;
  assign n7192 = ~n7183 & ~n7191;
  assign n7193 = ~n7189 & ~n7192;
  assign n7194 = n7089 & ~n7090;
  assign n7195 = n7144 & n7173;
  assign n7196 = n7182 & n7195;
  assign n7197 = n7144 & ~n7173;
  assign n7198 = n7143 & n7197;
  assign n7199 = n7178 & n7197;
  assign n7200 = ~n7198 & ~n7199;
  assign n7201 = n7143 & n7177;
  assign n7202 = n7125 & ~n7142;
  assign n7203 = n7174 & n7202;
  assign n7204 = ~n7201 & ~n7203;
  assign n7205 = n7200 & n7204;
  assign n7206 = ~n7179 & n7205;
  assign n7207 = ~n7196 & n7206;
  assign n7208 = ~n7175 & n7207;
  assign n7209 = n7194 & ~n7208;
  assign n7210 = n7195 & n7202;
  assign n7211 = n7143 & n7195;
  assign n7212 = n7200 & ~n7211;
  assign n7213 = ~n7210 & n7212;
  assign n7214 = n7188 & ~n7213;
  assign n7215 = n7211 ^ n7090;
  assign n7217 = n7197 & n7202;
  assign n7220 = n7178 & n7195;
  assign n7221 = ~n7217 & ~n7220;
  assign n7222 = ~n7196 & n7221;
  assign n7216 = n7182 & n7197;
  assign n7218 = ~n7216 & ~n7217;
  assign n7219 = ~n7210 & n7218;
  assign n7223 = n7222 ^ n7219;
  assign n7224 = n7222 ^ n7089;
  assign n7225 = n7224 ^ n7222;
  assign n7226 = n7223 & n7225;
  assign n7227 = n7226 ^ n7222;
  assign n7228 = n7227 ^ n7211;
  assign n7229 = ~n7215 & ~n7228;
  assign n7230 = n7229 ^ n7226;
  assign n7231 = n7230 ^ n7222;
  assign n7232 = n7231 ^ n7090;
  assign n7233 = ~n7211 & n7232;
  assign n7234 = n7233 ^ n7211;
  assign n7235 = n7234 ^ n7090;
  assign n7236 = ~n7214 & n7235;
  assign n7237 = ~n7209 & n7236;
  assign n7238 = ~n7193 & n7237;
  assign n7239 = ~n7186 & n7238;
  assign n7240 = n7175 ^ n7089;
  assign n7241 = n7240 ^ n7175;
  assign n7242 = n7210 ^ n7175;
  assign n7243 = n7241 & n7242;
  assign n7244 = n7243 ^ n7175;
  assign n7245 = ~n7090 & n7244;
  assign n7246 = n7239 & ~n7245;
  assign n7247 = n7181 & n7246;
  assign n7248 = n7247 ^ n5451;
  assign n7249 = n7248 ^ x122;
  assign n7250 = n5961 & ~n7249;
  assign n7251 = n6434 & n6629;
  assign n7252 = n6892 & ~n7048;
  assign n7253 = n7251 & n7252;
  assign n7254 = n7250 & n7253;
  assign n7255 = ~n7051 & ~n7254;
  assign n7256 = n6892 & n7048;
  assign n7257 = n6630 & n7256;
  assign n7258 = n7250 & n7257;
  assign n7259 = ~n5961 & n7249;
  assign n7260 = n6630 & n7252;
  assign n7261 = ~n6434 & n6629;
  assign n7262 = n7048 ^ n6892;
  assign n7263 = n7261 & ~n7262;
  assign n7264 = ~n7253 & ~n7257;
  assign n7265 = ~n7263 & n7264;
  assign n7266 = ~n6434 & ~n6629;
  assign n7267 = n7256 & n7266;
  assign n7268 = ~n6892 & n7048;
  assign n7269 = n6630 & n7268;
  assign n7270 = n7049 & n7251;
  assign n7271 = ~n7269 & ~n7270;
  assign n7272 = ~n7267 & n7271;
  assign n7273 = n7265 & n7272;
  assign n7274 = ~n7260 & n7273;
  assign n7275 = n7259 & ~n7274;
  assign n7276 = ~n7258 & ~n7275;
  assign n7277 = n7251 & n7256;
  assign n7278 = n5961 & n7277;
  assign n7279 = ~n5961 & ~n7249;
  assign n7280 = ~n7270 & ~n7277;
  assign n7281 = ~n7260 & n7280;
  assign n7282 = n7279 & ~n7281;
  assign n7283 = n7249 ^ n5961;
  assign n7284 = n7251 & n7268;
  assign n7285 = ~n7283 & n7284;
  assign n7286 = n7252 & n7266;
  assign n7287 = n7266 & n7268;
  assign n7288 = ~n7267 & ~n7287;
  assign n7290 = n7261 & n7268;
  assign n7289 = n7252 & n7261;
  assign n7291 = n7290 ^ n7289;
  assign n7292 = n7289 ^ n7250;
  assign n7293 = n7292 ^ n7250;
  assign n7294 = n7279 ^ n7250;
  assign n7295 = n7293 & ~n7294;
  assign n7296 = n7295 ^ n7250;
  assign n7297 = n7291 & ~n7296;
  assign n7298 = n7297 ^ n7290;
  assign n7299 = n7288 & ~n7298;
  assign n7300 = ~n7286 & n7299;
  assign n7301 = n7300 ^ n5961;
  assign n7302 = n7301 ^ n7300;
  assign n7303 = n7256 & n7261;
  assign n7304 = n7049 & n7266;
  assign n7305 = ~n7303 & ~n7304;
  assign n7306 = ~n7287 & n7305;
  assign n7307 = ~n7286 & n7306;
  assign n7308 = ~n7253 & n7307;
  assign n7309 = n7308 ^ n7300;
  assign n7310 = n7309 ^ n7300;
  assign n7311 = n7302 & ~n7310;
  assign n7312 = n7311 ^ n7300;
  assign n7313 = n7249 & ~n7312;
  assign n7314 = n7313 ^ n7300;
  assign n7315 = ~n7285 & n7314;
  assign n7316 = ~n7282 & n7315;
  assign n7317 = ~n7278 & n7316;
  assign n7318 = n7276 & n7317;
  assign n7319 = n7255 & n7318;
  assign n7320 = n7319 ^ n6282;
  assign n7321 = n7320 ^ x65;
  assign n7922 = ~n7089 & n7220;
  assign n7923 = n7188 & n7211;
  assign n7924 = n7177 & n7202;
  assign n7925 = ~n7183 & ~n7924;
  assign n7926 = n7194 & ~n7925;
  assign n7927 = ~n7923 & ~n7926;
  assign n7928 = ~n7922 & n7927;
  assign n8431 = n7188 & n7196;
  assign n8432 = ~n7179 & ~n7201;
  assign n8433 = n7194 & ~n8432;
  assign n8434 = ~n8431 & ~n8433;
  assign n8435 = n7091 & ~n7212;
  assign n8436 = ~n7189 & n7199;
  assign n8437 = ~n7198 & ~n7210;
  assign n8438 = ~n7188 & n8432;
  assign n8439 = n8437 & n8438;
  assign n8440 = ~n7216 & n8439;
  assign n8441 = n7187 & ~n8440;
  assign n8442 = ~n7175 & n7192;
  assign n8443 = n7091 & ~n8442;
  assign n8444 = n7218 & n8437;
  assign n8445 = n7194 & ~n8444;
  assign n8446 = ~n8443 & ~n8445;
  assign n8447 = n7177 & n7182;
  assign n8448 = ~n7203 & ~n8447;
  assign n7935 = ~n7175 & ~n7184;
  assign n8449 = ~n7935 & ~n8438;
  assign n8450 = n8448 & ~n8449;
  assign n8451 = ~n7189 & ~n8450;
  assign n8452 = n8446 & ~n8451;
  assign n8453 = ~n8441 & n8452;
  assign n8454 = ~n8436 & n8453;
  assign n8455 = ~n8435 & n8454;
  assign n8456 = n8434 & n8455;
  assign n8457 = n7928 & n8456;
  assign n8458 = n8457 ^ n6313;
  assign n8459 = n8458 ^ x101;
  assign n7995 = n6037 ^ n6004;
  assign n7996 = n6072 ^ n6004;
  assign n7997 = n7996 ^ n6037;
  assign n7998 = n7997 ^ n6004;
  assign n7999 = n7998 ^ n6004;
  assign n8000 = n7995 & ~n7999;
  assign n8001 = n8000 ^ n6004;
  assign n8002 = n6114 & n8001;
  assign n8003 = n8002 ^ n7997;
  assign n8460 = n6415 & ~n8003;
  assign n8005 = n6392 & n6396;
  assign n8006 = ~n6037 & ~n6114;
  assign n8007 = ~n6072 & n8006;
  assign n8008 = ~n6394 & ~n8007;
  assign n8009 = ~n8005 & n8008;
  assign n8010 = n6407 & n8009;
  assign n8011 = ~n6391 & n8010;
  assign n8461 = n6403 & ~n8011;
  assign n8462 = ~n8460 & ~n8461;
  assign n8014 = n6072 & n6117;
  assign n8015 = n6425 & ~n8014;
  assign n8016 = ~n6116 & n8008;
  assign n8017 = n8015 & n8016;
  assign n8018 = n8017 ^ n6385;
  assign n8019 = n8018 ^ n8017;
  assign n8020 = n6392 & ~n7995;
  assign n8021 = ~n6114 & n6387;
  assign n8022 = ~n8020 & ~n8021;
  assign n8023 = n8016 & n8022;
  assign n8024 = n8023 ^ n8017;
  assign n8025 = n8019 & ~n8024;
  assign n8026 = n8025 ^ n8017;
  assign n8463 = n6283 & n8026;
  assign n8464 = n8462 & ~n8463;
  assign n8465 = n8464 ^ n6291;
  assign n8466 = n8465 ^ x76;
  assign n7323 = n6700 & n6862;
  assign n7324 = n6844 & n6851;
  assign n7325 = ~n7323 & ~n7324;
  assign n8210 = n6700 & n6836;
  assign n7326 = ~n6843 & ~n6868;
  assign n8211 = n6854 & n7326;
  assign n8212 = n6828 & ~n8211;
  assign n8213 = ~n6843 & ~n6852;
  assign n8214 = ~n6861 & n8213;
  assign n8215 = n6700 & ~n8214;
  assign n8216 = ~n6837 & n6856;
  assign n8217 = ~n6827 & n8216;
  assign n8218 = n6844 & ~n8217;
  assign n8219 = ~n8215 & ~n8218;
  assign n7337 = n6826 & n6831;
  assign n8036 = ~n6872 & ~n7337;
  assign n8220 = n6699 & ~n8036;
  assign n8221 = ~n6823 & ~n6836;
  assign n8222 = n6828 & ~n8221;
  assign n7322 = n6828 & n6837;
  assign n8039 = ~n6848 & ~n6861;
  assign n8223 = ~n6862 & n8039;
  assign n8224 = ~n6832 & n8223;
  assign n8225 = n6846 & ~n8224;
  assign n8226 = ~n7322 & ~n8225;
  assign n8227 = n6830 & n8226;
  assign n8228 = ~n8222 & n8227;
  assign n8229 = ~n8220 & n8228;
  assign n8230 = n8219 & n8229;
  assign n8231 = ~n8212 & n8230;
  assign n8232 = ~n8210 & n8231;
  assign n8233 = n6850 ^ n6846;
  assign n8234 = n6851 ^ n6850;
  assign n8235 = n8234 ^ n6851;
  assign n8236 = n6851 ^ n6844;
  assign n8237 = n8235 & ~n8236;
  assign n8238 = n8237 ^ n6851;
  assign n8239 = n8233 & ~n8238;
  assign n8240 = n8239 ^ n6846;
  assign n8241 = n8232 & ~n8240;
  assign n8242 = n7325 & n8241;
  assign n8243 = n8242 ^ n5724;
  assign n8467 = n8243 ^ x116;
  assign n8468 = ~n8466 & n8467;
  assign n7359 = n6578 & n6596;
  assign n7360 = n6562 & n6591;
  assign n7361 = ~n7359 & ~n7360;
  assign n7362 = n6517 & n6586;
  assign n7363 = n7361 & ~n7362;
  assign n8469 = ~n6581 & ~n6584;
  assign n8470 = n6585 & ~n8469;
  assign n8471 = n6562 & ~n6616;
  assign n8472 = ~n6576 & ~n6586;
  assign n8473 = ~n8471 & ~n8472;
  assign n7377 = ~n6590 & ~n6614;
  assign n8474 = ~n6596 & n7377;
  assign n8475 = ~n6589 & n8474;
  assign n8476 = n6585 & ~n8475;
  assign n8477 = n6571 & ~n6598;
  assign n8478 = ~n8476 & ~n8477;
  assign n7364 = ~n6575 & ~n6584;
  assign n7365 = ~n6603 & n7364;
  assign n7366 = ~n6581 & n7365;
  assign n8479 = n6615 & n7366;
  assign n8480 = n8479 ^ n6605;
  assign n8481 = n8480 ^ n6605;
  assign n8482 = n6605 ^ n6561;
  assign n8483 = n8482 ^ n6605;
  assign n8484 = ~n8481 & n8483;
  assign n8485 = n8484 ^ n6605;
  assign n8486 = ~n6518 & ~n8485;
  assign n8487 = n8486 ^ n6605;
  assign n8488 = n8478 & n8487;
  assign n8489 = n8473 & n8488;
  assign n8490 = ~n8470 & n8489;
  assign n8491 = ~n6572 & n8490;
  assign n8492 = n7363 & n8491;
  assign n8493 = ~n6595 & n8492;
  assign n8494 = n8493 ^ n3669;
  assign n8495 = n8494 ^ x94;
  assign n8496 = n8468 & n8495;
  assign n8497 = ~n8459 & n8496;
  assign n8498 = ~n8466 & ~n8467;
  assign n8499 = n8459 & n8495;
  assign n8500 = n8498 & n8499;
  assign n8501 = ~n8497 & ~n8500;
  assign n7674 = n6036 ^ x114;
  assign n7675 = n6820 ^ x88;
  assign n7741 = n7674 & ~n7675;
  assign n7677 = n5651 & ~n7078;
  assign n7678 = n7066 ^ n5564;
  assign n7679 = n7678 ^ n7066;
  assign n7680 = n7083 ^ n7066;
  assign n7681 = n7679 & n7680;
  assign n7682 = n7681 ^ n7066;
  assign n7683 = n5565 & ~n7682;
  assign n7684 = ~n7677 & ~n7683;
  assign n7685 = n7060 ^ n7053;
  assign n7686 = n7685 ^ n7053;
  assign n7687 = n7053 ^ n5564;
  assign n7688 = n7687 ^ n7053;
  assign n7689 = ~n7686 & ~n7688;
  assign n7690 = n7689 ^ n7053;
  assign n7691 = ~n5565 & n7690;
  assign n7692 = n7691 ^ n7053;
  assign n7693 = n7684 & ~n7692;
  assign n7694 = n7693 ^ n3738;
  assign n7695 = n7694 ^ x82;
  assign n7696 = n4549 & ~n4557;
  assign n7697 = ~n4560 & ~n4593;
  assign n7698 = n3265 & ~n7697;
  assign n7699 = ~n7696 & ~n7698;
  assign n7700 = n4551 & n4581;
  assign n7701 = ~n4566 & ~n4578;
  assign n7702 = ~n4590 & n7701;
  assign n7703 = n4556 & ~n7702;
  assign n7704 = ~n7700 & ~n7703;
  assign n7705 = n7699 & n7704;
  assign n7706 = n6678 ^ n3670;
  assign n7707 = n7706 ^ n6678;
  assign n7708 = n6678 ^ n6454;
  assign n7709 = n7707 & n7708;
  assign n7710 = n7709 ^ n6678;
  assign n7711 = ~n3265 & ~n7710;
  assign n7712 = n7705 & ~n7711;
  assign n7713 = ~n6436 & n7712;
  assign n7714 = n6662 & n7713;
  assign n7715 = n4577 & n7714;
  assign n7716 = ~n4614 & n7715;
  assign n7717 = n6444 & n7716;
  assign n7718 = ~n4546 & n7717;
  assign n7719 = n7718 ^ n3774;
  assign n7720 = n7719 ^ x81;
  assign n7721 = n7695 & n7720;
  assign n7722 = n6384 ^ x64;
  assign n7723 = n6658 ^ x120;
  assign n7724 = ~n7722 & ~n7723;
  assign n7725 = n7721 & n7724;
  assign n7728 = ~n7695 & ~n7720;
  assign n7729 = n7722 & ~n7723;
  assign n7730 = n7728 & n7729;
  assign n7742 = ~n7725 & ~n7730;
  assign n7743 = n7741 & ~n7742;
  assign n7727 = ~n7674 & n7675;
  assign n7731 = n7727 & n7730;
  assign n7732 = n7674 & n7675;
  assign n7733 = n7695 & ~n7720;
  assign n7734 = ~n7722 & n7723;
  assign n7735 = n7733 & n7734;
  assign n7736 = n7722 & n7723;
  assign n7737 = n7728 & n7736;
  assign n7738 = ~n7735 & ~n7737;
  assign n7739 = n7732 & ~n7738;
  assign n7740 = ~n7731 & ~n7739;
  assign n7676 = ~n7674 & ~n7675;
  assign n8286 = n7676 & n7730;
  assign n8287 = n7740 & ~n8286;
  assign n7780 = n7721 & n7729;
  assign n8502 = ~n7674 & n7780;
  assign n7752 = ~n7727 & ~n7741;
  assign n7749 = ~n7695 & n7720;
  assign n7765 = n7724 & n7749;
  assign n8503 = ~n7752 & n7765;
  assign n8504 = ~n8502 & ~n8503;
  assign n7766 = n7729 & n7733;
  assign n8505 = n7741 & n7766;
  assign n7759 = n7729 & n7749;
  assign n8506 = n7727 & n7759;
  assign n7750 = n7736 & n7749;
  assign n7953 = n7750 & ~n7752;
  assign n7746 = n7724 & n7728;
  assign n7777 = n7675 ^ n7674;
  assign n8507 = n7746 & ~n7777;
  assign n7754 = n7734 & n7749;
  assign n7755 = n7721 & n7736;
  assign n7756 = ~n7754 & ~n7755;
  assign n7758 = n7724 & n7733;
  assign n8508 = n7738 & ~n7758;
  assign n8509 = n7756 & n8508;
  assign n8510 = n7676 & ~n8509;
  assign n8511 = ~n8507 & ~n8510;
  assign n7744 = n7721 & n7734;
  assign n7753 = n7733 & n7736;
  assign n7764 = n7728 & n7734;
  assign n8512 = ~n7753 & ~n7764;
  assign n8513 = ~n7744 & n8512;
  assign n8514 = ~n7752 & ~n8513;
  assign n7760 = ~n7758 & ~n7759;
  assign n7956 = n7760 & ~n7780;
  assign n7971 = ~n7744 & ~n7765;
  assign n8515 = n7956 & n7971;
  assign n8516 = n7732 & ~n8515;
  assign n8517 = ~n8514 & ~n8516;
  assign n8518 = n8511 & n8517;
  assign n8519 = ~n7953 & n8518;
  assign n8520 = ~n8506 & n8519;
  assign n8521 = ~n8505 & n8520;
  assign n8522 = n8504 & n8521;
  assign n8523 = n8287 & n8522;
  assign n8524 = ~n7743 & n8523;
  assign n8525 = n8524 ^ n3885;
  assign n8526 = n8525 ^ x67;
  assign n8102 = n6895 & n7011;
  assign n8103 = n6975 & ~n7007;
  assign n8104 = ~n8102 & ~n8103;
  assign n7568 = n6895 & ~n6981;
  assign n7569 = ~n7018 & ~n7021;
  assign n7570 = n6895 & ~n7569;
  assign n7571 = ~n7568 & ~n7570;
  assign n7572 = n6893 & n7022;
  assign n7573 = n6997 & ~n7572;
  assign n8322 = n6999 & n7010;
  assign n7576 = ~n6973 & ~n6993;
  assign n8323 = n7023 & n7576;
  assign n8324 = n6975 & ~n8323;
  assign n8325 = ~n8322 & ~n8324;
  assign n8326 = n6998 & ~n7019;
  assign n8327 = ~n6973 & ~n8326;
  assign n8328 = ~n6978 & n8327;
  assign n8329 = n8328 ^ n6894;
  assign n8330 = n8329 ^ n8328;
  assign n8331 = n8328 ^ n7006;
  assign n8332 = n8331 ^ n8328;
  assign n8333 = n8330 & n8332;
  assign n8334 = n8333 ^ n8328;
  assign n8335 = ~n6893 & ~n8334;
  assign n8336 = n8335 ^ n8328;
  assign n8337 = n8325 & n8336;
  assign n8338 = n7026 ^ n6998;
  assign n8339 = n7026 ^ n6895;
  assign n8340 = n8339 ^ n6895;
  assign n8341 = n7000 ^ n6895;
  assign n8342 = n8340 & ~n8341;
  assign n8343 = n8342 ^ n6895;
  assign n8344 = ~n8338 & n8343;
  assign n8345 = n8344 ^ n6998;
  assign n8346 = n8337 & ~n8345;
  assign n8347 = n7573 & n8346;
  assign n8348 = n7571 & n8347;
  assign n8349 = ~n6988 & n8348;
  assign n8350 = n8104 & n8349;
  assign n8351 = n8350 ^ n5822;
  assign n8527 = n8351 ^ x125;
  assign n8528 = n8526 & n8527;
  assign n8529 = ~n8501 & n8528;
  assign n8530 = n8466 & n8467;
  assign n8531 = n8495 & n8530;
  assign n8532 = ~n8459 & n8531;
  assign n8533 = ~n8459 & ~n8467;
  assign n8534 = ~n8466 & n8533;
  assign n8535 = n8495 & n8534;
  assign n8536 = ~n8532 & ~n8535;
  assign n8537 = ~n8526 & n8527;
  assign n8538 = ~n8536 & n8537;
  assign n8539 = ~n8529 & ~n8538;
  assign n8540 = ~n8495 & n8498;
  assign n8541 = n8459 & n8540;
  assign n8542 = n8537 & n8541;
  assign n8543 = n8466 & n8533;
  assign n8544 = n8495 & n8543;
  assign n8545 = n8526 & ~n8527;
  assign n8546 = ~n8537 & ~n8545;
  assign n8547 = n8544 & n8546;
  assign n8548 = ~n8542 & ~n8547;
  assign n8549 = n8468 & ~n8495;
  assign n8550 = n8459 & n8549;
  assign n8551 = n8466 & ~n8495;
  assign n8552 = n8467 & n8551;
  assign n8553 = ~n8459 & n8552;
  assign n8554 = ~n8550 & ~n8553;
  assign n8555 = ~n8459 & n8549;
  assign n8556 = ~n8467 & n8551;
  assign n8557 = n8459 & n8556;
  assign n8558 = ~n8555 & ~n8557;
  assign n8559 = ~n8500 & n8558;
  assign n8560 = n8554 & n8559;
  assign n8561 = n8537 & ~n8560;
  assign n8562 = ~n8467 & n8499;
  assign n8563 = n8466 & n8562;
  assign n8564 = n8528 & n8563;
  assign n8565 = ~n8526 & ~n8527;
  assign n8566 = n8468 & n8499;
  assign n8567 = ~n8563 & ~n8566;
  assign n8568 = ~n8497 & ~n8553;
  assign n8569 = ~n8541 & n8558;
  assign n8570 = n8568 & n8569;
  assign n8571 = n8567 & n8570;
  assign n8572 = n8565 & ~n8571;
  assign n8573 = ~n8564 & ~n8572;
  assign n8574 = ~n8561 & n8573;
  assign n8575 = ~n8495 & n8534;
  assign n8576 = ~n8552 & ~n8575;
  assign n8577 = ~n8541 & n8576;
  assign n8578 = n8577 ^ n8527;
  assign n8579 = n8578 ^ n8577;
  assign n8580 = ~n8532 & ~n8563;
  assign n8581 = ~n8550 & n8580;
  assign n8582 = n8577 & n8581;
  assign n8583 = ~n8497 & n8582;
  assign n8584 = n8583 ^ n8577;
  assign n8585 = ~n8579 & ~n8584;
  assign n8586 = n8585 ^ n8577;
  assign n8587 = n8526 & ~n8586;
  assign n8588 = n8574 & ~n8587;
  assign n8589 = n8548 & n8588;
  assign n8590 = n8539 & n8589;
  assign n8591 = n8590 ^ n6384;
  assign n8592 = n8591 ^ x112;
  assign n7327 = ~n6852 & n7326;
  assign n7328 = ~n6850 & n7327;
  assign n7329 = n6700 & ~n7328;
  assign n7330 = ~n6700 & ~n6823;
  assign n7331 = ~n6845 & n7330;
  assign n7332 = n6854 & n7331;
  assign n7333 = ~n6867 & ~n7332;
  assign n7334 = ~n7329 & ~n7333;
  assign n7335 = ~n6861 & ~n6872;
  assign n7336 = n6846 & ~n7335;
  assign n7338 = n6863 & ~n7337;
  assign n7339 = ~n6867 & ~n7338;
  assign n7340 = n6821 ^ n6789;
  assign n7341 = n6750 ^ n6723;
  assign n7342 = n7341 ^ n6821;
  assign n7343 = n7342 ^ n7341;
  assign n7344 = n7341 ^ n6750;
  assign n7345 = n7344 ^ n7341;
  assign n7346 = n7343 & n7345;
  assign n7347 = n7346 ^ n7341;
  assign n7348 = n7340 & n7347;
  assign n7349 = n7348 ^ n7341;
  assign n7350 = n6828 & n7349;
  assign n7351 = ~n7339 & ~n7350;
  assign n7352 = ~n7336 & n7351;
  assign n7353 = n7334 & n7352;
  assign n7354 = n7325 & n7353;
  assign n7355 = n6841 & n7354;
  assign n7356 = ~n7322 & n7355;
  assign n7357 = n7356 ^ n5009;
  assign n7358 = n7357 ^ x98;
  assign n7367 = ~n6614 & n7366;
  assign n7368 = ~n6597 & n7367;
  assign n7369 = n6562 & ~n7368;
  assign n7370 = ~n6569 & ~n6604;
  assign n7371 = ~n6581 & n7370;
  assign n7372 = n6616 & n7371;
  assign n7373 = ~n6590 & n7372;
  assign n7374 = ~n6574 & n7373;
  assign n7375 = n6585 & ~n7374;
  assign n7376 = ~n7369 & ~n7375;
  assign n7378 = n6578 & ~n7377;
  assign n7379 = n6592 & ~n6604;
  assign n7380 = n6571 & ~n7379;
  assign n7381 = ~n6578 & n7364;
  assign n7382 = ~n6566 & n6599;
  assign n7383 = ~n6589 & n7382;
  assign n7384 = ~n6571 & n7383;
  assign n7385 = ~n7381 & ~n7384;
  assign n7386 = n6586 & n7385;
  assign n7387 = ~n7380 & ~n7386;
  assign n7388 = ~n7378 & n7387;
  assign n7389 = n7376 & n7388;
  assign n7390 = n6573 & n7389;
  assign n7391 = n7363 & n7390;
  assign n7392 = n7391 ^ n5050;
  assign n7393 = n7392 ^ x72;
  assign n7394 = n7358 & ~n7393;
  assign n7395 = ~n4620 & ~n5133;
  assign n7396 = n5895 & n5906;
  assign n7397 = n7395 & n7396;
  assign n7398 = ~n5892 & ~n5920;
  assign n7399 = n5894 & ~n7398;
  assign n7400 = ~n7397 & ~n7399;
  assign n7401 = ~n5917 & n7395;
  assign n7402 = ~n5914 & ~n7401;
  assign n7403 = n5902 & n7395;
  assign n7404 = n5134 & n5944;
  assign n7405 = ~n7403 & ~n7404;
  assign n7406 = ~n5928 & ~n7396;
  assign n7407 = n5894 & ~n7406;
  assign n7408 = ~n5899 & ~n5925;
  assign n7409 = n5905 & ~n7408;
  assign n7410 = n5563 & n5896;
  assign n7411 = ~n5946 & n7398;
  assign n7412 = ~n7410 & n7411;
  assign n7413 = ~n5133 & ~n7412;
  assign n7414 = ~n7409 & ~n7413;
  assign n7415 = ~n7407 & n7414;
  assign n7416 = n7405 & n7415;
  assign n7417 = n7402 & n7416;
  assign n7418 = n5912 & n7417;
  assign n7419 = n7400 & n7418;
  assign n7420 = n7419 ^ n4649;
  assign n7421 = n7420 ^ x113;
  assign n7422 = n6722 ^ x73;
  assign n7423 = n7141 ^ x66;
  assign n7424 = n7422 & ~n7423;
  assign n7425 = n7088 ^ x107;
  assign n7426 = n6698 ^ x105;
  assign n7427 = ~n7425 & n7426;
  assign n7428 = ~n5325 & n5329;
  assign n7429 = n5300 & ~n5315;
  assign n7430 = ~n7428 & ~n7429;
  assign n7431 = ~n5304 & ~n5322;
  assign n7432 = n5312 & ~n7431;
  assign n7433 = ~n5328 & n6808;
  assign n7434 = n5291 & ~n7433;
  assign n7435 = ~n7432 & ~n7434;
  assign n7436 = n5340 & n6790;
  assign n7437 = ~n5289 & n7436;
  assign n7438 = n7437 ^ n5309;
  assign n7439 = n7438 ^ n5309;
  assign n7440 = n5309 ^ n5180;
  assign n7441 = n7440 ^ n5309;
  assign n7442 = ~n7439 & ~n7441;
  assign n7443 = n7442 ^ n5309;
  assign n7444 = n5179 & n7443;
  assign n7445 = n7444 ^ n5309;
  assign n7446 = n7435 & ~n7445;
  assign n7447 = n7430 & n7446;
  assign n7448 = n5321 & n7447;
  assign n7449 = n6800 & n7448;
  assign n7450 = n6794 & n7449;
  assign n7451 = n6041 & n7450;
  assign n7452 = ~n6791 & n7451;
  assign n7453 = ~n5306 & n7452;
  assign n7454 = n7453 ^ n3982;
  assign n7455 = n7454 ^ x80;
  assign n7456 = ~n5503 & n6024;
  assign n7457 = n5399 & ~n7456;
  assign n7458 = n5500 & n5538;
  assign n7459 = ~n5486 & n7458;
  assign n7460 = n5488 & ~n7459;
  assign n7461 = ~n7457 & ~n7460;
  assign n7462 = n5492 & n5507;
  assign n7463 = ~n5536 & n6022;
  assign n7464 = ~n5492 & n7463;
  assign n7465 = ~n5509 & n5539;
  assign n7466 = ~n5505 & n7465;
  assign n7467 = ~n7464 & ~n7466;
  assign n7468 = ~n5496 & ~n7467;
  assign n7469 = ~n5529 & n7468;
  assign n7470 = ~n6019 & ~n7469;
  assign n7471 = ~n7462 & ~n7470;
  assign n7472 = n7461 & n7471;
  assign n7473 = n5526 & n7472;
  assign n7474 = n6013 & n7473;
  assign n7475 = n5514 & n7474;
  assign n7476 = n6007 & n7475;
  assign n7477 = ~n5487 & n7476;
  assign n7478 = n7477 ^ n4076;
  assign n7479 = n7478 ^ x90;
  assign n7480 = ~n7455 & n7479;
  assign n7481 = n7427 & n7480;
  assign n7482 = ~n7425 & ~n7426;
  assign n7483 = n7455 & ~n7479;
  assign n7484 = n7482 & n7483;
  assign n7485 = ~n7481 & ~n7484;
  assign n7486 = n7424 & ~n7485;
  assign n7487 = ~n7422 & n7423;
  assign n7488 = n7427 & n7483;
  assign n7489 = ~n7484 & ~n7488;
  assign n7490 = n7487 & ~n7489;
  assign n7491 = n7425 & n7426;
  assign n7492 = n7455 & n7479;
  assign n7493 = n7491 & n7492;
  assign n7494 = n7483 & n7491;
  assign n7495 = ~n7493 & ~n7494;
  assign n7496 = n7427 & n7492;
  assign n7497 = ~n7455 & ~n7479;
  assign n7498 = n7482 & n7497;
  assign n7499 = n7427 & n7497;
  assign n7500 = ~n7498 & ~n7499;
  assign n7501 = ~n7496 & n7500;
  assign n7502 = n7495 & n7501;
  assign n7503 = n7424 & ~n7502;
  assign n7504 = n7425 & ~n7426;
  assign n7505 = n7480 & n7504;
  assign n7506 = n7422 & n7423;
  assign n7507 = n7483 & n7504;
  assign n7508 = n7497 & n7504;
  assign n7509 = ~n7493 & ~n7508;
  assign n7510 = ~n7507 & n7509;
  assign n7511 = n7506 & ~n7510;
  assign n7512 = ~n7422 & ~n7423;
  assign n7513 = n7480 & n7491;
  assign n7514 = n7492 & n7504;
  assign n7515 = ~n7508 & ~n7514;
  assign n7516 = ~n7513 & n7515;
  assign n7517 = n7512 & ~n7516;
  assign n7518 = ~n7511 & ~n7517;
  assign n7519 = ~n7505 & n7518;
  assign n7520 = ~n7503 & n7519;
  assign n7521 = ~n7488 & ~n7507;
  assign n7522 = n7521 ^ n7423;
  assign n7523 = n7522 ^ n7521;
  assign n7524 = n7480 & n7482;
  assign n7525 = n7491 & n7497;
  assign n7526 = ~n7496 & ~n7513;
  assign n7527 = ~n7525 & n7526;
  assign n7528 = ~n7524 & n7527;
  assign n7529 = ~n7514 & n7528;
  assign n7530 = n7529 ^ n7521;
  assign n7531 = n7523 & n7530;
  assign n7532 = n7531 ^ n7521;
  assign n7533 = ~n7422 & ~n7532;
  assign n7534 = n7520 & ~n7533;
  assign n7535 = n7482 & n7492;
  assign n7536 = ~n7499 & ~n7535;
  assign n7537 = n7536 ^ n7506;
  assign n7538 = n7536 ^ n7512;
  assign n7539 = n7538 ^ n7512;
  assign n7540 = ~n7481 & ~n7524;
  assign n7541 = n7540 ^ n7512;
  assign n7542 = n7539 & n7541;
  assign n7543 = n7542 ^ n7512;
  assign n7544 = ~n7537 & n7543;
  assign n7545 = n7544 ^ n7506;
  assign n7546 = n7534 & ~n7545;
  assign n7547 = ~n7490 & n7546;
  assign n7548 = ~n7486 & n7547;
  assign n7549 = n7548 ^ n4680;
  assign n7550 = n7549 ^ x104;
  assign n7551 = ~n7421 & n7550;
  assign n7552 = n6386 & ~n6412;
  assign n7553 = n6427 ^ n6283;
  assign n7554 = n7553 ^ n6283;
  assign n7555 = n6415 ^ n6283;
  assign n7556 = n7555 ^ n6283;
  assign n7557 = n7554 & n7556;
  assign n7558 = n7557 ^ n6283;
  assign n7559 = n6120 & n7558;
  assign n7560 = n7559 ^ n6283;
  assign n7561 = ~n7552 & ~n7560;
  assign n7562 = ~n6421 & n6423;
  assign n7563 = ~n6401 & n6403;
  assign n7564 = ~n7562 & ~n7563;
  assign n7565 = n7561 & n7564;
  assign n7566 = n7565 ^ n4715;
  assign n7567 = n7566 ^ x66;
  assign n7574 = ~n7000 & ~n7010;
  assign n7575 = n6895 & ~n7574;
  assign n7577 = ~n6999 & ~n7576;
  assign n7578 = ~n7575 & ~n7577;
  assign n7579 = ~n6894 & n6994;
  assign n7580 = ~n6980 & ~n7002;
  assign n7581 = n7007 & n7580;
  assign n7582 = ~n7021 & n7581;
  assign n7583 = n6975 & ~n7582;
  assign n7584 = ~n7579 & ~n7583;
  assign n7585 = n6999 & n7011;
  assign n7586 = ~n7000 & n7028;
  assign n7587 = ~n7006 & n7574;
  assign n7588 = ~n6978 & n7587;
  assign n7589 = ~n6984 & n7588;
  assign n7590 = ~n7586 & ~n7589;
  assign n7591 = n6893 & n7590;
  assign n7592 = ~n7585 & ~n7591;
  assign n7593 = n7584 & n7592;
  assign n7594 = n7578 & n7593;
  assign n7595 = n7573 & n7594;
  assign n7596 = n7571 & n7595;
  assign n7597 = n7596 ^ n4875;
  assign n7598 = n7597 ^ x65;
  assign n7599 = n7567 & n7598;
  assign n7600 = n7551 & n7599;
  assign n7601 = ~n7421 & ~n7550;
  assign n7602 = n7567 & ~n7598;
  assign n7603 = n7601 & n7602;
  assign n7604 = ~n7600 & ~n7603;
  assign n7605 = n7394 & ~n7604;
  assign n7606 = ~n7358 & n7393;
  assign n7607 = n7421 & ~n7550;
  assign n7608 = n7602 & n7607;
  assign n7609 = ~n7567 & ~n7598;
  assign n7610 = n7601 & n7609;
  assign n7611 = n7607 & n7609;
  assign n7612 = ~n7610 & ~n7611;
  assign n7613 = ~n7608 & n7612;
  assign n7614 = n7606 & ~n7613;
  assign n7615 = ~n7605 & ~n7614;
  assign n7616 = ~n7358 & ~n7393;
  assign n7617 = n7599 & n7607;
  assign n7618 = n7599 & n7601;
  assign n7619 = ~n7567 & n7598;
  assign n7620 = n7607 & n7619;
  assign n7621 = ~n7603 & ~n7620;
  assign n7622 = ~n7618 & n7621;
  assign n7623 = ~n7617 & n7622;
  assign n7624 = n7616 & ~n7623;
  assign n7625 = n7421 & n7550;
  assign n7626 = n7619 & n7625;
  assign n7627 = n7394 & n7626;
  assign n7628 = n7599 & n7625;
  assign n7629 = n7606 & n7628;
  assign n7630 = ~n7627 & ~n7629;
  assign n7631 = n7609 & n7625;
  assign n7632 = n7616 & n7631;
  assign n7633 = ~n7394 & ~n7606;
  assign n7634 = n7551 & n7602;
  assign n7635 = ~n7631 & ~n7634;
  assign n7636 = ~n7628 & n7635;
  assign n7637 = ~n7606 & n7636;
  assign n7638 = n7602 & n7625;
  assign n7639 = ~n7626 & ~n7634;
  assign n7640 = ~n7638 & n7639;
  assign n7641 = ~n7394 & n7640;
  assign n7642 = ~n7637 & ~n7641;
  assign n7643 = ~n7633 & n7642;
  assign n7644 = ~n7632 & ~n7643;
  assign n7645 = n7393 ^ n7358;
  assign n7646 = n7551 & n7609;
  assign n7647 = n7551 & n7619;
  assign n7648 = ~n7638 & ~n7647;
  assign n7649 = ~n7646 & n7648;
  assign n7650 = ~n7645 & ~n7649;
  assign n7651 = n7358 & n7393;
  assign n7652 = ~n7610 & ~n7620;
  assign n7653 = ~n7634 & n7652;
  assign n7654 = ~n7618 & n7653;
  assign n7655 = ~n7617 & n7654;
  assign n7656 = n7651 & ~n7655;
  assign n7657 = ~n7650 & ~n7656;
  assign n7658 = n7644 & n7657;
  assign n7659 = n7630 & n7658;
  assign n7660 = ~n7624 & n7659;
  assign n7661 = n7615 & n7660;
  assign n7662 = n7601 & n7619;
  assign n7663 = n7662 ^ n7394;
  assign n7664 = n7662 ^ n7606;
  assign n7665 = n7664 ^ n7606;
  assign n7666 = n7611 ^ n7606;
  assign n7667 = ~n7665 & ~n7666;
  assign n7668 = n7667 ^ n7606;
  assign n7669 = n7663 & n7668;
  assign n7670 = n7669 ^ n7394;
  assign n7671 = n7661 & ~n7670;
  assign n7672 = n7671 ^ n6003;
  assign n7673 = n7672 ^ x107;
  assign n7726 = n7676 & n7725;
  assign n7745 = n7727 & n7744;
  assign n7747 = ~n7674 & n7746;
  assign n7748 = ~n7745 & ~n7747;
  assign n7751 = n7674 & n7750;
  assign n7757 = ~n7753 & n7756;
  assign n7761 = n7757 & n7760;
  assign n7762 = ~n7752 & ~n7761;
  assign n7763 = ~n7751 & ~n7762;
  assign n7767 = ~n7765 & ~n7766;
  assign n7768 = ~n7764 & n7767;
  assign n7769 = n7732 & ~n7768;
  assign n7770 = ~n7759 & ~n7766;
  assign n7771 = n7756 & n7770;
  assign n7772 = ~n7744 & n7771;
  assign n7773 = n7676 & ~n7772;
  assign n7774 = ~n7769 & ~n7773;
  assign n7775 = n7763 & n7774;
  assign n7776 = n7748 & n7775;
  assign n7778 = n7737 ^ n7675;
  assign n7779 = n7778 ^ n7737;
  assign n7781 = ~n7725 & ~n7780;
  assign n7782 = n7781 ^ n7737;
  assign n7783 = n7779 & ~n7782;
  assign n7784 = n7783 ^ n7737;
  assign n7785 = ~n7777 & n7784;
  assign n7786 = n7776 & ~n7785;
  assign n7787 = ~n7743 & n7786;
  assign n7788 = n7740 & n7787;
  assign n7789 = ~n7726 & n7788;
  assign n7790 = n7789 ^ n5422;
  assign n7791 = n7790 ^ x107;
  assign n7792 = n7392 ^ x88;
  assign n7793 = ~n7791 & n7792;
  assign n7794 = n7248 ^ x97;
  assign n7795 = n5896 & n5900;
  assign n7796 = n7395 & n7795;
  assign n7797 = n7410 ^ n5133;
  assign n7798 = n7797 ^ n7410;
  assign n7799 = n7410 ^ n5925;
  assign n7800 = n7799 ^ n7410;
  assign n7801 = n7798 & n7800;
  assign n7802 = n7801 ^ n7410;
  assign n7803 = ~n5915 & n7802;
  assign n7804 = n7803 ^ n7410;
  assign n7805 = ~n7796 & ~n7804;
  assign n7806 = n5905 & n5942;
  assign n7807 = ~n5928 & n5947;
  assign n7808 = n5915 & ~n7807;
  assign n7809 = ~n7806 & ~n7808;
  assign n7810 = n5908 & n7395;
  assign n7811 = ~n5920 & ~n7410;
  assign n7812 = n5894 & ~n7811;
  assign n7813 = n5929 & ~n7396;
  assign n7814 = ~n5925 & n7813;
  assign n7815 = n7395 & ~n7814;
  assign n7816 = n5134 & n5902;
  assign n7817 = ~n7396 & ~n7795;
  assign n7818 = n5894 & ~n7817;
  assign n7819 = ~n7816 & ~n7818;
  assign n7820 = ~n5899 & n7819;
  assign n7821 = ~n5907 & n7820;
  assign n7822 = n5133 & ~n7821;
  assign n7823 = ~n7815 & ~n7822;
  assign n7824 = ~n7812 & n7823;
  assign n7825 = ~n7810 & n7824;
  assign n7826 = n7809 & n7825;
  assign n7827 = n7402 & n7826;
  assign n7828 = n7805 & n7827;
  assign n7829 = ~n5893 & n7828;
  assign n7830 = n7829 ^ n5482;
  assign n7831 = n7830 ^ x114;
  assign n7832 = ~n7794 & ~n7831;
  assign n7833 = n7793 & n7832;
  assign n7834 = n7549 ^ x82;
  assign n7835 = n7047 ^ x73;
  assign n7836 = n7834 & n7835;
  assign n7837 = n7833 & n7836;
  assign n7838 = ~n7792 & n7832;
  assign n7839 = ~n7791 & n7838;
  assign n7840 = ~n7834 & ~n7835;
  assign n7841 = n7839 & n7840;
  assign n7842 = ~n7837 & ~n7841;
  assign n7843 = n7793 & n7794;
  assign n7844 = ~n7831 & n7843;
  assign n7845 = ~n7834 & n7835;
  assign n7846 = n7844 & n7845;
  assign n7847 = n7791 & n7792;
  assign n7848 = n7831 & n7847;
  assign n7849 = ~n7794 & n7848;
  assign n7850 = ~n7791 & n7831;
  assign n7851 = ~n7792 & n7850;
  assign n7852 = ~n7794 & n7851;
  assign n7853 = ~n7849 & ~n7852;
  assign n7854 = n7834 & ~n7835;
  assign n7855 = ~n7853 & n7854;
  assign n7856 = ~n7846 & ~n7855;
  assign n7857 = n7794 & n7848;
  assign n7858 = n7845 & n7857;
  assign n7859 = n7840 & n7844;
  assign n7860 = ~n7858 & ~n7859;
  assign n7861 = n7792 & n7850;
  assign n7862 = n7794 & n7861;
  assign n7863 = n7836 & n7862;
  assign n7864 = ~n7792 & n7794;
  assign n7865 = n7850 & n7864;
  assign n7866 = n7845 & n7865;
  assign n7867 = ~n7863 & ~n7866;
  assign n7868 = n7791 & ~n7792;
  assign n7869 = n7832 & n7868;
  assign n7870 = n7832 & n7847;
  assign n7871 = ~n7869 & ~n7870;
  assign n7872 = n7854 & ~n7871;
  assign n7873 = ~n7791 & n7864;
  assign n7874 = ~n7831 & n7873;
  assign n7875 = n7854 & n7874;
  assign n7876 = n7845 & ~n7853;
  assign n7877 = ~n7875 & ~n7876;
  assign n7878 = n7845 & n7870;
  assign n7879 = ~n7831 & n7847;
  assign n7880 = n7794 & n7879;
  assign n7881 = n7791 & n7864;
  assign n7882 = n7831 & n7881;
  assign n7883 = ~n7862 & ~n7882;
  assign n7884 = ~n7880 & n7883;
  assign n7885 = n7884 ^ n7839;
  assign n7886 = n7885 ^ n7839;
  assign n7887 = n7839 ^ n7834;
  assign n7888 = n7887 ^ n7839;
  assign n7889 = ~n7886 & n7888;
  assign n7890 = n7889 ^ n7839;
  assign n7891 = ~n7835 & n7890;
  assign n7892 = n7891 ^ n7839;
  assign n7893 = ~n7878 & ~n7892;
  assign n7894 = n7877 & n7893;
  assign n7895 = ~n7872 & n7894;
  assign n7896 = ~n7831 & n7881;
  assign n7897 = n7845 & n7896;
  assign n7898 = ~n7836 & ~n7840;
  assign n7899 = ~n7794 & n7861;
  assign n7900 = ~n7865 & ~n7880;
  assign n7901 = ~n7882 & n7900;
  assign n7902 = ~n7794 & n7868;
  assign n7903 = n7831 & n7902;
  assign n7904 = ~n7833 & ~n7903;
  assign n7905 = ~n7836 & n7904;
  assign n7906 = ~n7840 & ~n7869;
  assign n7907 = ~n7905 & ~n7906;
  assign n7908 = n7901 & ~n7907;
  assign n7909 = ~n7899 & n7908;
  assign n7910 = ~n7898 & ~n7909;
  assign n7911 = ~n7897 & ~n7910;
  assign n7912 = n7895 & n7911;
  assign n7913 = n7867 & n7912;
  assign n7914 = n7860 & n7913;
  assign n7915 = n7856 & n7914;
  assign n7916 = n7842 & n7915;
  assign n7917 = n7916 ^ n6036;
  assign n7918 = n7917 ^ x90;
  assign n7919 = n7188 & n7191;
  assign n7920 = n7194 & ~n7212;
  assign n7921 = ~n7919 & ~n7920;
  assign n7929 = n7187 & n7203;
  assign n7930 = ~n7210 & ~n7220;
  assign n7931 = ~n7175 & n7930;
  assign n7932 = n7194 & ~n7931;
  assign n7933 = ~n7929 & ~n7932;
  assign n7934 = n7090 & n7196;
  assign n7936 = n7205 & n7935;
  assign n7937 = n7091 & ~n7936;
  assign n7938 = n7185 & ~n7187;
  assign n7939 = ~n7142 & n7177;
  assign n7940 = ~n7184 & ~n7939;
  assign n7941 = ~n7201 & n7940;
  assign n7942 = ~n7188 & n7941;
  assign n7943 = ~n7938 & ~n7942;
  assign n7944 = n7218 & ~n7943;
  assign n7945 = ~n7189 & ~n7944;
  assign n7946 = ~n7937 & ~n7945;
  assign n7947 = ~n7934 & n7946;
  assign n7948 = n7933 & n7947;
  assign n7949 = n7928 & n7948;
  assign n7950 = n7921 & n7949;
  assign n7951 = n7950 ^ n4356;
  assign n7952 = n7951 ^ x109;
  assign n7954 = ~n7754 & ~n7764;
  assign n7955 = ~n7777 & ~n7954;
  assign n7957 = n7676 & ~n7956;
  assign n7958 = ~n7955 & ~n7957;
  assign n7959 = n7723 ^ n7695;
  assign n7960 = n7723 ^ n7720;
  assign n7961 = n7960 ^ n7720;
  assign n7962 = n7722 ^ n7720;
  assign n7963 = n7962 ^ n7720;
  assign n7964 = ~n7961 & n7963;
  assign n7965 = n7964 ^ n7720;
  assign n7966 = ~n7959 & ~n7965;
  assign n7967 = n7732 & n7966;
  assign n7968 = ~n7735 & ~n7755;
  assign n7969 = ~n7746 & n7767;
  assign n7970 = ~n7741 & n7969;
  assign n7972 = ~n7758 & n7971;
  assign n7973 = ~n7727 & n7972;
  assign n7974 = ~n7970 & ~n7973;
  assign n7975 = n7968 & ~n7974;
  assign n7976 = ~n7730 & n7975;
  assign n7977 = ~n7752 & ~n7976;
  assign n7978 = ~n7967 & ~n7977;
  assign n7979 = n7753 ^ n7737;
  assign n7980 = n7979 ^ n7753;
  assign n7981 = n7753 ^ n7675;
  assign n7982 = n7981 ^ n7753;
  assign n7983 = n7980 & ~n7982;
  assign n7984 = n7983 ^ n7753;
  assign n7985 = n7674 & n7984;
  assign n7986 = n7985 ^ n7753;
  assign n7987 = n7978 & ~n7986;
  assign n7988 = n7958 & n7987;
  assign n7989 = ~n7785 & n7988;
  assign n7990 = ~n7726 & n7989;
  assign n7991 = ~n7953 & n7990;
  assign n7992 = n7991 ^ n5178;
  assign n7993 = n7992 ^ x91;
  assign n7994 = ~n7952 & ~n7993;
  assign n8004 = n6423 & ~n8003;
  assign n8012 = n6386 & ~n8011;
  assign n8013 = ~n8004 & ~n8012;
  assign n8027 = ~n6283 & ~n8026;
  assign n8028 = n8013 & ~n8027;
  assign n8029 = n8028 ^ n3264;
  assign n8030 = n8029 ^ x110;
  assign n8031 = n6700 & n7337;
  assign n8032 = ~n6832 & n6869;
  assign n8033 = n6828 & ~n8032;
  assign n8034 = ~n8031 & ~n8033;
  assign n8035 = n6699 & n6851;
  assign n8037 = n6870 & n8036;
  assign n8038 = n6844 & ~n8037;
  assign n8040 = n6854 & n8039;
  assign n8041 = n6844 & ~n8040;
  assign n8042 = ~n6850 & n6863;
  assign n8043 = n6846 & ~n8042;
  assign n8044 = ~n8041 & ~n8043;
  assign n8045 = ~n6846 & ~n6853;
  assign n8046 = ~n6861 & n7330;
  assign n8047 = ~n8045 & ~n8046;
  assign n8048 = n7326 & ~n8047;
  assign n8049 = n8048 ^ n6659;
  assign n8050 = n8049 ^ n8048;
  assign n8051 = n8048 ^ n6870;
  assign n8052 = n8051 ^ n8048;
  assign n8053 = n8050 & ~n8052;
  assign n8054 = n8053 ^ n8048;
  assign n8055 = ~n6699 & ~n8054;
  assign n8056 = n8055 ^ n8048;
  assign n8057 = n8044 & n8056;
  assign n8058 = ~n7322 & n8057;
  assign n8059 = n6830 & n8058;
  assign n8060 = ~n8038 & n8059;
  assign n8061 = ~n8035 & n8060;
  assign n8062 = n8034 & n8061;
  assign n8063 = n6840 & n8062;
  assign n8064 = n8063 ^ n5243;
  assign n8065 = n8064 ^ x77;
  assign n8066 = n8030 & n8065;
  assign n8067 = ~n7501 & n7506;
  assign n8068 = ~n7505 & ~n7525;
  assign n8069 = n7526 & n8068;
  assign n8070 = ~n7507 & n8069;
  assign n8071 = n7424 & ~n8070;
  assign n8072 = ~n7505 & n7536;
  assign n8073 = n7495 & n7540;
  assign n8074 = n8072 & n8073;
  assign n8075 = ~n7507 & n8074;
  assign n8076 = n7512 & ~n8075;
  assign n8077 = ~n7494 & ~n7508;
  assign n8078 = ~n7493 & n8077;
  assign n8079 = ~n7514 & n8078;
  assign n8080 = n7506 & ~n8079;
  assign n8081 = ~n7481 & ~n7488;
  assign n8082 = ~n7493 & ~n7513;
  assign n8083 = ~n7499 & n8082;
  assign n8084 = ~n7524 & n8083;
  assign n8085 = n7515 & n8084;
  assign n8086 = n8081 & n8085;
  assign n8087 = n7487 & ~n8086;
  assign n8088 = ~n8080 & ~n8087;
  assign n8089 = ~n8076 & n8088;
  assign n8090 = ~n8071 & n8089;
  assign n8091 = ~n8067 & n8090;
  assign n8092 = ~n7486 & n8091;
  assign n8093 = n7514 ^ n7423;
  assign n8094 = n8093 ^ n7514;
  assign n8095 = n7524 ^ n7514;
  assign n8096 = n8094 & n8095;
  assign n8097 = n8096 ^ n7514;
  assign n8098 = n7422 & n8097;
  assign n8099 = n8092 & ~n8098;
  assign n8100 = n8099 ^ n5286;
  assign n8101 = n8100 ^ x70;
  assign n8105 = ~n6978 & n7580;
  assign n8106 = n6998 & ~n8105;
  assign n8107 = ~n6993 & ~n7022;
  assign n8108 = n6895 & ~n8107;
  assign n8109 = ~n8106 & ~n8108;
  assign n8110 = n6893 & n7010;
  assign n8111 = ~n7000 & n7007;
  assign n8112 = n6984 & ~n8111;
  assign n8113 = ~n6986 & ~n7005;
  assign n8114 = n6895 & ~n8113;
  assign n8115 = n7023 & n7569;
  assign n8116 = n6998 & ~n8115;
  assign n8117 = ~n8114 & ~n8116;
  assign n8118 = n6894 ^ n6893;
  assign n8119 = ~n6990 & ~n7011;
  assign n8120 = n8119 ^ n6894;
  assign n8121 = n8120 ^ n8119;
  assign n8122 = ~n7005 & ~n7021;
  assign n8123 = n8122 ^ n8119;
  assign n8124 = ~n8121 & n8123;
  assign n8125 = n8124 ^ n8119;
  assign n8126 = ~n8118 & ~n8125;
  assign n8127 = n7576 & ~n8126;
  assign n8128 = n6999 & ~n8127;
  assign n8129 = n8117 & ~n8128;
  assign n8130 = ~n7568 & n8129;
  assign n8131 = ~n8112 & n8130;
  assign n8132 = ~n8110 & n8131;
  assign n8133 = n8109 & n8132;
  assign n8134 = n8104 & n8133;
  assign n8135 = n6983 & n8134;
  assign n8136 = n8135 ^ n5206;
  assign n8137 = n8136 ^ x92;
  assign n8138 = ~n8101 & n8137;
  assign n8139 = n8066 & n8138;
  assign n8140 = n7994 & n8139;
  assign n8141 = n7952 & n7993;
  assign n8142 = n8139 & n8141;
  assign n8143 = n8030 & ~n8065;
  assign n8144 = n8101 & ~n8137;
  assign n8145 = n8143 & n8144;
  assign n8146 = n7994 & n8145;
  assign n8147 = ~n8142 & ~n8146;
  assign n8148 = ~n8030 & n8065;
  assign n8149 = n8138 & n8148;
  assign n8150 = ~n8101 & ~n8137;
  assign n8151 = n8143 & n8150;
  assign n8152 = ~n8149 & ~n8151;
  assign n8153 = n8141 & ~n8152;
  assign n8154 = ~n7952 & n7993;
  assign n8155 = n8144 & n8148;
  assign n8156 = ~n8145 & ~n8155;
  assign n8157 = n8154 & ~n8156;
  assign n8158 = ~n8153 & ~n8157;
  assign n8159 = n8101 & n8137;
  assign n8160 = n8148 & n8159;
  assign n8161 = ~n7952 & n8160;
  assign n8162 = n7952 & ~n7993;
  assign n8163 = ~n8030 & ~n8065;
  assign n8164 = n8150 & n8163;
  assign n8165 = n8159 & n8163;
  assign n8166 = n8066 & n8159;
  assign n8167 = ~n8165 & ~n8166;
  assign n8168 = ~n8155 & n8167;
  assign n8169 = ~n8164 & n8168;
  assign n8170 = n8162 & ~n8169;
  assign n8171 = ~n8161 & ~n8170;
  assign n8172 = n8158 & n8171;
  assign n8173 = ~n8154 & ~n8162;
  assign n8183 = n8138 & n8163;
  assign n8184 = n8148 & n8150;
  assign n8185 = ~n8183 & ~n8184;
  assign n8186 = n8144 & n8163;
  assign n8187 = n8066 & n8144;
  assign n8188 = ~n8165 & ~n8187;
  assign n8189 = ~n8186 & n8188;
  assign n8190 = n8185 & n8189;
  assign n8174 = n8066 & n8150;
  assign n8175 = n8138 & n8143;
  assign n8176 = ~n8149 & ~n8175;
  assign n8177 = ~n8164 & n8176;
  assign n8178 = ~n8162 & n8177;
  assign n8179 = ~n8139 & ~n8151;
  assign n8180 = ~n8154 & n8179;
  assign n8181 = ~n8178 & ~n8180;
  assign n8182 = ~n8174 & ~n8181;
  assign n8191 = n8190 ^ n8182;
  assign n8192 = n8191 ^ n8190;
  assign n8193 = n8143 & n8159;
  assign n8194 = n8193 ^ n8190;
  assign n8195 = n8194 ^ n8190;
  assign n8196 = n8192 & ~n8195;
  assign n8197 = n8196 ^ n8190;
  assign n8198 = ~n8173 & n8197;
  assign n8199 = n8198 ^ n8190;
  assign n8200 = n8172 & n8199;
  assign n8201 = n8147 & n8200;
  assign n8202 = ~n8140 & n8201;
  assign n8203 = n8202 ^ n6071;
  assign n8204 = n8203 ^ x89;
  assign n8205 = n7918 & n8204;
  assign n8206 = ~n7918 & ~n8204;
  assign n8207 = ~n8205 & ~n8206;
  assign n8208 = ~n7673 & n8207;
  assign n8209 = n6433 ^ x69;
  assign n8244 = n8243 ^ x118;
  assign n8245 = ~n8209 & n8244;
  assign n8246 = n5960 ^ x93;
  assign n8247 = ~n7506 & ~n7512;
  assign n8248 = n7507 & ~n8247;
  assign n8249 = ~n7498 & n8081;
  assign n8250 = ~n7524 & n8249;
  assign n8251 = n7424 & ~n8250;
  assign n8252 = ~n8248 & ~n8251;
  assign n8253 = ~n7513 & n8077;
  assign n8254 = n7506 & ~n8253;
  assign n8255 = ~n7514 & n8082;
  assign n8256 = n7512 & ~n8255;
  assign n8257 = n7485 & ~n7512;
  assign n8258 = n7500 & ~n7506;
  assign n8259 = ~n7524 & n8258;
  assign n8260 = ~n8257 & ~n8259;
  assign n8261 = ~n7496 & ~n8260;
  assign n8262 = ~n8247 & ~n8261;
  assign n8263 = ~n7493 & n8068;
  assign n8264 = n7424 & ~n8263;
  assign n8267 = n7515 & n8068;
  assign n8265 = ~n7535 & n8081;
  assign n8266 = ~n7507 & n8265;
  assign n8268 = n8267 ^ n8266;
  assign n8269 = n8267 ^ n7487;
  assign n8270 = n8267 & n8269;
  assign n8271 = n8270 ^ n8267;
  assign n8272 = n8268 & n8271;
  assign n8273 = n8272 ^ n8270;
  assign n8274 = n8273 ^ n8267;
  assign n8275 = n8274 ^ n7487;
  assign n8276 = ~n8264 & n8275;
  assign n8277 = n8276 ^ n8264;
  assign n8278 = ~n8262 & ~n8277;
  assign n8279 = ~n8098 & n8278;
  assign n8280 = ~n8256 & n8279;
  assign n8281 = ~n8254 & n8280;
  assign n8282 = n8252 & n8281;
  assign n8283 = n8282 ^ n5797;
  assign n8284 = n8283 ^ x100;
  assign n8285 = n8246 & ~n8284;
  assign n8288 = ~n7744 & ~n7746;
  assign n8289 = n7741 & ~n8288;
  assign n8290 = n7737 & ~n7752;
  assign n8291 = n7760 & ~n7766;
  assign n8292 = ~n7725 & n8291;
  assign n8293 = n7674 & ~n8292;
  assign n8294 = ~n8290 & ~n8293;
  assign n8295 = n7756 ^ n7676;
  assign n8296 = n7756 ^ n7732;
  assign n8297 = n8296 ^ n7732;
  assign n8298 = n7753 ^ n7732;
  assign n8299 = n8297 & ~n8298;
  assign n8300 = n8299 ^ n7732;
  assign n8301 = ~n8295 & n8300;
  assign n8302 = n8301 ^ n7676;
  assign n8303 = n8294 & ~n8302;
  assign n8304 = ~n8289 & n8303;
  assign n8305 = ~n7744 & ~n7780;
  assign n8306 = ~n7676 & n8305;
  assign n8307 = n8306 ^ n7727;
  assign n8308 = n8306 ^ n7968;
  assign n8309 = n8308 ^ n7968;
  assign n8310 = n7968 ^ n7767;
  assign n8311 = ~n8309 & ~n8310;
  assign n8312 = n8311 ^ n7968;
  assign n8313 = ~n8307 & n8312;
  assign n8314 = n8313 ^ n7727;
  assign n8315 = n8304 & ~n8314;
  assign n8316 = n8287 & n8315;
  assign n8317 = ~n7726 & n8316;
  assign n8318 = ~n7953 & n8317;
  assign n8319 = ~n7758 & n8318;
  assign n8320 = n8319 ^ n5749;
  assign n8321 = n8320 ^ x86;
  assign n8352 = n8351 ^ x83;
  assign n8353 = n8321 & ~n8352;
  assign n8354 = n8285 & n8353;
  assign n8355 = n8245 & n8354;
  assign n8356 = n8209 & n8244;
  assign n8357 = ~n8246 & n8284;
  assign n8358 = ~n8321 & ~n8352;
  assign n8359 = n8357 & n8358;
  assign n8360 = n8246 & n8284;
  assign n8361 = n8353 & n8360;
  assign n8362 = ~n8359 & ~n8361;
  assign n8363 = n8356 & ~n8362;
  assign n8364 = ~n8355 & ~n8363;
  assign n8365 = n8209 & ~n8244;
  assign n8366 = n8321 & n8352;
  assign n8367 = n8360 & n8366;
  assign n8368 = ~n8321 & n8352;
  assign n8369 = n8285 & n8368;
  assign n8370 = ~n8246 & ~n8284;
  assign n8371 = n8368 & n8370;
  assign n8372 = n8285 & n8366;
  assign n8373 = ~n8371 & ~n8372;
  assign n8374 = ~n8369 & n8373;
  assign n8375 = ~n8367 & n8374;
  assign n8376 = n8365 & ~n8375;
  assign n8377 = n8353 & n8370;
  assign n8378 = n8358 & n8360;
  assign n8379 = ~n8377 & ~n8378;
  assign n8380 = ~n8359 & n8379;
  assign n8381 = n8245 & ~n8380;
  assign n8382 = ~n8376 & ~n8381;
  assign n8383 = ~n8209 & ~n8244;
  assign n8384 = ~n8361 & ~n8377;
  assign n8385 = n8353 & n8357;
  assign n8386 = ~n8378 & ~n8385;
  assign n8387 = n8384 & n8386;
  assign n8388 = n8383 & ~n8387;
  assign n8389 = n8285 & n8358;
  assign n8390 = n8358 & n8370;
  assign n8391 = ~n8389 & ~n8390;
  assign n8392 = n8356 & ~n8391;
  assign n8393 = n8365 & ~n8387;
  assign n8394 = n8357 & n8366;
  assign n8395 = n8360 & n8368;
  assign n8396 = ~n8371 & ~n8395;
  assign n8397 = ~n8394 & n8396;
  assign n8398 = ~n8367 & n8397;
  assign n8399 = n8245 & ~n8398;
  assign n8400 = ~n8356 & ~n8383;
  assign n8401 = n8357 & n8368;
  assign n8402 = n8366 & n8370;
  assign n8403 = ~n8372 & ~n8402;
  assign n8404 = ~n8394 & n8403;
  assign n8405 = n8404 ^ n8374;
  assign n8406 = n8244 ^ n8209;
  assign n8407 = n8374 ^ n8244;
  assign n8408 = n8406 & ~n8407;
  assign n8409 = n8408 ^ n8244;
  assign n8410 = n8405 & ~n8409;
  assign n8411 = n8410 ^ n8404;
  assign n8412 = ~n8401 & n8411;
  assign n8413 = ~n8400 & ~n8412;
  assign n8414 = ~n8399 & ~n8413;
  assign n8415 = ~n8393 & n8414;
  assign n8416 = ~n8392 & n8415;
  assign n8417 = ~n8388 & n8416;
  assign n8418 = n8382 & n8417;
  assign n8419 = n8364 & n8418;
  assign n8420 = n8419 ^ n6113;
  assign n8421 = n8420 ^ x80;
  assign n8422 = n7918 & n8421;
  assign n8423 = ~n8204 & n8422;
  assign n8424 = ~n7673 & n8421;
  assign n8425 = n7918 & n8424;
  assign n8426 = ~n8423 & ~n8425;
  assign n8427 = n7673 & ~n8421;
  assign n8428 = ~n8207 & n8427;
  assign n8429 = n8426 & ~n8428;
  assign n8430 = ~n8208 & n8429;
  assign n8593 = n8592 ^ n8430;
  assign n8594 = n8593 ^ n8430;
  assign n8595 = n8204 & n8421;
  assign n8596 = ~n8204 & n8427;
  assign n8597 = ~n8595 & ~n8596;
  assign n8598 = n7918 & ~n8597;
  assign n8599 = ~n7673 & ~n8421;
  assign n8600 = n8204 & n8599;
  assign n8601 = n7673 & n8204;
  assign n8602 = ~n8206 & ~n8601;
  assign n8603 = n8421 & ~n8602;
  assign n8604 = ~n8600 & ~n8603;
  assign n8605 = ~n8598 & n8604;
  assign n8606 = n8605 ^ n8430;
  assign n8607 = n8594 & n8606;
  assign n8608 = n8607 ^ n8430;
  assign n8609 = ~n7321 & n8608;
  assign n8610 = ~n7918 & n8204;
  assign n8611 = n8610 ^ n8424;
  assign n8612 = n7918 & n8427;
  assign n8613 = ~n8611 & ~n8612;
  assign n8614 = n8613 ^ n8592;
  assign n8615 = n8614 ^ n8613;
  assign n8616 = n8205 & n8424;
  assign n8617 = n7673 & n8422;
  assign n8618 = ~n7918 & n8599;
  assign n8619 = n7673 & ~n8207;
  assign n8620 = ~n8618 & ~n8619;
  assign n8621 = ~n8617 & n8620;
  assign n8622 = ~n8616 & n8621;
  assign n8623 = n8622 ^ n8613;
  assign n8624 = n8615 & n8623;
  assign n8625 = n8624 ^ n8613;
  assign n8626 = n7321 & ~n8625;
  assign n8627 = ~n8609 & ~n8626;
  assign n8628 = n8627 ^ n7566;
  assign n8629 = n8628 ^ x107;
  assign n8630 = n8565 & n8583;
  assign n8631 = n8533 & n8551;
  assign n8632 = ~n8555 & ~n8631;
  assign n8633 = ~n8575 & n8581;
  assign n8634 = n8632 & n8633;
  assign n8635 = n8528 & ~n8634;
  assign n8636 = n8495 ^ n8466;
  assign n8637 = n8467 ^ n8459;
  assign n8638 = n8495 ^ n8467;
  assign n8639 = n8638 ^ n8467;
  assign n8640 = n8637 & n8639;
  assign n8641 = n8640 ^ n8467;
  assign n8642 = ~n8636 & ~n8641;
  assign n8643 = n8642 ^ n8459;
  assign n8644 = n8545 & ~n8643;
  assign n8645 = ~n8635 & ~n8644;
  assign n8646 = ~n8630 & n8645;
  assign n8647 = n8567 ^ n8537;
  assign n8648 = n8576 ^ n8537;
  assign n8649 = n8648 ^ n8576;
  assign n8650 = n8576 ^ n8545;
  assign n8651 = ~n8649 & n8650;
  assign n8652 = n8651 ^ n8576;
  assign n8653 = ~n8647 & ~n8652;
  assign n8654 = n8653 ^ n8567;
  assign n8655 = n8646 & n8654;
  assign n8656 = ~n8542 & n8655;
  assign n8657 = n8539 & n8656;
  assign n8658 = n8657 ^ n7141;
  assign n8659 = n8658 ^ x99;
  assign n8660 = n8383 & ~n8386;
  assign n8661 = ~n8354 & ~n8390;
  assign n8662 = n8245 & ~n8661;
  assign n8663 = ~n8660 & ~n8662;
  assign n8664 = n8356 & ~n8386;
  assign n8665 = n8354 & n8383;
  assign n8666 = n8373 & ~n8394;
  assign n8667 = ~n8367 & n8666;
  assign n8668 = n8383 & ~n8667;
  assign n8669 = ~n8367 & ~n8401;
  assign n8670 = ~n8402 & n8669;
  assign n8671 = n8245 & ~n8670;
  assign n8672 = ~n8369 & ~n8402;
  assign n8673 = ~n8394 & n8672;
  assign n8674 = ~n8367 & n8673;
  assign n8675 = n8356 & ~n8674;
  assign n8676 = ~n8671 & ~n8675;
  assign n8677 = ~n8668 & n8676;
  assign n8678 = n8395 & n8406;
  assign n8679 = n8384 & n8666;
  assign n8680 = ~n8359 & n8679;
  assign n8681 = ~n8354 & n8680;
  assign n8682 = n8365 & ~n8681;
  assign n8683 = ~n8678 & ~n8682;
  assign n8684 = n8677 & n8683;
  assign n8685 = ~n8665 & n8684;
  assign n8686 = ~n8664 & n8685;
  assign n8687 = n8389 ^ n8244;
  assign n8688 = n8389 ^ n8209;
  assign n8689 = n8688 ^ n8209;
  assign n8690 = n8359 ^ n8209;
  assign n8691 = ~n8689 & n8690;
  assign n8692 = n8691 ^ n8209;
  assign n8693 = n8687 & ~n8692;
  assign n8694 = n8693 ^ n8244;
  assign n8695 = n8686 & ~n8694;
  assign n8696 = n8663 & n8695;
  assign n8697 = n8696 ^ n6722;
  assign n8698 = n8697 ^ x106;
  assign n8699 = ~n8659 & n8698;
  assign n8700 = n7194 & n7216;
  assign n8701 = ~n7189 & n7201;
  assign n8702 = ~n8700 & ~n8701;
  assign n8703 = n7200 & ~n7216;
  assign n8704 = ~n7220 & n8703;
  assign n8705 = ~n7203 & n8704;
  assign n8706 = n7188 & ~n8705;
  assign n8707 = ~n7191 & n7204;
  assign n8708 = n7194 & ~n8707;
  assign n8709 = n7221 & n8437;
  assign n8710 = n7187 & ~n8709;
  assign n8711 = ~n8708 & ~n8710;
  assign n8712 = ~n8706 & n8711;
  assign n8713 = ~n7185 & n7187;
  assign n8714 = n7144 ^ n7125;
  assign n8715 = n8714 ^ n7142;
  assign n8716 = n7173 ^ n7142;
  assign n8717 = n8716 ^ n7142;
  assign n8718 = n8716 ^ n7125;
  assign n8719 = n8717 & ~n8718;
  assign n8720 = n8719 ^ n8716;
  assign n8721 = ~n8715 & ~n8720;
  assign n8722 = n8721 ^ n8716;
  assign n8723 = n7091 & ~n8722;
  assign n8724 = ~n8713 & ~n8723;
  assign n8725 = n8712 & n8724;
  assign n8726 = n8702 & n8725;
  assign n8727 = n7181 & n8726;
  assign n8728 = n7921 & n8727;
  assign n8729 = n8728 ^ n5588;
  assign n8730 = n8729 ^ x96;
  assign n8731 = n7357 ^ x106;
  assign n8732 = ~n8730 & n8731;
  assign n8733 = n8730 & ~n8731;
  assign n8734 = ~n8732 & ~n8733;
  assign n8735 = ~n6561 & n6566;
  assign n8736 = n6571 & ~n7364;
  assign n8737 = ~n8735 & ~n8736;
  assign n8738 = n6576 & n6605;
  assign n8739 = n6578 & ~n8738;
  assign n8740 = ~n6590 & n6598;
  assign n8741 = ~n6589 & n8740;
  assign n8742 = n6578 & ~n8741;
  assign n8743 = n6515 ^ n6479;
  assign n8744 = n8743 ^ n6469;
  assign n8745 = ~n6435 & ~n8744;
  assign n8746 = n6571 & n8745;
  assign n8747 = ~n8742 & ~n8746;
  assign n8748 = n7371 & n7377;
  assign n8749 = ~n6591 & n8748;
  assign n8750 = n8749 ^ n6562;
  assign n8751 = n8749 ^ n6611;
  assign n8752 = n8751 ^ n6611;
  assign n8753 = n6611 ^ n6585;
  assign n8754 = ~n8752 & n8753;
  assign n8755 = n8754 ^ n6611;
  assign n8756 = ~n8750 & n8755;
  assign n8757 = n8756 ^ n6562;
  assign n8758 = n8747 & ~n8757;
  assign n8759 = ~n8739 & n8758;
  assign n8760 = n8737 & n8759;
  assign n8761 = ~n8470 & n8760;
  assign n8762 = ~n6595 & n8761;
  assign n8763 = n8762 ^ n5624;
  assign n8764 = n8763 ^ x105;
  assign n8765 = n7992 ^ x123;
  assign n8766 = ~n8764 & n8765;
  assign n8767 = ~n8734 & n8766;
  assign n8768 = n7420 ^ x99;
  assign n8769 = n8100 ^ x81;
  assign n8770 = n8768 & n8769;
  assign n8771 = n8765 ^ n8731;
  assign n8772 = n8765 ^ n8764;
  assign n8773 = n8772 ^ n8764;
  assign n8774 = n8731 ^ n8730;
  assign n8775 = n8774 ^ n8764;
  assign n8776 = n8775 ^ n8764;
  assign n8777 = n8776 ^ n8764;
  assign n8778 = n8773 & n8777;
  assign n8779 = n8778 ^ n8764;
  assign n8780 = ~n8771 & ~n8779;
  assign n8781 = n8780 ^ n8775;
  assign n8782 = n8770 & n8781;
  assign n8783 = ~n8768 & ~n8769;
  assign n8784 = n8764 & n8765;
  assign n8785 = ~n8730 & n8784;
  assign n8786 = n8730 & n8731;
  assign n8787 = ~n8765 & n8786;
  assign n8788 = ~n8764 & ~n8765;
  assign n8789 = ~n8731 & n8788;
  assign n8790 = ~n8787 & ~n8789;
  assign n8791 = ~n8785 & n8790;
  assign n8792 = n8783 & ~n8791;
  assign n8793 = ~n8782 & ~n8792;
  assign n8794 = n8768 & ~n8769;
  assign n8795 = n8764 & ~n8765;
  assign n8796 = ~n8730 & n8795;
  assign n8797 = n8788 ^ n8730;
  assign n8798 = n8797 ^ n8788;
  assign n8799 = n8788 ^ n8764;
  assign n8800 = n8799 ^ n8788;
  assign n8801 = n8798 & n8800;
  assign n8802 = n8801 ^ n8788;
  assign n8803 = ~n8731 & n8802;
  assign n8804 = n8803 ^ n8788;
  assign n8805 = ~n8796 & ~n8804;
  assign n8806 = n8794 & ~n8805;
  assign n8807 = ~n8768 & n8769;
  assign n8808 = ~n8730 & ~n8731;
  assign n8809 = ~n8765 & n8808;
  assign n8810 = ~n8786 & n8788;
  assign n8811 = ~n8809 & ~n8810;
  assign n8812 = ~n8731 & n8784;
  assign n8813 = ~n8766 & ~n8795;
  assign n8814 = n8786 & ~n8813;
  assign n8815 = ~n8812 & ~n8814;
  assign n8816 = n8811 & n8815;
  assign n8817 = n8807 & n8816;
  assign n8818 = ~n8806 & ~n8817;
  assign n8819 = n8793 & n8818;
  assign n8820 = ~n8767 & n8819;
  assign n8821 = n8820 ^ n7088;
  assign n8822 = n8821 ^ x104;
  assign n8823 = n8029 ^ x85;
  assign n8824 = n8494 ^ x102;
  assign n8825 = n8823 & n8824;
  assign n8826 = n5915 & n5925;
  assign n8827 = ~n5133 & n5902;
  assign n8828 = ~n8826 & ~n8827;
  assign n8829 = n5134 & n5946;
  assign n8830 = ~n5945 & ~n7795;
  assign n8831 = ~n5908 & n8830;
  assign n8832 = n5894 & ~n8831;
  assign n8833 = ~n8829 & ~n8832;
  assign n8834 = n8828 & n8833;
  assign n8835 = n5899 & n7395;
  assign n8836 = ~n5916 & n7406;
  assign n8837 = n5905 & ~n8836;
  assign n8838 = ~n5907 & n5917;
  assign n8839 = ~n7396 & n8838;
  assign n8840 = n5134 & ~n8839;
  assign n8841 = n5930 & ~n7410;
  assign n8842 = n7395 & ~n8841;
  assign n8843 = ~n8840 & ~n8842;
  assign n8844 = ~n8837 & n8843;
  assign n8845 = ~n8835 & n8844;
  assign n8846 = n8834 & n8845;
  assign n8847 = n5911 & n8846;
  assign n8848 = n7805 & n8847;
  assign n8849 = n7400 & n8848;
  assign n8850 = ~n5893 & n8849;
  assign n8851 = n8850 ^ n4538;
  assign n8852 = n8851 ^ x78;
  assign n8853 = n8525 ^ x124;
  assign n8854 = n8852 & ~n8853;
  assign n8855 = n7951 ^ x68;
  assign n8856 = ~n7507 & n8082;
  assign n8857 = n7506 & ~n8856;
  assign n8858 = ~n7508 & n8084;
  assign n8859 = n7424 & ~n8858;
  assign n8860 = ~n8857 & ~n8859;
  assign n8861 = ~n7514 & n8263;
  assign n8862 = n7512 & ~n8861;
  assign n8863 = n8072 & n8253;
  assign n8864 = n7487 & ~n8863;
  assign n8865 = ~n7488 & ~n7496;
  assign n8866 = ~n7482 & n8865;
  assign n8867 = ~n7512 & n8866;
  assign n8868 = n8081 & n8258;
  assign n8869 = n7501 & n8265;
  assign n8870 = ~n8868 & ~n8869;
  assign n8871 = ~n8867 & n8870;
  assign n8872 = ~n8247 & n8871;
  assign n8873 = ~n8864 & ~n8872;
  assign n8874 = ~n8862 & n8873;
  assign n8875 = n8860 & n8874;
  assign n8876 = ~n7490 & n8875;
  assign n8877 = ~n7486 & n8876;
  assign n8878 = ~n8098 & n8877;
  assign n8879 = n8878 ^ n4146;
  assign n8880 = n8879 ^ x126;
  assign n8881 = ~n8855 & n8880;
  assign n8882 = n8854 & n8881;
  assign n8883 = n8852 & n8853;
  assign n8884 = ~n8855 & ~n8880;
  assign n8885 = n8883 & n8884;
  assign n8886 = ~n8882 & ~n8885;
  assign n8887 = n8825 & ~n8886;
  assign n8888 = n8855 & n8880;
  assign n8889 = n8883 & n8888;
  assign n8890 = n8825 & n8889;
  assign n8891 = ~n8823 & n8824;
  assign n8892 = ~n8852 & n8853;
  assign n8893 = n8881 & n8892;
  assign n8894 = ~n8852 & ~n8853;
  assign n8895 = n8884 & n8894;
  assign n8896 = ~n8893 & ~n8895;
  assign n8897 = n8891 & ~n8896;
  assign n8898 = ~n8890 & ~n8897;
  assign n8899 = n8823 & ~n8824;
  assign n8900 = n8855 & ~n8880;
  assign n8901 = n8894 & n8900;
  assign n8902 = n8899 & n8901;
  assign n8903 = ~n8823 & ~n8824;
  assign n8904 = n8888 & n8894;
  assign n8905 = n8892 & n8900;
  assign n8906 = ~n8904 & ~n8905;
  assign n8907 = n8903 & ~n8906;
  assign n8908 = ~n8902 & ~n8907;
  assign n8909 = n8824 ^ n8823;
  assign n8910 = n8854 & n8888;
  assign n8911 = ~n8909 & n8910;
  assign n8912 = n8881 & n8883;
  assign n8913 = ~n8882 & ~n8912;
  assign n8914 = n8891 & ~n8913;
  assign n8915 = ~n8911 & ~n8914;
  assign n8916 = n8854 & n8884;
  assign n8917 = n8884 & n8892;
  assign n8918 = ~n8916 & ~n8917;
  assign n8919 = ~n8901 & n8918;
  assign n8920 = ~n8905 & n8919;
  assign n8921 = n8825 & ~n8920;
  assign n8922 = n8855 ^ n8853;
  assign n8923 = n8922 ^ n8880;
  assign n8924 = n8880 ^ n8855;
  assign n8925 = n8855 ^ n8852;
  assign n8926 = n8925 ^ n8855;
  assign n8927 = n8924 & n8926;
  assign n8928 = n8927 ^ n8855;
  assign n8929 = n8923 & ~n8928;
  assign n8930 = ~n8889 & ~n8929;
  assign n8931 = n8903 & ~n8930;
  assign n8932 = ~n8921 & ~n8931;
  assign n8933 = n8883 & n8900;
  assign n8934 = n8888 & n8892;
  assign n8935 = ~n8910 & ~n8934;
  assign n8936 = ~n8933 & n8935;
  assign n8937 = n8899 & ~n8936;
  assign n8938 = n8854 & n8900;
  assign n8939 = ~n8901 & ~n8933;
  assign n8940 = ~n8938 & n8939;
  assign n8941 = ~n8899 & n8940;
  assign n8942 = ~n8904 & n8941;
  assign n8943 = n8896 & ~n8912;
  assign n8944 = ~n8938 & n8943;
  assign n8945 = n8899 & ~n8944;
  assign n8946 = ~n8891 & ~n8945;
  assign n8947 = ~n8942 & ~n8946;
  assign n8948 = ~n8937 & ~n8947;
  assign n8949 = n8932 & n8948;
  assign n8950 = n8915 & n8949;
  assign n8951 = n8908 & n8950;
  assign n8952 = n8898 & n8951;
  assign n8953 = ~n8887 & n8952;
  assign n8954 = n8953 ^ n6698;
  assign n8955 = n8954 ^ x73;
  assign n8956 = ~n8822 & n8955;
  assign n8957 = n7833 & n7854;
  assign n8958 = n7845 & ~n7883;
  assign n8959 = ~n8957 & ~n8958;
  assign n8960 = n7845 & n7880;
  assign n8961 = ~n7870 & ~n7903;
  assign n8962 = ~n7857 & n8961;
  assign n8963 = n7854 & ~n8962;
  assign n8964 = ~n8960 & ~n8963;
  assign n8965 = n7836 & n7874;
  assign n8966 = ~n7865 & ~n7896;
  assign n8967 = ~n7862 & n8966;
  assign n8968 = ~n7898 & ~n8967;
  assign n8969 = n7854 & ~n7901;
  assign n8970 = ~n7833 & ~n7839;
  assign n8971 = n7845 & ~n8970;
  assign n8972 = ~n8969 & ~n8971;
  assign n8973 = n7877 & n8972;
  assign n8974 = ~n7849 & n7906;
  assign n8975 = ~n7903 & n8974;
  assign n8976 = ~n8962 & ~n8975;
  assign n8977 = n8976 ^ n7836;
  assign n8978 = ~n7849 & ~n7869;
  assign n8979 = n8978 ^ n8976;
  assign n8980 = n8979 ^ n8978;
  assign n8981 = n8978 ^ n7840;
  assign n8982 = n8980 & n8981;
  assign n8983 = n8982 ^ n8978;
  assign n8984 = n8977 & n8983;
  assign n8985 = n8984 ^ n7836;
  assign n8986 = n8973 & ~n8985;
  assign n8987 = n7842 & n8986;
  assign n8988 = ~n8968 & n8987;
  assign n8989 = ~n8965 & n8988;
  assign n8990 = n8964 & n8989;
  assign n8991 = n7860 & n8990;
  assign n8992 = n8959 & n8991;
  assign n8993 = n8992 ^ n7478;
  assign n8994 = n8993 ^ x123;
  assign n8995 = n8956 & n8994;
  assign n8996 = n8162 & n8183;
  assign n8997 = ~n8140 & ~n8996;
  assign n8998 = n8154 & n8160;
  assign n8999 = n8141 & n8175;
  assign n9000 = ~n8998 & ~n8999;
  assign n9001 = n7994 & n8193;
  assign n9002 = n8141 & n8184;
  assign n9003 = ~n9001 & ~n9002;
  assign n9004 = n8141 & n8174;
  assign n9005 = n7994 & ~n8167;
  assign n9006 = ~n9004 & ~n9005;
  assign n9007 = ~n8173 & n8187;
  assign n9008 = n8152 & ~n8174;
  assign n9009 = ~n8193 & n9008;
  assign n9010 = n8156 & n9009;
  assign n9011 = n8162 & ~n9010;
  assign n9012 = ~n9007 & ~n9011;
  assign n9013 = ~n8145 & ~n8186;
  assign n9014 = n8154 & ~n9013;
  assign n9015 = n7994 & n8164;
  assign n9016 = n8152 & ~n8193;
  assign n9017 = ~n8151 & ~n8164;
  assign n9018 = ~n8154 & n9017;
  assign n9019 = ~n9016 & ~n9018;
  assign n9020 = ~n9015 & ~n9019;
  assign n9021 = ~n8184 & n9020;
  assign n9022 = n9021 ^ n7993;
  assign n9023 = n9022 ^ n9021;
  assign n9024 = ~n8160 & n8167;
  assign n9025 = ~n8186 & n9024;
  assign n9026 = n9025 ^ n9021;
  assign n9027 = n9026 ^ n9021;
  assign n9028 = n9023 & ~n9027;
  assign n9029 = n9028 ^ n9021;
  assign n9030 = n7952 & ~n9029;
  assign n9031 = n9030 ^ n9021;
  assign n9032 = ~n9014 & n9031;
  assign n9033 = n9012 & n9032;
  assign n9034 = n9006 & n9033;
  assign n9035 = n9003 & n9034;
  assign n9036 = n8147 & n9035;
  assign n9037 = n9000 & n9036;
  assign n9038 = n8997 & n9037;
  assign n9039 = n9038 ^ n7454;
  assign n9040 = n9039 ^ x113;
  assign n9041 = n8995 & n9040;
  assign n9042 = n8699 & n9041;
  assign n9043 = n8659 & ~n8698;
  assign n9044 = n8822 & n8994;
  assign n9045 = n8955 & n9044;
  assign n9046 = n9040 & n9045;
  assign n9047 = n9043 & n9046;
  assign n9048 = ~n8955 & ~n9040;
  assign n9049 = ~n8822 & n9048;
  assign n9050 = ~n8994 & n9049;
  assign n9051 = n8699 & n9050;
  assign n9052 = ~n9047 & ~n9051;
  assign n9053 = ~n9042 & n9052;
  assign n9054 = ~n9040 & n9045;
  assign n9055 = n8699 & n9054;
  assign n9056 = n9043 & n9050;
  assign n9057 = ~n9055 & ~n9056;
  assign n9058 = n8659 & n8698;
  assign n9059 = ~n8659 & ~n8698;
  assign n9060 = ~n9058 & ~n9059;
  assign n9061 = ~n8994 & n9040;
  assign n9062 = n8956 & n9061;
  assign n9063 = n8994 & n9049;
  assign n9064 = ~n9062 & ~n9063;
  assign n9065 = ~n9060 & ~n9064;
  assign n9066 = ~n8955 & n9044;
  assign n9067 = n9040 & n9066;
  assign n9068 = ~n9058 & ~n9067;
  assign n9069 = n8822 & n9061;
  assign n9070 = ~n8955 & n9069;
  assign n9071 = n8822 & n9048;
  assign n9072 = ~n8994 & n9071;
  assign n9073 = ~n9054 & ~n9072;
  assign n9074 = ~n9067 & n9073;
  assign n9075 = ~n9070 & n9074;
  assign n9076 = ~n9068 & ~n9075;
  assign n9077 = ~n9065 & ~n9076;
  assign n9078 = n8956 & ~n8994;
  assign n9079 = ~n9040 & n9078;
  assign n9080 = ~n9072 & ~n9079;
  assign n9081 = n9044 & n9048;
  assign n9082 = ~n9046 & ~n9081;
  assign n9083 = ~n9070 & n9082;
  assign n9084 = n9080 & n9083;
  assign n9085 = n9059 & ~n9084;
  assign n9086 = n9041 & n9058;
  assign n9087 = ~n8822 & ~n8955;
  assign n9088 = n8994 & n9087;
  assign n9089 = n9040 & n9088;
  assign n9090 = n8659 & n9089;
  assign n9091 = ~n9086 & ~n9090;
  assign n9092 = n8822 & n8955;
  assign n9093 = ~n8994 & n9092;
  assign n9094 = ~n9040 & n9093;
  assign n9095 = n8995 & ~n9040;
  assign n9096 = n9061 & n9087;
  assign n9097 = ~n9062 & ~n9096;
  assign n9098 = ~n9095 & n9097;
  assign n9099 = ~n9094 & n9098;
  assign n9100 = n8699 & ~n9099;
  assign n9101 = n9061 & n9092;
  assign n9102 = ~n9081 & ~n9101;
  assign n9103 = ~n9095 & n9102;
  assign n9104 = ~n9079 & n9103;
  assign n9105 = n9043 & ~n9104;
  assign n9106 = ~n9100 & ~n9105;
  assign n9107 = n9091 & n9106;
  assign n9108 = ~n9085 & n9107;
  assign n9109 = n9077 & n9108;
  assign n9110 = n9057 & n9109;
  assign n9111 = n9053 & n9110;
  assign n9112 = n9111 ^ n7549;
  assign n9113 = n9112 ^ x80;
  assign n9114 = n8629 & n9113;
  assign n9115 = n7606 & n7620;
  assign n9116 = ~n7608 & ~n7618;
  assign n9117 = n7394 & ~n9116;
  assign n9118 = ~n9115 & ~n9117;
  assign n9119 = ~n7611 & ~n7617;
  assign n9120 = ~n7358 & ~n9119;
  assign n9121 = ~n7603 & ~n7610;
  assign n9122 = n7616 & ~n9121;
  assign n9123 = ~n7628 & ~n7647;
  assign n9124 = n7616 & ~n9123;
  assign n9125 = ~n7635 & ~n7645;
  assign n9126 = n7567 ^ n7421;
  assign n9127 = n9126 ^ n7598;
  assign n9128 = n7550 & ~n9127;
  assign n9129 = ~n7633 & n9128;
  assign n9130 = ~n7617 & ~n7662;
  assign n9131 = ~n7600 & ~n7610;
  assign n9132 = n9130 & n9131;
  assign n9133 = n7621 & n9132;
  assign n9134 = n7651 & ~n9133;
  assign n9135 = ~n9129 & ~n9134;
  assign n9136 = ~n9125 & n9135;
  assign n9137 = ~n9124 & n9136;
  assign n9138 = ~n9122 & n9137;
  assign n9139 = ~n9120 & n9138;
  assign n9140 = n9118 & n9139;
  assign n9141 = ~n7670 & n9140;
  assign n9142 = n9141 ^ n5132;
  assign n9143 = n9142 ^ x118;
  assign n9144 = n8891 & n8916;
  assign n9145 = n8903 & ~n8935;
  assign n9146 = ~n9144 & ~n9145;
  assign n9147 = n8903 & n8917;
  assign n9148 = n8899 ^ n8893;
  assign n9149 = n8893 ^ n8825;
  assign n9150 = n9149 ^ n8825;
  assign n9151 = n8895 ^ n8825;
  assign n9152 = ~n9150 & ~n9151;
  assign n9153 = n9152 ^ n8825;
  assign n9154 = n9148 & n9153;
  assign n9155 = n9154 ^ n8899;
  assign n9156 = ~n9147 & ~n9155;
  assign n9157 = n8895 & ~n8909;
  assign n9158 = n8881 & n8894;
  assign n9159 = n8906 & ~n9158;
  assign n9160 = n8891 & ~n9159;
  assign n9161 = ~n9157 & ~n9160;
  assign n9162 = n8899 & ~n8919;
  assign n9163 = n8886 & ~n8893;
  assign n9164 = ~n8938 & n9163;
  assign n9165 = n8903 & ~n9164;
  assign n9166 = ~n8912 & ~n8933;
  assign n9167 = ~n8934 & n9166;
  assign n9168 = ~n8901 & n9167;
  assign n9169 = n8891 & ~n9168;
  assign n9170 = ~n8889 & ~n8904;
  assign n9171 = ~n8825 & n9170;
  assign n9172 = ~n8933 & n9171;
  assign n9173 = n8906 & ~n8938;
  assign n9174 = ~n8910 & n9173;
  assign n9175 = n8825 & ~n9174;
  assign n9176 = ~n8899 & ~n9175;
  assign n9177 = ~n9172 & ~n9176;
  assign n9178 = ~n9169 & ~n9177;
  assign n9179 = ~n9165 & n9178;
  assign n9180 = ~n9162 & n9179;
  assign n9181 = n9161 & n9180;
  assign n9182 = n9156 & n9181;
  assign n9183 = n9146 & n9182;
  assign n9184 = ~n8887 & n9183;
  assign n9185 = n9184 ^ n4619;
  assign n9186 = n9185 ^ x109;
  assign n9187 = n9143 & n9186;
  assign n9188 = n8245 & ~n8373;
  assign n9189 = n8383 & ~n8669;
  assign n9190 = ~n8385 & ~n8389;
  assign n9191 = n8365 & ~n9190;
  assign n9192 = ~n9189 & ~n9191;
  assign n9193 = ~n9188 & n9192;
  assign n9194 = n8362 & n8673;
  assign n9195 = ~n8372 & n9194;
  assign n9196 = n8365 & ~n9195;
  assign n9197 = n8386 & n8669;
  assign n9198 = ~n8389 & n9197;
  assign n9199 = n8245 & ~n9198;
  assign n9200 = ~n9196 & ~n9199;
  assign n9201 = ~n8379 & ~n8400;
  assign n9202 = ~n8369 & n8666;
  assign n9203 = n8356 & ~n9202;
  assign n9204 = n8396 & n8661;
  assign n9205 = n8383 & ~n9204;
  assign n9206 = ~n9203 & ~n9205;
  assign n9207 = ~n9201 & n9206;
  assign n9208 = n9200 & n9207;
  assign n9209 = n9193 & n9208;
  assign n9210 = n8364 & n9209;
  assign n9211 = n9210 ^ n5889;
  assign n9212 = n9211 ^ x85;
  assign n9213 = n7836 & n7839;
  assign n9214 = n7840 & n7870;
  assign n9215 = ~n9213 & ~n9214;
  assign n9216 = ~n7835 & ~n7900;
  assign n9217 = ~n7869 & ~n7899;
  assign n9218 = ~n7849 & n9217;
  assign n9219 = ~n7839 & n9218;
  assign n9220 = n7845 & ~n9219;
  assign n9221 = ~n7844 & ~n7882;
  assign n9222 = ~n7896 & n9221;
  assign n9223 = n7854 & ~n9222;
  assign n9224 = n8961 & n9217;
  assign n9225 = ~n7840 & n9224;
  assign n9226 = ~n7852 & n7905;
  assign n9227 = ~n9225 & ~n9226;
  assign n9228 = ~n7857 & ~n9227;
  assign n9229 = ~n7874 & n9228;
  assign n9230 = ~n7898 & ~n9229;
  assign n9231 = ~n9223 & ~n9230;
  assign n9232 = ~n9220 & n9231;
  assign n9233 = ~n9216 & n9232;
  assign n9234 = n7867 & n9233;
  assign n9235 = n7856 & n9234;
  assign n9236 = n8959 & n9235;
  assign n9237 = n9215 & n9236;
  assign n9238 = n9237 ^ n5561;
  assign n9239 = n9238 ^ x100;
  assign n9240 = ~n9212 & ~n9239;
  assign n9241 = n8734 & ~n8764;
  assign n9242 = ~n8785 & ~n9241;
  assign n9243 = n8732 & n8788;
  assign n9244 = n8733 & n8795;
  assign n9245 = ~n9243 & ~n9244;
  assign n9246 = n9242 & n9245;
  assign n9247 = n8783 & ~n9246;
  assign n9248 = n8733 & n8766;
  assign n9249 = n8784 & n8786;
  assign n9250 = n8732 & n8795;
  assign n9251 = ~n9249 & ~n9250;
  assign n9252 = ~n9248 & n9251;
  assign n9253 = n8732 & n8766;
  assign n9254 = ~n8731 & n8813;
  assign n9255 = ~n9253 & ~n9254;
  assign n9256 = n9252 & n9255;
  assign n9257 = n8794 & ~n9256;
  assign n9258 = ~n9247 & ~n9257;
  assign n9259 = ~n8764 & n8808;
  assign n9260 = n8766 & n8786;
  assign n9261 = ~n9259 & ~n9260;
  assign n9262 = n8764 & n8786;
  assign n9263 = n8731 & n8784;
  assign n9264 = ~n9262 & ~n9263;
  assign n9265 = ~n8809 & n9264;
  assign n9266 = ~n9248 & n9265;
  assign n9267 = n9261 & n9266;
  assign n9268 = n9267 ^ n8768;
  assign n9269 = n9268 ^ n9267;
  assign n9270 = n9252 & n9261;
  assign n9271 = n9245 & n9270;
  assign n9272 = n9271 ^ n9267;
  assign n9273 = n9269 & ~n9272;
  assign n9274 = n9273 ^ n9267;
  assign n9275 = n8769 & n9274;
  assign n9276 = n9258 & ~n9275;
  assign n9277 = n9276 ^ n5671;
  assign n9278 = n9277 ^ x91;
  assign n9279 = ~n7993 & n8174;
  assign n9280 = ~n8164 & ~n8183;
  assign n9281 = n7994 & ~n9280;
  assign n9282 = ~n8165 & n9017;
  assign n9283 = n8154 & ~n9282;
  assign n9284 = n8168 & n9009;
  assign n9285 = n8141 & ~n9284;
  assign n9286 = ~n9283 & ~n9285;
  assign n9287 = n8149 & n8162;
  assign n9288 = n8065 ^ n8030;
  assign n9289 = n8137 ^ n8030;
  assign n9290 = n9288 & n9289;
  assign n9291 = n9290 ^ n8030;
  assign n9292 = n8101 & n9291;
  assign n9293 = n7993 & ~n9292;
  assign n9294 = n8156 & ~n8186;
  assign n9295 = n8173 & n9294;
  assign n9296 = ~n8166 & n9294;
  assign n9297 = ~n8154 & n9296;
  assign n9298 = ~n9295 & ~n9297;
  assign n9299 = ~n9293 & n9298;
  assign n9300 = ~n9287 & ~n9299;
  assign n9301 = n9286 & n9300;
  assign n9302 = ~n9281 & n9301;
  assign n9303 = ~n9279 & n9302;
  assign n9304 = n9003 & n9303;
  assign n9305 = n8175 ^ n8162;
  assign n9306 = n8175 ^ n8154;
  assign n9307 = n9306 ^ n8154;
  assign n9308 = n8164 ^ n8154;
  assign n9309 = ~n9307 & ~n9308;
  assign n9310 = n9309 ^ n8154;
  assign n9311 = n9305 & n9310;
  assign n9312 = n9311 ^ n8162;
  assign n9313 = n9304 & ~n9312;
  assign n9314 = ~n8140 & n9313;
  assign n9315 = n9314 ^ n5355;
  assign n9316 = n9315 ^ x78;
  assign n9317 = ~n9278 & n9316;
  assign n9318 = n9240 & n9317;
  assign n9319 = n9187 & n9318;
  assign n9320 = ~n9143 & n9186;
  assign n9321 = ~n9212 & n9239;
  assign n9322 = n9317 & n9321;
  assign n9323 = n9320 & n9322;
  assign n9324 = n9212 & ~n9239;
  assign n9325 = n9278 & n9316;
  assign n9326 = n9324 & n9325;
  assign n9327 = n9187 & n9326;
  assign n9328 = ~n9323 & ~n9327;
  assign n9329 = ~n9319 & n9328;
  assign n9330 = n9278 & ~n9316;
  assign n9331 = n9321 & n9330;
  assign n9332 = ~n9278 & ~n9316;
  assign n9333 = n9324 & n9332;
  assign n9334 = ~n9331 & ~n9333;
  assign n9335 = n9320 & ~n9334;
  assign n9336 = ~n9143 & ~n9186;
  assign n9337 = n9321 & n9332;
  assign n9338 = ~n9318 & ~n9337;
  assign n9339 = n9336 & ~n9338;
  assign n9340 = n9240 & n9330;
  assign n9341 = n9212 & n9239;
  assign n9342 = n9332 & n9341;
  assign n9343 = n9321 & n9325;
  assign n9344 = n9317 & n9324;
  assign n9345 = ~n9343 & ~n9344;
  assign n9346 = ~n9342 & n9345;
  assign n9347 = ~n9340 & n9346;
  assign n9348 = n9187 & ~n9347;
  assign n9349 = n9325 & n9341;
  assign n9350 = n9324 & n9330;
  assign n9351 = ~n9331 & ~n9350;
  assign n9352 = ~n9349 & n9351;
  assign n9353 = n9345 & n9352;
  assign n9354 = n9336 & ~n9353;
  assign n9355 = ~n9348 & ~n9354;
  assign n9356 = n9186 ^ n9143;
  assign n9357 = ~n9337 & ~n9350;
  assign n9358 = n9240 & n9325;
  assign n9359 = n9330 & n9341;
  assign n9360 = ~n9358 & ~n9359;
  assign n9361 = ~n9326 & n9360;
  assign n9362 = n9357 & n9361;
  assign n9363 = n9362 ^ n9186;
  assign n9364 = n9363 ^ n9362;
  assign n9365 = ~n9340 & ~n9359;
  assign n9366 = n9345 & n9365;
  assign n9367 = ~n9322 & n9366;
  assign n9368 = n9357 & n9367;
  assign n9369 = ~n9342 & n9368;
  assign n9370 = n9369 ^ n9362;
  assign n9371 = ~n9364 & ~n9370;
  assign n9372 = n9371 ^ n9362;
  assign n9373 = n9356 & ~n9372;
  assign n9374 = n9355 & ~n9373;
  assign n9375 = ~n9339 & n9374;
  assign n9376 = ~n9335 & n9375;
  assign n9377 = n9333 ^ n9186;
  assign n9378 = n9377 ^ n9333;
  assign n9379 = n9357 ^ n9333;
  assign n9380 = n9378 & ~n9379;
  assign n9381 = n9380 ^ n9333;
  assign n9382 = ~n9356 & n9381;
  assign n9383 = n9376 & ~n9382;
  assign n9384 = n9329 & n9383;
  assign n9385 = n9384 ^ n7420;
  assign n9386 = n9385 ^ x89;
  assign n9387 = n8807 & ~n9246;
  assign n9388 = n8770 & ~n9256;
  assign n9389 = ~n9387 & ~n9388;
  assign n9390 = ~n8769 & ~n9274;
  assign n9391 = n9389 & ~n9390;
  assign n9392 = n9391 ^ n6478;
  assign n9393 = n9392 ^ x69;
  assign n9394 = n9315 ^ x86;
  assign n9395 = n9393 & ~n9394;
  assign n9396 = n5961 & n7249;
  assign n9397 = ~n7280 & n9396;
  assign n9398 = n7049 & n7261;
  assign n9399 = ~n7287 & ~n9398;
  assign n9400 = n7259 & ~n9399;
  assign n9401 = ~n9397 & ~n9400;
  assign n9402 = n7250 & n7290;
  assign n9403 = n7250 & n7289;
  assign n9404 = ~n9402 & ~n9403;
  assign n9405 = n7259 & n7267;
  assign n9406 = n7249 & n7286;
  assign n9407 = ~n9405 & ~n9406;
  assign n9408 = n5961 & n7257;
  assign n9409 = n6629 ^ n6434;
  assign n9410 = n9409 ^ n7048;
  assign n9411 = ~n6892 & n9410;
  assign n9412 = n7250 & n9411;
  assign n9413 = ~n9408 & ~n9412;
  assign n9414 = ~n7269 & ~n7304;
  assign n9415 = ~n7290 & n9414;
  assign n9416 = ~n7260 & n9415;
  assign n9417 = n7288 & n9416;
  assign n9418 = n7279 & ~n9417;
  assign n9419 = ~n7050 & n7264;
  assign n9420 = ~n7277 & n9419;
  assign n9421 = n7259 & ~n9420;
  assign n9422 = ~n7289 & n7305;
  assign n9423 = ~n7290 & n9422;
  assign n9424 = n9396 & ~n9423;
  assign n9425 = ~n9421 & ~n9424;
  assign n9426 = ~n9418 & n9425;
  assign n9427 = n9413 & n9426;
  assign n9428 = n9407 & n9427;
  assign n9429 = n7260 ^ n5961;
  assign n9430 = n9429 ^ n7260;
  assign n9431 = ~n7253 & ~n7277;
  assign n9432 = n9431 ^ n7260;
  assign n9433 = ~n9430 & ~n9432;
  assign n9434 = n9433 ^ n7260;
  assign n9435 = ~n7249 & n9434;
  assign n9436 = n9428 & ~n9435;
  assign n9437 = n9404 & n9436;
  assign n9438 = n9401 & n9437;
  assign n9439 = n9438 ^ n6933;
  assign n9440 = n9439 ^ x110;
  assign n9441 = n8528 & ~n8554;
  assign n9442 = n8499 & n8530;
  assign n9443 = n8565 & n9442;
  assign n9444 = ~n9441 & ~n9443;
  assign n9445 = ~n8541 & ~n8631;
  assign n9446 = n8528 & ~n9445;
  assign n9447 = ~n8550 & n8569;
  assign n9448 = n8545 & ~n9447;
  assign n9449 = ~n8535 & ~n9442;
  assign n9450 = n8528 & ~n9449;
  assign n9451 = ~n8557 & n8576;
  assign n9452 = n8565 & ~n9451;
  assign n9453 = ~n9450 & ~n9452;
  assign n9454 = ~n9448 & n9453;
  assign n9455 = ~n8544 & n8580;
  assign n9456 = ~n8537 & n9455;
  assign n9457 = ~n8497 & ~n8545;
  assign n9458 = ~n9456 & ~n9457;
  assign n9459 = ~n8566 & ~n9458;
  assign n9460 = ~n8546 & ~n9459;
  assign n9461 = n9454 & ~n9460;
  assign n9462 = n8539 & n9461;
  assign n9463 = ~n9446 & n9462;
  assign n9464 = n8501 & ~n8544;
  assign n9465 = n9464 ^ n8527;
  assign n9466 = n9465 ^ n9464;
  assign n9467 = n8459 & n8552;
  assign n9468 = ~n8557 & ~n9467;
  assign n9469 = ~n8550 & n9468;
  assign n9470 = ~n8544 & n9469;
  assign n9471 = n9470 ^ n9464;
  assign n9472 = n9466 & n9471;
  assign n9473 = n9472 ^ n9464;
  assign n9474 = ~n8526 & ~n9473;
  assign n9475 = n9463 & ~n9474;
  assign n9476 = n9444 & n9475;
  assign n9477 = n9476 ^ n6967;
  assign n9478 = n9477 ^ x125;
  assign n9479 = ~n9440 & n9478;
  assign n9480 = n9142 ^ x108;
  assign n9481 = n8244 & n8395;
  assign n9482 = n8365 & ~n8667;
  assign n9483 = ~n9481 & ~n9482;
  assign n9484 = ~n8390 & n8672;
  assign n9485 = ~n8400 & ~n9484;
  assign n9486 = n8354 & n8365;
  assign n9487 = n8245 & ~n8384;
  assign n9488 = ~n9486 & ~n9487;
  assign n9489 = n8401 & n8406;
  assign n9490 = n8383 & n8389;
  assign n9491 = ~n8377 & ~n8385;
  assign n9492 = n8356 & ~n9491;
  assign n9493 = ~n9490 & ~n9492;
  assign n9494 = ~n9489 & n9493;
  assign n9495 = n9488 & n9494;
  assign n9496 = ~n9485 & n9495;
  assign n9497 = n9483 & n9496;
  assign n9498 = ~n8363 & n9497;
  assign n9499 = n9193 & n9498;
  assign n9500 = n8663 & n9499;
  assign n9501 = n9500 ^ n6560;
  assign n9502 = n9501 ^ x83;
  assign n9503 = ~n9480 & ~n9502;
  assign n9504 = n9479 & n9503;
  assign n9505 = n9440 & n9478;
  assign n9506 = n9480 & ~n9502;
  assign n9507 = n9505 & n9506;
  assign n9508 = ~n9504 & ~n9507;
  assign n9509 = n9395 & ~n9508;
  assign n9510 = ~n9393 & n9394;
  assign n9511 = n9480 & n9502;
  assign n9512 = n9479 & n9511;
  assign n9513 = ~n9480 & n9502;
  assign n9514 = n9505 & n9513;
  assign n9515 = ~n9512 & ~n9514;
  assign n9516 = n9510 & ~n9515;
  assign n9517 = n9395 & n9514;
  assign n9518 = n9505 & n9511;
  assign n9519 = ~n9393 & ~n9394;
  assign n9520 = n9518 & n9519;
  assign n9521 = ~n9517 & ~n9520;
  assign n9522 = n9440 & ~n9478;
  assign n9523 = n9513 & n9522;
  assign n9524 = n9519 & n9523;
  assign n9525 = ~n9440 & ~n9478;
  assign n9526 = n9503 & n9525;
  assign n9527 = n9506 & n9522;
  assign n9528 = ~n9526 & ~n9527;
  assign n9529 = n9510 & ~n9528;
  assign n9530 = ~n9524 & ~n9529;
  assign n9531 = n9513 & n9525;
  assign n9532 = n9511 & n9522;
  assign n9533 = ~n9531 & ~n9532;
  assign n9534 = ~n9519 & ~n9533;
  assign n9535 = n9506 & n9525;
  assign n9536 = ~n9504 & ~n9535;
  assign n9537 = n9510 & ~n9536;
  assign n9538 = ~n9534 & ~n9537;
  assign n9539 = n9393 & n9394;
  assign n9540 = n9479 & n9513;
  assign n9541 = n9511 & n9525;
  assign n9542 = ~n9540 & ~n9541;
  assign n9543 = n9539 & ~n9542;
  assign n9544 = n9503 & n9522;
  assign n9545 = ~n9535 & ~n9544;
  assign n9546 = ~n9518 & n9545;
  assign n9547 = n9395 & ~n9546;
  assign n9548 = ~n9543 & ~n9547;
  assign n9549 = n9503 & n9505;
  assign n9550 = n9479 & n9506;
  assign n9551 = ~n9544 & ~n9550;
  assign n9552 = ~n9527 & n9551;
  assign n9553 = ~n9539 & n9552;
  assign n9554 = ~n9507 & n9545;
  assign n9555 = ~n9519 & n9554;
  assign n9556 = ~n9553 & ~n9555;
  assign n9557 = ~n9549 & ~n9556;
  assign n9558 = n9557 ^ n9519;
  assign n9559 = ~n9512 & ~n9540;
  assign n9560 = n9559 ^ n9557;
  assign n9561 = n9560 ^ n9559;
  assign n9562 = n9559 ^ n9539;
  assign n9563 = ~n9561 & n9562;
  assign n9564 = n9563 ^ n9559;
  assign n9565 = ~n9558 & n9564;
  assign n9566 = n9565 ^ n9519;
  assign n9567 = n9548 & ~n9566;
  assign n9568 = n9538 & n9567;
  assign n9569 = n9530 & n9568;
  assign n9570 = n9521 & n9569;
  assign n9571 = ~n9516 & n9570;
  assign n9572 = ~n9509 & n9571;
  assign n9573 = n9572 ^ n7597;
  assign n9574 = n9573 ^ x106;
  assign n9575 = n9386 & ~n9574;
  assign n9576 = n9114 & n9575;
  assign n9577 = n7672 ^ x75;
  assign n9578 = n9501 ^ x93;
  assign n9579 = ~n9577 & n9578;
  assign n9580 = n9392 ^ x94;
  assign n9581 = n7840 & ~n9217;
  assign n9582 = n7836 & ~n8961;
  assign n9583 = ~n9581 & ~n9582;
  assign n9584 = n7853 & ~n7899;
  assign n9585 = ~n7903 & n9584;
  assign n9586 = n7845 & ~n9585;
  assign n9587 = ~n7857 & n7883;
  assign n9588 = ~n7896 & n9587;
  assign n9589 = n7854 & ~n9588;
  assign n9590 = ~n7874 & n7900;
  assign n9591 = ~n7862 & n9590;
  assign n9592 = n7840 & ~n9591;
  assign n9593 = ~n9589 & ~n9592;
  assign n9594 = ~n7880 & n9222;
  assign n9595 = n7845 & ~n9594;
  assign n9596 = ~n7862 & n9222;
  assign n9597 = n7836 & ~n9596;
  assign n9598 = ~n7852 & n8970;
  assign n9599 = ~n7870 & n9598;
  assign n9600 = n7854 & ~n9599;
  assign n9601 = ~n9597 & ~n9600;
  assign n9602 = ~n9595 & n9601;
  assign n9603 = n9593 & n9602;
  assign n9604 = ~n9586 & n9603;
  assign n9605 = n9583 & n9604;
  assign n9606 = n9215 & n9605;
  assign n9607 = n7842 & n9606;
  assign n9608 = n9607 ^ n6514;
  assign n9609 = n9608 ^ x124;
  assign n9610 = ~n9580 & ~n9609;
  assign n9611 = n8825 & n8929;
  assign n9612 = ~n8885 & ~n8910;
  assign n9613 = ~n8933 & n9612;
  assign n9614 = n8891 & ~n9613;
  assign n9615 = ~n8885 & n9166;
  assign n9616 = n8903 & ~n9615;
  assign n9617 = ~n9614 & ~n9616;
  assign n9618 = ~n9611 & n9617;
  assign n9619 = ~n8909 & ~n8935;
  assign n9620 = ~n8916 & n9173;
  assign n9621 = n8913 & n9620;
  assign n9622 = ~n8893 & n9621;
  assign n9623 = n8899 & ~n9622;
  assign n9624 = ~n9619 & ~n9623;
  assign n9625 = n9618 & n9624;
  assign n9626 = n8908 & n9625;
  assign n9627 = n9161 & n9626;
  assign n9628 = n8898 & n9627;
  assign n9629 = n9628 ^ n6468;
  assign n9630 = n9629 ^ x76;
  assign n9631 = n7320 ^ x117;
  assign n9632 = ~n9630 & ~n9631;
  assign n9633 = n9610 & n9632;
  assign n9634 = n9579 & n9633;
  assign n9635 = n9577 & ~n9578;
  assign n9636 = n9630 & n9631;
  assign n9637 = n9610 & n9636;
  assign n9638 = n9580 & n9609;
  assign n9639 = n9636 & n9638;
  assign n9640 = ~n9637 & ~n9639;
  assign n9641 = n9635 & ~n9640;
  assign n9642 = ~n9634 & ~n9641;
  assign n9643 = ~n9630 & n9631;
  assign n9644 = n9610 & n9643;
  assign n9645 = n9635 & n9644;
  assign n9646 = n9580 & ~n9609;
  assign n9647 = n9632 & n9646;
  assign n9648 = n9579 & n9647;
  assign n9649 = ~n9645 & ~n9648;
  assign n9650 = ~n9577 & ~n9578;
  assign n9651 = n9639 & n9650;
  assign n9652 = ~n9580 & n9609;
  assign n9653 = n9630 & ~n9631;
  assign n9654 = n9652 & n9653;
  assign n9655 = n9579 & n9654;
  assign n9656 = ~n9651 & ~n9655;
  assign n9657 = n9638 & n9643;
  assign n9658 = ~n9637 & ~n9657;
  assign n9659 = n9579 & ~n9658;
  assign n9660 = n9636 & n9646;
  assign n9661 = n9636 & n9652;
  assign n9662 = ~n9660 & ~n9661;
  assign n9663 = n9579 & ~n9662;
  assign n9664 = n9638 & n9653;
  assign n9665 = n9632 & n9638;
  assign n9666 = ~n9664 & ~n9665;
  assign n9667 = n9632 & n9652;
  assign n9668 = n9646 & n9653;
  assign n9669 = ~n9667 & ~n9668;
  assign n9670 = n9666 & n9669;
  assign n9671 = n9635 & ~n9670;
  assign n9672 = ~n9663 & ~n9671;
  assign n9673 = n9577 & n9578;
  assign n9674 = ~n9650 & ~n9673;
  assign n9675 = n9643 & n9652;
  assign n9676 = ~n9660 & ~n9675;
  assign n9677 = ~n9644 & ~n9647;
  assign n9678 = ~n9665 & n9677;
  assign n9679 = ~n9654 & n9678;
  assign n9680 = ~n9673 & n9679;
  assign n9681 = n9610 & n9653;
  assign n9682 = ~n9665 & ~n9681;
  assign n9683 = ~n9633 & n9682;
  assign n9684 = ~n9647 & n9683;
  assign n9685 = ~n9650 & n9684;
  assign n9686 = ~n9680 & ~n9685;
  assign n9687 = n9676 & ~n9686;
  assign n9688 = ~n9674 & ~n9687;
  assign n9689 = n9672 & ~n9688;
  assign n9690 = n9643 & n9646;
  assign n9691 = n9690 ^ n9668;
  assign n9692 = n9691 ^ n9690;
  assign n9693 = n9690 ^ n9578;
  assign n9694 = n9693 ^ n9690;
  assign n9695 = n9692 & n9694;
  assign n9696 = n9695 ^ n9690;
  assign n9697 = ~n9577 & n9696;
  assign n9698 = n9697 ^ n9690;
  assign n9699 = n9689 & ~n9698;
  assign n9700 = n9578 ^ n9577;
  assign n9701 = n9661 ^ n9578;
  assign n9702 = n9701 ^ n9661;
  assign n9703 = n9664 ^ n9661;
  assign n9704 = n9702 & n9703;
  assign n9705 = n9704 ^ n9661;
  assign n9706 = ~n9700 & n9705;
  assign n9707 = n9699 & ~n9706;
  assign n9708 = ~n9659 & n9707;
  assign n9709 = n9656 & n9708;
  assign n9710 = n9649 & n9709;
  assign n9711 = n9642 & n9710;
  assign n9712 = n9711 ^ n7392;
  assign n9713 = n9712 ^ x113;
  assign n9714 = n8954 ^ x122;
  assign n9715 = n7267 & n9396;
  assign n9716 = n7259 & n7277;
  assign n9717 = ~n9715 & ~n9716;
  assign n9718 = n7050 & ~n7283;
  assign n9719 = n7264 & ~n7270;
  assign n9720 = ~n7290 & n9719;
  assign n9721 = n7279 & ~n9720;
  assign n9722 = ~n9718 & ~n9721;
  assign n9723 = n5961 & n7286;
  assign n9724 = n7265 & ~n7269;
  assign n9725 = n7250 & ~n9724;
  assign n9728 = ~n7287 & ~n7289;
  assign n9726 = ~n7284 & n7305;
  assign n9727 = ~n7267 & n9726;
  assign n9729 = n9728 ^ n9727;
  assign n9730 = n9729 ^ n9728;
  assign n9731 = n9728 ^ n7249;
  assign n9732 = n9731 ^ n9728;
  assign n9733 = ~n9730 & n9732;
  assign n9734 = n9733 ^ n9728;
  assign n9735 = n7283 & ~n9734;
  assign n9736 = n9735 ^ n9728;
  assign n9737 = ~n9725 & n9736;
  assign n9738 = ~n9723 & n9737;
  assign n9739 = n9722 & n9738;
  assign n9740 = n9717 & n9739;
  assign n9741 = n9401 & n9740;
  assign n9742 = ~n9402 & n9741;
  assign n9743 = ~n7260 & n9742;
  assign n9744 = n9743 ^ n6658;
  assign n9745 = n9744 ^ x66;
  assign n9746 = ~n9714 & n9745;
  assign n9747 = n7651 & ~n9116;
  assign n9748 = ~n9124 & ~n9747;
  assign n9749 = ~n7633 & ~n7648;
  assign n9750 = ~n7358 & n7600;
  assign n9752 = n7612 & n7621;
  assign n9751 = n7652 & n9116;
  assign n9753 = n9752 ^ n9751;
  assign n9754 = n9752 ^ n7393;
  assign n9755 = n9754 ^ n9752;
  assign n9756 = n9753 & ~n9755;
  assign n9757 = n9756 ^ n9752;
  assign n9758 = ~n7358 & ~n9757;
  assign n9759 = ~n7626 & ~n7646;
  assign n9760 = n9130 & n9759;
  assign n9761 = n7635 & n9760;
  assign n9762 = n9761 ^ n7393;
  assign n9763 = n9762 ^ n9761;
  assign n9764 = n7622 & ~n7628;
  assign n9765 = ~n7611 & n9764;
  assign n9766 = n9765 ^ n9761;
  assign n9767 = ~n9763 & n9766;
  assign n9768 = n9767 ^ n9761;
  assign n9769 = n7358 & ~n9768;
  assign n9770 = ~n9758 & ~n9769;
  assign n9771 = ~n7632 & n9770;
  assign n9772 = ~n9750 & n9771;
  assign n9773 = ~n9749 & n9772;
  assign n9774 = n9748 & n9773;
  assign n9775 = n7630 & n9774;
  assign n9776 = n9775 ^ n6749;
  assign n9777 = n9776 ^ x120;
  assign n9778 = n8528 & n8557;
  assign n9779 = ~n8535 & n8567;
  assign n9780 = n8565 & ~n9779;
  assign n9781 = ~n9778 & ~n9780;
  assign n9787 = ~n8500 & ~n9442;
  assign n9788 = ~n8532 & n9787;
  assign n9789 = n8528 & ~n9788;
  assign n9790 = n8554 & ~n9789;
  assign n9791 = ~n8575 & n9790;
  assign n9782 = n8501 & ~n8532;
  assign n9783 = ~n8541 & n9782;
  assign n9784 = ~n8537 & n9783;
  assign n9785 = n8580 & n9457;
  assign n9786 = ~n9784 & ~n9785;
  assign n9792 = n9791 ^ n9786;
  assign n9793 = n9792 ^ n9791;
  assign n9794 = n8632 & n9468;
  assign n9795 = n9794 ^ n9791;
  assign n9796 = n9795 ^ n9791;
  assign n9797 = ~n9793 & n9796;
  assign n9798 = n9797 ^ n9791;
  assign n9799 = ~n8546 & n9798;
  assign n9800 = n9799 ^ n9791;
  assign n9801 = n9781 & n9800;
  assign n9802 = n8548 & n9801;
  assign n9803 = n9444 & n9802;
  assign n9804 = n9803 ^ n6788;
  assign n9805 = n9804 ^ x98;
  assign n9806 = n9777 & ~n9805;
  assign n9807 = n8697 ^ x81;
  assign n9808 = n8139 & ~n8173;
  assign n9809 = n7994 & ~n9008;
  assign n9810 = ~n9808 & ~n9809;
  assign n9811 = n8141 & ~n9296;
  assign n9812 = ~n8165 & ~n8184;
  assign n9813 = n8154 & ~n9812;
  assign n9814 = ~n8151 & n8185;
  assign n9815 = n8141 & ~n9814;
  assign n9816 = n8156 & ~n8187;
  assign n9817 = n8154 & ~n9816;
  assign n9818 = n8193 ^ n7993;
  assign n9819 = ~n8145 & ~n8160;
  assign n9820 = ~n8174 & n9819;
  assign n9821 = n9820 ^ n8189;
  assign n9822 = n8189 ^ n7952;
  assign n9823 = n9822 ^ n8189;
  assign n9824 = n9821 & n9823;
  assign n9825 = n9824 ^ n8189;
  assign n9826 = n9825 ^ n8193;
  assign n9827 = n9818 & ~n9826;
  assign n9828 = n9827 ^ n9824;
  assign n9829 = n9828 ^ n8189;
  assign n9830 = n9829 ^ n7993;
  assign n9831 = ~n8193 & ~n9830;
  assign n9832 = n9831 ^ n8193;
  assign n9833 = n9832 ^ n7993;
  assign n9834 = ~n9817 & ~n9833;
  assign n9835 = ~n9815 & n9834;
  assign n9836 = n9000 & n9835;
  assign n9837 = ~n9813 & n9836;
  assign n9838 = ~n9811 & n9837;
  assign n9839 = n9810 & n9838;
  assign n9840 = ~n9312 & n9839;
  assign n9841 = n8997 & n9840;
  assign n9842 = n9841 ^ n6820;
  assign n9843 = n9842 ^ x72;
  assign n9844 = ~n9807 & n9843;
  assign n9845 = n9806 & n9844;
  assign n9846 = n9746 & n9845;
  assign n9847 = ~n9714 & ~n9745;
  assign n9848 = ~n9777 & n9805;
  assign n9849 = n9807 & ~n9843;
  assign n9850 = n9848 & n9849;
  assign n9851 = n9847 & n9850;
  assign n9852 = n9714 & n9745;
  assign n9853 = n9777 & n9805;
  assign n9854 = n9844 & n9853;
  assign n9855 = n9806 & n9849;
  assign n9856 = ~n9854 & ~n9855;
  assign n9857 = n9852 & ~n9856;
  assign n9858 = ~n9851 & ~n9857;
  assign n9859 = ~n9846 & n9858;
  assign n9860 = ~n9807 & ~n9843;
  assign n9861 = n9853 & n9860;
  assign n9862 = n9852 & n9861;
  assign n9863 = n9714 & ~n9745;
  assign n9864 = ~n9777 & ~n9805;
  assign n9865 = n9860 & n9864;
  assign n9866 = ~n9845 & ~n9865;
  assign n9867 = n9863 & ~n9866;
  assign n9868 = ~n9862 & ~n9867;
  assign n9869 = n9807 & n9843;
  assign n9870 = n9806 & n9869;
  assign n9871 = n9847 & n9870;
  assign n9872 = n9746 & n9865;
  assign n9873 = ~n9871 & ~n9872;
  assign n9874 = n9854 & n9863;
  assign n9875 = n9844 & n9848;
  assign n9876 = n9852 & n9875;
  assign n9877 = n9746 & n9850;
  assign n9878 = ~n9876 & ~n9877;
  assign n9879 = ~n9874 & n9878;
  assign n9880 = n9806 & n9860;
  assign n9881 = n9847 & n9880;
  assign n9882 = n9864 & n9869;
  assign n9883 = ~n9855 & ~n9882;
  assign n9884 = n9746 & ~n9883;
  assign n9885 = ~n9881 & ~n9884;
  assign n9886 = n9852 & n9880;
  assign n9887 = n9848 & n9860;
  assign n9888 = n9853 & n9869;
  assign n9889 = ~n9875 & ~n9888;
  assign n9890 = ~n9887 & n9889;
  assign n9891 = n9746 & ~n9890;
  assign n9892 = ~n9886 & ~n9891;
  assign n9893 = n9863 & n9887;
  assign n9894 = n9844 & n9864;
  assign n9895 = n9849 & n9853;
  assign n9896 = ~n9861 & ~n9882;
  assign n9897 = ~n9854 & n9896;
  assign n9898 = ~n9895 & n9897;
  assign n9899 = ~n9894 & n9898;
  assign n9900 = n9847 & ~n9899;
  assign n9901 = ~n9893 & ~n9900;
  assign n9907 = ~n9870 & ~n9882;
  assign n9908 = ~n9850 & n9907;
  assign n9902 = n9849 & n9864;
  assign n9903 = n9848 & n9869;
  assign n9904 = ~n9895 & ~n9903;
  assign n9905 = ~n9870 & n9904;
  assign n9906 = ~n9902 & n9905;
  assign n9909 = n9908 ^ n9906;
  assign n9910 = n9908 ^ n9745;
  assign n9911 = n9910 ^ n9908;
  assign n9912 = n9909 & ~n9911;
  assign n9913 = n9912 ^ n9908;
  assign n9914 = n9714 & ~n9913;
  assign n9915 = n9901 & ~n9914;
  assign n9916 = n9892 & n9915;
  assign n9917 = n9885 & n9916;
  assign n9918 = n9879 & n9917;
  assign n9919 = n9873 & n9918;
  assign n9920 = n9868 & n9919;
  assign n9921 = n9859 & n9920;
  assign n9922 = n9921 ^ n7357;
  assign n9923 = n9922 ^ x74;
  assign n9924 = n9713 & n9923;
  assign n9925 = ~n9713 & ~n9923;
  assign n9926 = ~n9924 & ~n9925;
  assign n9927 = n9576 & ~n9926;
  assign n9928 = n9923 ^ n9713;
  assign n9929 = ~n8629 & ~n9113;
  assign n9930 = n9575 & n9929;
  assign n9931 = n9930 ^ n9923;
  assign n9932 = n9931 ^ n9930;
  assign n9933 = ~n9386 & ~n9574;
  assign n9934 = n9114 & n9933;
  assign n9935 = n9386 & n9574;
  assign n9936 = n9114 & n9935;
  assign n9937 = ~n9934 & ~n9936;
  assign n9938 = n9937 ^ n9930;
  assign n9939 = ~n9932 & ~n9938;
  assign n9940 = n9939 ^ n9930;
  assign n9941 = n9928 & n9940;
  assign n9942 = ~n9927 & ~n9941;
  assign n9943 = ~n9386 & n9574;
  assign n9944 = n9114 & n9943;
  assign n9945 = n9713 & ~n9923;
  assign n9946 = n9944 & n9945;
  assign n9947 = ~n8629 & n9113;
  assign n9948 = n9575 & n9947;
  assign n9949 = n9943 & n9947;
  assign n9950 = ~n9948 & ~n9949;
  assign n9951 = ~n9926 & ~n9950;
  assign n9952 = ~n9946 & ~n9951;
  assign n9953 = ~n9713 & n9923;
  assign n9954 = n9929 & n9933;
  assign n9955 = n8629 & ~n9113;
  assign n9956 = n9943 & n9955;
  assign n9957 = n9575 & n9955;
  assign n9958 = ~n9956 & ~n9957;
  assign n9959 = ~n9954 & n9958;
  assign n9960 = n9953 & ~n9959;
  assign n9961 = n9933 & n9955;
  assign n9962 = n9929 & n9935;
  assign n9963 = n9935 & n9955;
  assign n9964 = ~n9956 & ~n9963;
  assign n9965 = ~n9962 & n9964;
  assign n9966 = ~n9961 & n9965;
  assign n9967 = n9925 & ~n9966;
  assign n9968 = n9574 ^ n9386;
  assign n9969 = n9386 ^ n8629;
  assign n9970 = n9969 ^ n9386;
  assign n9971 = ~n9968 & ~n9970;
  assign n9972 = n9971 ^ n9386;
  assign n9973 = n9113 & ~n9972;
  assign n9974 = n9953 & n9973;
  assign n9975 = n9933 & n9947;
  assign n9976 = n9929 & n9943;
  assign n9977 = ~n9975 & ~n9976;
  assign n9978 = ~n9963 & n9977;
  assign n9979 = ~n9945 & n9978;
  assign n9980 = ~n9961 & n9979;
  assign n9981 = ~n9957 & ~n9976;
  assign n9982 = ~n9954 & n9981;
  assign n9983 = ~n9930 & n9982;
  assign n9984 = n9945 & ~n9983;
  assign n9985 = ~n9924 & ~n9984;
  assign n9986 = ~n9980 & ~n9985;
  assign n9987 = ~n9974 & ~n9986;
  assign n9988 = ~n9967 & n9987;
  assign n9989 = ~n9960 & n9988;
  assign n9990 = n9935 & n9947;
  assign n9991 = n9990 ^ n9713;
  assign n9992 = n9991 ^ n9990;
  assign n9993 = n9990 ^ n9936;
  assign n9994 = n9993 ^ n9990;
  assign n9995 = n9992 & n9994;
  assign n9996 = n9995 ^ n9990;
  assign n9997 = n9923 & n9996;
  assign n9998 = n9997 ^ n9990;
  assign n9999 = n9989 & ~n9998;
  assign n10000 = n9952 & n9999;
  assign n10001 = n9942 & n10000;
  assign n10002 = n10001 ^ n7672;
  assign n10003 = n10002 ^ x118;
  assign n10004 = n7321 & ~n8592;
  assign n10005 = ~n8430 & n10004;
  assign n10006 = n7321 & n8592;
  assign n10007 = ~n8605 & n10006;
  assign n10008 = ~n10005 & ~n10007;
  assign n10009 = ~n7321 & n8592;
  assign n10010 = ~n8621 & n10009;
  assign n10011 = ~n7321 & ~n8592;
  assign n10012 = ~n8610 & ~n8612;
  assign n10013 = n10012 ^ n8204;
  assign n10014 = ~n8424 & n10013;
  assign n10015 = n10014 ^ n8204;
  assign n10016 = n10011 & ~n10015;
  assign n10017 = ~n10010 & ~n10016;
  assign n10018 = n10008 & n10017;
  assign n10019 = ~n8616 & n10018;
  assign n10020 = n10019 ^ n6433;
  assign n10021 = n10020 ^ x108;
  assign n10022 = ~n9847 & ~n9852;
  assign n10023 = ~n9887 & ~n9894;
  assign n10024 = ~n10022 & ~n10023;
  assign n10025 = n9746 & ~n9905;
  assign n10026 = ~n10024 & ~n10025;
  assign n10027 = n9714 & n9880;
  assign n10028 = ~n9845 & ~n9861;
  assign n10029 = n9847 & ~n10028;
  assign n10030 = ~n10027 & ~n10029;
  assign n10031 = ~n9865 & ~n9875;
  assign n10032 = n9863 & ~n10031;
  assign n10033 = n9746 & ~n9896;
  assign n10034 = ~n9888 & ~n9902;
  assign n10035 = ~n10022 & ~n10034;
  assign n10036 = ~n9895 & n9907;
  assign n10037 = ~n9855 & n10036;
  assign n10038 = n9863 & ~n10037;
  assign n10039 = ~n10035 & ~n10038;
  assign n10040 = ~n10033 & n10039;
  assign n10041 = n9873 & n10040;
  assign n10042 = n9859 & n10041;
  assign n10043 = ~n10032 & n10042;
  assign n10044 = n10030 & n10043;
  assign n10045 = n10026 & n10044;
  assign n10046 = n9879 & n10045;
  assign n10047 = n10046 ^ n8243;
  assign n10048 = n10047 ^ x94;
  assign n10049 = ~n10021 & n10048;
  assign n10050 = ~n8781 & n8794;
  assign n10051 = n8770 & ~n8805;
  assign n10052 = ~n10050 & ~n10051;
  assign n10053 = n8767 & n8769;
  assign n10054 = ~n8791 & n8807;
  assign n10055 = ~n10053 & ~n10054;
  assign n10056 = n8783 & ~n8816;
  assign n10057 = n10055 & ~n10056;
  assign n10058 = n10052 & n10057;
  assign n10059 = n10058 ^ n7694;
  assign n10060 = n10059 ^ x115;
  assign n10061 = ~n8895 & n9173;
  assign n10062 = ~n8889 & n10061;
  assign n10063 = ~n8912 & n10062;
  assign n10064 = ~n8885 & n10063;
  assign n10065 = n8891 & ~n10064;
  assign n10066 = ~n8934 & n9171;
  assign n10067 = ~n8938 & n10066;
  assign n10068 = ~n8941 & ~n10067;
  assign n10069 = n10068 ^ n8824;
  assign n10070 = n10069 ^ n10068;
  assign n10071 = ~n8905 & n8913;
  assign n10072 = ~n8901 & n10071;
  assign n10073 = n10072 ^ n10068;
  assign n10074 = n10073 ^ n10068;
  assign n10075 = ~n10070 & ~n10074;
  assign n10076 = n10075 ^ n10068;
  assign n10077 = ~n8823 & n10076;
  assign n10078 = n10077 ^ n10068;
  assign n10079 = ~n10065 & ~n10078;
  assign n10080 = n9158 ^ n8886;
  assign n10081 = n10080 ^ n9158;
  assign n10082 = n9158 ^ n8824;
  assign n10083 = n10082 ^ n9158;
  assign n10084 = ~n10081 & ~n10083;
  assign n10085 = n10084 ^ n9158;
  assign n10086 = n8909 & n10085;
  assign n10087 = n10086 ^ n9158;
  assign n10088 = n10079 & ~n10087;
  assign n10089 = ~n8890 & n10088;
  assign n10090 = n9156 & n10089;
  assign n10091 = n9146 & n10090;
  assign n10092 = ~n8887 & n10091;
  assign n10093 = n10092 ^ n7719;
  assign n10094 = n10093 ^ x114;
  assign n10095 = ~n10060 & ~n10094;
  assign n10096 = n8591 ^ x97;
  assign n10097 = n9744 ^ x88;
  assign n10098 = ~n10096 & n10097;
  assign n10099 = n10095 & n10098;
  assign n10100 = n10060 & n10094;
  assign n10101 = ~n10096 & ~n10097;
  assign n10102 = n10100 & n10101;
  assign n10103 = ~n10099 & ~n10102;
  assign n10104 = n7917 ^ x82;
  assign n10105 = n9842 ^ x121;
  assign n10106 = n10104 & n10105;
  assign n10107 = ~n10103 & n10106;
  assign n10108 = n10060 & ~n10094;
  assign n10109 = n10096 & ~n10097;
  assign n10110 = n10108 & n10109;
  assign n10111 = ~n10060 & n10094;
  assign n10112 = n10101 & n10111;
  assign n10113 = ~n10110 & ~n10112;
  assign n10114 = n10109 & n10111;
  assign n10115 = n10095 & n10101;
  assign n10116 = ~n10114 & ~n10115;
  assign n10117 = n10113 & n10116;
  assign n10118 = n10104 & ~n10105;
  assign n10119 = ~n10117 & n10118;
  assign n10120 = ~n10107 & ~n10119;
  assign n10121 = n10100 & n10109;
  assign n10122 = n10096 & n10097;
  assign n10123 = n10111 & n10122;
  assign n10124 = n10095 & n10122;
  assign n10125 = n10098 & n10108;
  assign n10126 = ~n10124 & ~n10125;
  assign n10127 = ~n10123 & n10126;
  assign n10128 = ~n10121 & n10127;
  assign n10129 = ~n10104 & n10105;
  assign n10130 = ~n10128 & n10129;
  assign n10131 = n10098 & n10111;
  assign n10132 = ~n10124 & ~n10131;
  assign n10133 = ~n10104 & ~n10105;
  assign n10134 = ~n10132 & n10133;
  assign n10135 = ~n10130 & ~n10134;
  assign n10136 = n10100 & n10122;
  assign n10137 = n10108 & n10122;
  assign n10138 = ~n10136 & ~n10137;
  assign n10139 = n10105 ^ n10104;
  assign n10140 = ~n10138 & ~n10139;
  assign n10141 = ~n10131 & ~n10136;
  assign n10142 = n10118 & ~n10141;
  assign n10143 = n10121 & n10133;
  assign n10144 = ~n10142 & ~n10143;
  assign n10145 = n10106 & ~n10117;
  assign n10146 = n10118 & ~n10126;
  assign n10147 = ~n10145 & ~n10146;
  assign n10148 = n10101 & n10108;
  assign n10149 = ~n10112 & ~n10148;
  assign n10150 = n10116 & n10149;
  assign n10151 = n10129 & ~n10150;
  assign n10152 = n10095 & n10109;
  assign n10153 = ~n10099 & ~n10112;
  assign n10154 = ~n10152 & n10153;
  assign n10155 = n10133 & ~n10154;
  assign n10156 = ~n10151 & ~n10155;
  assign n10157 = n10147 & n10156;
  assign n10158 = n10144 & n10157;
  assign n10159 = ~n10140 & n10158;
  assign n10160 = n10135 & n10159;
  assign n10161 = n10120 & n10160;
  assign n10162 = n10161 ^ n8320;
  assign n10163 = n10162 ^ x125;
  assign n10164 = n9143 & ~n9186;
  assign n10165 = ~n9351 & n10164;
  assign n10166 = n9240 & n9332;
  assign n10167 = n9187 & n10166;
  assign n10168 = n9320 & n9342;
  assign n10169 = ~n10167 & ~n10168;
  assign n10170 = ~n9187 & ~n9336;
  assign n10171 = ~n9349 & ~n9358;
  assign n10172 = n10170 & ~n10171;
  assign n10173 = n9345 & ~n10166;
  assign n10174 = ~n9337 & n10173;
  assign n10175 = n10164 & ~n10174;
  assign n10176 = ~n10172 & ~n10175;
  assign n10177 = n9336 & n9369;
  assign n10178 = ~n9340 & n9357;
  assign n10179 = ~n9344 & n10178;
  assign n10180 = n9320 & ~n10179;
  assign n10181 = ~n9331 & n9367;
  assign n10182 = n9187 & ~n10181;
  assign n10183 = ~n10180 & ~n10182;
  assign n10184 = ~n10177 & n10183;
  assign n10185 = n10176 & n10184;
  assign n10186 = n10169 & n10185;
  assign n10187 = n9328 & n10186;
  assign n10188 = ~n10165 & n10187;
  assign n10189 = n10188 ^ n5960;
  assign n10190 = n10189 ^ x69;
  assign n10191 = ~n10163 & n10190;
  assign n10192 = n9531 & n9539;
  assign n10193 = n9521 & ~n10192;
  assign n10194 = n9519 & ~n9536;
  assign n10195 = ~n9516 & ~n10194;
  assign n10196 = n9539 & ~n9545;
  assign n10197 = ~n9531 & ~n9550;
  assign n10198 = n9519 & ~n10197;
  assign n10199 = ~n10196 & ~n10198;
  assign n10200 = n9515 & ~n9523;
  assign n10201 = n9508 & n10200;
  assign n10202 = n9539 & ~n10201;
  assign n10203 = ~n9541 & ~n9549;
  assign n10204 = n9510 & ~n10203;
  assign n10205 = ~n9507 & ~n9544;
  assign n10206 = n9519 & ~n10205;
  assign n10207 = ~n10204 & ~n10206;
  assign n10208 = n9530 & n10207;
  assign n10209 = ~n10202 & n10208;
  assign n10210 = n9394 ^ n9393;
  assign n10211 = ~n9518 & ~n9540;
  assign n10212 = n10211 ^ n9394;
  assign n10213 = n10212 ^ n10211;
  assign n10214 = ~n9526 & ~n9550;
  assign n10215 = n9542 & n10214;
  assign n10216 = ~n9532 & n10215;
  assign n10217 = n10216 ^ n10211;
  assign n10218 = ~n10213 & n10217;
  assign n10219 = n10218 ^ n10211;
  assign n10220 = n10210 & ~n10219;
  assign n10221 = n10209 & ~n10220;
  assign n10222 = n10199 & n10221;
  assign n10223 = n10195 & n10222;
  assign n10224 = n10193 & n10223;
  assign n10225 = ~n9509 & n10224;
  assign n10226 = n10225 ^ n8351;
  assign n10227 = n10226 ^ x126;
  assign n10228 = n9043 & n9067;
  assign n10229 = ~n9041 & ~n9089;
  assign n10230 = n8699 & ~n10229;
  assign n10231 = ~n10228 & ~n10230;
  assign n10232 = n9058 & n9094;
  assign n10233 = n8659 & n9070;
  assign n10234 = ~n10232 & ~n10233;
  assign n10235 = n9043 & ~n9102;
  assign n10236 = ~n9046 & ~n9072;
  assign n10237 = ~n9060 & ~n10236;
  assign n10238 = ~n10235 & ~n10237;
  assign n10239 = n10234 & n10238;
  assign n10240 = ~n9054 & ~n9081;
  assign n10241 = n9059 & ~n10240;
  assign n10242 = ~n9079 & ~n9096;
  assign n10243 = n8699 & ~n10242;
  assign n10244 = ~n9089 & n9098;
  assign n10245 = n9059 & ~n10244;
  assign n10246 = ~n9054 & n9102;
  assign n10247 = ~n9067 & n10246;
  assign n10248 = n8699 & ~n10247;
  assign n10249 = ~n9050 & n10229;
  assign n10250 = ~n9095 & n10249;
  assign n10251 = ~n9043 & n10250;
  assign n10252 = ~n9063 & n9080;
  assign n10253 = ~n9041 & n10252;
  assign n10254 = ~n9058 & n10253;
  assign n10255 = n8659 & ~n10254;
  assign n10256 = ~n10251 & n10255;
  assign n10257 = ~n10248 & ~n10256;
  assign n10258 = ~n10245 & n10257;
  assign n10259 = ~n10243 & n10258;
  assign n10260 = ~n10241 & n10259;
  assign n10261 = n10239 & n10260;
  assign n10262 = n10231 & n10261;
  assign n10263 = n10262 ^ n8283;
  assign n10264 = n10263 ^ x76;
  assign n10265 = n10227 & ~n10264;
  assign n10266 = n10191 & n10265;
  assign n10267 = n10049 & n10266;
  assign n10268 = n10021 & ~n10048;
  assign n10269 = n10163 & ~n10190;
  assign n10270 = n10265 & n10269;
  assign n10271 = n10163 & n10190;
  assign n10272 = n10227 & n10264;
  assign n10273 = n10271 & n10272;
  assign n10274 = ~n10163 & ~n10190;
  assign n10275 = n10272 & n10274;
  assign n10276 = ~n10273 & ~n10275;
  assign n10277 = ~n10270 & n10276;
  assign n10278 = n10268 & ~n10277;
  assign n10279 = ~n10021 & ~n10048;
  assign n10280 = ~n10227 & ~n10264;
  assign n10281 = n10191 & n10280;
  assign n10282 = ~n10227 & n10264;
  assign n10283 = n10191 & n10282;
  assign n10284 = n10269 & n10280;
  assign n10285 = ~n10283 & ~n10284;
  assign n10286 = ~n10281 & n10285;
  assign n10287 = n10279 & ~n10286;
  assign n10288 = ~n10278 & ~n10287;
  assign n10289 = n10021 & n10048;
  assign n10290 = n10274 & n10280;
  assign n10291 = n10271 & n10280;
  assign n10292 = ~n10290 & ~n10291;
  assign n10293 = n10289 & ~n10292;
  assign n10294 = n10274 & n10282;
  assign n10295 = n10289 & n10294;
  assign n10296 = n10265 & n10271;
  assign n10297 = n10268 & n10296;
  assign n10298 = ~n10295 & ~n10297;
  assign n10299 = ~n10021 & n10294;
  assign n10300 = n10048 ^ n10021;
  assign n10301 = n10191 & n10272;
  assign n10302 = n10269 & n10272;
  assign n10303 = ~n10301 & ~n10302;
  assign n10304 = ~n10300 & ~n10303;
  assign n10305 = ~n10299 & ~n10304;
  assign n10306 = n10265 & n10274;
  assign n10307 = ~n10296 & ~n10306;
  assign n10308 = n10279 & ~n10307;
  assign n10309 = n10269 & n10282;
  assign n10310 = ~n10266 & ~n10284;
  assign n10311 = ~n10309 & n10310;
  assign n10312 = n10289 & ~n10311;
  assign n10313 = n10276 & ~n10306;
  assign n10314 = n10049 & ~n10313;
  assign n10315 = n10271 & n10282;
  assign n10316 = n10300 & n10315;
  assign n10317 = ~n10291 & ~n10309;
  assign n10318 = n10049 & ~n10317;
  assign n10319 = n10285 & n10313;
  assign n10320 = n10268 & ~n10319;
  assign n10321 = ~n10318 & ~n10320;
  assign n10322 = ~n10316 & n10321;
  assign n10323 = ~n10314 & n10322;
  assign n10324 = ~n10312 & n10323;
  assign n10325 = ~n10308 & n10324;
  assign n10326 = n10305 & n10325;
  assign n10327 = n10298 & n10326;
  assign n10328 = ~n10293 & n10327;
  assign n10329 = n10288 & n10328;
  assign n10330 = ~n10267 & n10329;
  assign n10331 = n10330 ^ n9501;
  assign n10332 = n10331 ^ x69;
  assign n10333 = n10003 & n10332;
  assign n10334 = n10189 ^ x120;
  assign n10335 = n8821 ^ x116;
  assign n10336 = n9238 ^ x102;
  assign n10337 = ~n10335 & n10336;
  assign n10338 = n8658 ^ x77;
  assign n10339 = ~n7263 & ~n7284;
  assign n10340 = n9396 & ~n10339;
  assign n10341 = n7250 & ~n7272;
  assign n10342 = ~n10340 & ~n10341;
  assign n10343 = n7279 & ~n7307;
  assign n10344 = ~n7257 & ~n7270;
  assign n10345 = ~n7283 & ~n10344;
  assign n10346 = ~n7253 & n9416;
  assign n10347 = n7259 & ~n10346;
  assign n10348 = ~n10345 & ~n10347;
  assign n10349 = ~n10343 & n10348;
  assign n10350 = n10342 & n10349;
  assign n10351 = n9407 & n10350;
  assign n10352 = ~n9435 & n10351;
  assign n10353 = n7255 & n10352;
  assign n10354 = n9717 & n10353;
  assign n10355 = n9404 & n10354;
  assign n10356 = n10355 ^ n7172;
  assign n10357 = n10356 ^ x84;
  assign n10358 = n10338 & n10357;
  assign n10359 = n9185 ^ x67;
  assign n10360 = ~n7621 & n7651;
  assign n10361 = ~n7631 & n9131;
  assign n10362 = n7394 & ~n10361;
  assign n10363 = ~n7611 & ~n7638;
  assign n10364 = n7616 & ~n10363;
  assign n10365 = n7621 & n9116;
  assign n10366 = n7394 & ~n10365;
  assign n10367 = ~n10364 & ~n10366;
  assign n10368 = ~n7626 & n7635;
  assign n10369 = n7606 & ~n10368;
  assign n10370 = n7635 & n9123;
  assign n10371 = n7651 & ~n10370;
  assign n10372 = n7616 ^ n7606;
  assign n10374 = ~n7603 & ~n7662;
  assign n10375 = n9116 & n10374;
  assign n10373 = n7604 & n9119;
  assign n10376 = n10375 ^ n10373;
  assign n10377 = n10375 ^ n7616;
  assign n10378 = n10377 ^ n10375;
  assign n10379 = ~n10376 & ~n10378;
  assign n10380 = n10379 ^ n10375;
  assign n10381 = n10372 & ~n10380;
  assign n10382 = n10381 ^ n7606;
  assign n10383 = ~n10371 & ~n10382;
  assign n10384 = ~n10369 & n10383;
  assign n10385 = n10367 & n10384;
  assign n10386 = ~n10362 & n10385;
  assign n10387 = ~n10360 & n10386;
  assign n10388 = n9748 & n10387;
  assign n10389 = n7630 & n10388;
  assign n10390 = n10389 ^ n7124;
  assign n10391 = n10390 ^ x70;
  assign n10392 = ~n10359 & n10391;
  assign n10393 = n10358 & n10392;
  assign n10394 = ~n10359 & ~n10391;
  assign n10395 = n10358 & n10394;
  assign n10396 = ~n10393 & ~n10395;
  assign n10397 = n10359 & n10391;
  assign n10398 = n10338 & ~n10357;
  assign n10399 = n10397 & n10398;
  assign n10400 = n10359 & ~n10391;
  assign n10401 = ~n10338 & ~n10357;
  assign n10402 = n10400 & n10401;
  assign n10403 = ~n10399 & ~n10402;
  assign n10404 = n10396 & n10403;
  assign n10405 = n10337 & ~n10404;
  assign n10406 = n10398 & n10400;
  assign n10407 = n10337 & n10406;
  assign n10408 = n10335 & ~n10336;
  assign n10409 = ~n10338 & n10357;
  assign n10410 = n10392 & n10409;
  assign n10411 = n10392 & n10398;
  assign n10412 = ~n10410 & ~n10411;
  assign n10413 = n10408 & ~n10412;
  assign n10414 = ~n10407 & ~n10413;
  assign n10415 = n10335 & n10336;
  assign n10416 = n10397 & n10409;
  assign n10417 = n10415 & n10416;
  assign n10418 = ~n10335 & ~n10336;
  assign n10419 = n10400 & n10409;
  assign n10420 = n10358 & n10397;
  assign n10421 = ~n10419 & ~n10420;
  assign n10422 = n10418 & ~n10421;
  assign n10423 = ~n10417 & ~n10422;
  assign n10424 = n10357 ^ n10338;
  assign n10425 = n10397 & ~n10424;
  assign n10426 = n10408 & n10425;
  assign n10427 = n10358 & n10400;
  assign n10428 = n10415 & n10427;
  assign n10429 = ~n10426 & ~n10428;
  assign n10430 = ~n10338 & n10394;
  assign n10431 = ~n10416 & ~n10430;
  assign n10432 = n10337 & ~n10431;
  assign n10433 = n10394 & n10401;
  assign n10434 = ~n10393 & ~n10419;
  assign n10435 = ~n10433 & n10434;
  assign n10436 = ~n10406 & n10435;
  assign n10437 = n10408 & ~n10436;
  assign n10438 = ~n10432 & ~n10437;
  assign n10439 = n10392 & n10401;
  assign n10440 = n10394 & n10398;
  assign n10441 = ~n10439 & ~n10440;
  assign n10442 = n10418 & ~n10441;
  assign n10443 = ~n10415 & ~n10418;
  assign n10444 = ~n10357 & n10397;
  assign n10445 = n10396 & ~n10415;
  assign n10446 = ~n10433 & n10441;
  assign n10447 = ~n10395 & n10446;
  assign n10448 = ~n10418 & n10447;
  assign n10449 = ~n10445 & ~n10448;
  assign n10450 = ~n10444 & ~n10449;
  assign n10451 = ~n10443 & ~n10450;
  assign n10452 = ~n10442 & ~n10451;
  assign n10453 = n10438 & n10452;
  assign n10454 = n10429 & n10453;
  assign n10455 = n10423 & n10454;
  assign n10456 = n10414 & n10455;
  assign n10457 = ~n10405 & n10456;
  assign n10458 = n10457 ^ n7248;
  assign n10459 = n10458 ^ x98;
  assign n10460 = ~n10334 & n10459;
  assign n10461 = ~n9527 & ~n9531;
  assign n10462 = n9395 & ~n10461;
  assign n10463 = ~n9514 & n9542;
  assign n10464 = ~n9531 & n10463;
  assign n10465 = n9510 & ~n10464;
  assign n10466 = ~n10462 & ~n10465;
  assign n10467 = n9539 & ~n10214;
  assign n10468 = ~n9535 & ~n9549;
  assign n10469 = n9519 & ~n10468;
  assign n10470 = ~n9523 & n9559;
  assign n10471 = n9539 & ~n10470;
  assign n10472 = ~n9518 & ~n9523;
  assign n10473 = n9542 & n10472;
  assign n10474 = n9395 & ~n10473;
  assign n10475 = ~n10471 & ~n10474;
  assign n10476 = n9519 & n9532;
  assign n10477 = ~n9504 & n10205;
  assign n10478 = ~n9527 & n10477;
  assign n10479 = n9510 & ~n10478;
  assign n10480 = ~n10476 & ~n10479;
  assign n10481 = n10475 & n10480;
  assign n10482 = n9532 ^ n9394;
  assign n10483 = n10482 ^ n9532;
  assign n10484 = n10200 ^ n9532;
  assign n10485 = ~n10483 & ~n10484;
  assign n10486 = n10485 ^ n9532;
  assign n10487 = ~n10210 & n10486;
  assign n10488 = n10481 & ~n10487;
  assign n10489 = ~n10469 & n10488;
  assign n10490 = ~n10467 & n10489;
  assign n10491 = n10466 & n10490;
  assign n10492 = n10199 & n10491;
  assign n10493 = ~n9509 & n10492;
  assign n10494 = n10493 ^ n7047;
  assign n10495 = n10494 ^ x65;
  assign n10496 = n10020 ^ x96;
  assign n10497 = ~n10495 & n10496;
  assign n10498 = ~n9644 & ~n9675;
  assign n10499 = n9579 & ~n10498;
  assign n10500 = n9640 & n9676;
  assign n10501 = n9650 & ~n10500;
  assign n10502 = ~n10499 & ~n10501;
  assign n10503 = ~n9654 & ~n9690;
  assign n10504 = n9650 & ~n10503;
  assign n10505 = ~n9668 & n9682;
  assign n10506 = ~n9654 & n10505;
  assign n10507 = n9635 & ~n10506;
  assign n10508 = ~n10504 & ~n10507;
  assign n10509 = ~n9657 & ~n9660;
  assign n10510 = ~n9690 & n10509;
  assign n10511 = n9635 & ~n10510;
  assign n10512 = ~n9654 & n9666;
  assign n10513 = n9579 & ~n10512;
  assign n10514 = ~n10511 & ~n10513;
  assign n10515 = n9649 & n10514;
  assign n10516 = n10508 & n10515;
  assign n10517 = n10502 & n10516;
  assign n10518 = n9673 ^ n9669;
  assign n10519 = n9669 ^ n9650;
  assign n10520 = n10519 ^ n9650;
  assign n10521 = n9630 ^ n9609;
  assign n10522 = n10521 ^ n9580;
  assign n10523 = n10522 ^ n9609;
  assign n10524 = n10523 ^ n9631;
  assign n10525 = n10521 ^ n9631;
  assign n10526 = n10525 ^ n10521;
  assign n10527 = n10521 ^ n9609;
  assign n10528 = n10526 & n10527;
  assign n10529 = n10528 ^ n10521;
  assign n10530 = n10524 & ~n10529;
  assign n10531 = n10530 ^ n10521;
  assign n10532 = n10531 ^ n9650;
  assign n10533 = n10520 & n10532;
  assign n10534 = n10533 ^ n9650;
  assign n10535 = ~n10518 & n10534;
  assign n10536 = n10535 ^ n9673;
  assign n10537 = n10517 & ~n10536;
  assign n10538 = ~n9659 & n10537;
  assign n10539 = n10538 ^ n6628;
  assign n10540 = n10539 ^ x105;
  assign n10541 = n9847 & n9855;
  assign n10542 = n9850 & n9863;
  assign n10543 = n9746 & n9861;
  assign n10544 = ~n10542 & ~n10543;
  assign n10545 = ~n10541 & n10544;
  assign n10546 = ~n9871 & n10545;
  assign n10547 = ~n9887 & ~n9902;
  assign n10548 = n9746 & ~n10547;
  assign n10549 = n9897 & ~n9902;
  assign n10550 = n9863 & ~n10549;
  assign n10551 = ~n9888 & n9907;
  assign n10552 = n9746 & ~n10551;
  assign n10553 = ~n9902 & n10023;
  assign n10554 = ~n9854 & n10553;
  assign n10555 = n9847 & ~n10554;
  assign n10556 = ~n10552 & ~n10555;
  assign n10557 = ~n10550 & n10556;
  assign n10558 = n9894 ^ n9852;
  assign n10559 = n9894 ^ n9746;
  assign n10560 = n10559 ^ n9746;
  assign n10561 = n9843 ^ n9807;
  assign n10562 = n9843 ^ n9805;
  assign n10563 = n10562 ^ n9843;
  assign n10564 = n9843 ^ n9777;
  assign n10565 = n10564 ^ n9843;
  assign n10566 = ~n10563 & ~n10565;
  assign n10567 = n10566 ^ n9843;
  assign n10568 = ~n10561 & n10567;
  assign n10569 = n10568 ^ n9746;
  assign n10570 = ~n10560 & ~n10569;
  assign n10571 = n10570 ^ n9746;
  assign n10572 = n10558 & n10571;
  assign n10573 = n10572 ^ n9852;
  assign n10574 = n10557 & ~n10573;
  assign n10575 = n9904 ^ n9855;
  assign n10576 = n10575 ^ n9855;
  assign n10577 = n9855 ^ n9745;
  assign n10578 = n10577 ^ n9855;
  assign n10579 = ~n10576 & ~n10578;
  assign n10580 = n10579 ^ n9855;
  assign n10581 = ~n9714 & n10580;
  assign n10582 = n10581 ^ n9855;
  assign n10583 = n10574 & ~n10582;
  assign n10584 = ~n10548 & n10583;
  assign n10585 = n9878 & n10584;
  assign n10586 = n10546 & n10585;
  assign n10587 = n9868 & n10586;
  assign n10588 = n10587 ^ n6891;
  assign n10589 = n10588 ^ x115;
  assign n10590 = n10540 & n10589;
  assign n10591 = n10497 & n10590;
  assign n10592 = n10495 & n10496;
  assign n10593 = n10540 & ~n10589;
  assign n10594 = n10592 & n10593;
  assign n10595 = ~n10591 & ~n10594;
  assign n10596 = n10460 & ~n10595;
  assign n10597 = n10459 ^ n10334;
  assign n10598 = ~n10540 & n10589;
  assign n10599 = n10497 & n10598;
  assign n10600 = n10599 ^ n10459;
  assign n10601 = n10600 ^ n10599;
  assign n10602 = n10495 & ~n10496;
  assign n10603 = ~n10540 & ~n10589;
  assign n10604 = n10602 & n10603;
  assign n10605 = n10604 ^ n10599;
  assign n10606 = ~n10601 & n10605;
  assign n10607 = n10606 ^ n10599;
  assign n10608 = n10597 & n10607;
  assign n10609 = ~n10596 & ~n10608;
  assign n10610 = n10334 & n10459;
  assign n10611 = n10592 & n10603;
  assign n10612 = n10610 & n10611;
  assign n10613 = n10590 & n10602;
  assign n10614 = n10460 & n10613;
  assign n10615 = n10497 & n10593;
  assign n10616 = n10610 & n10615;
  assign n10617 = ~n10614 & ~n10616;
  assign n10618 = ~n10612 & n10617;
  assign n10619 = ~n10334 & ~n10459;
  assign n10620 = ~n10495 & ~n10496;
  assign n10621 = n10598 & n10620;
  assign n10622 = n10619 & n10621;
  assign n10623 = n10593 & n10602;
  assign n10624 = n10610 & n10623;
  assign n10625 = ~n10622 & ~n10624;
  assign n10626 = n10590 & n10592;
  assign n10627 = n10460 & n10626;
  assign n10628 = n10598 & n10602;
  assign n10629 = n10593 & n10620;
  assign n10630 = ~n10628 & ~n10629;
  assign n10631 = n10610 & ~n10630;
  assign n10632 = ~n10627 & ~n10631;
  assign n10633 = n10497 & n10603;
  assign n10634 = n10603 & n10620;
  assign n10635 = ~n10628 & ~n10634;
  assign n10636 = ~n10633 & n10635;
  assign n10637 = n10460 & ~n10636;
  assign n10638 = n10334 & ~n10459;
  assign n10639 = n10592 & n10598;
  assign n10640 = ~n10599 & ~n10626;
  assign n10641 = ~n10639 & n10640;
  assign n10642 = n10638 & ~n10641;
  assign n10643 = ~n10591 & ~n10611;
  assign n10644 = n10619 & ~n10643;
  assign n10645 = ~n10642 & ~n10644;
  assign n10646 = n10615 & n10638;
  assign n10647 = ~n10633 & ~n10639;
  assign n10648 = n10619 & ~n10647;
  assign n10649 = ~n10646 & ~n10648;
  assign n10650 = n10645 & n10649;
  assign n10651 = ~n10637 & n10650;
  assign n10652 = n10590 & n10620;
  assign n10655 = ~n10613 & ~n10652;
  assign n10656 = ~n10623 & n10655;
  assign n10653 = ~n10599 & ~n10639;
  assign n10654 = ~n10652 & n10653;
  assign n10657 = n10656 ^ n10654;
  assign n10658 = n10657 ^ n10656;
  assign n10659 = n10656 ^ n10334;
  assign n10660 = n10659 ^ n10656;
  assign n10661 = ~n10658 & n10660;
  assign n10662 = n10661 ^ n10656;
  assign n10663 = n10459 & ~n10662;
  assign n10664 = n10663 ^ n10656;
  assign n10665 = n10651 & n10664;
  assign n10666 = n10632 & n10665;
  assign n10667 = n10625 & n10666;
  assign n10668 = n10618 & n10667;
  assign n10669 = n10609 & n10668;
  assign n10670 = n10669 ^ n7320;
  assign n10671 = n10670 ^ x93;
  assign n10672 = n10494 ^ x114;
  assign n10673 = n9112 ^ x123;
  assign n10674 = ~n10672 & ~n10673;
  assign n10675 = ~n10126 & n10129;
  assign n10676 = n10118 & n10148;
  assign n10677 = ~n10675 & ~n10676;
  assign n10678 = n10129 & n10136;
  assign n10679 = n10102 & n10133;
  assign n10680 = ~n10678 & ~n10679;
  assign n10681 = n10106 & n10137;
  assign n10682 = n10118 & n10152;
  assign n10683 = ~n10681 & ~n10682;
  assign n10684 = n10680 & n10683;
  assign n10685 = n10102 & n10129;
  assign n10686 = n10106 & n10121;
  assign n10687 = ~n10685 & ~n10686;
  assign n10688 = ~n10116 & n10139;
  assign n10689 = n10098 & n10100;
  assign n10690 = ~n10137 & ~n10689;
  assign n10691 = n10118 & ~n10690;
  assign n10692 = ~n10688 & ~n10691;
  assign n10693 = ~n10113 & ~n10139;
  assign n10694 = ~n10099 & ~n10110;
  assign n10695 = n10129 & ~n10694;
  assign n10696 = n10106 & n10115;
  assign n10697 = ~n10127 & ~n10139;
  assign n10698 = n10099 & n10133;
  assign n10699 = ~n10697 & ~n10698;
  assign n10700 = ~n10696 & n10699;
  assign n10701 = ~n10695 & n10700;
  assign n10702 = ~n10693 & n10701;
  assign n10703 = n10692 & n10702;
  assign n10704 = n10687 & n10703;
  assign n10705 = n10684 & n10704;
  assign n10706 = n10677 & n10705;
  assign n10707 = n10144 & n10706;
  assign n10708 = n10707 ^ n7790;
  assign n10709 = n10708 ^ x112;
  assign n10710 = n9322 & n10164;
  assign n10711 = ~n9339 & ~n10710;
  assign n10712 = n9320 & ~n9346;
  assign n10713 = ~n9326 & ~n9343;
  assign n10714 = ~n9331 & n10713;
  assign n10715 = n10164 & ~n10714;
  assign n10716 = n9317 & n9341;
  assign n10717 = n10171 & ~n10716;
  assign n10718 = ~n9344 & n10717;
  assign n10719 = n9336 & ~n10718;
  assign n10720 = n10170 ^ n9365;
  assign n10721 = n10720 ^ n9365;
  assign n10722 = ~n9333 & ~n10166;
  assign n10723 = ~n9342 & n10722;
  assign n10724 = n10723 ^ n9365;
  assign n10725 = n10721 & n10724;
  assign n10726 = n10725 ^ n9365;
  assign n10727 = ~n10719 & n10726;
  assign n10728 = ~n10715 & n10727;
  assign n10729 = ~n10712 & n10728;
  assign n10730 = n9239 ^ n9212;
  assign n10731 = n10730 ^ n9239;
  assign n10732 = n9316 ^ n9239;
  assign n10733 = n10732 ^ n9239;
  assign n10734 = n10731 & ~n10733;
  assign n10735 = n10734 ^ n9239;
  assign n10736 = ~n9278 & n10735;
  assign n10737 = n10736 ^ n9336;
  assign n10738 = n10737 ^ n10736;
  assign n10739 = n10736 ^ n9350;
  assign n10740 = n10739 ^ n10736;
  assign n10741 = ~n10738 & n10740;
  assign n10742 = n10741 ^ n10736;
  assign n10743 = ~n9187 & n10742;
  assign n10744 = n10743 ^ n10736;
  assign n10745 = n10729 & ~n10744;
  assign n10746 = ~n9335 & n10745;
  assign n10747 = n9329 & n10746;
  assign n10748 = n10711 & n10747;
  assign n10749 = n10748 ^ n7830;
  assign n10750 = n10749 ^ x90;
  assign n10751 = n10709 & ~n10750;
  assign n10752 = n10458 ^ x73;
  assign n10753 = n9712 ^ x64;
  assign n10754 = n10752 & n10753;
  assign n10755 = n10751 & n10754;
  assign n10756 = n10674 & n10755;
  assign n10757 = n10752 & ~n10753;
  assign n10758 = n10751 & n10757;
  assign n10759 = n10674 & n10758;
  assign n10760 = ~n10756 & ~n10759;
  assign n10761 = ~n10672 & n10673;
  assign n10762 = n10709 & n10750;
  assign n10763 = ~n10752 & ~n10753;
  assign n10764 = n10762 & n10763;
  assign n10765 = n10761 & n10764;
  assign n10766 = ~n10752 & n10753;
  assign n10767 = n10751 & n10766;
  assign n10768 = n10761 & n10767;
  assign n10769 = ~n10709 & n10750;
  assign n10770 = n10757 & n10769;
  assign n10771 = n10674 & n10770;
  assign n10772 = ~n10768 & ~n10771;
  assign n10773 = ~n10765 & n10772;
  assign n10774 = n10672 & n10673;
  assign n10775 = n10762 & n10766;
  assign n10776 = n10774 & n10775;
  assign n10777 = ~n10709 & ~n10750;
  assign n10778 = n10754 & n10777;
  assign n10779 = ~n10758 & ~n10778;
  assign n10780 = n10761 & ~n10779;
  assign n10781 = ~n10776 & ~n10780;
  assign n10782 = n10672 & ~n10673;
  assign n10783 = n10763 & n10777;
  assign n10784 = ~n10767 & ~n10783;
  assign n10785 = n10782 & ~n10784;
  assign n10786 = n10757 & n10777;
  assign n10787 = n10786 ^ n10672;
  assign n10788 = n10787 ^ n10786;
  assign n10789 = n10766 & n10777;
  assign n10790 = ~n10764 & ~n10789;
  assign n10791 = n10790 ^ n10786;
  assign n10792 = n10788 & ~n10791;
  assign n10793 = n10792 ^ n10786;
  assign n10794 = n10673 & n10793;
  assign n10795 = ~n10785 & ~n10794;
  assign n10796 = n10782 & n10789;
  assign n10797 = n10750 & n10754;
  assign n10798 = ~n10709 & n10797;
  assign n10799 = n10763 & n10769;
  assign n10800 = ~n10775 & ~n10799;
  assign n10801 = ~n10798 & n10800;
  assign n10802 = n10761 & ~n10801;
  assign n10803 = n10757 & n10762;
  assign n10804 = ~n10798 & ~n10803;
  assign n10805 = n10770 & n10782;
  assign n10806 = n10758 & n10774;
  assign n10807 = ~n10805 & ~n10806;
  assign n10808 = n10804 & n10807;
  assign n10809 = ~n10778 & n10808;
  assign n10810 = n10809 ^ n10673;
  assign n10811 = n10810 ^ n10809;
  assign n10812 = n10709 & n10797;
  assign n10813 = n10766 & n10769;
  assign n10814 = n10751 & n10763;
  assign n10815 = ~n10775 & ~n10814;
  assign n10816 = ~n10813 & n10815;
  assign n10817 = ~n10812 & n10816;
  assign n10818 = n10817 ^ n10809;
  assign n10819 = n10818 ^ n10809;
  assign n10820 = ~n10811 & ~n10819;
  assign n10821 = n10820 ^ n10809;
  assign n10822 = ~n10672 & ~n10821;
  assign n10823 = n10822 ^ n10809;
  assign n10824 = ~n10802 & n10823;
  assign n10825 = ~n10796 & n10824;
  assign n10826 = n10795 & n10825;
  assign n10827 = n10673 ^ n10672;
  assign n10828 = n10814 ^ n10799;
  assign n10829 = n10828 ^ n10799;
  assign n10830 = n10799 ^ n10673;
  assign n10831 = n10830 ^ n10799;
  assign n10832 = n10829 & ~n10831;
  assign n10833 = n10832 ^ n10799;
  assign n10834 = n10827 & n10833;
  assign n10835 = n10834 ^ n10799;
  assign n10836 = n10826 & ~n10835;
  assign n10837 = n10781 & n10836;
  assign n10838 = n10773 & n10837;
  assign n10839 = n10760 & n10838;
  assign n10840 = n10839 ^ n9608;
  assign n10841 = n10840 ^ x100;
  assign n10842 = ~n10671 & n10841;
  assign n10843 = n9385 ^ x104;
  assign n10844 = ~n9062 & ~n9079;
  assign n10845 = n9043 & ~n10844;
  assign n10846 = n9059 & ~n9074;
  assign n10847 = n9103 & n10236;
  assign n10848 = ~n9067 & n10847;
  assign n10849 = n8699 & ~n10848;
  assign n10850 = ~n10846 & ~n10849;
  assign n10851 = ~n9060 & n9094;
  assign n10852 = ~n9095 & ~n9096;
  assign n10853 = n9058 & ~n10852;
  assign n10854 = n9064 & ~n10853;
  assign n10855 = n10229 & n10854;
  assign n10856 = n9098 & n10229;
  assign n10857 = ~n9043 & n10244;
  assign n10858 = ~n10856 & ~n10857;
  assign n10859 = ~n9059 & ~n10858;
  assign n10860 = ~n10855 & ~n10859;
  assign n10861 = n10860 ^ n8659;
  assign n10862 = n10860 ^ n8698;
  assign n10863 = n10862 ^ n8698;
  assign n10864 = ~n9070 & n10240;
  assign n10865 = n10864 ^ n8698;
  assign n10866 = ~n10863 & ~n10865;
  assign n10867 = n10866 ^ n8698;
  assign n10868 = n10861 & ~n10867;
  assign n10869 = n10868 ^ n8659;
  assign n10870 = ~n10851 & ~n10869;
  assign n10871 = n10850 & n10870;
  assign n10872 = ~n10845 & n10871;
  assign n10873 = n9053 & n10872;
  assign n10874 = n10873 ^ n8100;
  assign n10875 = n10874 ^ x122;
  assign n10876 = n10843 & ~n10875;
  assign n10877 = n10113 & ~n10152;
  assign n10878 = n10129 & ~n10877;
  assign n10879 = ~n10100 & ~n10108;
  assign n10880 = n10098 & ~n10879;
  assign n10881 = ~n10123 & ~n10880;
  assign n10882 = ~n10131 & n10881;
  assign n10883 = ~n10110 & n10882;
  assign n10884 = ~n10102 & n10883;
  assign n10885 = n10118 & ~n10884;
  assign n10886 = ~n10878 & ~n10885;
  assign n10887 = n10115 & n10139;
  assign n10888 = ~n10121 & ~n10148;
  assign n10889 = n10153 & n10888;
  assign n10890 = n10106 & ~n10889;
  assign n10891 = n10132 ^ n10105;
  assign n10892 = n10891 ^ n10132;
  assign n10893 = n10881 ^ n10132;
  assign n10894 = n10893 ^ n10132;
  assign n10895 = n10892 & ~n10894;
  assign n10896 = n10895 ^ n10132;
  assign n10897 = n10139 & ~n10896;
  assign n10898 = n10897 ^ n10132;
  assign n10899 = n10136 ^ n10105;
  assign n10900 = n10899 ^ n10136;
  assign n10901 = ~n10114 & n10888;
  assign n10902 = ~n10123 & n10901;
  assign n10903 = ~n10137 & n10902;
  assign n10904 = n10903 ^ n10136;
  assign n10905 = ~n10900 & ~n10904;
  assign n10906 = n10905 ^ n10136;
  assign n10907 = ~n10139 & n10906;
  assign n10908 = n10898 & ~n10907;
  assign n10909 = ~n10890 & n10908;
  assign n10910 = ~n10887 & n10909;
  assign n10911 = n10886 & n10910;
  assign n10912 = n10684 & n10911;
  assign n10913 = n10912 ^ n7992;
  assign n10914 = n10913 ^ x99;
  assign n10915 = n10399 & n10408;
  assign n10916 = ~n10442 & ~n10915;
  assign n10917 = n10408 & n10427;
  assign n10918 = ~n10411 & ~n10433;
  assign n10919 = ~n10425 & n10918;
  assign n10920 = n10415 & ~n10919;
  assign n10921 = ~n10917 & ~n10920;
  assign n10922 = n10402 & ~n10443;
  assign n10923 = ~n10410 & ~n10440;
  assign n10924 = ~n10444 & n10923;
  assign n10925 = n10435 & n10924;
  assign n10926 = n10337 & ~n10925;
  assign n10927 = ~n10922 & ~n10926;
  assign n10928 = n10421 & n10441;
  assign n10929 = n10408 & ~n10928;
  assign n10930 = n10394 & n10409;
  assign n10931 = ~n10395 & ~n10930;
  assign n10932 = n10415 & ~n10931;
  assign n10933 = n10412 & ~n10427;
  assign n10934 = n10418 & ~n10933;
  assign n10935 = ~n10932 & ~n10934;
  assign n10936 = ~n10929 & n10935;
  assign n10937 = n10927 & n10936;
  assign n10938 = n10921 & n10937;
  assign n10939 = n10423 & n10938;
  assign n10940 = n10414 & n10939;
  assign n10941 = n10916 & n10940;
  assign n10942 = n10941 ^ n8729;
  assign n10943 = n10942 ^ x72;
  assign n10944 = n9922 ^ x82;
  assign n10945 = n10943 & n10944;
  assign n10946 = n10914 & n10945;
  assign n10947 = n9668 & n9673;
  assign n10948 = n9579 & ~n9640;
  assign n10949 = ~n10947 & ~n10948;
  assign n10950 = ~n9647 & ~n9667;
  assign n10951 = n9650 & ~n10950;
  assign n10952 = ~n9664 & ~n9681;
  assign n10953 = ~n9674 & ~n10952;
  assign n10954 = ~n9577 & ~n9579;
  assign n10955 = n9665 & ~n10954;
  assign n10956 = ~n9633 & n9676;
  assign n10957 = n9635 & ~n10956;
  assign n10958 = ~n10955 & ~n10957;
  assign n10959 = n9579 & ~n9669;
  assign n10967 = ~n9644 & ~n9654;
  assign n10960 = ~n9661 & ~n9690;
  assign n10961 = n9676 & n10960;
  assign n10962 = ~n9673 & n10961;
  assign n10963 = ~n9657 & n10960;
  assign n10964 = ~n9644 & n10963;
  assign n10965 = ~n9650 & n10964;
  assign n10966 = ~n10962 & ~n10965;
  assign n10968 = n10967 ^ n10966;
  assign n10969 = ~n9674 & ~n10968;
  assign n10970 = n10969 ^ n10967;
  assign n10971 = ~n10959 & n10970;
  assign n10972 = n10958 & n10971;
  assign n10973 = n9642 & n10972;
  assign n10974 = ~n10953 & n10973;
  assign n10975 = ~n10951 & n10974;
  assign n10976 = n10949 & n10975;
  assign n10977 = n10976 ^ n8763;
  assign n10978 = n10977 ^ x81;
  assign n10979 = n10914 & n10978;
  assign n10980 = ~n10914 & ~n10978;
  assign n10981 = ~n10979 & ~n10980;
  assign n10982 = ~n10943 & ~n10944;
  assign n10983 = n10981 & n10982;
  assign n10984 = ~n10943 & n10944;
  assign n10985 = ~n10914 & n10984;
  assign n10986 = n10943 & ~n10944;
  assign n10987 = n10978 & n10986;
  assign n10988 = ~n10985 & ~n10987;
  assign n10989 = ~n10983 & n10988;
  assign n10990 = ~n10946 & n10989;
  assign n10991 = n10876 & n10990;
  assign n10992 = ~n10843 & n10875;
  assign n10993 = n10943 ^ n10914;
  assign n10994 = n10993 ^ n10978;
  assign n10995 = n10994 ^ n10943;
  assign n10996 = n10995 ^ n10978;
  assign n10997 = n10996 ^ n10944;
  assign n10998 = n10978 ^ n10943;
  assign n10999 = n10944 ^ n10943;
  assign n11000 = n10999 ^ n10943;
  assign n11001 = ~n10998 & ~n11000;
  assign n11002 = n11001 ^ n10943;
  assign n11003 = ~n10997 & ~n11002;
  assign n11004 = n11003 ^ n10994;
  assign n11005 = n10992 & n11004;
  assign n11006 = ~n10991 & ~n11005;
  assign n11007 = n10843 & n10875;
  assign n11008 = n10945 & n10981;
  assign n11009 = n10914 & ~n10978;
  assign n11010 = n10982 & ~n11009;
  assign n11011 = ~n11008 & ~n11010;
  assign n11012 = n10980 & n10984;
  assign n11013 = ~n10981 & n10986;
  assign n11014 = ~n11012 & ~n11013;
  assign n11015 = n11011 & n11014;
  assign n11016 = n11007 & ~n11015;
  assign n11017 = ~n10843 & ~n10875;
  assign n11018 = ~n10979 & n10984;
  assign n11019 = n10945 & n10980;
  assign n11020 = ~n11018 & ~n11019;
  assign n11021 = ~n10980 & n10986;
  assign n11022 = ~n10914 & n10978;
  assign n11023 = n10982 & n11022;
  assign n11024 = ~n11021 & ~n11023;
  assign n11025 = n11020 & n11024;
  assign n11026 = n11017 & ~n11025;
  assign n11027 = ~n11016 & ~n11026;
  assign n11028 = n11006 & n11027;
  assign n11029 = n11028 ^ n9392;
  assign n11030 = n11029 ^ x70;
  assign n11031 = n8422 ^ n7673;
  assign n11032 = ~n8204 & ~n11031;
  assign n11033 = n8424 ^ n8205;
  assign n11034 = n11033 ^ n8205;
  assign n11035 = n8610 ^ n8205;
  assign n11036 = ~n11034 & n11035;
  assign n11037 = n11036 ^ n8205;
  assign n11038 = ~n11032 & ~n11037;
  assign n11039 = n10006 & ~n11038;
  assign n11040 = n8421 ^ n8204;
  assign n11041 = n8421 ^ n7673;
  assign n11042 = n11041 ^ n7673;
  assign n11043 = n8204 ^ n7918;
  assign n11044 = n11043 ^ n7673;
  assign n11045 = n11044 ^ n7673;
  assign n11046 = ~n11042 & ~n11045;
  assign n11047 = n11046 ^ n7673;
  assign n11048 = n11040 & n11047;
  assign n11049 = n11048 ^ n11043;
  assign n11050 = n10011 & n11049;
  assign n11051 = ~n11039 & ~n11050;
  assign n11052 = ~n7918 & ~n11040;
  assign n11053 = n11052 ^ n8599;
  assign n11054 = ~n8617 & ~n11053;
  assign n11055 = n10009 & n11054;
  assign n11056 = ~n8204 & n8424;
  assign n11057 = n8205 & ~n8424;
  assign n11058 = ~n7918 & ~n8597;
  assign n11059 = ~n11057 & ~n11058;
  assign n11060 = ~n11056 & n11059;
  assign n11061 = n10004 & ~n11060;
  assign n11062 = ~n11055 & ~n11061;
  assign n11063 = n11051 & n11062;
  assign n11064 = n11063 ^ n8029;
  assign n11065 = n11064 ^ x124;
  assign n11066 = n9657 & ~n9674;
  assign n11067 = n9635 & ~n10960;
  assign n11068 = ~n11066 & ~n11067;
  assign n11069 = n9661 & n9673;
  assign n11070 = n9669 & n10964;
  assign n11071 = ~n9664 & n11070;
  assign n11072 = n9579 & ~n11071;
  assign n11073 = n10950 & n10952;
  assign n11074 = ~n9635 & n11073;
  assign n11075 = ~n9633 & ~n9664;
  assign n11076 = n9682 & n11075;
  assign n11077 = ~n9673 & n11076;
  assign n11078 = ~n11074 & ~n11077;
  assign n11079 = ~n9637 & ~n11078;
  assign n11080 = ~n9660 & n11079;
  assign n11081 = n9577 & ~n11080;
  assign n11082 = ~n11072 & ~n11081;
  assign n11085 = ~n9675 & ~n9690;
  assign n11083 = n9677 & ~n9681;
  assign n11084 = ~n9668 & n11083;
  assign n11086 = n11085 ^ n11084;
  assign n11087 = n11085 ^ n9650;
  assign n11088 = n11085 & n11087;
  assign n11089 = n11088 ^ n11085;
  assign n11090 = n11086 & n11089;
  assign n11091 = n11090 ^ n11088;
  assign n11092 = n11091 ^ n11085;
  assign n11093 = n11092 ^ n9650;
  assign n11094 = n11082 & n11093;
  assign n11095 = n11094 ^ n11082;
  assign n11096 = ~n11069 & n11095;
  assign n11097 = n11068 & n11096;
  assign n11098 = n9656 & n11097;
  assign n11099 = n11098 ^ n8494;
  assign n11100 = n11099 ^ x78;
  assign n11101 = n11065 & n11100;
  assign n11102 = ~n10139 & n10148;
  assign n11103 = n10110 & n10133;
  assign n11104 = ~n11102 & ~n11103;
  assign n11105 = n10106 & ~n10116;
  assign n11106 = ~n10103 & n10118;
  assign n11107 = n10122 ^ n10098;
  assign n11108 = n10094 ^ n10060;
  assign n11109 = n11107 & n11108;
  assign n11110 = n11109 ^ n10098;
  assign n11111 = ~n10139 & n11110;
  assign n11112 = ~n10112 & n10141;
  assign n11113 = ~n10121 & n11112;
  assign n11114 = n10129 & ~n11113;
  assign n11115 = ~n11111 & ~n11114;
  assign n11116 = n10152 ^ n10105;
  assign n11117 = n11116 ^ n10152;
  assign n11118 = n10152 ^ n10113;
  assign n11119 = n11118 ^ n10152;
  assign n11120 = ~n11117 & ~n11119;
  assign n11121 = n11120 ^ n10152;
  assign n11122 = n10104 & n11121;
  assign n11123 = n11122 ^ n10152;
  assign n11124 = n11115 & ~n11123;
  assign n11125 = n10683 & n11124;
  assign n11126 = n10677 & n11125;
  assign n11127 = ~n11106 & n11126;
  assign n11128 = ~n11105 & n11127;
  assign n11129 = n11104 & n11128;
  assign n11130 = n10687 & n11129;
  assign n11131 = n10144 & n11130;
  assign n11132 = n11131 ^ n8525;
  assign n11133 = n11132 ^ x100;
  assign n11134 = ~n10439 & n10918;
  assign n11135 = n10415 & ~n11134;
  assign n11136 = ~n10419 & ~n10425;
  assign n11137 = n10408 & ~n11136;
  assign n11138 = ~n10393 & ~n10930;
  assign n11139 = n10412 & n11138;
  assign n11140 = n10337 & ~n11139;
  assign n11141 = n10406 ^ n10336;
  assign n11144 = ~n10402 & n10421;
  assign n11142 = ~n10416 & ~n10427;
  assign n11143 = ~n10410 & n11142;
  assign n11145 = n11144 ^ n11143;
  assign n11146 = n11144 ^ n10335;
  assign n11147 = n11146 ^ n11144;
  assign n11148 = n11145 & n11147;
  assign n11149 = n11148 ^ n11144;
  assign n11150 = n11149 ^ n10406;
  assign n11151 = ~n11141 & ~n11150;
  assign n11152 = n11151 ^ n11148;
  assign n11153 = n11152 ^ n11144;
  assign n11154 = n11153 ^ n10336;
  assign n11155 = ~n10406 & n11154;
  assign n11156 = n11155 ^ n10406;
  assign n11157 = n11156 ^ n10336;
  assign n11158 = ~n11140 & n11157;
  assign n11159 = n10396 & ~n10439;
  assign n11160 = ~n10402 & n11159;
  assign n11161 = n11160 ^ n10335;
  assign n11162 = n11161 ^ n11160;
  assign n11163 = n10403 & n11142;
  assign n11164 = n11163 ^ n11160;
  assign n11165 = ~n11162 & n11164;
  assign n11166 = n11165 ^ n11160;
  assign n11167 = ~n10336 & ~n11166;
  assign n11168 = n11158 & ~n11167;
  assign n11169 = ~n11137 & n11168;
  assign n11170 = ~n11135 & n11169;
  assign n11171 = n10930 ^ n10418;
  assign n11172 = n10418 ^ n10415;
  assign n11173 = n11172 ^ n10415;
  assign n11174 = n10415 ^ n10395;
  assign n11175 = n11173 & ~n11174;
  assign n11176 = n11175 ^ n10415;
  assign n11177 = n11171 & ~n11176;
  assign n11178 = n11177 ^ n10930;
  assign n11179 = n11170 & ~n11178;
  assign n11180 = n10916 & n11179;
  assign n11181 = n11180 ^ n7951;
  assign n11182 = n11181 ^ x75;
  assign n11183 = ~n11133 & ~n11182;
  assign n11184 = ~n9344 & ~n9349;
  assign n11185 = n10164 & ~n11184;
  assign n11186 = n9187 & ~n9360;
  assign n11187 = ~n11185 & ~n11186;
  assign n11188 = ~n9340 & ~n9342;
  assign n11189 = n9336 & ~n11188;
  assign n11190 = ~n9343 & n10171;
  assign n11191 = ~n9322 & n11190;
  assign n11192 = n9320 & ~n11191;
  assign n11193 = ~n11189 & ~n11192;
  assign n11194 = n10713 & ~n10716;
  assign n11195 = n11194 ^ n10170;
  assign n11196 = n11195 ^ n11194;
  assign n11197 = ~n9318 & ~n9359;
  assign n11198 = ~n9333 & n11197;
  assign n11199 = n11198 ^ n11194;
  assign n11200 = n11196 & n11199;
  assign n11201 = n11200 ^ n11194;
  assign n11202 = n11193 & n11201;
  assign n11203 = n11187 & n11202;
  assign n11204 = n10169 & n11203;
  assign n11205 = ~n9382 & n11204;
  assign n11206 = n10711 & n11205;
  assign n11207 = ~n10165 & n11206;
  assign n11208 = n11207 ^ n8851;
  assign n11209 = n11208 ^ x117;
  assign n11210 = ~n9060 & n9079;
  assign n11211 = n8659 & n9063;
  assign n11212 = ~n11210 & ~n11211;
  assign n11213 = ~n9070 & ~n9094;
  assign n11214 = n9043 & ~n11213;
  assign n11215 = ~n9062 & n9083;
  assign n11216 = n8699 & ~n11215;
  assign n11217 = ~n11214 & ~n11216;
  assign n11218 = ~n9041 & n9097;
  assign n11219 = n9059 & ~n11218;
  assign n11220 = n8698 ^ n8659;
  assign n11221 = ~n9089 & n10236;
  assign n11222 = ~n9054 & n11221;
  assign n11223 = n11222 ^ n10247;
  assign n11224 = n10247 ^ n8698;
  assign n11225 = n11224 ^ n10247;
  assign n11226 = n11223 & n11225;
  assign n11227 = n11226 ^ n10247;
  assign n11228 = ~n11220 & ~n11227;
  assign n11229 = ~n11219 & ~n11228;
  assign n11230 = n11217 & n11229;
  assign n11231 = n11212 & n11230;
  assign n11232 = ~n10853 & n11231;
  assign n11233 = n9052 & n11232;
  assign n11234 = ~n10845 & n11233;
  assign n11235 = n10231 & n11234;
  assign n11236 = n9057 & n11235;
  assign n11237 = n11236 ^ n8879;
  assign n11238 = n11237 ^ x102;
  assign n11239 = n11209 & n11238;
  assign n11240 = n11183 & n11239;
  assign n11241 = n11101 & n11240;
  assign n11242 = ~n11065 & n11100;
  assign n11243 = ~n11133 & n11182;
  assign n11244 = n11239 & n11243;
  assign n11245 = n11133 & n11182;
  assign n11246 = n11209 & ~n11238;
  assign n11247 = n11245 & n11246;
  assign n11248 = ~n11244 & ~n11247;
  assign n11249 = n11242 & ~n11248;
  assign n11250 = ~n11241 & ~n11249;
  assign n11251 = ~n11065 & ~n11100;
  assign n11252 = ~n11209 & ~n11238;
  assign n11253 = n11245 & n11252;
  assign n11254 = n11251 & n11253;
  assign n11255 = n11065 & ~n11100;
  assign n11256 = n11183 & n11252;
  assign n11257 = n11133 & ~n11182;
  assign n11258 = n11239 & n11257;
  assign n11259 = ~n11209 & n11238;
  assign n11260 = n11183 & n11259;
  assign n11261 = ~n11258 & ~n11260;
  assign n11262 = ~n11256 & n11261;
  assign n11263 = n11255 & ~n11262;
  assign n11264 = ~n11254 & ~n11263;
  assign n11266 = n11257 & n11259;
  assign n11265 = n11246 & n11257;
  assign n11267 = n11266 ^ n11265;
  assign n11268 = n11267 ^ n11266;
  assign n11269 = n11266 ^ n11065;
  assign n11270 = n11269 ^ n11266;
  assign n11271 = n11268 & n11270;
  assign n11272 = n11271 ^ n11266;
  assign n11273 = n11100 & n11272;
  assign n11274 = n11273 ^ n11266;
  assign n11275 = n11264 & ~n11274;
  assign n11276 = ~n11101 & ~n11251;
  assign n11277 = n11183 & n11246;
  assign n11278 = n11252 & n11257;
  assign n11279 = ~n11277 & ~n11278;
  assign n11280 = ~n11276 & ~n11279;
  assign n11281 = n11243 & n11259;
  assign n11282 = ~n11253 & ~n11281;
  assign n11283 = n11242 & ~n11282;
  assign n11284 = n11239 & n11245;
  assign n11285 = ~n11281 & ~n11284;
  assign n11286 = n11251 & ~n11285;
  assign n11287 = ~n11258 & n11279;
  assign n11288 = ~n11240 & n11287;
  assign n11289 = n11242 & ~n11288;
  assign n11290 = n11245 & n11259;
  assign n11291 = n11243 & n11252;
  assign n11292 = ~n11290 & ~n11291;
  assign n11293 = n11285 & n11292;
  assign n11294 = n11101 & ~n11293;
  assign n11295 = n11243 & n11246;
  assign n11296 = ~n11291 & ~n11295;
  assign n11297 = n11255 & ~n11296;
  assign n11298 = n11248 & ~n11297;
  assign n11299 = ~n11100 & ~n11298;
  assign n11300 = ~n11294 & ~n11299;
  assign n11301 = ~n11289 & n11300;
  assign n11302 = ~n11286 & n11301;
  assign n11303 = ~n11283 & n11302;
  assign n11304 = ~n11280 & n11303;
  assign n11305 = n11275 & n11304;
  assign n11306 = n11250 & n11305;
  assign n11307 = n11306 ^ n9629;
  assign n11308 = n11307 ^ x83;
  assign n11309 = ~n11030 & ~n11308;
  assign n11310 = n10842 & n11309;
  assign n11311 = n10333 & n11310;
  assign n11312 = n10003 & ~n10332;
  assign n11313 = n10671 & n10841;
  assign n11314 = ~n11030 & n11308;
  assign n11315 = n11313 & n11314;
  assign n11316 = n11030 & ~n11308;
  assign n11317 = n11313 & n11316;
  assign n11318 = ~n11315 & ~n11317;
  assign n11319 = n11312 & ~n11318;
  assign n11320 = ~n11311 & ~n11319;
  assign n11321 = ~n10003 & ~n10332;
  assign n11322 = n11030 & n11308;
  assign n11323 = n10842 & n11322;
  assign n11324 = n11321 & n11323;
  assign n11325 = ~n10003 & n10332;
  assign n11326 = ~n11321 & ~n11325;
  assign n11327 = n10842 & n11316;
  assign n11328 = ~n11326 & n11327;
  assign n11329 = ~n10671 & ~n10841;
  assign n11330 = n11322 & n11329;
  assign n11331 = n10333 & n11330;
  assign n11332 = n10671 & ~n10841;
  assign n11333 = n11322 & n11332;
  assign n11334 = n11325 & n11333;
  assign n11335 = ~n11331 & ~n11334;
  assign n11336 = ~n10671 & n11314;
  assign n11337 = ~n10841 & n11336;
  assign n11338 = n11316 & n11329;
  assign n11339 = n11313 & n11322;
  assign n11340 = n11309 & n11332;
  assign n11341 = n11309 & n11313;
  assign n11342 = n11316 & n11332;
  assign n11343 = ~n11341 & ~n11342;
  assign n11344 = ~n11340 & n11343;
  assign n11345 = ~n11339 & n11344;
  assign n11346 = ~n11338 & n11345;
  assign n11347 = ~n11337 & n11346;
  assign n11348 = n10333 & ~n11347;
  assign n11349 = n11314 & n11332;
  assign n11350 = n10841 & n11336;
  assign n11351 = ~n11338 & ~n11350;
  assign n11352 = ~n11317 & n11351;
  assign n11353 = ~n11340 & n11352;
  assign n11354 = ~n11349 & n11353;
  assign n11355 = ~n11333 & n11354;
  assign n11356 = n11321 & ~n11355;
  assign n11357 = n11030 ^ n10671;
  assign n11358 = n11357 ^ n10841;
  assign n11359 = n11308 ^ n10841;
  assign n11360 = n11359 ^ n10841;
  assign n11361 = n10841 ^ n10671;
  assign n11362 = n11361 ^ n10841;
  assign n11363 = n11360 & n11362;
  assign n11364 = n11363 ^ n10841;
  assign n11365 = ~n11358 & ~n11364;
  assign n11366 = n11325 & n11365;
  assign n11367 = ~n11312 & ~n11325;
  assign n11368 = ~n11323 & ~n11330;
  assign n11369 = ~n11367 & ~n11368;
  assign n11370 = ~n11310 & ~n11349;
  assign n11371 = n11343 & n11370;
  assign n11372 = n11312 & ~n11371;
  assign n11373 = ~n11369 & ~n11372;
  assign n11374 = ~n11366 & n11373;
  assign n11375 = ~n11356 & n11374;
  assign n11376 = ~n11348 & n11375;
  assign n11377 = n11335 & n11376;
  assign n11378 = ~n11328 & n11377;
  assign n11379 = ~n11324 & n11378;
  assign n11380 = n11320 & n11379;
  assign n11381 = n11380 ^ n9712;
  assign n11382 = n11381 ^ x81;
  assign n11383 = ~n9936 & ~n9949;
  assign n11384 = n9953 & ~n11383;
  assign n11385 = ~n9926 & ~n9981;
  assign n11386 = ~n9954 & ~n9963;
  assign n11387 = n9924 & ~n11386;
  assign n11388 = ~n9954 & ~n9962;
  assign n11389 = ~n9948 & n9958;
  assign n11390 = n11388 & n11389;
  assign n11391 = n9945 & ~n11390;
  assign n11392 = ~n9961 & n11388;
  assign n11393 = ~n9944 & n11392;
  assign n11394 = n9953 & ~n11393;
  assign n11395 = ~n11391 & ~n11394;
  assign n11396 = ~n9923 & n9975;
  assign n11397 = ~n9934 & ~n9948;
  assign n11398 = ~n9990 & n11397;
  assign n11399 = ~n9926 & ~n11398;
  assign n11400 = ~n11396 & ~n11399;
  assign n11401 = n11395 & n11400;
  assign n11402 = ~n11387 & n11401;
  assign n11403 = ~n11385 & n11402;
  assign n11404 = n9964 ^ n9576;
  assign n11405 = n11404 ^ n9576;
  assign n11406 = n9713 ^ n9576;
  assign n11407 = n11406 ^ n9576;
  assign n11408 = ~n11405 & ~n11407;
  assign n11409 = n11408 ^ n9576;
  assign n11410 = ~n9923 & n11409;
  assign n11411 = n11410 ^ n9576;
  assign n11412 = n11403 & ~n11411;
  assign n11413 = ~n9941 & n11412;
  assign n11414 = ~n11384 & n11413;
  assign n11415 = n11414 ^ n9776;
  assign n11416 = n11415 ^ x96;
  assign n11417 = n10296 & ~n10300;
  assign n11418 = ~n10277 & n10279;
  assign n11419 = ~n11417 & ~n11418;
  assign n11420 = ~n10270 & n10303;
  assign n11421 = n10289 & ~n11420;
  assign n11422 = ~n10309 & ~n10315;
  assign n11423 = n10268 & ~n11422;
  assign n11424 = n10279 & n10315;
  assign n11425 = n10266 & n10268;
  assign n11426 = ~n11424 & ~n11425;
  assign n11427 = n10227 ^ n10190;
  assign n11429 = n11427 ^ n10227;
  assign n11430 = ~n10163 & ~n11429;
  assign n11428 = n10264 & n11427;
  assign n11431 = n11430 ^ n11428;
  assign n11432 = n10049 & n11431;
  assign n11433 = n10286 & ~n10290;
  assign n11434 = n10289 & ~n11433;
  assign n11435 = ~n11432 & ~n11434;
  assign n11436 = n11426 & n11435;
  assign n11437 = n10288 & n11436;
  assign n11438 = ~n11423 & n11437;
  assign n11439 = ~n11421 & n11438;
  assign n11440 = n11419 & n11439;
  assign n11441 = n10296 ^ n10048;
  assign n11442 = n11441 ^ n10296;
  assign n11443 = n10296 ^ n10292;
  assign n11444 = ~n11442 & ~n11443;
  assign n11445 = n11444 ^ n10296;
  assign n11446 = n10300 & n11445;
  assign n11447 = n11440 & ~n11446;
  assign n11448 = ~n10267 & n11447;
  assign n11449 = n11448 ^ n8697;
  assign n11450 = n11449 ^ x122;
  assign n11451 = ~n11416 & ~n11450;
  assign n11452 = n10226 ^ x101;
  assign n11453 = n11132 ^ x110;
  assign n11454 = n11452 & ~n11453;
  assign n11455 = n10337 & ~n10928;
  assign n11456 = n10403 & n11138;
  assign n11457 = ~n10406 & n11456;
  assign n11458 = n10418 & ~n11457;
  assign n11459 = ~n11455 & ~n11458;
  assign n11460 = ~n10419 & n10923;
  assign n11461 = ~n10443 & ~n11460;
  assign n11462 = ~n10416 & n11134;
  assign n11463 = ~n10395 & n11462;
  assign n11464 = n10408 & ~n11463;
  assign n11465 = ~n11461 & ~n11464;
  assign n11466 = n11459 & n11465;
  assign n11467 = n10429 & n11466;
  assign n11468 = n10921 & n11467;
  assign n11469 = ~n10405 & n11468;
  assign n11470 = n11469 ^ n8458;
  assign n11471 = n11470 ^ x77;
  assign n11472 = n10047 ^ x92;
  assign n11473 = n11471 & n11472;
  assign n11474 = n10004 & ~n11049;
  assign n11475 = n10011 & ~n11060;
  assign n11476 = ~n11474 & ~n11475;
  assign n11477 = n10009 & ~n11038;
  assign n11478 = n10006 & ~n11054;
  assign n11479 = ~n11477 & ~n11478;
  assign n11480 = n11476 & n11479;
  assign n11481 = n11480 ^ n8465;
  assign n11482 = n11481 ^ x83;
  assign n11483 = n11099 ^ x70;
  assign n11484 = ~n11482 & ~n11483;
  assign n11485 = n11473 & n11484;
  assign n11486 = n11454 & n11485;
  assign n11487 = n11471 & ~n11472;
  assign n11488 = n11484 & n11487;
  assign n11489 = n11454 & n11488;
  assign n11490 = ~n11452 & ~n11453;
  assign n11491 = n11482 & n11483;
  assign n11492 = n11473 & n11491;
  assign n11493 = ~n11482 & n11483;
  assign n11494 = n11487 & n11493;
  assign n11495 = ~n11492 & ~n11494;
  assign n11496 = n11473 & n11493;
  assign n11497 = ~n11471 & ~n11472;
  assign n11498 = n11491 & n11497;
  assign n11499 = ~n11496 & ~n11498;
  assign n11500 = n11482 & ~n11483;
  assign n11501 = n11473 & n11500;
  assign n11502 = ~n11471 & n11472;
  assign n11503 = n11484 & n11502;
  assign n11504 = n11497 & n11500;
  assign n11505 = ~n11503 & ~n11504;
  assign n11506 = ~n11501 & n11505;
  assign n11507 = n11499 & n11506;
  assign n11508 = n11495 & n11507;
  assign n11509 = n11490 & ~n11508;
  assign n11510 = n11452 & n11453;
  assign n11511 = ~n11488 & n11506;
  assign n11512 = n11510 & ~n11511;
  assign n11513 = n11487 & n11491;
  assign n11514 = ~n11496 & ~n11513;
  assign n11515 = n11510 & ~n11514;
  assign n11516 = n11493 & n11502;
  assign n11517 = n11491 & n11502;
  assign n11518 = ~n11494 & ~n11517;
  assign n11519 = n11500 & n11502;
  assign n11520 = n11484 & n11497;
  assign n11521 = ~n11519 & ~n11520;
  assign n11522 = n11518 & n11521;
  assign n11523 = ~n11516 & n11522;
  assign n11524 = n11454 & ~n11523;
  assign n11525 = ~n11515 & ~n11524;
  assign n11526 = n11453 & n11516;
  assign n11527 = ~n11452 & n11453;
  assign n11528 = ~n11513 & ~n11517;
  assign n11529 = ~n11485 & ~n11488;
  assign n11530 = n11521 & n11529;
  assign n11531 = n11528 & n11530;
  assign n11532 = n11527 & ~n11531;
  assign n11533 = ~n11526 & ~n11532;
  assign n11534 = n11525 & n11533;
  assign n11535 = ~n11512 & n11534;
  assign n11536 = ~n11509 & n11535;
  assign n11537 = n11487 & n11500;
  assign n11538 = n11537 ^ n11453;
  assign n11539 = n11538 ^ n11537;
  assign n11540 = n11493 & n11497;
  assign n11541 = n11540 ^ n11537;
  assign n11542 = ~n11539 & n11541;
  assign n11543 = n11542 ^ n11537;
  assign n11544 = ~n11452 & n11543;
  assign n11545 = n11536 & ~n11544;
  assign n11546 = n11539 & n11541;
  assign n11547 = n11546 ^ n11537;
  assign n11548 = n11452 & n11547;
  assign n11549 = n11545 & ~n11548;
  assign n11550 = ~n11489 & n11549;
  assign n11551 = ~n11486 & n11550;
  assign n11552 = n11551 ^ n9804;
  assign n11553 = n11552 ^ x74;
  assign n11554 = n10913 ^ x67;
  assign n11555 = n11181 ^ x85;
  assign n11556 = n11554 & ~n11555;
  assign n11557 = ~n9393 & n9541;
  assign n11558 = n9510 & n9523;
  assign n11559 = ~n11557 & ~n11558;
  assign n11560 = n9519 & n9527;
  assign n11561 = n9528 & n10205;
  assign n11562 = n9395 & ~n11561;
  assign n11563 = ~n11560 & ~n11562;
  assign n11564 = n9536 & ~n9549;
  assign n11565 = ~n9550 & n11564;
  assign n11566 = n9539 & ~n11565;
  assign n11567 = n9539 & ~n10472;
  assign n11568 = ~n9531 & n9559;
  assign n11569 = n9395 & ~n11568;
  assign n11570 = ~n9507 & n11564;
  assign n11571 = n9510 & ~n11570;
  assign n11572 = ~n11569 & ~n11571;
  assign n11573 = ~n11567 & n11572;
  assign n11574 = n10193 & n11573;
  assign n11575 = ~n10487 & n11574;
  assign n11576 = ~n11566 & n11575;
  assign n11577 = n11563 & n11576;
  assign n11578 = n11559 & n11577;
  assign n11579 = n10195 & n11578;
  assign n11580 = n11579 ^ n8136;
  assign n11581 = n11580 ^ x68;
  assign n11582 = n9847 & ~n9890;
  assign n11583 = n9852 & ~n10023;
  assign n11584 = ~n11582 & ~n11583;
  assign n11585 = ~n9880 & ~n9894;
  assign n11586 = n9863 & ~n11585;
  assign n11587 = ~n9882 & n9904;
  assign n11588 = n9714 & ~n11587;
  assign n11589 = ~n11586 & ~n11588;
  assign n11590 = n9854 ^ n9746;
  assign n11591 = n9854 ^ n9847;
  assign n11592 = n11591 ^ n9847;
  assign n11593 = n9903 ^ n9847;
  assign n11594 = ~n11592 & ~n11593;
  assign n11595 = n11594 ^ n9847;
  assign n11596 = n11590 & n11595;
  assign n11597 = n11596 ^ n9746;
  assign n11598 = n11589 & ~n11597;
  assign n11599 = n11584 & n11598;
  assign n11600 = ~n10548 & n11599;
  assign n11601 = n9885 & n11600;
  assign n11602 = n10546 & n11601;
  assign n11603 = n9868 & n11602;
  assign n11604 = n9859 & n11603;
  assign n11605 = n11604 ^ n8064;
  assign n11606 = n11605 ^ x116;
  assign n11607 = ~n11581 & n11606;
  assign n11608 = n11064 ^ x86;
  assign n11609 = n10874 ^ x109;
  assign n11610 = n11608 & ~n11609;
  assign n11611 = n11607 & n11610;
  assign n11612 = n11556 & n11611;
  assign n11613 = n11554 & n11555;
  assign n11614 = n11581 & n11610;
  assign n11615 = n11606 & n11614;
  assign n11616 = n11613 & n11615;
  assign n11617 = ~n11612 & ~n11616;
  assign n11618 = ~n11554 & ~n11555;
  assign n11619 = n11581 & ~n11608;
  assign n11620 = n11609 & n11619;
  assign n11621 = n11606 & n11620;
  assign n11622 = n11607 & ~n11608;
  assign n11623 = n11609 & n11622;
  assign n11624 = n11608 & n11609;
  assign n11625 = ~n11606 & n11624;
  assign n11626 = n11581 & n11625;
  assign n11627 = ~n11623 & ~n11626;
  assign n11628 = ~n11621 & n11627;
  assign n11629 = n11618 & ~n11628;
  assign n11630 = ~n11554 & n11555;
  assign n11631 = ~n11581 & ~n11606;
  assign n11632 = ~n11608 & ~n11609;
  assign n11633 = n11631 & n11632;
  assign n11634 = n11610 & n11631;
  assign n11635 = ~n11606 & n11614;
  assign n11636 = ~n11634 & ~n11635;
  assign n11637 = n11608 ^ n11581;
  assign n11638 = n11637 ^ n11581;
  assign n11639 = n11606 ^ n11581;
  assign n11640 = n11639 ^ n11581;
  assign n11641 = n11638 & n11640;
  assign n11642 = n11641 ^ n11581;
  assign n11643 = n11609 & n11642;
  assign n11644 = n11636 & ~n11643;
  assign n11645 = ~n11633 & n11644;
  assign n11646 = n11630 & ~n11645;
  assign n11647 = ~n11608 & n11631;
  assign n11648 = n11609 & n11647;
  assign n11649 = ~n11609 & n11619;
  assign n11650 = n11606 & n11649;
  assign n11651 = ~n11611 & ~n11634;
  assign n11652 = ~n11650 & n11651;
  assign n11653 = ~n11648 & n11652;
  assign n11654 = n11618 & ~n11653;
  assign n11655 = n11581 & n11624;
  assign n11656 = n11606 & n11655;
  assign n11657 = ~n11606 & n11620;
  assign n11658 = ~n11648 & ~n11657;
  assign n11659 = ~n11656 & n11658;
  assign n11660 = ~n11581 & n11625;
  assign n11661 = n11607 & n11632;
  assign n11662 = ~n11635 & ~n11661;
  assign n11663 = ~n11660 & n11662;
  assign n11664 = ~n11615 & n11663;
  assign n11665 = n11659 & n11664;
  assign n11666 = n11556 & ~n11665;
  assign n11667 = ~n11654 & ~n11666;
  assign n11672 = ~n11623 & ~n11625;
  assign n11668 = ~n11606 & n11649;
  assign n11669 = ~n11611 & ~n11633;
  assign n11670 = ~n11668 & n11669;
  assign n11671 = ~n11634 & n11670;
  assign n11673 = n11672 ^ n11671;
  assign n11674 = n11672 ^ n11613;
  assign n11675 = n11672 & n11674;
  assign n11676 = n11675 ^ n11672;
  assign n11677 = n11673 & n11676;
  assign n11678 = n11677 ^ n11675;
  assign n11679 = n11678 ^ n11672;
  assign n11680 = n11679 ^ n11613;
  assign n11681 = n11667 & n11680;
  assign n11682 = n11681 ^ n11667;
  assign n11683 = ~n11646 & n11682;
  assign n11684 = ~n11629 & n11683;
  assign n11685 = n11656 ^ n11555;
  assign n11686 = n11685 ^ n11656;
  assign n11687 = n11656 ^ n11650;
  assign n11688 = n11686 & n11687;
  assign n11689 = n11688 ^ n11656;
  assign n11690 = ~n11554 & n11689;
  assign n11691 = n11684 & ~n11690;
  assign n11692 = n11617 & n11691;
  assign n11693 = n11692 ^ n9842;
  assign n11694 = n11693 ^ x113;
  assign n11695 = ~n11553 & ~n11694;
  assign n11696 = n11451 & n11695;
  assign n11697 = n10610 & n10621;
  assign n11698 = n10460 & n10639;
  assign n11699 = n10619 & n10623;
  assign n11700 = ~n11698 & ~n11699;
  assign n11701 = ~n11697 & n11700;
  assign n11702 = ~n10459 & n10604;
  assign n11703 = ~n10615 & n10640;
  assign n11704 = ~n10633 & n11703;
  assign n11705 = n10619 & ~n11704;
  assign n11706 = ~n11702 & ~n11705;
  assign n11707 = ~n10623 & ~n10634;
  assign n11708 = ~n10611 & n10630;
  assign n11709 = n11707 & n11708;
  assign n11710 = n10460 & ~n11709;
  assign n11711 = n10647 & n10655;
  assign n11712 = n10610 & ~n11711;
  assign n11713 = ~n10594 & n10635;
  assign n11714 = n10640 & n11713;
  assign n11715 = ~n10652 & n11714;
  assign n11716 = n10638 & ~n11715;
  assign n11717 = ~n11712 & ~n11716;
  assign n11718 = ~n11710 & n11717;
  assign n11719 = n11706 & n11718;
  assign n11720 = n10617 & n11719;
  assign n11721 = n10625 & n11720;
  assign n11722 = n11701 & n11721;
  assign n11723 = ~n10591 & n11722;
  assign n11724 = n11723 ^ n9744;
  assign n11725 = n11724 ^ x107;
  assign n11726 = n11242 & n11266;
  assign n11727 = ~n11253 & ~n11295;
  assign n11728 = n11255 & ~n11727;
  assign n11729 = ~n11726 & ~n11728;
  assign n11730 = ~n11290 & ~n11295;
  assign n11731 = n11101 & ~n11730;
  assign n11732 = n11255 & ~n11285;
  assign n11733 = n11242 & ~n11261;
  assign n11734 = ~n11732 & ~n11733;
  assign n11735 = ~n11244 & ~n11290;
  assign n11736 = n11251 & ~n11735;
  assign n11747 = ~n11258 & ~n11277;
  assign n11748 = ~n11244 & n11727;
  assign n11749 = n11242 & ~n11748;
  assign n11750 = n11747 & ~n11749;
  assign n11751 = ~n11266 & n11750;
  assign n11752 = ~n11291 & n11751;
  assign n11737 = ~n11260 & ~n11265;
  assign n11738 = ~n11256 & n11737;
  assign n11739 = ~n11251 & n11738;
  assign n11740 = ~n11240 & ~n11265;
  assign n11741 = ~n11291 & n11740;
  assign n11742 = ~n11101 & n11741;
  assign n11743 = ~n11739 & ~n11742;
  assign n11744 = ~n11278 & ~n11743;
  assign n11745 = ~n11247 & n11744;
  assign n11746 = ~n11281 & n11745;
  assign n11753 = n11752 ^ n11746;
  assign n11754 = ~n11276 & n11753;
  assign n11755 = n11754 ^ n11752;
  assign n11756 = ~n11736 & n11755;
  assign n11757 = n11734 & n11756;
  assign n11758 = ~n11731 & n11757;
  assign n11759 = n11729 & n11758;
  assign n11760 = n11759 ^ n8954;
  assign n11761 = n11760 ^ x98;
  assign n11762 = ~n11725 & n11761;
  assign n11763 = n11696 & n11762;
  assign n11764 = n11553 & ~n11694;
  assign n11765 = n11451 & n11764;
  assign n11766 = n11762 & n11765;
  assign n11767 = ~n11725 & ~n11761;
  assign n11768 = n11696 & n11767;
  assign n11769 = ~n11766 & ~n11768;
  assign n11770 = n11725 & ~n11761;
  assign n11771 = ~n11416 & n11450;
  assign n11772 = n11695 & n11771;
  assign n11773 = n11416 & n11450;
  assign n11774 = ~n11553 & n11694;
  assign n11775 = n11773 & n11774;
  assign n11776 = n11764 & n11773;
  assign n11777 = ~n11775 & ~n11776;
  assign n11778 = ~n11772 & n11777;
  assign n11779 = n11770 & ~n11778;
  assign n11780 = n11769 & ~n11779;
  assign n11781 = n11725 & n11761;
  assign n11782 = n11696 & n11781;
  assign n11783 = n11451 & n11774;
  assign n11784 = n11553 & n11694;
  assign n11785 = n11451 & n11784;
  assign n11786 = ~n11783 & ~n11785;
  assign n11787 = ~n11767 & ~n11781;
  assign n11788 = ~n11786 & ~n11787;
  assign n11789 = n11695 & n11773;
  assign n11790 = n11762 & n11789;
  assign n11791 = n11416 & ~n11450;
  assign n11792 = n11774 & n11791;
  assign n11793 = n11770 & n11792;
  assign n11794 = ~n11790 & ~n11793;
  assign n11795 = n11784 & n11791;
  assign n11796 = n11770 & n11795;
  assign n11797 = n11764 & n11771;
  assign n11798 = ~n11775 & ~n11797;
  assign n11799 = n11767 & ~n11798;
  assign n11800 = n11771 & n11784;
  assign n11801 = n11781 & n11800;
  assign n11802 = n11765 & n11770;
  assign n11803 = ~n11801 & ~n11802;
  assign n11804 = ~n11799 & n11803;
  assign n11805 = ~n11796 & n11804;
  assign n11806 = n11771 & n11774;
  assign n11807 = n11762 & n11806;
  assign n11808 = ~n11776 & ~n11806;
  assign n11809 = n11767 & ~n11808;
  assign n11810 = n11773 & n11784;
  assign n11811 = n11762 & n11810;
  assign n11812 = n11695 & n11791;
  assign n11813 = n11770 & n11812;
  assign n11814 = ~n11811 & ~n11813;
  assign n11815 = ~n11809 & n11814;
  assign n11816 = ~n11777 & n11781;
  assign n11817 = ~n11762 & ~n11781;
  assign n11818 = n11797 & ~n11817;
  assign n11819 = ~n11816 & ~n11818;
  assign n11820 = n11815 & n11819;
  assign n11821 = ~n11807 & n11820;
  assign n11822 = n11805 & n11821;
  assign n11823 = n11794 & n11822;
  assign n11824 = ~n11788 & n11823;
  assign n11825 = n11761 ^ n11725;
  assign n11826 = n11800 ^ n11761;
  assign n11827 = n11826 ^ n11800;
  assign n11828 = ~n11792 & ~n11795;
  assign n11829 = n11828 ^ n11800;
  assign n11830 = n11827 & ~n11829;
  assign n11831 = n11830 ^ n11800;
  assign n11832 = n11825 & n11831;
  assign n11833 = n11824 & ~n11832;
  assign n11834 = ~n11782 & n11833;
  assign n11835 = n11812 ^ n11761;
  assign n11836 = n11835 ^ n11812;
  assign n11837 = n11764 & n11791;
  assign n11838 = n11837 ^ n11812;
  assign n11839 = ~n11836 & n11838;
  assign n11840 = n11839 ^ n11812;
  assign n11841 = ~n11825 & n11840;
  assign n11842 = n11834 & ~n11841;
  assign n11843 = n11780 & n11842;
  assign n11844 = ~n11763 & n11843;
  assign n11845 = n11844 ^ n9922;
  assign n11846 = n11845 ^ x107;
  assign n11847 = n11382 & n11846;
  assign n11848 = ~n9923 & n9930;
  assign n11849 = n9925 & n9957;
  assign n11850 = ~n11848 & ~n11849;
  assign n11851 = n9924 & ~n11388;
  assign n11852 = ~n9961 & ~n9963;
  assign n11853 = ~n9926 & ~n11852;
  assign n11854 = n9950 & n9964;
  assign n11855 = ~n9976 & n11854;
  assign n11856 = n9945 & ~n11855;
  assign n11857 = ~n9956 & ~n9975;
  assign n11858 = n9981 & n11857;
  assign n11859 = ~n9961 & n11858;
  assign n11860 = n9953 & ~n11859;
  assign n11861 = ~n9944 & ~n9990;
  assign n11862 = ~n9975 & n11861;
  assign n11863 = ~n9926 & ~n11862;
  assign n11864 = ~n11860 & ~n11863;
  assign n11865 = ~n11856 & n11864;
  assign n11866 = n9942 & n11865;
  assign n11867 = ~n11853 & n11866;
  assign n11868 = ~n11851 & n11867;
  assign n11869 = n11850 & n11868;
  assign n11870 = ~n11384 & n11869;
  assign n11871 = n11870 ^ n9142;
  assign n11872 = n11871 ^ x94;
  assign n11873 = ~n11276 & n11291;
  assign n11874 = ~n11256 & n11747;
  assign n11875 = ~n11265 & n11874;
  assign n11876 = ~n11290 & n11875;
  assign n11877 = n11255 & ~n11876;
  assign n11878 = ~n11873 & ~n11877;
  assign n11879 = n11261 & n11279;
  assign n11880 = n11248 & n11879;
  assign n11881 = ~n11281 & n11880;
  assign n11882 = n11101 & ~n11881;
  assign n11883 = n11287 & n11737;
  assign n11884 = n11251 & ~n11883;
  assign n11885 = ~n11284 & n11727;
  assign n11886 = ~n11240 & n11885;
  assign n11887 = n11242 & ~n11886;
  assign n11888 = ~n11884 & ~n11887;
  assign n11889 = ~n11882 & n11888;
  assign n11890 = n11878 & n11889;
  assign n11891 = ~n11249 & n11890;
  assign n11892 = n11100 ^ n11065;
  assign n11893 = n11244 ^ n11100;
  assign n11894 = n11893 ^ n11244;
  assign n11895 = n11256 ^ n11244;
  assign n11896 = n11894 & n11895;
  assign n11897 = n11896 ^ n11244;
  assign n11898 = n11892 & n11897;
  assign n11899 = n11891 & ~n11898;
  assign n11900 = n11729 & n11899;
  assign n11901 = ~n11286 & n11900;
  assign n11902 = n11901 ^ n9185;
  assign n11903 = n11902 ^ x85;
  assign n11904 = ~n11872 & ~n11903;
  assign n11905 = n11004 & n11017;
  assign n11906 = n10876 & ~n11015;
  assign n11907 = ~n11905 & ~n11906;
  assign n11908 = n11025 ^ n10843;
  assign n11909 = n11908 ^ n11025;
  assign n11910 = n11025 ^ n10990;
  assign n11911 = n11909 & ~n11910;
  assign n11912 = n11911 ^ n11025;
  assign n11913 = n10875 & n11912;
  assign n11914 = n11907 & ~n11913;
  assign n11915 = n11914 ^ n9277;
  assign n11916 = n11915 ^ x67;
  assign n11917 = n10774 & n10814;
  assign n11918 = n10774 & n10813;
  assign n11919 = n10775 & n10782;
  assign n11920 = n10761 & n10770;
  assign n11921 = ~n11919 & ~n11920;
  assign n11922 = ~n11918 & n11921;
  assign n11923 = ~n11917 & n11922;
  assign n11924 = n10774 & n10789;
  assign n11925 = ~n10755 & n10804;
  assign n11926 = n10761 & ~n11925;
  assign n11927 = ~n11924 & ~n11926;
  assign n11928 = ~n10767 & n10790;
  assign n11929 = n10674 & ~n11928;
  assign n11930 = ~n10786 & ~n10812;
  assign n11931 = ~n10827 & ~n11930;
  assign n11932 = ~n10778 & ~n10783;
  assign n11933 = n10761 & ~n11932;
  assign n11934 = ~n11931 & ~n11933;
  assign n11935 = n10753 ^ n10750;
  assign n11936 = n11935 ^ n10753;
  assign n11937 = n10753 ^ n10752;
  assign n11938 = n11937 ^ n10753;
  assign n11939 = n11936 & ~n11938;
  assign n11940 = n11939 ^ n10753;
  assign n11941 = n10752 ^ n10709;
  assign n11942 = n11941 ^ n10750;
  assign n11943 = n11942 ^ n10752;
  assign n11944 = n11943 ^ n10753;
  assign n11945 = n11940 & n11944;
  assign n11946 = n11945 ^ n11941;
  assign n11947 = n10782 & ~n11946;
  assign n11948 = n11934 & ~n11947;
  assign n11949 = ~n10776 & n11948;
  assign n11950 = n10773 & n11949;
  assign n11951 = ~n10756 & n11950;
  assign n11952 = ~n10806 & n11951;
  assign n11953 = ~n11929 & n11952;
  assign n11954 = n11927 & n11953;
  assign n11955 = ~n10835 & n11954;
  assign n11956 = n11923 & n11955;
  assign n11957 = n11956 ^ n9238;
  assign n11958 = n11957 ^ x76;
  assign n11959 = n11916 & ~n11958;
  assign n11960 = ~n10021 & n10281;
  assign n11961 = ~n10293 & ~n11960;
  assign n11962 = ~n10300 & n10309;
  assign n11963 = ~n10021 & n10315;
  assign n11964 = ~n11962 & ~n11963;
  assign n11965 = n10279 & n10294;
  assign n11966 = n10281 & n10289;
  assign n11967 = ~n11965 & ~n11966;
  assign n11968 = n11964 & n11967;
  assign n11969 = ~n10285 & n10300;
  assign n11970 = ~n10273 & n11420;
  assign n11971 = n10268 & ~n11970;
  assign n11972 = n10277 & ~n10301;
  assign n11973 = n10021 & n11972;
  assign n11974 = ~n10275 & ~n10289;
  assign n11975 = n10307 & n11974;
  assign n11976 = ~n10266 & n11975;
  assign n11977 = ~n10300 & ~n11976;
  assign n11978 = ~n10314 & ~n11977;
  assign n11979 = ~n11973 & ~n11978;
  assign n11980 = ~n11971 & ~n11979;
  assign n11981 = ~n11969 & n11980;
  assign n11982 = n11968 & n11981;
  assign n11983 = n11961 & n11982;
  assign n11984 = ~n11446 & n11983;
  assign n11985 = n11984 ^ n9211;
  assign n11986 = n11985 ^ x124;
  assign n11987 = n11618 & n11660;
  assign n11988 = n11613 & n11668;
  assign n11989 = n11556 & ~n11669;
  assign n11990 = ~n11988 & ~n11989;
  assign n11991 = n11618 & n11668;
  assign n11992 = ~n11616 & ~n11991;
  assign n11993 = n11556 & n11668;
  assign n11994 = n11607 & n11624;
  assign n11995 = ~n11648 & ~n11994;
  assign n11996 = n11630 & ~n11995;
  assign n11997 = ~n11993 & ~n11996;
  assign n11998 = n11630 & ~n11664;
  assign n11999 = n11636 & n11995;
  assign n12000 = ~n11623 & n11999;
  assign n12001 = n11618 & ~n12000;
  assign n12002 = ~n11998 & ~n12001;
  assign n12003 = ~n11556 & ~n11630;
  assign n12004 = n11621 & ~n12003;
  assign n12005 = ~n11625 & ~n11657;
  assign n12006 = ~n11615 & n12005;
  assign n12007 = n11556 & ~n12006;
  assign n12008 = ~n11634 & ~n11661;
  assign n12009 = ~n11643 & n12008;
  assign n12010 = n11613 & ~n12009;
  assign n12011 = ~n12007 & ~n12010;
  assign n12012 = ~n12004 & n12011;
  assign n12013 = n12002 & n12012;
  assign n12014 = n11997 & n12013;
  assign n12015 = n11992 & n12014;
  assign n12016 = ~n11690 & n12015;
  assign n12017 = n11990 & n12016;
  assign n12018 = ~n11987 & n12017;
  assign n12019 = n12018 ^ n9315;
  assign n12020 = n12019 ^ x117;
  assign n12021 = ~n11986 & n12020;
  assign n12022 = n11959 & n12021;
  assign n12023 = n11904 & n12022;
  assign n12024 = n11872 & n11903;
  assign n12025 = n11916 & n11958;
  assign n12026 = ~n11986 & ~n12020;
  assign n12027 = n12025 & n12026;
  assign n12028 = n12024 & n12027;
  assign n12029 = ~n12023 & ~n12028;
  assign n12030 = n11904 & n12027;
  assign n12031 = ~n11872 & n11903;
  assign n12032 = n11986 & ~n12020;
  assign n12033 = n11959 & n12032;
  assign n12034 = n12031 & n12033;
  assign n12035 = ~n11916 & n11958;
  assign n12036 = n11986 & n12020;
  assign n12037 = n12035 & n12036;
  assign n12038 = n11959 & n12036;
  assign n12039 = ~n12037 & ~n12038;
  assign n12040 = n11904 & ~n12039;
  assign n12041 = ~n12034 & ~n12040;
  assign n12042 = n11904 & n12033;
  assign n12043 = ~n11916 & ~n11958;
  assign n12044 = n12036 & n12043;
  assign n12045 = n12021 & n12035;
  assign n12046 = ~n12044 & ~n12045;
  assign n12047 = n12024 & ~n12046;
  assign n12048 = ~n12042 & ~n12047;
  assign n12049 = n12024 & n12038;
  assign n12050 = n12021 & n12025;
  assign n12051 = n12021 & n12043;
  assign n12052 = ~n12050 & ~n12051;
  assign n12053 = n12031 & ~n12052;
  assign n12054 = ~n12049 & ~n12053;
  assign n12055 = n12032 & n12043;
  assign n12056 = n12025 & n12032;
  assign n12057 = n12026 & n12043;
  assign n12058 = ~n12056 & ~n12057;
  assign n12059 = ~n12022 & n12058;
  assign n12060 = ~n12055 & n12059;
  assign n12061 = n12024 & ~n12060;
  assign n12062 = n11872 & ~n11903;
  assign n12063 = n12032 & n12035;
  assign n12064 = ~n12038 & ~n12045;
  assign n12065 = ~n12050 & n12064;
  assign n12066 = ~n12055 & n12065;
  assign n12067 = ~n12063 & n12066;
  assign n12068 = n12058 & n12067;
  assign n12069 = ~n12027 & n12068;
  assign n12070 = n12062 & n12069;
  assign n12071 = ~n12061 & ~n12070;
  assign n12072 = n12026 & n12035;
  assign n12073 = ~n12055 & ~n12072;
  assign n12074 = ~n12045 & n12073;
  assign n12075 = n11904 & ~n12074;
  assign n12076 = ~n12063 & n12073;
  assign n12077 = ~n12044 & n12076;
  assign n12078 = ~n12027 & n12077;
  assign n12079 = n12031 & ~n12078;
  assign n12080 = ~n12075 & ~n12079;
  assign n12081 = n12071 & n12080;
  assign n12082 = n12054 & n12081;
  assign n12083 = n12048 & n12082;
  assign n12084 = n12041 & n12083;
  assign n12085 = ~n12030 & n12084;
  assign n12086 = n12029 & n12085;
  assign n12087 = n12086 ^ n9385;
  assign n12088 = n12087 ^ x122;
  assign n12089 = n10670 ^ x106;
  assign n12090 = ~n11498 & ~n11516;
  assign n12091 = n11454 & ~n12090;
  assign n12092 = n11454 & n11503;
  assign n12093 = ~n11494 & n11528;
  assign n12094 = n11510 & ~n12093;
  assign n12095 = ~n12092 & ~n12094;
  assign n12096 = n11454 & n11501;
  assign n12097 = ~n11503 & ~n11537;
  assign n12098 = n11510 & ~n12097;
  assign n12099 = ~n12096 & ~n12098;
  assign n12100 = ~n11513 & ~n11519;
  assign n12101 = n11454 & ~n12100;
  assign n12102 = ~n11485 & ~n11504;
  assign n12103 = n11510 & ~n12102;
  assign n12104 = ~n12101 & ~n12103;
  assign n12105 = n11483 ^ n11471;
  assign n12106 = n12105 ^ n11472;
  assign n12107 = n12106 ^ n11482;
  assign n12108 = n12107 ^ n11483;
  assign n12109 = n12108 ^ n11472;
  assign n12110 = n11483 ^ n11472;
  assign n12111 = n11483 ^ n11482;
  assign n12112 = n12111 ^ n11483;
  assign n12113 = n12110 & n12112;
  assign n12114 = n12113 ^ n11483;
  assign n12115 = ~n12109 & ~n12114;
  assign n12116 = n12115 ^ n12106;
  assign n12117 = n11527 & n12116;
  assign n12118 = ~n11488 & ~n11519;
  assign n12119 = ~n11492 & n12097;
  assign n12120 = n11518 & n12119;
  assign n12121 = n12118 & n12120;
  assign n12122 = ~n11540 & n12121;
  assign n12123 = n11490 & ~n12122;
  assign n12124 = ~n12117 & ~n12123;
  assign n12125 = n12104 & n12124;
  assign n12126 = ~n11548 & n12125;
  assign n12127 = n12099 & n12126;
  assign n12128 = n12095 & n12127;
  assign n12129 = ~n11489 & n12128;
  assign n12130 = ~n12091 & n12129;
  assign n12131 = n12130 ^ n8591;
  assign n12132 = n12131 ^ x88;
  assign n12133 = ~n12089 & ~n12132;
  assign n12134 = n10283 & n10289;
  assign n12135 = ~n10284 & ~n10291;
  assign n12136 = n10279 & ~n12135;
  assign n12137 = ~n12134 & ~n12136;
  assign n12138 = ~n10021 & n10309;
  assign n12139 = ~n10290 & ~n10315;
  assign n12140 = ~n10296 & n12139;
  assign n12141 = n10049 & ~n12140;
  assign n12142 = ~n12138 & ~n12141;
  assign n12143 = ~n10302 & ~n10306;
  assign n12144 = ~n10273 & n12143;
  assign n12145 = ~n10049 & n12144;
  assign n12146 = ~n11974 & ~n12145;
  assign n12147 = ~n10270 & ~n12146;
  assign n12148 = n12147 ^ n10021;
  assign n12149 = n12148 ^ n12147;
  assign n12150 = ~n10301 & n10313;
  assign n12151 = n12150 ^ n12147;
  assign n12152 = n12151 ^ n12147;
  assign n12153 = ~n12149 & ~n12152;
  assign n12154 = n12153 ^ n12147;
  assign n12155 = ~n10048 & ~n12154;
  assign n12156 = n12155 ^ n12147;
  assign n12159 = n10276 & ~n10301;
  assign n12157 = ~n10281 & n12135;
  assign n12158 = ~n10309 & n12157;
  assign n12160 = n12159 ^ n12158;
  assign n12161 = n12159 ^ n10268;
  assign n12162 = n12159 & n12161;
  assign n12163 = n12162 ^ n12159;
  assign n12164 = n12160 & n12163;
  assign n12165 = n12164 ^ n12162;
  assign n12166 = n12165 ^ n12159;
  assign n12167 = n12166 ^ n10268;
  assign n12168 = n12156 & n12167;
  assign n12169 = n12168 ^ n12156;
  assign n12170 = n12142 & n12169;
  assign n12171 = n12137 & n12170;
  assign n12172 = n10298 & n12171;
  assign n12173 = n11961 & n12172;
  assign n12174 = ~n10267 & n12173;
  assign n12175 = n12174 ^ n8420;
  assign n12176 = n12175 ^ x121;
  assign n12213 = n10761 & n10799;
  assign n12214 = ~n10806 & ~n12213;
  assign n12215 = n10755 & n10774;
  assign n12216 = n10782 & n10786;
  assign n12217 = ~n12215 & ~n12216;
  assign n12218 = n10674 & n10803;
  assign n12219 = ~n10764 & ~n10770;
  assign n12220 = n10774 & ~n12219;
  assign n12221 = n10778 & ~n10827;
  assign n12222 = n10790 & n10815;
  assign n12223 = n10674 & ~n12222;
  assign n12224 = ~n12221 & ~n12223;
  assign n12225 = ~n10783 & ~n10813;
  assign n12226 = ~n10812 & n12225;
  assign n12227 = n10761 & ~n12226;
  assign n12228 = ~n10799 & n11925;
  assign n12229 = n10782 & ~n12228;
  assign n12230 = ~n12227 & ~n12229;
  assign n12231 = n12224 & n12230;
  assign n12232 = ~n12220 & n12231;
  assign n12233 = ~n12218 & n12232;
  assign n12234 = n10772 & n12233;
  assign n12235 = ~n10785 & n12234;
  assign n12236 = n12217 & n12235;
  assign n12237 = n11923 & n12236;
  assign n12238 = n10781 & n12237;
  assign n12239 = n12214 & n12238;
  assign n12240 = ~n10756 & n12239;
  assign n12241 = n12240 ^ n7917;
  assign n12242 = n12241 ^ x66;
  assign n12211 = n10002 ^ x112;
  assign n12177 = n11556 & n11648;
  assign n12178 = ~n11611 & ~n11635;
  assign n12179 = n11613 & ~n12178;
  assign n12180 = ~n11623 & ~n11657;
  assign n12181 = ~n11626 & n12180;
  assign n12182 = ~n11656 & n12181;
  assign n12183 = n11556 & ~n12182;
  assign n12184 = ~n11660 & n11995;
  assign n12185 = ~n11621 & n12184;
  assign n12186 = n11613 & ~n12185;
  assign n12187 = ~n12183 & ~n12186;
  assign n12188 = ~n11615 & n12008;
  assign n12189 = n11618 & ~n12188;
  assign n12190 = n11662 & n11669;
  assign n12191 = n11630 & ~n12190;
  assign n12192 = ~n12189 & ~n12191;
  assign n12193 = n12187 & n12192;
  assign n12194 = ~n11629 & n12193;
  assign n12195 = ~n11987 & n12194;
  assign n12196 = ~n12179 & n12195;
  assign n12197 = ~n12177 & n12196;
  assign n12198 = n11650 ^ n11630;
  assign n12199 = n11650 ^ n11556;
  assign n12200 = n12199 ^ n11556;
  assign n12201 = n11659 ^ n11556;
  assign n12202 = ~n12200 & n12201;
  assign n12203 = n12202 ^ n11556;
  assign n12204 = n12198 & n12203;
  assign n12205 = n12204 ^ n11630;
  assign n12206 = n12197 & ~n12205;
  assign n12207 = n11992 & n12206;
  assign n12208 = n11990 & n12207;
  assign n12209 = n12208 ^ n8203;
  assign n12210 = n12209 ^ x65;
  assign n12212 = n12211 ^ n12210;
  assign n12243 = n12242 ^ n12212;
  assign n12244 = n12176 & n12243;
  assign n12245 = ~n12176 & n12210;
  assign n12246 = n12242 & n12245;
  assign n12247 = ~n12176 & ~n12210;
  assign n12248 = n12211 & n12247;
  assign n12249 = ~n12246 & ~n12248;
  assign n12250 = ~n12244 & n12249;
  assign n12251 = n12133 & n12250;
  assign n12252 = n12089 & ~n12132;
  assign n12253 = ~n12176 & ~n12242;
  assign n12254 = ~n12212 & n12253;
  assign n12255 = n12176 & ~n12210;
  assign n12256 = n12255 ^ n12242;
  assign n12257 = n12256 ^ n12255;
  assign n12258 = n12211 ^ n12176;
  assign n12259 = n12258 ^ n12255;
  assign n12260 = n12257 & n12259;
  assign n12261 = n12260 ^ n12255;
  assign n12262 = ~n12254 & ~n12261;
  assign n12263 = n12252 & ~n12262;
  assign n12264 = ~n12251 & ~n12263;
  assign n12265 = ~n12089 & n12132;
  assign n12266 = n12176 & n12210;
  assign n12267 = ~n12211 & n12266;
  assign n12268 = n12242 & n12267;
  assign n12269 = n12253 ^ n12210;
  assign n12270 = n12269 ^ n12253;
  assign n12271 = n12211 & n12242;
  assign n12272 = n12258 & ~n12271;
  assign n12273 = n12272 ^ n12253;
  assign n12274 = ~n12270 & ~n12273;
  assign n12275 = n12274 ^ n12253;
  assign n12276 = ~n12268 & ~n12275;
  assign n12277 = n12265 & n12276;
  assign n12278 = n12089 & n12132;
  assign n12279 = n12242 & n12247;
  assign n12283 = ~n12211 & ~n12266;
  assign n12280 = n12210 ^ n12176;
  assign n12281 = n12211 & n12280;
  assign n12282 = n12281 ^ n12210;
  assign n12284 = n12283 ^ n12282;
  assign n12285 = n12242 & n12284;
  assign n12286 = n12285 ^ n12282;
  assign n12287 = ~n12279 & ~n12286;
  assign n12288 = n12278 & ~n12287;
  assign n12289 = ~n12277 & ~n12288;
  assign n12290 = n12264 & n12289;
  assign n12291 = n12290 ^ n8628;
  assign n12292 = n12291 ^ x104;
  assign n12293 = n10331 ^ x126;
  assign n12294 = n10604 & n10610;
  assign n12295 = n10589 ^ n10495;
  assign n12296 = n10540 ^ n10495;
  assign n12297 = n12296 ^ n10496;
  assign n12298 = n12297 ^ n10589;
  assign n12299 = n12297 ^ n10496;
  assign n12300 = ~n12298 & ~n12299;
  assign n12301 = n12300 ^ n12297;
  assign n12302 = ~n12295 & ~n12301;
  assign n12303 = n12302 ^ n12297;
  assign n12304 = ~n10615 & n12303;
  assign n12305 = n10638 & ~n12304;
  assign n12306 = ~n10604 & ~n10629;
  assign n12307 = n10595 & ~n10599;
  assign n12308 = n12306 & n12307;
  assign n12309 = ~n10639 & n12308;
  assign n12310 = ~n10613 & n12309;
  assign n12311 = n10619 & ~n12310;
  assign n12312 = ~n10613 & ~n10615;
  assign n12313 = n10460 & ~n12312;
  assign n12314 = n10610 ^ n10460;
  assign n12317 = ~n10652 & n11707;
  assign n12315 = ~n10626 & n10647;
  assign n12316 = ~n10652 & n12315;
  assign n12318 = n12317 ^ n12316;
  assign n12319 = n12317 ^ n10610;
  assign n12320 = n12319 ^ n12317;
  assign n12321 = ~n12318 & n12320;
  assign n12322 = n12321 ^ n12317;
  assign n12323 = n12314 & n12322;
  assign n12324 = n12323 ^ n10460;
  assign n12325 = ~n12313 & ~n12324;
  assign n12326 = ~n12311 & n12325;
  assign n12327 = ~n12305 & n12326;
  assign n12328 = ~n12294 & n12327;
  assign n12329 = ~n10608 & n12328;
  assign n12330 = n10632 & n12329;
  assign n12331 = n11701 & n12330;
  assign n12332 = n12331 ^ n9439;
  assign n12333 = n12332 ^ x86;
  assign n12334 = n12293 & n12333;
  assign n12335 = n11871 ^ x84;
  assign n12336 = n11453 & n11501;
  assign n12337 = n11527 & ~n12118;
  assign n12338 = ~n12336 & ~n12337;
  assign n12339 = n11454 & n11540;
  assign n12340 = ~n11496 & n11528;
  assign n12341 = n11490 & ~n12340;
  assign n12342 = ~n12339 & ~n12341;
  assign n12343 = n11510 & n11520;
  assign n12344 = ~n11492 & ~n11517;
  assign n12345 = n11454 & ~n12344;
  assign n12346 = n11499 & n11528;
  assign n12347 = n11510 & ~n12346;
  assign n12348 = ~n12345 & ~n12347;
  assign n12349 = n11505 & n11529;
  assign n12350 = n11490 & ~n12349;
  assign n12351 = n11495 & ~n11516;
  assign n12352 = ~n11540 & n12351;
  assign n12353 = n11527 & ~n12352;
  assign n12354 = ~n12350 & ~n12353;
  assign n12355 = n12348 & n12354;
  assign n12356 = ~n12091 & n12355;
  assign n12357 = ~n12343 & n12356;
  assign n12358 = n12342 & n12357;
  assign n12359 = n12338 & n12358;
  assign n12360 = ~n11544 & n12359;
  assign n12361 = n12099 & n12360;
  assign n12362 = ~n11489 & n12361;
  assign n12363 = ~n11486 & n12362;
  assign n12364 = n12363 ^ n9477;
  assign n12365 = n12364 ^ x101;
  assign n12366 = n12335 & ~n12365;
  assign n12367 = n12334 & n12366;
  assign n12368 = n11029 ^ x108;
  assign n12369 = n12019 ^ x125;
  assign n12370 = ~n12368 & ~n12369;
  assign n12371 = n12367 & n12370;
  assign n12372 = ~n12368 & n12369;
  assign n12373 = ~n12335 & ~n12365;
  assign n12374 = n12334 & n12373;
  assign n12375 = n12293 & ~n12333;
  assign n12376 = n12366 & n12375;
  assign n12377 = ~n12374 & ~n12376;
  assign n12378 = n12372 & ~n12377;
  assign n12379 = ~n12371 & ~n12378;
  assign n12380 = ~n12293 & ~n12333;
  assign n12381 = n12373 & n12380;
  assign n12382 = n12335 & n12365;
  assign n12383 = n12380 & n12382;
  assign n12384 = ~n12381 & ~n12383;
  assign n12385 = n12372 & ~n12384;
  assign n12386 = ~n12335 & n12365;
  assign n12387 = n12334 & n12386;
  assign n12388 = ~n12376 & ~n12387;
  assign n12389 = n12370 & ~n12388;
  assign n12390 = n12368 & n12369;
  assign n12391 = n12334 & n12382;
  assign n12392 = n12375 & n12386;
  assign n12393 = ~n12391 & ~n12392;
  assign n12394 = n12390 & ~n12393;
  assign n12395 = ~n12389 & ~n12394;
  assign n12396 = ~n12385 & n12395;
  assign n12397 = ~n12293 & n12333;
  assign n12398 = n12382 & n12397;
  assign n12399 = n12380 & n12386;
  assign n12400 = ~n12398 & ~n12399;
  assign n12401 = n12372 & ~n12400;
  assign n12402 = n12368 & ~n12369;
  assign n12403 = n12366 & n12397;
  assign n12404 = ~n12381 & ~n12403;
  assign n12405 = n12402 & ~n12404;
  assign n12406 = ~n12401 & ~n12405;
  assign n12407 = n12370 & n12398;
  assign n12408 = n12373 & n12397;
  assign n12409 = n12390 & n12408;
  assign n12410 = ~n12407 & ~n12409;
  assign n12411 = n12370 & n12408;
  assign n12412 = n12383 & n12390;
  assign n12413 = ~n12411 & ~n12412;
  assign n12414 = ~n12372 & ~n12402;
  assign n12415 = n12392 & ~n12414;
  assign n12416 = n12413 & ~n12415;
  assign n12417 = n12369 ^ n12368;
  assign n12418 = n12403 ^ n12369;
  assign n12419 = n12418 ^ n12403;
  assign n12420 = n12366 & n12380;
  assign n12421 = n12420 ^ n12403;
  assign n12422 = ~n12419 & n12421;
  assign n12423 = n12422 ^ n12403;
  assign n12424 = ~n12417 & n12423;
  assign n12425 = n12374 ^ n12372;
  assign n12426 = n12425 ^ n12374;
  assign n12427 = n12386 & n12397;
  assign n12428 = n12427 ^ n12374;
  assign n12429 = n12428 ^ n12374;
  assign n12430 = ~n12426 & n12429;
  assign n12431 = n12430 ^ n12374;
  assign n12432 = ~n12402 & n12431;
  assign n12433 = n12432 ^ n12374;
  assign n12434 = ~n12424 & ~n12433;
  assign n12435 = n12391 & ~n12414;
  assign n12436 = ~n12383 & ~n12427;
  assign n12437 = ~n12367 & n12436;
  assign n12438 = n12402 & ~n12437;
  assign n12439 = ~n12435 & ~n12438;
  assign n12440 = n12373 & n12375;
  assign n12441 = n12440 ^ n12390;
  assign n12442 = n12375 & n12382;
  assign n12443 = n12442 ^ n12440;
  assign n12444 = n12443 ^ n12442;
  assign n12445 = n12442 ^ n12370;
  assign n12446 = n12444 & ~n12445;
  assign n12447 = n12446 ^ n12442;
  assign n12448 = n12441 & ~n12447;
  assign n12449 = n12448 ^ n12390;
  assign n12450 = n12439 & ~n12449;
  assign n12451 = n12434 & n12450;
  assign n12452 = n12416 & n12451;
  assign n12453 = n12410 & n12452;
  assign n12454 = n12406 & n12453;
  assign n12455 = n12396 & n12454;
  assign n12456 = n12379 & n12455;
  assign n12457 = n12456 ^ n9573;
  assign n12458 = n12457 ^ x74;
  assign n12459 = n10945 & n11022;
  assign n12460 = n10945 & n10978;
  assign n12461 = n10981 & n10984;
  assign n12462 = ~n12460 & ~n12461;
  assign n12463 = n10986 ^ n10982;
  assign n12464 = n11022 ^ n10982;
  assign n12465 = n12464 ^ n10982;
  assign n12466 = n12463 & ~n12465;
  assign n12467 = n12466 ^ n10982;
  assign n12468 = n12462 & ~n12467;
  assign n12469 = n11007 & ~n12468;
  assign n12470 = n10986 & n11009;
  assign n12471 = n10984 ^ n10979;
  assign n12472 = n12471 ^ n10984;
  assign n12473 = n10984 ^ n10982;
  assign n12474 = ~n12472 & n12473;
  assign n12475 = n12474 ^ n10984;
  assign n12476 = ~n12470 & ~n12475;
  assign n12477 = ~n10946 & n12476;
  assign n12478 = n10876 & ~n12477;
  assign n12479 = ~n12469 & ~n12478;
  assign n12480 = n10945 & ~n10979;
  assign n12481 = ~n10983 & ~n12480;
  assign n12482 = ~n10981 & n10984;
  assign n12483 = n10986 & n11022;
  assign n12484 = ~n12482 & ~n12483;
  assign n12485 = n12481 & n12484;
  assign n12486 = n10992 & ~n12485;
  assign n12487 = n10914 & n10984;
  assign n12488 = n10978 & n10982;
  assign n12489 = ~n12487 & ~n12488;
  assign n12490 = ~n11013 & n12489;
  assign n12491 = ~n11019 & n12490;
  assign n12492 = n11017 & ~n12491;
  assign n12493 = ~n12486 & ~n12492;
  assign n12494 = n12479 & n12493;
  assign n12495 = ~n12459 & n12494;
  assign n12496 = n12495 ^ n8821;
  assign n12497 = n12496 ^ x80;
  assign n12498 = ~n11555 & n11650;
  assign n12499 = n11556 & n11635;
  assign n12500 = ~n12498 & ~n12499;
  assign n12501 = n11613 & n11633;
  assign n12502 = n11555 ^ n11554;
  assign n12503 = ~n11662 & ~n12502;
  assign n12504 = n11630 & ~n12180;
  assign n12505 = n11618 & ~n12182;
  assign n12506 = ~n11615 & n11652;
  assign n12507 = n11630 & ~n12506;
  assign n12508 = ~n12505 & ~n12507;
  assign n12509 = n11625 ^ n11554;
  assign n12510 = ~n11621 & ~n11656;
  assign n12511 = n12510 ^ n11995;
  assign n12512 = n11995 ^ n11555;
  assign n12513 = n12512 ^ n11995;
  assign n12514 = n12511 & n12513;
  assign n12515 = n12514 ^ n11995;
  assign n12516 = n12515 ^ n11625;
  assign n12517 = ~n12509 & ~n12516;
  assign n12518 = n12517 ^ n12514;
  assign n12519 = n12518 ^ n11995;
  assign n12520 = n12519 ^ n11554;
  assign n12521 = ~n11625 & n12520;
  assign n12522 = n12521 ^ n11625;
  assign n12523 = n12522 ^ n11554;
  assign n12524 = n12508 & n12523;
  assign n12525 = ~n12504 & n12524;
  assign n12526 = ~n12503 & n12525;
  assign n12527 = ~n12501 & n12526;
  assign n12528 = n12500 & n12527;
  assign n12529 = n11997 & n12528;
  assign n12530 = n11617 & n12529;
  assign n12531 = ~n11987 & n12530;
  assign n12532 = n12531 ^ n9039;
  assign n12533 = n12532 ^ x89;
  assign n12534 = n12497 & ~n12533;
  assign n12535 = n10674 & ~n10804;
  assign n12536 = n10790 & ~n10812;
  assign n12537 = ~n10778 & n12536;
  assign n12538 = ~n10755 & n12537;
  assign n12539 = n10761 & ~n12538;
  assign n12540 = ~n12535 & ~n12539;
  assign n12541 = ~n10783 & ~n10797;
  assign n12542 = n10774 & ~n12541;
  assign n12543 = n10779 & n12219;
  assign n12544 = n10782 & ~n12543;
  assign n12545 = ~n10789 & n10800;
  assign n12546 = ~n10786 & n12545;
  assign n12547 = n10674 & ~n12546;
  assign n12548 = ~n12544 & ~n12547;
  assign n12549 = ~n12542 & n12548;
  assign n12550 = n12540 & n12549;
  assign n12551 = n10795 & n12550;
  assign n12552 = n12217 & n12551;
  assign n12553 = n11922 & n12552;
  assign n12554 = n12214 & n12553;
  assign n12555 = n10760 & n12554;
  assign n12556 = n12555 ^ n8993;
  assign n12557 = n12556 ^ x99;
  assign n12558 = n11760 ^ x114;
  assign n12559 = n12557 & ~n12558;
  assign n12560 = n12534 & n12559;
  assign n12561 = ~n11501 & ~n11504;
  assign n12562 = ~n11516 & n12561;
  assign n12563 = n11510 & ~n12562;
  assign n12564 = n11490 & n12116;
  assign n12565 = ~n12563 & ~n12564;
  assign n12566 = n11453 & ~n11521;
  assign n12567 = n11495 & ~n11537;
  assign n12568 = ~n11504 & n12567;
  assign n12569 = n11454 & ~n12568;
  assign n12570 = ~n11498 & n12120;
  assign n12571 = n11527 & ~n12570;
  assign n12572 = ~n12569 & ~n12571;
  assign n12573 = ~n12566 & n12572;
  assign n12574 = n12565 & n12573;
  assign n12575 = n12095 & n12574;
  assign n12576 = ~n11486 & n12575;
  assign n12577 = ~n12091 & n12576;
  assign n12578 = n12577 ^ n8658;
  assign n12579 = n12578 ^ x104;
  assign n12580 = n11449 ^ x82;
  assign n12581 = ~n12579 & n12580;
  assign n12582 = n12497 & n12533;
  assign n12583 = n12557 & n12558;
  assign n12584 = n12582 & n12583;
  assign n12585 = n12581 & n12584;
  assign n12586 = ~n12579 & ~n12580;
  assign n12587 = ~n12557 & n12558;
  assign n12588 = ~n12497 & ~n12533;
  assign n12589 = n12587 & n12588;
  assign n12590 = n12586 & n12589;
  assign n12591 = ~n12585 & ~n12590;
  assign n12592 = n12583 & n12588;
  assign n12593 = ~n12497 & n12533;
  assign n12594 = n12583 & n12593;
  assign n12595 = ~n12557 & ~n12558;
  assign n12596 = n12593 & n12595;
  assign n12597 = ~n12594 & ~n12596;
  assign n12598 = ~n12592 & n12597;
  assign n12599 = n12581 & ~n12598;
  assign n12600 = n12579 & n12580;
  assign n12601 = n12534 & n12595;
  assign n12602 = n12600 & n12601;
  assign n12603 = n12579 & ~n12580;
  assign n12604 = n12587 & n12593;
  assign n12605 = n12559 & n12588;
  assign n12606 = ~n12604 & ~n12605;
  assign n12607 = n12603 & ~n12606;
  assign n12608 = ~n12602 & ~n12607;
  assign n12609 = ~n12599 & n12608;
  assign n12610 = ~n12586 & ~n12600;
  assign n12611 = n12559 & n12593;
  assign n12612 = ~n12610 & n12611;
  assign n12613 = n12534 & n12583;
  assign n12614 = n12534 & n12587;
  assign n12615 = n12559 & n12582;
  assign n12616 = ~n12614 & ~n12615;
  assign n12617 = ~n12613 & n12616;
  assign n12618 = n12597 & n12617;
  assign n12619 = n12603 & ~n12618;
  assign n12620 = ~n12612 & ~n12619;
  assign n12621 = n12588 & n12595;
  assign n12622 = n12582 & n12587;
  assign n12623 = ~n12589 & ~n12622;
  assign n12624 = ~n12621 & n12623;
  assign n12625 = n12581 & ~n12624;
  assign n12626 = n12582 & n12595;
  assign n12627 = ~n12604 & ~n12626;
  assign n12628 = ~n12601 & ~n12613;
  assign n12629 = ~n12615 & n12628;
  assign n12630 = n12627 & n12629;
  assign n12631 = n12586 & ~n12630;
  assign n12632 = ~n12584 & ~n12626;
  assign n12633 = ~n12589 & ~n12605;
  assign n12634 = ~n12592 & n12633;
  assign n12635 = n12632 & n12634;
  assign n12636 = n12600 & ~n12635;
  assign n12637 = ~n12631 & ~n12636;
  assign n12638 = ~n12625 & n12637;
  assign n12639 = n12620 & n12638;
  assign n12640 = n12609 & n12639;
  assign n12641 = n12591 & n12640;
  assign n12642 = ~n12560 & n12641;
  assign n12643 = n12642 ^ n9112;
  assign n12644 = n12643 ^ x113;
  assign n12645 = n12458 & ~n12644;
  assign n12646 = n12292 & n12645;
  assign n12647 = n12088 & n12646;
  assign n12648 = n11847 & n12647;
  assign n12649 = n12088 & ~n12292;
  assign n12650 = n12458 & n12644;
  assign n12651 = n12649 & n12650;
  assign n12652 = n11846 ^ n11382;
  assign n12653 = n12651 & n12652;
  assign n12654 = n12088 & n12292;
  assign n12655 = n12650 & n12654;
  assign n12656 = n11382 & ~n11846;
  assign n12657 = n12655 & n12656;
  assign n12658 = ~n12088 & n12646;
  assign n12659 = n11847 & n12658;
  assign n12660 = ~n12657 & ~n12659;
  assign n12661 = ~n12653 & n12660;
  assign n12662 = ~n11382 & n11846;
  assign n12663 = n12655 & n12662;
  assign n12664 = ~n12458 & n12644;
  assign n12665 = n12649 & n12664;
  assign n12666 = ~n11382 & ~n11846;
  assign n12667 = n12665 & n12666;
  assign n12668 = ~n12088 & ~n12292;
  assign n12669 = ~n12458 & ~n12644;
  assign n12670 = n12668 & n12669;
  assign n12671 = n12649 & n12669;
  assign n12672 = ~n12670 & ~n12671;
  assign n12673 = n12656 & ~n12672;
  assign n12674 = ~n12667 & ~n12673;
  assign n12675 = ~n12663 & n12674;
  assign n12676 = ~n12088 & n12292;
  assign n12677 = n12664 & n12676;
  assign n12678 = n12652 & n12677;
  assign n12679 = n12662 & n12665;
  assign n12680 = ~n12678 & ~n12679;
  assign n12681 = n12654 & n12664;
  assign n12682 = ~n11846 & n12681;
  assign n12683 = n12645 & n12649;
  assign n12684 = ~n12670 & ~n12683;
  assign n12685 = n11847 & ~n12684;
  assign n12686 = n12645 & n12668;
  assign n12687 = n12654 & n12669;
  assign n12688 = ~n12686 & ~n12687;
  assign n12689 = n12656 & ~n12688;
  assign n12690 = n12650 & n12668;
  assign n12691 = n12664 & n12668;
  assign n12692 = ~n12681 & ~n12691;
  assign n12693 = ~n12690 & n12692;
  assign n12694 = ~n12677 & n12693;
  assign n12695 = n11847 & ~n12694;
  assign n12696 = ~n12689 & ~n12695;
  assign n12697 = n12650 & n12676;
  assign n12698 = n12669 & n12676;
  assign n12699 = ~n12671 & ~n12698;
  assign n12700 = ~n12697 & n12699;
  assign n12701 = ~n12686 & n12700;
  assign n12702 = n12662 & ~n12701;
  assign n12703 = ~n12683 & ~n12698;
  assign n12704 = ~n12690 & n12703;
  assign n12705 = ~n12691 & n12704;
  assign n12706 = ~n12646 & n12705;
  assign n12707 = n12666 & ~n12706;
  assign n12708 = ~n12702 & ~n12707;
  assign n12709 = n12696 & n12708;
  assign n12710 = ~n12685 & n12709;
  assign n12711 = ~n12682 & n12710;
  assign n12712 = n12680 & n12711;
  assign n12713 = n12675 & n12712;
  assign n12714 = n12661 & n12713;
  assign n12715 = ~n12648 & n12714;
  assign n12716 = n12715 ^ n10002;
  assign n12717 = n12716 ^ x80;
  assign n12718 = n12241 ^ x123;
  assign n12719 = n11693 ^ x97;
  assign n12720 = n12718 & ~n12719;
  assign n12721 = n10945 & ~n10980;
  assign n12722 = n12476 & ~n12721;
  assign n12723 = n11007 & ~n12722;
  assign n12724 = ~n12459 & n12491;
  assign n12725 = n10992 & ~n12724;
  assign n12726 = ~n12723 & ~n12725;
  assign n12727 = n12468 ^ n10843;
  assign n12728 = n12727 ^ n12468;
  assign n12729 = n12485 ^ n12468;
  assign n12730 = ~n12728 & n12729;
  assign n12731 = n12730 ^ n12468;
  assign n12732 = ~n10875 & n12731;
  assign n12733 = n12726 & ~n12732;
  assign n12734 = n12733 ^ n10059;
  assign n12735 = n12734 ^ x120;
  assign n12736 = n11724 ^ x64;
  assign n12737 = ~n12735 & n12736;
  assign n12738 = n12131 ^ x73;
  assign n12739 = n11276 & ~n11292;
  assign n12740 = n11255 & ~n11879;
  assign n12741 = ~n12739 & ~n12740;
  assign n12742 = ~n11266 & n11737;
  assign n12743 = ~n11240 & n12742;
  assign n12744 = n11251 & ~n12743;
  assign n12745 = ~n11247 & ~n11295;
  assign n12746 = n11251 & ~n12745;
  assign n12747 = ~n11266 & n11279;
  assign n12748 = n11242 & ~n12747;
  assign n12749 = ~n12746 & ~n12748;
  assign n12750 = n11255 & n11284;
  assign n12751 = n11101 & n11261;
  assign n12752 = n11261 ^ n11252;
  assign n12753 = n12751 ^ n11183;
  assign n12754 = n12752 & n12753;
  assign n12755 = n12754 ^ n11183;
  assign n12756 = n12751 & n12755;
  assign n12757 = n12756 ^ n11101;
  assign n12758 = ~n12750 & ~n12757;
  assign n12759 = n12749 & n12758;
  assign n12760 = ~n12744 & n12759;
  assign n12761 = n12741 & n12760;
  assign n12762 = ~n11731 & n12761;
  assign n12763 = ~n11898 & n12762;
  assign n12764 = n11250 & n12763;
  assign n12765 = ~n11286 & n12764;
  assign n12766 = n12765 ^ n10093;
  assign n12767 = n12766 ^ x90;
  assign n12768 = n12738 & n12767;
  assign n12769 = n12737 & n12768;
  assign n12770 = n12738 & ~n12767;
  assign n12771 = n12737 & n12770;
  assign n12772 = ~n12769 & ~n12771;
  assign n12773 = n12720 & ~n12772;
  assign n12774 = n12718 & n12719;
  assign n12775 = n12735 & ~n12736;
  assign n12776 = n12768 & n12775;
  assign n12777 = n12774 & n12776;
  assign n12778 = ~n12718 & ~n12719;
  assign n12779 = n12771 & n12778;
  assign n12780 = ~n12777 & ~n12779;
  assign n12781 = ~n12738 & ~n12767;
  assign n12782 = n12775 & n12781;
  assign n12783 = ~n12735 & ~n12736;
  assign n12784 = n12768 & n12783;
  assign n12785 = ~n12776 & ~n12784;
  assign n12786 = ~n12782 & n12785;
  assign n12787 = n12778 & ~n12786;
  assign n12788 = n12781 & n12783;
  assign n12789 = n12735 & n12736;
  assign n12790 = n12770 & n12789;
  assign n12791 = n12781 & n12789;
  assign n12792 = ~n12790 & ~n12791;
  assign n12793 = ~n12788 & n12792;
  assign n12794 = n12774 & ~n12793;
  assign n12795 = ~n12787 & ~n12794;
  assign n12796 = ~n12718 & n12790;
  assign n12797 = n12770 & n12783;
  assign n12798 = ~n12718 & n12719;
  assign n12799 = ~n12720 & ~n12798;
  assign n12800 = n12797 & ~n12799;
  assign n12801 = ~n12796 & ~n12800;
  assign n12802 = ~n12738 & n12767;
  assign n12803 = n12783 & n12802;
  assign n12804 = n12770 & n12775;
  assign n12805 = ~n12803 & ~n12804;
  assign n12806 = ~n12788 & n12805;
  assign n12807 = n12798 & ~n12806;
  assign n12808 = n12789 & n12802;
  assign n12809 = ~n12782 & ~n12803;
  assign n12810 = ~n12808 & n12809;
  assign n12811 = n12720 & ~n12810;
  assign n12812 = ~n12807 & ~n12811;
  assign n12813 = n12801 & n12812;
  assign n12814 = n12768 & n12789;
  assign n12815 = ~n12791 & ~n12814;
  assign n12816 = n12815 ^ n12799;
  assign n12817 = n12816 ^ n12815;
  assign n12818 = n12775 & n12802;
  assign n12819 = n12737 & n12802;
  assign n12820 = n12737 & n12781;
  assign n12821 = ~n12819 & ~n12820;
  assign n12822 = ~n12818 & n12821;
  assign n12823 = n12822 ^ n12815;
  assign n12824 = n12817 & n12823;
  assign n12825 = n12824 ^ n12815;
  assign n12826 = n12813 & n12825;
  assign n12827 = n12795 & n12826;
  assign n12828 = n12780 & n12827;
  assign n12829 = ~n12773 & n12828;
  assign n12830 = n12769 ^ n12718;
  assign n12831 = n12830 ^ n12769;
  assign n12832 = n12784 ^ n12769;
  assign n12833 = n12831 & n12832;
  assign n12834 = n12833 ^ n12769;
  assign n12835 = n12719 & n12834;
  assign n12836 = n12829 & ~n12835;
  assign n12837 = n12836 ^ n10913;
  assign n12838 = n12837 ^ x102;
  assign n12839 = n12496 ^ x92;
  assign n12840 = n11957 ^ x78;
  assign n12841 = n12839 & ~n12840;
  assign n12842 = n9925 & ~n9950;
  assign n12843 = n9924 & ~n11857;
  assign n12844 = ~n12842 & ~n12843;
  assign n12845 = n9953 & ~n11397;
  assign n12846 = ~n9963 & n11398;
  assign n12847 = n9945 & ~n12846;
  assign n12848 = ~n12845 & ~n12847;
  assign n12849 = n9981 & n11388;
  assign n12850 = n9923 & ~n12849;
  assign n12851 = ~n9576 & ~n9936;
  assign n12852 = ~n9926 & ~n12851;
  assign n12853 = ~n9930 & n9979;
  assign n12854 = ~n9976 & n11392;
  assign n12855 = ~n9925 & n12854;
  assign n12856 = ~n12853 & ~n12855;
  assign n12857 = ~n12852 & ~n12856;
  assign n12858 = ~n12850 & n12857;
  assign n12859 = n12848 & n12858;
  assign n12860 = n12844 & n12859;
  assign n12861 = ~n11384 & n12860;
  assign n12862 = n12861 ^ n10390;
  assign n12863 = n12862 ^ x109;
  assign n12864 = n12578 ^ x116;
  assign n12865 = n12863 & n12864;
  assign n12866 = n10619 & ~n10640;
  assign n12867 = ~n10626 & ~n10633;
  assign n12868 = n10610 & ~n12867;
  assign n12869 = ~n12866 & ~n12868;
  assign n12870 = n10638 & ~n12307;
  assign n12871 = ~n10652 & n12306;
  assign n12872 = n10460 & ~n12871;
  assign n12873 = ~n10613 & ~n10621;
  assign n12874 = ~n10633 & n12873;
  assign n12875 = n10638 & ~n12874;
  assign n12876 = n10635 & n10655;
  assign n12877 = n10610 & ~n12876;
  assign n12878 = n10630 & ~n10652;
  assign n12879 = n10619 & ~n12878;
  assign n12880 = ~n12877 & ~n12879;
  assign n12881 = ~n12875 & n12880;
  assign n12882 = n10609 & n12881;
  assign n12883 = n11700 & n12882;
  assign n12884 = ~n12872 & n12883;
  assign n12885 = ~n12870 & n12884;
  assign n12886 = n12869 & n12885;
  assign n12887 = n10618 & n12886;
  assign n12888 = n10649 & n12887;
  assign n12889 = n12888 ^ n10356;
  assign n12890 = n12889 ^ x91;
  assign n12891 = n11902 ^ x110;
  assign n12892 = ~n12890 & n12891;
  assign n12893 = n12865 & n12892;
  assign n12894 = n12863 & ~n12864;
  assign n12895 = n12890 & n12891;
  assign n12896 = n12894 & n12895;
  assign n12897 = ~n12863 & ~n12864;
  assign n12898 = n12892 & n12897;
  assign n12899 = ~n12896 & ~n12898;
  assign n12900 = ~n12893 & n12899;
  assign n12901 = n12841 & ~n12900;
  assign n12902 = n12839 & n12840;
  assign n12903 = n12890 & ~n12891;
  assign n12904 = n12894 & n12903;
  assign n12905 = n12902 & n12904;
  assign n12906 = ~n12839 & ~n12840;
  assign n12907 = ~n12863 & n12864;
  assign n12908 = n12903 & n12907;
  assign n12909 = ~n12890 & ~n12891;
  assign n12910 = n12907 & n12909;
  assign n12911 = ~n12904 & ~n12910;
  assign n12912 = ~n12908 & n12911;
  assign n12913 = n12906 & ~n12912;
  assign n12914 = ~n12905 & ~n12913;
  assign n12915 = ~n12901 & n12914;
  assign n12916 = n12897 & n12903;
  assign n12917 = n12902 & n12916;
  assign n12918 = ~n12839 & n12840;
  assign n12919 = n12865 & n12909;
  assign n12920 = n12894 & n12909;
  assign n12921 = ~n12919 & ~n12920;
  assign n12922 = n12918 & ~n12921;
  assign n12923 = ~n12917 & ~n12922;
  assign n12924 = n12865 & n12895;
  assign n12925 = n12841 & n12924;
  assign n12926 = n12865 & n12903;
  assign n12927 = n12840 & n12926;
  assign n12928 = n12898 & n12918;
  assign n12929 = n12841 & ~n12911;
  assign n12930 = ~n12928 & ~n12929;
  assign n12931 = n12895 & n12897;
  assign n12932 = ~n12919 & ~n12931;
  assign n12933 = n12841 & ~n12932;
  assign n12934 = n12892 & n12907;
  assign n12935 = n12892 & n12894;
  assign n12936 = ~n12934 & ~n12935;
  assign n12937 = n12895 & n12907;
  assign n12938 = ~n12920 & ~n12937;
  assign n12939 = n12936 & n12938;
  assign n12940 = n12902 & ~n12939;
  assign n12941 = ~n12933 & ~n12940;
  assign n12942 = n12897 & n12909;
  assign n12943 = n12942 ^ n12839;
  assign n12944 = n12942 ^ n12840;
  assign n12945 = n12944 ^ n12840;
  assign n12946 = ~n12893 & ~n12937;
  assign n12947 = ~n12931 & n12946;
  assign n12948 = ~n12906 & n12947;
  assign n12949 = ~n12924 & ~n12931;
  assign n12950 = n12918 & ~n12946;
  assign n12951 = n12949 & ~n12950;
  assign n12952 = n12936 & n12951;
  assign n12953 = ~n12948 & ~n12952;
  assign n12954 = n12953 ^ n12840;
  assign n12955 = ~n12945 & ~n12954;
  assign n12956 = n12955 ^ n12840;
  assign n12957 = ~n12943 & n12956;
  assign n12958 = n12957 ^ n12839;
  assign n12959 = n12941 & n12958;
  assign n12960 = n12930 & n12959;
  assign n12961 = ~n12927 & n12960;
  assign n12962 = ~n12925 & n12961;
  assign n12963 = n12923 & n12962;
  assign n12964 = n12915 & n12963;
  assign n12965 = n12964 ^ n11181;
  assign n12966 = n12965 ^ x116;
  assign n12967 = n12838 & n12966;
  assign n12968 = n12132 ^ n12089;
  assign n12969 = ~n12242 & n12255;
  assign n12970 = n12211 & n12266;
  assign n12971 = ~n12176 & ~n12243;
  assign n12972 = ~n12970 & ~n12971;
  assign n12973 = ~n12969 & n12972;
  assign n12974 = n12973 ^ n12132;
  assign n12975 = n12974 ^ n12973;
  assign n12976 = n12258 ^ n12211;
  assign n12977 = n12242 ^ n12210;
  assign n12978 = n12977 ^ n12211;
  assign n12979 = n12978 ^ n12211;
  assign n12980 = n12976 & n12979;
  assign n12981 = n12980 ^ n12211;
  assign n12982 = n12280 & ~n12981;
  assign n12983 = n12982 ^ n12977;
  assign n12984 = n12983 ^ n12973;
  assign n12985 = ~n12975 & n12984;
  assign n12986 = n12985 ^ n12973;
  assign n12987 = ~n12968 & ~n12986;
  assign n12988 = n12242 & n12255;
  assign n12989 = n12247 & ~n12271;
  assign n12990 = ~n12988 & ~n12989;
  assign n12991 = n12245 ^ n12242;
  assign n12992 = n12991 ^ n12245;
  assign n12993 = n12266 ^ n12245;
  assign n12994 = n12993 ^ n12245;
  assign n12995 = ~n12992 & n12994;
  assign n12996 = n12995 ^ n12245;
  assign n12997 = ~n12211 & n12996;
  assign n12998 = n12997 ^ n12245;
  assign n12999 = n12990 & ~n12998;
  assign n13000 = n12999 ^ n12132;
  assign n13001 = n13000 ^ n12999;
  assign n13002 = n12176 & n12212;
  assign n13003 = ~n12247 & ~n13002;
  assign n13004 = n13003 ^ n12258;
  assign n13005 = ~n12242 & n13004;
  assign n13006 = n13005 ^ n12258;
  assign n13007 = n13006 ^ n12999;
  assign n13008 = n13001 & ~n13007;
  assign n13009 = n13008 ^ n12999;
  assign n13010 = n12968 & ~n13009;
  assign n13011 = ~n12987 & ~n13010;
  assign n13012 = n13011 ^ n11064;
  assign n13013 = n13012 ^ x117;
  assign n13014 = n11770 & n11776;
  assign n13015 = ~n11782 & ~n13014;
  assign n13016 = ~n11785 & ~n11795;
  assign n13017 = n11762 & ~n13016;
  assign n13018 = n11770 & n11810;
  assign n13019 = n11767 & n11800;
  assign n13020 = ~n13018 & ~n13019;
  assign n13021 = n11762 & n11837;
  assign n13022 = ~n11785 & ~n11812;
  assign n13023 = ~n11772 & n13022;
  assign n13024 = n11767 & ~n13023;
  assign n13025 = ~n11783 & ~n11789;
  assign n13026 = n11770 & ~n13025;
  assign n13027 = ~n11807 & ~n13026;
  assign n13028 = ~n11696 & ~n11800;
  assign n13029 = n11770 & ~n13028;
  assign n13030 = n11762 & ~n11777;
  assign n13031 = ~n13029 & ~n13030;
  assign n13032 = n11794 & n13031;
  assign n13033 = n11804 & n13032;
  assign n13034 = n13027 & n13033;
  assign n13035 = ~n13024 & n13034;
  assign n13036 = ~n13021 & n13035;
  assign n13037 = n11792 ^ n11781;
  assign n13038 = n11781 ^ n11767;
  assign n13039 = n13038 ^ n11767;
  assign n13040 = ~n11783 & ~n11837;
  assign n13041 = n11808 & n13040;
  assign n13042 = ~n11789 & n13041;
  assign n13043 = n13042 ^ n11767;
  assign n13044 = n13039 & n13043;
  assign n13045 = n13044 ^ n11767;
  assign n13046 = n13037 & ~n13045;
  assign n13047 = n13046 ^ n11792;
  assign n13048 = n13036 & ~n13047;
  assign n13049 = n11769 & n13048;
  assign n13050 = n13020 & n13049;
  assign n13051 = ~n13017 & n13050;
  assign n13052 = n13015 & n13051;
  assign n13053 = n13052 ^ n11605;
  assign n13054 = n13053 ^ x84;
  assign n13055 = ~n13013 & n13054;
  assign n13056 = n12399 & n12402;
  assign n13057 = n12372 & n12408;
  assign n13058 = ~n12384 & n12414;
  assign n13059 = ~n13057 & ~n13058;
  assign n13060 = ~n13056 & n13059;
  assign n13061 = n12370 & n12374;
  assign n13062 = ~n12368 & n12442;
  assign n13063 = ~n12387 & ~n12403;
  assign n13064 = n12372 & ~n13063;
  assign n13065 = ~n13062 & ~n13064;
  assign n13066 = ~n13061 & n13065;
  assign n13067 = ~n12387 & ~n12420;
  assign n13068 = ~n12367 & n13067;
  assign n13069 = n12390 & ~n13068;
  assign n13070 = ~n12398 & ~n12427;
  assign n13071 = ~n12403 & n13070;
  assign n13072 = n12377 & n13071;
  assign n13073 = ~n12392 & n13072;
  assign n13074 = ~n12440 & n13073;
  assign n13075 = n12402 & ~n13074;
  assign n13076 = ~n13069 & ~n13075;
  assign n13077 = n13066 & n13076;
  assign n13078 = n12410 & n13077;
  assign n13079 = n13060 & n13078;
  assign n13080 = n12396 & n13079;
  assign n13081 = n12379 & n13080;
  assign n13082 = n13081 ^ n11580;
  assign n13083 = n13082 ^ x67;
  assign n13084 = n12592 & n12603;
  assign n13085 = ~n12611 & n12634;
  assign n13086 = n12586 & ~n13085;
  assign n13087 = ~n12594 & ~n12621;
  assign n13088 = ~n12605 & n13087;
  assign n13089 = ~n12622 & n13088;
  assign n13090 = n12600 & ~n13089;
  assign n13091 = n12610 & n12629;
  assign n13092 = ~n12584 & n13091;
  assign n13093 = n12580 ^ n12579;
  assign n13096 = ~n12584 & ~n12615;
  assign n13094 = ~n12622 & n12632;
  assign n13095 = ~n12560 & n13094;
  assign n13097 = n13096 ^ n13095;
  assign n13098 = n13096 ^ n12580;
  assign n13099 = n13098 ^ n13096;
  assign n13100 = ~n13097 & ~n13099;
  assign n13101 = n13100 ^ n13096;
  assign n13102 = ~n13093 & n13101;
  assign n13103 = n13102 ^ n12579;
  assign n13104 = ~n13092 & n13103;
  assign n13105 = ~n13090 & ~n13104;
  assign n13106 = ~n13086 & n13105;
  assign n13107 = ~n13084 & n13106;
  assign n13108 = n12617 & ~n12626;
  assign n13109 = ~n12560 & n13108;
  assign n13110 = n13109 ^ n12589;
  assign n13111 = n13110 ^ n12589;
  assign n13112 = n12589 ^ n12580;
  assign n13113 = n13112 ^ n12589;
  assign n13114 = ~n13111 & n13113;
  assign n13115 = n13114 ^ n12589;
  assign n13116 = ~n12579 & n13115;
  assign n13117 = n13116 ^ n12589;
  assign n13118 = n13107 & ~n13117;
  assign n13119 = n12609 & n13118;
  assign n13120 = n13119 ^ n10874;
  assign n13121 = n13120 ^ x77;
  assign n13122 = ~n13083 & ~n13121;
  assign n13123 = n13055 & n13122;
  assign n13124 = n12967 & n13123;
  assign n13125 = ~n12838 & n12966;
  assign n13126 = n13013 & n13054;
  assign n13127 = n13122 & n13126;
  assign n13128 = n13125 & n13127;
  assign n13129 = ~n13124 & ~n13128;
  assign n13130 = ~n13013 & ~n13054;
  assign n13131 = ~n13083 & n13121;
  assign n13132 = n13130 & n13131;
  assign n13133 = n13126 & n13131;
  assign n13134 = ~n13132 & ~n13133;
  assign n13135 = n12967 & ~n13134;
  assign n13136 = n12838 & ~n12966;
  assign n13137 = n13083 & ~n13121;
  assign n13138 = n13055 & n13137;
  assign n13139 = n13013 & ~n13054;
  assign n13140 = n13137 & n13139;
  assign n13141 = n13122 & n13130;
  assign n13142 = ~n13140 & ~n13141;
  assign n13143 = ~n13138 & n13142;
  assign n13144 = ~n13127 & n13143;
  assign n13145 = n13136 & ~n13144;
  assign n13146 = ~n13135 & ~n13145;
  assign n13147 = n13083 & n13121;
  assign n13148 = n13130 & n13147;
  assign n13149 = ~n12838 & ~n12966;
  assign n13150 = ~n12967 & ~n13149;
  assign n13151 = n13148 & ~n13150;
  assign n13152 = n13130 & n13137;
  assign n13153 = n13126 & n13137;
  assign n13154 = ~n13123 & ~n13153;
  assign n13155 = ~n13152 & n13154;
  assign n13156 = n13149 & ~n13155;
  assign n13157 = n13131 & n13139;
  assign n13158 = n13136 & n13157;
  assign n13159 = n12967 & n13152;
  assign n13160 = ~n13134 & n13149;
  assign n13161 = ~n13159 & ~n13160;
  assign n13162 = n13139 & n13147;
  assign n13163 = n13136 & n13162;
  assign n13164 = n13122 & n13139;
  assign n13165 = ~n13138 & ~n13164;
  assign n13166 = n12967 & ~n13165;
  assign n13167 = ~n13163 & ~n13166;
  assign n13168 = n13153 ^ n13125;
  assign n13169 = n13153 ^ n12967;
  assign n13170 = n13169 ^ n12967;
  assign n13171 = ~n13141 & ~n13164;
  assign n13172 = n13171 ^ n12967;
  assign n13173 = ~n13170 & n13172;
  assign n13174 = n13173 ^ n12967;
  assign n13175 = n13168 & n13174;
  assign n13176 = n13175 ^ n13125;
  assign n13178 = n13055 & n13147;
  assign n13188 = ~n13157 & ~n13178;
  assign n13177 = n13055 & n13131;
  assign n13179 = ~n13177 & ~n13178;
  assign n13180 = ~n13125 & n13179;
  assign n13181 = n13136 & n13178;
  assign n13182 = n13126 & n13147;
  assign n13183 = ~n13148 & ~n13182;
  assign n13184 = ~n13177 & n13183;
  assign n13185 = ~n13181 & n13184;
  assign n13186 = ~n13162 & n13185;
  assign n13187 = ~n13180 & ~n13186;
  assign n13189 = n13188 ^ n13187;
  assign n13190 = n13189 ^ n13188;
  assign n13191 = n13188 ^ n12967;
  assign n13192 = n13191 ^ n13188;
  assign n13193 = n13190 & ~n13192;
  assign n13194 = n13193 ^ n13188;
  assign n13195 = ~n13149 & ~n13194;
  assign n13196 = n13195 ^ n13188;
  assign n13197 = ~n13176 & n13196;
  assign n13198 = n13167 & n13197;
  assign n13199 = n13161 & n13198;
  assign n13200 = ~n13158 & n13199;
  assign n13201 = ~n13156 & n13200;
  assign n13202 = ~n13151 & n13201;
  assign n13203 = n13146 & n13202;
  assign n13204 = n13129 & n13203;
  assign n13205 = n13204 ^ n12209;
  assign n13206 = n13205 ^ x98;
  assign n13207 = ~n12717 & n13206;
  assign n13208 = ~n12839 & n12919;
  assign n13209 = ~n12910 & ~n12916;
  assign n13210 = n12840 & ~n13209;
  assign n13211 = ~n13208 & ~n13210;
  assign n13212 = n12918 & n12942;
  assign n13213 = ~n12896 & n12936;
  assign n13214 = ~n12908 & n13213;
  assign n13215 = n12902 & ~n13214;
  assign n13216 = ~n12935 & n12949;
  assign n13217 = ~n12937 & n13216;
  assign n13218 = n12918 & ~n13217;
  assign n13219 = ~n12916 & ~n12926;
  assign n13220 = n12938 & n13219;
  assign n13221 = ~n12919 & n13220;
  assign n13222 = n12841 & ~n13221;
  assign n13223 = ~n13218 & ~n13222;
  assign n13224 = n12924 ^ n12906;
  assign n13225 = n12924 ^ n12902;
  assign n13226 = n13225 ^ n12902;
  assign n13227 = n12902 ^ n12900;
  assign n13228 = ~n13226 & n13227;
  assign n13229 = n13228 ^ n12902;
  assign n13230 = n13224 & n13229;
  assign n13231 = n13230 ^ n12906;
  assign n13232 = n13223 & ~n13231;
  assign n13233 = ~n13215 & n13232;
  assign n13234 = ~n13212 & n13233;
  assign n13235 = n13211 & n13234;
  assign n13236 = n12915 & n13235;
  assign n13237 = n13236 ^ n10458;
  assign n13238 = n13237 ^ x106;
  assign n13239 = n11381 ^ x97;
  assign n13240 = ~n13238 & n13239;
  assign n13241 = n12025 & n12036;
  assign n13242 = ~n12051 & ~n13241;
  assign n13243 = n11904 & ~n13242;
  assign n13244 = ~n12031 & ~n12062;
  assign n13245 = n11959 & n12026;
  assign n13246 = ~n12072 & ~n13245;
  assign n13247 = ~n12056 & n13246;
  assign n13248 = ~n13244 & ~n13247;
  assign n13249 = ~n13243 & ~n13248;
  assign n13250 = n11872 & n12033;
  assign n13251 = n12031 & ~n12066;
  assign n13252 = ~n13250 & ~n13251;
  assign n13253 = ~n12057 & ~n12063;
  assign n13254 = n13244 & ~n13253;
  assign n13255 = n12046 & ~n12050;
  assign n13256 = ~n12055 & n13255;
  assign n13257 = n12062 & ~n13256;
  assign n13258 = n11958 ^ n11916;
  assign n13259 = n13258 ^ n11916;
  assign n13260 = n11986 ^ n11916;
  assign n13261 = n13260 ^ n11916;
  assign n13262 = ~n13259 & n13261;
  assign n13263 = n13262 ^ n11916;
  assign n13264 = n12020 & n13263;
  assign n13265 = n12024 & n13264;
  assign n13266 = ~n13257 & ~n13265;
  assign n13267 = ~n13254 & n13266;
  assign n13268 = n13252 & n13267;
  assign n13269 = n13249 & n13268;
  assign n13270 = n12041 & n13269;
  assign n13271 = ~n12030 & n13270;
  assign n13272 = n12029 & n13271;
  assign n13273 = n13272 ^ n10749;
  assign n13274 = n13273 ^ x123;
  assign n13275 = n12720 & n12769;
  assign n13276 = ~n12814 & ~n12819;
  assign n13277 = n12778 & ~n13276;
  assign n13278 = ~n13275 & ~n13277;
  assign n13279 = n12720 & n12818;
  assign n13280 = ~n12771 & ~n12791;
  assign n13281 = n12774 & ~n13280;
  assign n13282 = ~n13279 & ~n13281;
  assign n13283 = ~n12800 & n13282;
  assign n13284 = n12778 & n12818;
  assign n13285 = n12782 & ~n12799;
  assign n13286 = ~n13284 & ~n13285;
  assign n13287 = n12774 & n12818;
  assign n13288 = n12798 & n12808;
  assign n13289 = ~n13287 & ~n13288;
  assign n13290 = ~n12718 & n12788;
  assign n13291 = ~n12804 & ~n12808;
  assign n13292 = ~n12784 & n13291;
  assign n13293 = n12778 & ~n13292;
  assign n13294 = ~n13290 & ~n13293;
  assign n13295 = ~n12790 & n13276;
  assign n13296 = ~n12784 & n13295;
  assign n13297 = ~n12799 & ~n13296;
  assign n13298 = n12805 & ~n12820;
  assign n13299 = ~n12769 & n13298;
  assign n13300 = n12774 & ~n13299;
  assign n13301 = ~n13297 & ~n13300;
  assign n13302 = n13294 & n13301;
  assign n13303 = n12780 & n13302;
  assign n13304 = n13289 & n13303;
  assign n13305 = n13286 & n13304;
  assign n13306 = n13283 & n13305;
  assign n13307 = n13278 & n13306;
  assign n13308 = n13307 ^ n10708;
  assign n13309 = n13308 ^ x80;
  assign n13310 = ~n13274 & n13309;
  assign n13311 = n12398 & n12402;
  assign n13312 = n12414 & n12420;
  assign n13313 = ~n13311 & ~n13312;
  assign n13314 = n12388 & n12393;
  assign n13315 = ~n12383 & n13314;
  assign n13316 = n12370 & ~n13315;
  assign n13317 = ~n12440 & ~n12442;
  assign n13318 = ~n12381 & n13071;
  assign n13319 = n13317 & n13318;
  assign n13320 = n12372 & ~n13319;
  assign n13321 = ~n13316 & ~n13320;
  assign n13322 = n13313 & n13321;
  assign n13323 = ~n12368 & n12374;
  assign n13324 = ~n12399 & ~n12427;
  assign n13325 = n12390 & ~n13324;
  assign n13326 = n12388 & ~n12391;
  assign n13327 = ~n12440 & n13326;
  assign n13328 = n12390 & ~n13327;
  assign n13329 = ~n12402 & ~n13328;
  assign n13330 = ~n12387 & ~n12390;
  assign n13331 = ~n13326 & ~n13330;
  assign n13332 = n13317 & ~n13331;
  assign n13333 = ~n12367 & n13332;
  assign n13334 = ~n13329 & ~n13333;
  assign n13335 = ~n13325 & ~n13334;
  assign n13336 = ~n13323 & n13335;
  assign n13337 = n13322 & n13336;
  assign n13338 = ~n12405 & n13337;
  assign n13339 = n12416 & n13338;
  assign n13340 = n13339 ^ n10494;
  assign n13341 = n13340 ^ x82;
  assign n13342 = n12643 ^ x120;
  assign n13343 = ~n13341 & n13342;
  assign n13344 = n13310 & n13343;
  assign n13345 = n13240 & n13344;
  assign n13346 = n13341 & n13342;
  assign n13347 = n13274 & n13309;
  assign n13348 = n13238 & ~n13239;
  assign n13349 = n13347 & n13348;
  assign n13350 = n13346 & n13349;
  assign n13351 = n13349 ^ n13341;
  assign n13352 = n13351 ^ n13349;
  assign n13353 = n13274 & ~n13309;
  assign n13354 = n13238 & n13239;
  assign n13355 = n13353 & n13354;
  assign n13356 = ~n13274 & ~n13309;
  assign n13357 = ~n13238 & ~n13239;
  assign n13358 = n13356 & n13357;
  assign n13359 = ~n13355 & ~n13358;
  assign n13360 = n13359 ^ n13349;
  assign n13361 = n13352 & ~n13360;
  assign n13362 = n13361 ^ n13349;
  assign n13363 = n13342 & n13362;
  assign n13364 = ~n13350 & ~n13363;
  assign n13365 = n13344 & n13354;
  assign n13366 = n13240 & n13353;
  assign n13367 = n13310 & n13357;
  assign n13368 = ~n13366 & ~n13367;
  assign n13369 = n13346 & ~n13368;
  assign n13370 = ~n13365 & ~n13369;
  assign n13371 = ~n13341 & ~n13342;
  assign n13372 = n13310 & n13354;
  assign n13373 = n13348 & n13353;
  assign n13374 = ~n13372 & ~n13373;
  assign n13375 = n13371 & ~n13374;
  assign n13376 = n13240 & n13347;
  assign n13377 = n13353 & n13357;
  assign n13378 = ~n13376 & ~n13377;
  assign n13379 = n13343 & ~n13378;
  assign n13380 = ~n13375 & ~n13379;
  assign n13381 = n13240 & n13356;
  assign n13382 = n13346 & n13381;
  assign n13383 = n13343 & n13355;
  assign n13384 = n13341 & ~n13342;
  assign n13385 = ~n13378 & n13384;
  assign n13386 = ~n13383 & ~n13385;
  assign n13387 = ~n13382 & n13386;
  assign n13388 = n13348 & n13356;
  assign n13389 = n13343 & n13388;
  assign n13390 = n13346 & ~n13374;
  assign n13391 = ~n13389 & ~n13390;
  assign n13392 = n13344 & n13357;
  assign n13393 = n13347 & n13354;
  assign n13394 = n13240 & n13310;
  assign n13395 = ~n13393 & ~n13394;
  assign n13396 = ~n13358 & n13395;
  assign n13397 = n13354 & n13356;
  assign n13398 = n13310 & n13348;
  assign n13399 = ~n13397 & ~n13398;
  assign n13400 = ~n13373 & n13399;
  assign n13401 = n13396 & n13400;
  assign n13402 = n13384 & ~n13401;
  assign n13403 = ~n13358 & ~n13381;
  assign n13404 = n13347 & n13357;
  assign n13405 = ~n13366 & ~n13404;
  assign n13406 = ~n13349 & ~n13397;
  assign n13407 = n13405 & n13406;
  assign n13408 = n13403 & n13407;
  assign n13409 = n13371 & ~n13408;
  assign n13410 = ~n13402 & ~n13409;
  assign n13411 = ~n13392 & n13410;
  assign n13412 = n13391 & n13411;
  assign n13413 = n13387 & n13412;
  assign n13414 = n13380 & n13413;
  assign n13415 = n13370 & n13414;
  assign n13416 = n13364 & n13415;
  assign n13417 = ~n13345 & n13416;
  assign n13418 = n13417 ^ n12241;
  assign n13419 = n13418 ^ x99;
  assign n13420 = ~n12414 & ~n13317;
  assign n13421 = ~n12377 & n12390;
  assign n13422 = ~n13420 & ~n13421;
  assign n13423 = n12367 & n12372;
  assign n13424 = n12370 & n12403;
  assign n13425 = ~n13423 & ~n13424;
  assign n13426 = ~n12391 & ~n12420;
  assign n13427 = n12402 & ~n13426;
  assign n13428 = ~n12387 & ~n12392;
  assign n13429 = n12414 & ~n13428;
  assign n13430 = ~n13427 & ~n13429;
  assign n13431 = n13425 & n13430;
  assign n13432 = n13422 & n13431;
  assign n13433 = n12434 & n13432;
  assign n13434 = n12406 & n13433;
  assign n13435 = n13060 & n13434;
  assign n13436 = n12379 & n13435;
  assign n13437 = n13436 ^ n10226;
  assign n13438 = n13437 ^ x94;
  assign n13439 = ~n12045 & ~n12051;
  assign n13440 = n12062 & ~n13439;
  assign n13441 = n11872 & ~n13246;
  assign n13442 = ~n13440 & ~n13441;
  assign n13443 = ~n12027 & n12039;
  assign n13444 = ~n12055 & n13443;
  assign n13445 = ~n13244 & ~n13444;
  assign n13446 = n13253 & n13255;
  assign n13447 = n12024 & ~n13446;
  assign n13448 = ~n13445 & ~n13447;
  assign n13449 = n12031 & ~n12058;
  assign n13450 = n11904 & n12069;
  assign n13451 = ~n13449 & ~n13450;
  assign n13452 = n13448 & n13451;
  assign n13453 = n13442 & n13452;
  assign n13454 = n12054 & n13453;
  assign n13455 = n13454 ^ n10189;
  assign n13456 = n13455 ^ x100;
  assign n13457 = ~n13438 & n13456;
  assign n13458 = n12778 & ~n12809;
  assign n13459 = ~n12814 & n13280;
  assign n13460 = ~n12797 & n13459;
  assign n13461 = ~n12776 & n13460;
  assign n13462 = n12798 & ~n13461;
  assign n13463 = ~n13458 & ~n13462;
  assign n13464 = n12799 & n12804;
  assign n13465 = ~n12782 & n13276;
  assign n13466 = n12774 & ~n13465;
  assign n13467 = ~n12797 & n13295;
  assign n13468 = n12778 & ~n13467;
  assign n13469 = ~n12788 & n13292;
  assign n13470 = n12720 & ~n13469;
  assign n13471 = ~n13468 & ~n13470;
  assign n13472 = ~n13466 & n13471;
  assign n13473 = ~n13464 & n13472;
  assign n13474 = n13463 & n13473;
  assign n13475 = n13289 & n13474;
  assign n13476 = n13282 & n13475;
  assign n13477 = n13286 & n13476;
  assign n13478 = ~n12773 & n13477;
  assign n13479 = ~n12835 & n13478;
  assign n13480 = n13479 ^ n10162;
  assign n13481 = n13480 ^ x93;
  assign n13482 = n12579 & n12601;
  assign n13483 = n12586 & ~n13096;
  assign n13484 = ~n13482 & ~n13483;
  assign n13485 = n12600 & n12622;
  assign n13486 = n12606 & ~n12621;
  assign n13487 = ~n12592 & n13486;
  assign n13488 = n12581 & ~n13487;
  assign n13489 = ~n13485 & ~n13488;
  assign n13490 = n13484 & n13489;
  assign n13491 = ~n12560 & n12616;
  assign n13492 = n12603 & ~n13491;
  assign n13493 = ~n12613 & ~n12626;
  assign n13494 = ~n12610 & ~n13493;
  assign n13495 = n12581 & ~n13491;
  assign n13496 = n12586 & ~n13088;
  assign n13497 = n12598 & ~n12605;
  assign n13498 = ~n12603 & n13497;
  assign n13499 = ~n12611 & n12627;
  assign n13500 = ~n12592 & n13499;
  assign n13501 = ~n12600 & n13500;
  assign n13502 = ~n13498 & ~n13501;
  assign n13503 = n12579 & n13502;
  assign n13504 = ~n13496 & ~n13503;
  assign n13505 = ~n13495 & n13504;
  assign n13506 = n12591 & n13505;
  assign n13507 = ~n13494 & n13506;
  assign n13508 = ~n13492 & n13507;
  assign n13509 = n13490 & n13508;
  assign n13510 = n13509 ^ n10263;
  assign n13511 = n13510 ^ x75;
  assign n13512 = ~n13481 & n13511;
  assign n13513 = n13457 & n13512;
  assign n13514 = n13438 & ~n13456;
  assign n13515 = n13512 & n13514;
  assign n13516 = ~n13513 & ~n13515;
  assign n13517 = ~n12250 & n12252;
  assign n13518 = n12265 & n12286;
  assign n13519 = ~n13517 & ~n13518;
  assign n13520 = n12133 & ~n12262;
  assign n13521 = n12247 & n12271;
  assign n13522 = ~n12276 & n12278;
  assign n13523 = ~n13521 & ~n13522;
  assign n13524 = ~n13520 & n13523;
  assign n13525 = n13519 & n13524;
  assign n13526 = n13525 ^ n10020;
  assign n13527 = n13526 ^ x76;
  assign n13528 = n11553 ^ n11450;
  assign n13529 = n11694 ^ n11450;
  assign n13530 = n11450 ^ n11416;
  assign n13531 = n13530 ^ n11450;
  assign n13532 = ~n13529 & n13531;
  assign n13533 = n13532 ^ n11450;
  assign n13534 = ~n13528 & n13533;
  assign n13535 = n11762 & n13534;
  assign n13536 = n11798 & ~n11806;
  assign n13537 = n11770 & ~n13536;
  assign n13538 = ~n11792 & ~n11810;
  assign n13539 = ~n11765 & n13040;
  assign n13540 = n13539 ^ n13022;
  assign n13541 = n13539 ^ n11781;
  assign n13542 = n13541 ^ n11781;
  assign n13543 = ~n11767 & ~n11837;
  assign n13544 = n13543 ^ n11781;
  assign n13545 = ~n13542 & n13544;
  assign n13546 = n13545 ^ n11781;
  assign n13547 = n13540 & ~n13546;
  assign n13548 = n13547 ^ n13022;
  assign n13549 = n13538 & n13548;
  assign n13550 = ~n11772 & n13549;
  assign n13551 = ~n11787 & ~n13550;
  assign n13552 = ~n13537 & ~n13551;
  assign n13553 = ~n13535 & n13552;
  assign n13554 = ~n13017 & n13553;
  assign n13555 = n13015 & n13554;
  assign n13556 = n11805 & n13555;
  assign n13557 = n13027 & n13556;
  assign n13558 = ~n11763 & n13557;
  assign n13559 = n13558 ^ n10047;
  assign n13560 = n13559 ^ x125;
  assign n13561 = ~n13527 & ~n13560;
  assign n13562 = ~n13516 & n13561;
  assign n13563 = n13527 & n13560;
  assign n13564 = n13481 & n13511;
  assign n13565 = n13457 & n13564;
  assign n13566 = ~n13438 & ~n13456;
  assign n13567 = n13512 & n13566;
  assign n13568 = ~n13565 & ~n13567;
  assign n13569 = n13563 & ~n13568;
  assign n13570 = ~n13562 & ~n13569;
  assign n13571 = ~n13527 & n13560;
  assign n13572 = n13481 & ~n13511;
  assign n13573 = n13457 & n13572;
  assign n13574 = n13571 & n13573;
  assign n13575 = n13438 & n13456;
  assign n13576 = ~n13481 & ~n13511;
  assign n13577 = n13575 & n13576;
  assign n13578 = n13527 & ~n13560;
  assign n13579 = n13577 & n13578;
  assign n13580 = ~n13574 & ~n13579;
  assign n13581 = ~n13571 & ~n13578;
  assign n13582 = n13513 & ~n13581;
  assign n13583 = n13564 & n13575;
  assign n13584 = n13514 & n13564;
  assign n13585 = ~n13583 & ~n13584;
  assign n13586 = n13566 & n13572;
  assign n13587 = n13512 & n13575;
  assign n13588 = n13514 & n13576;
  assign n13589 = ~n13587 & ~n13588;
  assign n13590 = ~n13586 & n13589;
  assign n13591 = ~n13567 & n13590;
  assign n13592 = n13585 & n13591;
  assign n13593 = n13571 & ~n13592;
  assign n13594 = ~n13582 & ~n13593;
  assign n13595 = n13572 & n13575;
  assign n13596 = ~n13588 & ~n13595;
  assign n13597 = ~n13583 & n13596;
  assign n13598 = n13578 & ~n13597;
  assign n13599 = n13564 & n13566;
  assign n13600 = ~n13565 & ~n13586;
  assign n13601 = ~n13599 & n13600;
  assign n13602 = ~n13560 & ~n13601;
  assign n13603 = n13457 & n13576;
  assign n13604 = n13566 & n13576;
  assign n13605 = ~n13603 & ~n13604;
  assign n13606 = n13563 & ~n13605;
  assign n13607 = ~n13584 & ~n13595;
  assign n13608 = n13514 & n13572;
  assign n13609 = ~n13515 & ~n13608;
  assign n13610 = n13607 & n13609;
  assign n13611 = ~n13561 & n13610;
  assign n13612 = ~n13577 & n13596;
  assign n13613 = ~n13563 & n13612;
  assign n13614 = ~n13611 & ~n13613;
  assign n13615 = n13581 & n13614;
  assign n13616 = ~n13606 & ~n13615;
  assign n13617 = ~n13602 & n13616;
  assign n13618 = ~n13598 & n13617;
  assign n13619 = n13594 & n13618;
  assign n13620 = n13580 & n13619;
  assign n13621 = n13570 & n13620;
  assign n13622 = n13621 ^ n12175;
  assign n13623 = n13622 ^ x89;
  assign n13624 = n13419 & n13623;
  assign n13625 = ~n13419 & ~n13623;
  assign n13626 = ~n13624 & ~n13625;
  assign n13627 = n13207 & ~n13626;
  assign n13628 = n13455 ^ x88;
  assign n13629 = n13237 ^ x66;
  assign n13630 = n13628 & ~n13629;
  assign n13631 = n13526 ^ x64;
  assign n13632 = n11321 & n11333;
  assign n13633 = n10333 & n11327;
  assign n13634 = ~n13632 & ~n13633;
  assign n13635 = ~n11317 & n11343;
  assign n13636 = n11325 & ~n13635;
  assign n13637 = n11309 & n11329;
  assign n13638 = ~n11338 & ~n13637;
  assign n13639 = ~n11342 & n13638;
  assign n13640 = ~n11310 & n13639;
  assign n13641 = n11321 & ~n13640;
  assign n13642 = ~n13636 & ~n13641;
  assign n13643 = ~n11340 & ~n11342;
  assign n13644 = n11312 & ~n13643;
  assign n13645 = ~n11315 & ~n11340;
  assign n13646 = n10333 & ~n13645;
  assign n13647 = n11312 & n11333;
  assign n13648 = n11325 & n11327;
  assign n13649 = ~n13647 & ~n13648;
  assign n13650 = n11325 & n11337;
  assign n13651 = n11310 & n11312;
  assign n13652 = ~n13650 & ~n13651;
  assign n13653 = n10332 ^ n10003;
  assign n13654 = ~n11339 & ~n11349;
  assign n13655 = n13654 ^ n11351;
  assign n13656 = n13653 & n13655;
  assign n13657 = n13656 ^ n13654;
  assign n13658 = n13652 & n13657;
  assign n13659 = n13649 & n13658;
  assign n13660 = ~n13646 & n13659;
  assign n13661 = ~n13644 & n13660;
  assign n13662 = n13642 & n13661;
  assign n13663 = n13634 & n13662;
  assign n13664 = n11323 & ~n13653;
  assign n13665 = n13663 & ~n13664;
  assign n13666 = n11335 & n13665;
  assign n13667 = n11320 & n13666;
  assign n13668 = n13667 ^ n10539;
  assign n13669 = n13668 ^ x73;
  assign n13670 = n13631 & n13669;
  assign n13671 = n11772 & n11781;
  assign n13672 = n11767 & n11806;
  assign n13673 = ~n13671 & ~n13672;
  assign n13674 = n11777 & ~n11810;
  assign n13675 = n11762 & ~n13674;
  assign n13676 = ~n11792 & n13040;
  assign n13677 = n11770 & ~n13676;
  assign n13678 = ~n13675 & ~n13677;
  assign n13679 = n13673 & n13678;
  assign n13680 = n11800 & ~n11817;
  assign n13681 = ~n11789 & ~n11797;
  assign n13682 = ~n11787 & ~n13681;
  assign n13683 = n11762 & n11783;
  assign n13684 = n11770 & n11797;
  assign n13685 = ~n13683 & ~n13684;
  assign n13686 = n11795 & ~n11817;
  assign n13687 = n11767 & ~n13538;
  assign n13688 = n11781 & ~n13040;
  assign n13689 = ~n13687 & ~n13688;
  assign n13690 = ~n13686 & n13689;
  assign n13691 = n13685 & n13690;
  assign n13692 = ~n11841 & n13691;
  assign n13693 = n11780 & n13692;
  assign n13694 = ~n11763 & n13693;
  assign n13695 = ~n13682 & n13694;
  assign n13696 = ~n13680 & n13695;
  assign n13697 = n13679 & n13696;
  assign n13698 = n13020 & n13697;
  assign n13699 = n13698 ^ n10588;
  assign n13700 = n13699 ^ x112;
  assign n13701 = n13340 ^ x98;
  assign n13702 = n13700 & ~n13701;
  assign n13703 = n13670 & n13702;
  assign n13704 = n13630 & n13703;
  assign n13705 = n13628 & n13629;
  assign n13706 = ~n13700 & n13701;
  assign n13707 = n13670 & n13706;
  assign n13708 = ~n13700 & ~n13701;
  assign n13709 = n13631 & ~n13669;
  assign n13710 = n13708 & n13709;
  assign n13711 = ~n13707 & ~n13710;
  assign n13712 = n13705 & ~n13711;
  assign n13713 = ~n13631 & n13669;
  assign n13714 = n13706 & n13713;
  assign n13715 = n13630 & n13714;
  assign n13716 = n13629 ^ n13628;
  assign n13717 = n13700 & n13701;
  assign n13718 = n13713 & n13717;
  assign n13719 = n13718 ^ n13629;
  assign n13720 = n13719 ^ n13718;
  assign n13721 = ~n13631 & ~n13669;
  assign n13722 = n13706 & n13721;
  assign n13723 = n13722 ^ n13718;
  assign n13724 = ~n13720 & n13723;
  assign n13725 = n13724 ^ n13718;
  assign n13726 = ~n13716 & n13725;
  assign n13727 = ~n13715 & ~n13726;
  assign n13728 = n13628 & n13722;
  assign n13729 = n13717 & n13721;
  assign n13730 = n13702 & n13721;
  assign n13731 = ~n13729 & ~n13730;
  assign n13732 = ~n13629 & ~n13731;
  assign n13733 = ~n13728 & ~n13732;
  assign n13734 = ~n13628 & ~n13629;
  assign n13735 = n13702 & n13713;
  assign n13736 = n13734 & n13735;
  assign n13737 = ~n13628 & n13629;
  assign n13738 = n13670 & n13708;
  assign n13739 = n13709 & n13717;
  assign n13740 = ~n13738 & ~n13739;
  assign n13741 = n13708 & n13713;
  assign n13742 = ~n13718 & ~n13741;
  assign n13743 = ~n13729 & n13742;
  assign n13744 = n13701 ^ n13700;
  assign n13745 = n13709 & n13744;
  assign n13746 = ~n13703 & ~n13745;
  assign n13747 = n13743 & n13746;
  assign n13748 = n13740 & n13747;
  assign n13749 = n13737 & ~n13748;
  assign n13750 = ~n13736 & ~n13749;
  assign n13751 = n13708 & n13721;
  assign n13752 = ~n13730 & ~n13751;
  assign n13753 = n13705 & ~n13752;
  assign n13754 = ~n13705 & ~n13734;
  assign n13755 = ~n13703 & ~n13734;
  assign n13756 = n13702 & n13709;
  assign n13757 = ~n13707 & ~n13756;
  assign n13758 = ~n13705 & n13757;
  assign n13759 = ~n13738 & n13758;
  assign n13760 = ~n13755 & ~n13759;
  assign n13761 = ~n13754 & n13760;
  assign n13762 = n13670 & n13717;
  assign n13763 = n13762 ^ n13630;
  assign n13764 = n13762 ^ n13754;
  assign n13765 = n13764 ^ n13754;
  assign n13766 = ~n13710 & ~n13739;
  assign n13767 = n13766 ^ n13754;
  assign n13768 = ~n13765 & ~n13767;
  assign n13769 = n13768 ^ n13754;
  assign n13770 = n13763 & ~n13769;
  assign n13771 = n13770 ^ n13630;
  assign n13772 = ~n13761 & ~n13771;
  assign n13773 = ~n13753 & n13772;
  assign n13774 = n13750 & n13773;
  assign n13775 = n13733 & n13774;
  assign n13776 = n13727 & n13775;
  assign n13777 = ~n13712 & n13776;
  assign n13778 = ~n13704 & n13777;
  assign n13779 = n13778 ^ n10670;
  assign n13780 = n13779 ^ x74;
  assign n13781 = n13437 ^ x69;
  assign n13782 = n12774 & n12808;
  assign n13783 = n12788 & n12799;
  assign n13784 = ~n13782 & ~n13783;
  assign n13785 = ~n12782 & ~n12797;
  assign n13786 = n12778 & ~n13785;
  assign n13787 = n12778 & ~n13280;
  assign n13788 = ~n12790 & ~n12820;
  assign n13789 = ~n12808 & n13788;
  assign n13790 = ~n12799 & ~n13789;
  assign n13791 = ~n13787 & ~n13790;
  assign n13792 = ~n12784 & ~n12803;
  assign n13793 = n12798 & ~n13792;
  assign n13794 = ~n12776 & n12809;
  assign n13795 = n12774 & ~n13794;
  assign n13796 = ~n13793 & ~n13795;
  assign n13797 = n13791 & n13796;
  assign n13798 = n13278 & n13797;
  assign n13799 = ~n12835 & n13798;
  assign n13800 = ~n13786 & n13799;
  assign n13801 = n12776 ^ n12719;
  assign n13802 = n13801 ^ n12776;
  assign n13803 = n12805 ^ n12776;
  assign n13804 = n13803 ^ n12776;
  assign n13805 = ~n13802 & ~n13804;
  assign n13806 = n13805 ^ n12776;
  assign n13807 = n12718 & n13806;
  assign n13808 = n13807 ^ n12776;
  assign n13809 = n13800 & ~n13808;
  assign n13810 = n13784 & n13809;
  assign n13811 = n13283 & n13810;
  assign n13812 = n13811 ^ n11132;
  assign n13813 = n13812 ^ x78;
  assign n13814 = n13781 & ~n13813;
  assign n13815 = n12265 & ~n12973;
  assign n13816 = n12133 & ~n12999;
  assign n13817 = ~n13815 & ~n13816;
  assign n13818 = n12252 & n12983;
  assign n13819 = n12278 & ~n13006;
  assign n13820 = ~n13818 & ~n13819;
  assign n13821 = n13817 & n13820;
  assign n13822 = n13821 ^ n11481;
  assign n13823 = n13822 ^ x118;
  assign n13824 = n12893 & n12918;
  assign n13825 = n12841 & ~n13219;
  assign n13826 = ~n13824 & ~n13825;
  assign n13827 = ~n12839 & ~n12949;
  assign n13828 = ~n12898 & ~n12937;
  assign n13829 = n12906 & ~n13828;
  assign n13830 = ~n13827 & ~n13829;
  assign n13831 = n12900 & ~n12934;
  assign n13832 = n12902 & ~n13831;
  assign n13833 = ~n12893 & n13213;
  assign n13834 = n12841 & ~n13833;
  assign n13835 = ~n12908 & ~n12920;
  assign n13836 = ~n12918 & ~n12942;
  assign n13837 = ~n12919 & n13836;
  assign n13838 = ~n12839 & ~n13837;
  assign n13839 = n13835 & ~n13838;
  assign n13840 = n13219 & n13839;
  assign n13841 = n13835 & n13836;
  assign n13842 = ~n12906 & n12912;
  assign n13843 = ~n13841 & ~n13842;
  assign n13844 = ~n12919 & ~n13843;
  assign n13845 = n13844 ^ n12840;
  assign n13846 = ~n12839 & ~n13845;
  assign n13847 = n13846 ^ n12840;
  assign n13848 = ~n13840 & n13847;
  assign n13849 = ~n13834 & ~n13848;
  assign n13850 = ~n13832 & n13849;
  assign n13851 = n13830 & n13850;
  assign n13852 = n13826 & n13851;
  assign n13853 = n12930 & n13852;
  assign n13854 = n13853 ^ n11470;
  assign n13855 = n13854 ^ x108;
  assign n13856 = n13823 & n13855;
  assign n13857 = n11312 & n11330;
  assign n13858 = n11321 & n11337;
  assign n13859 = ~n13857 & ~n13858;
  assign n13860 = ~n11349 & n13638;
  assign n13861 = n11312 & ~n13860;
  assign n13862 = ~n11341 & n13654;
  assign n13863 = ~n11333 & n13862;
  assign n13864 = n11351 & n13863;
  assign n13865 = n10333 & ~n13864;
  assign n13866 = ~n13861 & ~n13865;
  assign n13867 = n11344 & ~n13637;
  assign n13868 = n11321 & ~n13867;
  assign n13869 = ~n11333 & ~n11339;
  assign n13870 = n11312 & ~n13869;
  assign n13871 = ~n11350 & ~n13637;
  assign n13872 = n11345 & n13871;
  assign n13873 = ~n11330 & n13872;
  assign n13874 = n11325 & ~n13873;
  assign n13875 = ~n13870 & ~n13874;
  assign n13876 = ~n13868 & n13875;
  assign n13877 = n13866 & n13876;
  assign n13878 = n13634 & n13877;
  assign n13879 = n13859 & n13878;
  assign n13880 = ~n11328 & n13879;
  assign n13881 = ~n11324 & n13880;
  assign n13882 = n11320 & n13881;
  assign n13883 = n13882 ^ n11099;
  assign n13884 = n13883 ^ x101;
  assign n13885 = n13559 ^ x91;
  assign n13886 = ~n13884 & ~n13885;
  assign n13887 = n13856 & n13886;
  assign n13888 = n13814 & n13887;
  assign n13889 = ~n13781 & ~n13813;
  assign n13890 = ~n13884 & n13885;
  assign n13891 = n13823 & ~n13855;
  assign n13892 = n13890 & n13891;
  assign n13893 = n13889 & n13892;
  assign n13894 = n13781 & n13813;
  assign n13895 = n13884 & n13885;
  assign n13896 = ~n13823 & ~n13855;
  assign n13897 = n13895 & n13896;
  assign n13898 = ~n13823 & n13855;
  assign n13899 = n13884 & ~n13885;
  assign n13900 = n13898 & n13899;
  assign n13901 = ~n13897 & ~n13900;
  assign n13902 = n13894 & ~n13901;
  assign n13903 = ~n13893 & ~n13902;
  assign n13904 = n13892 & n13894;
  assign n13905 = n13856 & n13899;
  assign n13906 = n13889 & n13905;
  assign n13907 = ~n13904 & ~n13906;
  assign n13908 = n13886 & n13898;
  assign n13909 = ~n13892 & ~n13908;
  assign n13910 = n13814 & ~n13909;
  assign n13911 = ~n13781 & n13813;
  assign n13912 = n13884 ^ n13823;
  assign n13913 = n13912 ^ n13885;
  assign n13914 = n13913 ^ n13884;
  assign n13915 = n13914 ^ n13855;
  assign n13916 = n13915 ^ n13885;
  assign n13917 = n13885 ^ n13884;
  assign n13918 = n13884 ^ n13855;
  assign n13919 = n13918 ^ n13884;
  assign n13920 = n13917 & n13919;
  assign n13921 = n13920 ^ n13884;
  assign n13922 = n13916 & n13921;
  assign n13923 = n13922 ^ n13913;
  assign n13924 = n13911 & n13923;
  assign n13925 = ~n13887 & ~n13908;
  assign n13926 = n13890 & n13896;
  assign n13927 = ~n13897 & ~n13926;
  assign n13928 = n13895 & n13898;
  assign n13929 = n13891 & n13899;
  assign n13930 = ~n13928 & ~n13929;
  assign n13931 = n13927 & n13930;
  assign n13932 = n13925 & n13931;
  assign n13933 = n13889 & ~n13932;
  assign n13934 = n13896 & n13899;
  assign n13935 = n13890 & n13898;
  assign n13936 = ~n13926 & ~n13935;
  assign n13937 = ~n13934 & n13936;
  assign n13938 = n13891 & n13895;
  assign n13939 = ~n13900 & ~n13938;
  assign n13940 = n13937 & n13939;
  assign n13941 = n13814 & ~n13940;
  assign n13942 = n13856 & n13890;
  assign n13943 = n13886 & n13896;
  assign n13944 = ~n13942 & ~n13943;
  assign n13945 = ~n13908 & n13944;
  assign n13946 = ~n13929 & n13945;
  assign n13947 = ~n13905 & n13946;
  assign n13948 = n13894 & ~n13947;
  assign n13949 = ~n13941 & ~n13948;
  assign n13950 = ~n13933 & n13949;
  assign n13951 = ~n13924 & n13950;
  assign n13952 = ~n13910 & n13951;
  assign n13953 = n13907 & n13952;
  assign n13954 = n13903 & n13953;
  assign n13955 = ~n13888 & n13954;
  assign n13956 = n13955 ^ n12131;
  assign n13957 = n13956 ^ x121;
  assign n13958 = n13780 & ~n13957;
  assign n13959 = ~n13419 & n13623;
  assign n13960 = n12717 & n13959;
  assign n13961 = n13419 & ~n13623;
  assign n13962 = n12717 & ~n13206;
  assign n13963 = n13961 & n13962;
  assign n13964 = ~n13960 & ~n13963;
  assign n13965 = n12717 & n13206;
  assign n13966 = ~n13961 & n13965;
  assign n13967 = ~n12717 & ~n13206;
  assign n13968 = n13625 & n13967;
  assign n13969 = ~n13966 & ~n13968;
  assign n13970 = n13207 & n13961;
  assign n13971 = n13959 & n13967;
  assign n13972 = ~n13970 & ~n13971;
  assign n13973 = n13969 & n13972;
  assign n13974 = n13964 & n13973;
  assign n13975 = n13958 & n13974;
  assign n13976 = ~n13780 & ~n13957;
  assign n13977 = ~n13419 & n13965;
  assign n13978 = ~n13963 & ~n13977;
  assign n13979 = n13961 & n13965;
  assign n13980 = n13624 & n13967;
  assign n13981 = ~n13979 & ~n13980;
  assign n13982 = n13978 & n13981;
  assign n13983 = ~n13971 & n13982;
  assign n13984 = n13976 & ~n13983;
  assign n13985 = ~n13975 & ~n13984;
  assign n13986 = ~n13780 & n13957;
  assign n13987 = n13419 ^ n12717;
  assign n13988 = n13987 ^ n13206;
  assign n13989 = n13623 ^ n12717;
  assign n13990 = n13206 ^ n12717;
  assign n13991 = n13990 ^ n12717;
  assign n13992 = ~n13989 & ~n13991;
  assign n13993 = n13992 ^ n12717;
  assign n13994 = ~n13988 & n13993;
  assign n13995 = n13994 ^ n12717;
  assign n13996 = n13986 & n13995;
  assign n13997 = n13780 & n13957;
  assign n13998 = n13624 & n13965;
  assign n13999 = n13964 & ~n13998;
  assign n14000 = n13972 & n13999;
  assign n14001 = n13997 & ~n14000;
  assign n14002 = ~n13996 & ~n14001;
  assign n14003 = n13985 & n14002;
  assign n14004 = ~n13627 & n14003;
  assign n14005 = n14004 ^ n13526;
  assign n14006 = n14005 ^ x97;
  assign n14007 = n12087 ^ x72;
  assign n14008 = n13120 ^ x90;
  assign n14009 = n14007 & ~n14008;
  assign n14010 = n12837 ^ x96;
  assign n14011 = n12840 & n12896;
  assign n14012 = ~n12924 & ~n12937;
  assign n14013 = n12918 & ~n14012;
  assign n14014 = ~n14011 & ~n14013;
  assign n14015 = ~n12898 & ~n12934;
  assign n14016 = ~n12893 & n14015;
  assign n14017 = n12906 & ~n14016;
  assign n14018 = n12863 & n12903;
  assign n14019 = n13835 & ~n14018;
  assign n14020 = n12841 & ~n14019;
  assign n14021 = ~n12924 & n14016;
  assign n14022 = n12841 & ~n14021;
  assign n14023 = n12891 ^ n12863;
  assign n14024 = n14023 ^ n12864;
  assign n14025 = n12891 ^ n12864;
  assign n14026 = n14025 ^ n12864;
  assign n14027 = ~n14024 & n14026;
  assign n14028 = n14027 ^ n12864;
  assign n14029 = n12890 & n14028;
  assign n14030 = n14029 ^ n14023;
  assign n14031 = n12902 & ~n14030;
  assign n14032 = ~n14022 & ~n14031;
  assign n14033 = ~n12902 & ~n12906;
  assign n14034 = n12931 & ~n14033;
  assign n14035 = n13835 ^ n12839;
  assign n14036 = ~n12916 & ~n12919;
  assign n14037 = n14036 ^ n14018;
  assign n14038 = n14018 ^ n12840;
  assign n14039 = n14038 ^ n14018;
  assign n14040 = ~n14037 & n14039;
  assign n14041 = n14040 ^ n14018;
  assign n14042 = n14041 ^ n13835;
  assign n14043 = ~n14035 & ~n14042;
  assign n14044 = n14043 ^ n14040;
  assign n14045 = n14044 ^ n14018;
  assign n14046 = n14045 ^ n12839;
  assign n14047 = n13835 & n14046;
  assign n14048 = n14047 ^ n13835;
  assign n14049 = n14048 ^ n12839;
  assign n14050 = ~n14034 & n14049;
  assign n14051 = n14032 & n14050;
  assign n14052 = ~n14020 & n14051;
  assign n14053 = ~n14017 & n14052;
  assign n14054 = n14014 & n14053;
  assign n14055 = ~n12928 & n14054;
  assign n14056 = n14055 ^ n10942;
  assign n14057 = n14056 ^ x105;
  assign n14058 = ~n14010 & n14057;
  assign n14059 = ~n11315 & n11343;
  assign n14060 = n11312 & ~n14059;
  assign n14061 = ~n11337 & n11353;
  assign n14062 = n10333 & ~n14061;
  assign n14063 = ~n14060 & ~n14062;
  assign n14064 = ~n11370 & ~n13653;
  assign n14065 = n11318 & n13643;
  assign n14066 = n11321 & ~n14065;
  assign n14067 = ~n11327 & n13871;
  assign n14068 = n11312 & ~n14067;
  assign n14069 = n13638 & n13863;
  assign n14070 = ~n11323 & n14069;
  assign n14071 = n11325 & ~n14070;
  assign n14072 = ~n14068 & ~n14071;
  assign n14073 = ~n14066 & n14072;
  assign n14074 = ~n14064 & n14073;
  assign n14075 = n14063 & n14074;
  assign n14076 = ~n13664 & n14075;
  assign n14077 = n13859 & n14076;
  assign n14078 = n13649 & n14077;
  assign n14079 = n14078 ^ n10977;
  assign n14080 = n14079 ^ x114;
  assign n14081 = n11845 ^ x115;
  assign n14082 = n14080 & ~n14081;
  assign n14083 = n14058 & n14082;
  assign n14084 = n14010 & n14057;
  assign n14085 = ~n14080 & n14081;
  assign n14086 = n14084 & n14085;
  assign n14087 = ~n14080 & ~n14081;
  assign n14088 = ~n14057 & n14087;
  assign n14089 = ~n14086 & ~n14088;
  assign n14090 = ~n14083 & n14089;
  assign n14091 = ~n14010 & ~n14057;
  assign n14092 = n14081 & n14091;
  assign n14093 = n14080 & n14081;
  assign n14094 = ~n14087 & ~n14093;
  assign n14095 = n14084 & ~n14094;
  assign n14096 = ~n14092 & ~n14095;
  assign n14097 = n14090 & n14096;
  assign n14098 = n14009 & n14097;
  assign n14099 = ~n14007 & n14008;
  assign n14100 = n14010 & ~n14057;
  assign n14101 = n14082 & n14100;
  assign n14102 = n14093 & n14100;
  assign n14103 = ~n14010 & n14085;
  assign n14104 = n14090 & ~n14103;
  assign n14105 = ~n14102 & n14104;
  assign n14106 = ~n14101 & n14105;
  assign n14107 = n14099 & ~n14106;
  assign n14108 = ~n14098 & ~n14107;
  assign n14109 = n14007 & n14008;
  assign n14110 = n14085 & n14100;
  assign n14111 = n14084 & n14087;
  assign n14112 = ~n14110 & ~n14111;
  assign n14113 = ~n14010 & n14087;
  assign n14114 = ~n14101 & ~n14113;
  assign n14115 = n14084 & n14093;
  assign n14116 = n14091 & n14093;
  assign n14117 = n14082 & n14084;
  assign n14118 = ~n14116 & ~n14117;
  assign n14119 = ~n14115 & n14118;
  assign n14120 = n14114 & n14119;
  assign n14121 = n14112 & n14120;
  assign n14122 = n14109 & ~n14121;
  assign n14123 = ~n14007 & ~n14008;
  assign n14124 = n14081 ^ n14057;
  assign n14125 = n14124 ^ n14080;
  assign n14126 = n14125 ^ n14081;
  assign n14127 = n14081 ^ n14010;
  assign n14128 = n14127 ^ n14010;
  assign n14129 = n14080 ^ n14010;
  assign n14130 = n14129 ^ n14010;
  assign n14131 = n14128 & ~n14130;
  assign n14132 = n14131 ^ n14010;
  assign n14133 = n14126 & n14132;
  assign n14134 = n14133 ^ n14124;
  assign n14135 = n14123 & ~n14134;
  assign n14136 = ~n14122 & ~n14135;
  assign n14137 = n14108 & n14136;
  assign n14138 = n14137 ^ n11029;
  assign n14139 = n14138 ^ x76;
  assign n14140 = n13133 & n13136;
  assign n14141 = ~n13181 & ~n14140;
  assign n14142 = n13129 & n14141;
  assign n14143 = ~n13150 & n13162;
  assign n14144 = ~n13132 & ~n13157;
  assign n14145 = ~n13177 & n14144;
  assign n14146 = ~n12838 & ~n14145;
  assign n14147 = ~n14143 & ~n14146;
  assign n14148 = ~n13127 & n13184;
  assign n14149 = n12967 & ~n14148;
  assign n14150 = n13142 & ~n13164;
  assign n14151 = ~n13148 & n14150;
  assign n14152 = n13136 & ~n14151;
  assign n14153 = ~n14149 & ~n14152;
  assign n14154 = n13150 & n13182;
  assign n14155 = ~n13127 & ~n13153;
  assign n14156 = ~n13141 & n14155;
  assign n14157 = ~n13152 & n14156;
  assign n14158 = n14157 ^ n13143;
  assign n14159 = n13143 ^ n12966;
  assign n14160 = n14159 ^ n13143;
  assign n14161 = n14158 & ~n14160;
  assign n14162 = n14161 ^ n13143;
  assign n14163 = ~n12838 & ~n14162;
  assign n14164 = ~n14154 & ~n14163;
  assign n14165 = n14153 & n14164;
  assign n14166 = n14147 & n14165;
  assign n14167 = n13167 & n14166;
  assign n14168 = n14142 & n14167;
  assign n14169 = n14168 ^ n12019;
  assign n14170 = n14169 ^ x93;
  assign n14171 = ~n14139 & n14170;
  assign n14172 = n13737 & n13762;
  assign n14173 = n13705 & n13730;
  assign n14174 = ~n14172 & ~n14173;
  assign n14175 = n13734 & n13762;
  assign n14176 = ~n13731 & n13737;
  assign n14177 = ~n14175 & ~n14176;
  assign n14178 = n13628 & n13735;
  assign n14179 = ~n13714 & ~n13751;
  assign n14180 = ~n13754 & ~n14179;
  assign n14181 = ~n14178 & ~n14180;
  assign n14182 = ~n13703 & n13766;
  assign n14183 = n13737 & ~n14182;
  assign n14184 = ~n13729 & n13746;
  assign n14185 = n13734 & ~n14184;
  assign n14186 = ~n13722 & ~n13741;
  assign n14187 = n13754 & ~n14186;
  assign n14188 = n13740 & ~n13762;
  assign n14189 = ~n13630 & n14188;
  assign n14190 = n13758 & n13766;
  assign n14191 = ~n14189 & ~n14190;
  assign n14192 = n13628 & n14191;
  assign n14193 = ~n14187 & ~n14192;
  assign n14194 = ~n14185 & n14193;
  assign n14195 = ~n14183 & n14194;
  assign n14196 = n14181 & n14195;
  assign n14197 = n13727 & n14196;
  assign n14198 = n14177 & n14197;
  assign n14199 = n14174 & n14198;
  assign n14200 = n14199 ^ n12332;
  assign n14201 = n14200 ^ x117;
  assign n14202 = n12658 & n12662;
  assign n14203 = ~n12665 & ~n12677;
  assign n14204 = n11847 & ~n14203;
  assign n14205 = ~n14202 & ~n14204;
  assign n14206 = n12662 & n12687;
  assign n14207 = n12656 & n12683;
  assign n14208 = ~n14206 & ~n14207;
  assign n14209 = ~n12670 & n12699;
  assign n14210 = n12666 & ~n14209;
  assign n14211 = ~n12655 & ~n12690;
  assign n14212 = n12666 & ~n14211;
  assign n14213 = n12666 & ~n14203;
  assign n14214 = ~n12686 & n12703;
  assign n14215 = n11847 & ~n14214;
  assign n14216 = n12458 ^ n12292;
  assign n14217 = n14216 ^ n12088;
  assign n14218 = n14217 ^ n12644;
  assign n14219 = n12458 ^ n12088;
  assign n14220 = ~n12644 & ~n14219;
  assign n14221 = n14218 & n14220;
  assign n14222 = n14221 ^ n14218;
  assign n14223 = n12652 & n14222;
  assign n14224 = ~n14215 & ~n14223;
  assign n14225 = ~n14213 & n14224;
  assign n14226 = ~n12648 & n14225;
  assign n14227 = ~n14212 & n14226;
  assign n14228 = ~n14210 & n14227;
  assign n14229 = ~n12670 & ~n12697;
  assign n14230 = n14229 ^ n12647;
  assign n14231 = n14230 ^ n12647;
  assign n14232 = n12647 ^ n11382;
  assign n14233 = n14232 ^ n12647;
  assign n14234 = ~n14231 & n14233;
  assign n14235 = n14234 ^ n12647;
  assign n14236 = n11846 & n14235;
  assign n14237 = n14236 ^ n12647;
  assign n14238 = n14228 & ~n14237;
  assign n14239 = n14208 & n14238;
  assign n14240 = n14205 & n14239;
  assign n14241 = n14240 ^ n11871;
  assign n14242 = n14241 ^ x83;
  assign n14243 = ~n14201 & n14242;
  assign n14244 = n13561 & n13583;
  assign n14245 = n13573 & n13578;
  assign n14246 = ~n14244 & ~n14245;
  assign n14247 = n13563 & n13586;
  assign n14248 = n13515 & n13571;
  assign n14249 = ~n14247 & ~n14248;
  assign n14250 = ~n13599 & ~n13603;
  assign n14251 = n13578 & ~n14250;
  assign n14252 = n14249 & ~n14251;
  assign n14253 = n13560 & n13587;
  assign n14254 = ~n13581 & ~n13596;
  assign n14255 = ~n14253 & ~n14254;
  assign n14256 = ~n13515 & n13585;
  assign n14257 = n13578 & ~n14256;
  assign n14258 = ~n13604 & n14250;
  assign n14259 = n13561 & ~n14258;
  assign n14260 = ~n14257 & ~n14259;
  assign n14261 = ~n13577 & ~n13608;
  assign n14262 = n13581 & ~n14261;
  assign n14265 = ~n13599 & ~n13604;
  assign n14263 = ~n13573 & ~n13604;
  assign n14264 = n13600 & n14263;
  assign n14266 = n14265 ^ n14264;
  assign n14267 = n14265 ^ n13527;
  assign n14268 = n14267 ^ n14265;
  assign n14269 = n14266 & ~n14268;
  assign n14270 = n14269 ^ n14265;
  assign n14271 = n13560 & ~n14270;
  assign n14272 = ~n14262 & ~n14271;
  assign n14273 = n14260 & n14272;
  assign n14274 = n14255 & n14273;
  assign n14275 = n14252 & n14274;
  assign n14276 = n14246 & n14275;
  assign n14277 = n13570 & n14276;
  assign n14278 = n14277 ^ n10331;
  assign n14279 = n14278 ^ x94;
  assign n14280 = ~n13928 & ~n13934;
  assign n14281 = ~n13938 & n14280;
  assign n14282 = n13814 & ~n14281;
  assign n14283 = n13856 & n13895;
  assign n14284 = ~n13934 & ~n14283;
  assign n14285 = n13894 & ~n14284;
  assign n14286 = ~n13887 & n13944;
  assign n14287 = n13889 & ~n14286;
  assign n14288 = ~n14285 & ~n14287;
  assign n14289 = n13814 & n13897;
  assign n14290 = ~n13905 & ~n13938;
  assign n14291 = n13930 & n14290;
  assign n14292 = n13911 & ~n14291;
  assign n14293 = n13814 & n13942;
  assign n14294 = ~n13929 & ~n14283;
  assign n14295 = n13901 & n14294;
  assign n14296 = n14295 ^ n13813;
  assign n14297 = n14296 ^ n14295;
  assign n14298 = n13925 & n13936;
  assign n14299 = n14298 ^ n14295;
  assign n14300 = n14297 & n14299;
  assign n14301 = n14300 ^ n14295;
  assign n14302 = ~n13781 & ~n14301;
  assign n14303 = n13935 ^ n13781;
  assign n14304 = ~n13884 & n13891;
  assign n14305 = ~n13908 & ~n14304;
  assign n14306 = n14305 ^ n13929;
  assign n14307 = n13929 ^ n13813;
  assign n14308 = n14307 ^ n13929;
  assign n14309 = ~n14306 & n14308;
  assign n14310 = n14309 ^ n13929;
  assign n14311 = n14310 ^ n13935;
  assign n14312 = ~n14303 & n14311;
  assign n14313 = n14312 ^ n14309;
  assign n14314 = n14313 ^ n13929;
  assign n14315 = n14314 ^ n13781;
  assign n14316 = ~n13935 & ~n14315;
  assign n14317 = n14316 ^ n13935;
  assign n14318 = n14317 ^ n13781;
  assign n14319 = ~n14302 & n14318;
  assign n14320 = ~n14293 & n14319;
  assign n14321 = ~n13888 & n14320;
  assign n14322 = ~n14292 & n14321;
  assign n14323 = ~n14289 & n14322;
  assign n14324 = n14288 & n14323;
  assign n14325 = n13903 & n14324;
  assign n14326 = ~n14282 & n14325;
  assign n14327 = n14326 ^ n12364;
  assign n14328 = n14327 ^ x69;
  assign n14329 = n14279 & ~n14328;
  assign n14330 = n14243 & n14329;
  assign n14331 = n14171 & n14330;
  assign n14332 = n14139 & ~n14170;
  assign n14333 = n14201 & n14242;
  assign n14334 = ~n14279 & n14328;
  assign n14335 = n14333 & n14334;
  assign n14336 = ~n14201 & ~n14242;
  assign n14337 = n14334 & n14336;
  assign n14338 = ~n14335 & ~n14337;
  assign n14339 = n14332 & ~n14338;
  assign n14340 = ~n14331 & ~n14339;
  assign n14341 = n14139 & n14170;
  assign n14342 = ~n14139 & ~n14170;
  assign n14343 = ~n14341 & ~n14342;
  assign n14344 = n14243 & n14334;
  assign n14345 = ~n14343 & n14344;
  assign n14346 = n14329 & n14336;
  assign n14347 = ~n14170 & n14346;
  assign n14348 = ~n14345 & ~n14347;
  assign n14349 = n14201 & ~n14242;
  assign n14350 = n14279 & n14328;
  assign n14351 = n14349 & n14350;
  assign n14352 = n14336 & n14350;
  assign n14353 = ~n14346 & ~n14352;
  assign n14354 = ~n14351 & n14353;
  assign n14355 = n14171 & ~n14354;
  assign n14356 = ~n14279 & ~n14328;
  assign n14357 = n14336 & n14356;
  assign n14358 = n14243 & n14356;
  assign n14359 = n14349 & n14356;
  assign n14360 = ~n14358 & ~n14359;
  assign n14361 = ~n14357 & n14360;
  assign n14362 = n14341 & ~n14361;
  assign n14363 = ~n14355 & ~n14362;
  assign n14364 = n14348 & n14363;
  assign n14365 = n14333 & n14356;
  assign n14366 = n14332 & n14365;
  assign n14367 = n14334 & n14349;
  assign n14368 = ~n14358 & ~n14367;
  assign n14369 = n14342 & ~n14368;
  assign n14370 = n14201 & n14329;
  assign n14371 = n14243 & n14350;
  assign n14372 = ~n14352 & ~n14371;
  assign n14373 = ~n14370 & n14372;
  assign n14374 = n14341 & ~n14373;
  assign n14375 = n14329 & n14333;
  assign n14376 = n14329 & n14349;
  assign n14377 = ~n14351 & ~n14371;
  assign n14378 = ~n14376 & n14377;
  assign n14379 = ~n14375 & n14378;
  assign n14380 = n14342 & ~n14379;
  assign n14381 = ~n14374 & ~n14380;
  assign n14382 = ~n14359 & ~n14365;
  assign n14383 = n14338 & n14382;
  assign n14384 = n14171 & ~n14383;
  assign n14385 = n14333 & n14350;
  assign n14386 = ~n14376 & ~n14385;
  assign n14387 = ~n14330 & ~n14341;
  assign n14388 = n14386 & n14387;
  assign n14389 = ~n14352 & n14388;
  assign n14390 = n14332 & ~n14389;
  assign n14391 = ~n14384 & ~n14390;
  assign n14392 = n14381 & n14391;
  assign n14393 = ~n14369 & n14392;
  assign n14394 = ~n14366 & n14393;
  assign n14395 = n14364 & n14394;
  assign n14396 = n14340 & n14395;
  assign n14397 = n14396 ^ n13340;
  assign n14398 = n14397 ^ x66;
  assign n14399 = n14006 & ~n14398;
  assign n14400 = n12716 ^ x86;
  assign n14401 = n14278 ^ x100;
  assign n14402 = n14400 & ~n14401;
  assign n14403 = n14138 ^ x101;
  assign n14404 = n13779 ^ x124;
  assign n14405 = n14403 & n14404;
  assign n14406 = n13342 ^ n13341;
  assign n14407 = n13394 & ~n14406;
  assign n14408 = n13346 & n13404;
  assign n14409 = ~n14407 & ~n14408;
  assign n14410 = n13343 & n13393;
  assign n14411 = n13355 ^ n13341;
  assign n14412 = n14411 ^ n13355;
  assign n14413 = ~n13349 & ~n13372;
  assign n14414 = n14413 ^ n13355;
  assign n14415 = n14412 & ~n14414;
  assign n14416 = n14415 ^ n13355;
  assign n14417 = ~n13342 & n14416;
  assign n14418 = ~n14410 & ~n14417;
  assign n14419 = n13344 & n13348;
  assign n14420 = n13384 & ~n13405;
  assign n14421 = ~n14419 & ~n14420;
  assign n14422 = n13341 & ~n13399;
  assign n14423 = ~n13377 & n13403;
  assign n14424 = n13343 & ~n14423;
  assign n14425 = n13374 & ~n13388;
  assign n14426 = ~n13358 & n13368;
  assign n14427 = n14425 & n14426;
  assign n14428 = n13371 & ~n14427;
  assign n14429 = ~n14424 & ~n14428;
  assign n14430 = ~n14422 & n14429;
  assign n14431 = n14421 & n14430;
  assign n14432 = n14418 & n14431;
  assign n14433 = n13387 & n14432;
  assign n14434 = n13364 & n14433;
  assign n14435 = n14409 & n14434;
  assign n14436 = ~n13345 & n14435;
  assign n14437 = n14436 ^ n10840;
  assign n14438 = n14437 ^ x68;
  assign n14439 = n13012 ^ x92;
  assign n14440 = n13883 ^ x109;
  assign n14441 = ~n14439 & n14440;
  assign n14442 = n13812 ^ x68;
  assign n14443 = n12050 & ~n13244;
  assign n14444 = n11904 & ~n12058;
  assign n14445 = ~n14443 & ~n14444;
  assign n14446 = n12024 & ~n13242;
  assign n14447 = ~n12022 & n12039;
  assign n14448 = n12062 & ~n14447;
  assign n14449 = ~n12037 & n13439;
  assign n14450 = n12031 & ~n14449;
  assign n14451 = n12063 ^ n11903;
  assign n14454 = ~n12055 & ~n13245;
  assign n14452 = ~n12033 & ~n12056;
  assign n14453 = ~n12022 & n14452;
  assign n14455 = n14454 ^ n14453;
  assign n14456 = n14454 ^ n11872;
  assign n14457 = n14456 ^ n14454;
  assign n14458 = n14455 & ~n14457;
  assign n14459 = n14458 ^ n14454;
  assign n14460 = n14459 ^ n12063;
  assign n14461 = ~n14451 & ~n14460;
  assign n14462 = n14461 ^ n14458;
  assign n14463 = n14462 ^ n14454;
  assign n14464 = n14463 ^ n11903;
  assign n14465 = ~n12063 & n14464;
  assign n14466 = n14465 ^ n12063;
  assign n14467 = n14466 ^ n11903;
  assign n14468 = ~n14450 & n14467;
  assign n14469 = n12046 & ~n13241;
  assign n14470 = n14469 ^ n11872;
  assign n14471 = n14470 ^ n14469;
  assign n14472 = ~n12033 & n12076;
  assign n14473 = n14472 ^ n14469;
  assign n14474 = n14471 & n14473;
  assign n14475 = n14474 ^ n14469;
  assign n14476 = ~n11903 & ~n14475;
  assign n14477 = n14468 & ~n14476;
  assign n14478 = n12029 & n14477;
  assign n14479 = ~n14448 & n14478;
  assign n14480 = ~n14446 & n14479;
  assign n14481 = n14445 & n14480;
  assign n14482 = n12048 & n14481;
  assign n14483 = ~n12030 & n14482;
  assign n14484 = n14483 ^ n11208;
  assign n14485 = n14484 ^ x85;
  assign n14486 = n14442 & n14485;
  assign n14487 = n12965 ^ x110;
  assign n14488 = n12586 & n12592;
  assign n14489 = n12579 & n12611;
  assign n14490 = ~n14488 & ~n14489;
  assign n14491 = n12581 & ~n12629;
  assign n14492 = n12594 & n12600;
  assign n14493 = ~n12603 & n12610;
  assign n14494 = n12604 & ~n14493;
  assign n14495 = n12533 ^ n12497;
  assign n14496 = n14495 ^ n12558;
  assign n14497 = n14496 ^ n12533;
  assign n14498 = n14497 ^ n14496;
  assign n14499 = n14496 ^ n12558;
  assign n14500 = ~n14498 & n14499;
  assign n14501 = n14500 ^ n14496;
  assign n14502 = n12557 & n14501;
  assign n14503 = n14502 ^ n14496;
  assign n14504 = n12603 & n14503;
  assign n14505 = ~n14494 & ~n14504;
  assign n14506 = ~n12596 & n12634;
  assign n14507 = n12581 & ~n14506;
  assign n14508 = ~n12584 & n13491;
  assign n14509 = ~n12600 & n14508;
  assign n14510 = ~n12613 & n12632;
  assign n14511 = ~n12605 & n14510;
  assign n14512 = ~n12586 & n14511;
  assign n14513 = ~n14509 & ~n14512;
  assign n14514 = ~n12621 & ~n14513;
  assign n14515 = ~n12610 & ~n14514;
  assign n14516 = ~n14507 & ~n14515;
  assign n14517 = n14505 & n14516;
  assign n14518 = ~n14492 & n14517;
  assign n14519 = ~n14491 & n14518;
  assign n14520 = n14490 & n14519;
  assign n14521 = n12591 & n14520;
  assign n14522 = n14521 ^ n11237;
  assign n14523 = n14522 ^ x70;
  assign n14524 = n14487 & ~n14523;
  assign n14525 = n14486 & n14524;
  assign n14526 = n14441 & n14525;
  assign n14527 = ~n14439 & ~n14440;
  assign n14528 = n14442 & ~n14485;
  assign n14529 = n14487 & n14523;
  assign n14530 = n14528 & n14529;
  assign n14531 = ~n14442 & n14485;
  assign n14532 = n14529 & n14531;
  assign n14533 = ~n14530 & ~n14532;
  assign n14534 = n14527 & ~n14533;
  assign n14535 = n14525 & n14527;
  assign n14536 = n14439 & n14440;
  assign n14537 = ~n14527 & ~n14536;
  assign n14538 = ~n14442 & ~n14485;
  assign n14539 = ~n14487 & ~n14523;
  assign n14540 = n14538 & n14539;
  assign n14541 = n14486 & n14539;
  assign n14542 = ~n14540 & ~n14541;
  assign n14543 = ~n14537 & ~n14542;
  assign n14544 = ~n14535 & ~n14543;
  assign n14549 = ~n14487 & n14523;
  assign n14550 = n14486 & n14549;
  assign n14545 = n14529 & n14538;
  assign n14546 = n14524 & n14528;
  assign n14547 = ~n14545 & ~n14546;
  assign n14548 = ~n14532 & n14547;
  assign n14551 = n14550 ^ n14548;
  assign n14552 = n14551 ^ n14550;
  assign n14553 = n14550 ^ n14439;
  assign n14554 = n14553 ^ n14550;
  assign n14555 = ~n14552 & ~n14554;
  assign n14556 = n14555 ^ n14550;
  assign n14557 = n14440 & n14556;
  assign n14558 = n14557 ^ n14550;
  assign n14559 = n14544 & ~n14558;
  assign n14560 = n14538 & n14549;
  assign n14561 = n14528 & n14539;
  assign n14562 = ~n14560 & ~n14561;
  assign n14563 = n14536 & ~n14562;
  assign n14564 = n14439 & ~n14440;
  assign n14565 = n14531 & n14539;
  assign n14566 = n14528 & n14549;
  assign n14567 = n14531 & n14549;
  assign n14568 = ~n14566 & ~n14567;
  assign n14569 = ~n14565 & n14568;
  assign n14570 = n14564 & ~n14569;
  assign n14571 = n14441 & ~n14542;
  assign n14572 = n14524 & n14531;
  assign n14573 = n14572 ^ n14536;
  assign n14574 = n14572 ^ n14564;
  assign n14575 = n14574 ^ n14564;
  assign n14576 = n14486 & n14529;
  assign n14577 = n14576 ^ n14564;
  assign n14578 = ~n14575 & ~n14577;
  assign n14579 = n14578 ^ n14564;
  assign n14580 = n14573 & n14579;
  assign n14581 = n14580 ^ n14536;
  assign n14582 = ~n14571 & ~n14581;
  assign n14583 = ~n14560 & ~n14566;
  assign n14584 = n14441 & ~n14583;
  assign n14585 = n14527 & ~n14547;
  assign n14586 = ~n14584 & ~n14585;
  assign n14587 = n14564 ^ n14536;
  assign n14588 = n14524 & n14538;
  assign n14589 = n14547 & ~n14588;
  assign n14590 = n14589 ^ n14533;
  assign n14591 = n14564 ^ n14533;
  assign n14592 = n14591 ^ n14533;
  assign n14593 = ~n14590 & n14592;
  assign n14594 = n14593 ^ n14533;
  assign n14595 = n14587 & n14594;
  assign n14596 = n14595 ^ n14536;
  assign n14597 = n14586 & ~n14596;
  assign n14598 = n14582 & n14597;
  assign n14599 = ~n14570 & n14598;
  assign n14600 = ~n14563 & n14599;
  assign n14601 = n14559 & n14600;
  assign n14602 = ~n14534 & n14601;
  assign n14603 = ~n14526 & n14602;
  assign n14604 = n14603 ^ n11307;
  assign n14605 = n14604 ^ x118;
  assign n14606 = ~n14438 & n14605;
  assign n14607 = n14405 & n14606;
  assign n14608 = n14402 & n14607;
  assign n14609 = ~n14400 & ~n14401;
  assign n14610 = ~n14403 & n14404;
  assign n14611 = n14438 & ~n14605;
  assign n14612 = n14610 & n14611;
  assign n14613 = ~n14438 & ~n14605;
  assign n14614 = n14405 & n14613;
  assign n14615 = ~n14612 & ~n14614;
  assign n14616 = n14609 & ~n14615;
  assign n14617 = ~n14608 & ~n14616;
  assign n14618 = ~n14403 & ~n14404;
  assign n14619 = n14402 & n14618;
  assign n14620 = n14438 & n14605;
  assign n14621 = n14619 & n14620;
  assign n14622 = n14400 & n14401;
  assign n14623 = ~n14609 & ~n14622;
  assign n14624 = n14403 & ~n14404;
  assign n14625 = n14611 & n14624;
  assign n14626 = n14623 & n14625;
  assign n14627 = ~n14400 & n14401;
  assign n14628 = n14610 & n14613;
  assign n14629 = n14627 & n14628;
  assign n14630 = ~n14626 & ~n14629;
  assign n14631 = ~n14621 & n14630;
  assign n14632 = n14620 & n14624;
  assign n14633 = n14627 & n14632;
  assign n14634 = n14622 & n14632;
  assign n14635 = n14618 & n14620;
  assign n14636 = n14627 & n14635;
  assign n14637 = ~n14634 & ~n14636;
  assign n14638 = ~n14633 & n14637;
  assign n14639 = n14613 & n14624;
  assign n14640 = n14627 & n14639;
  assign n14641 = n14605 ^ n14438;
  assign n14642 = n14622 ^ n14605;
  assign n14643 = n14642 ^ n14622;
  assign n14644 = n14622 ^ n14609;
  assign n14645 = n14643 & n14644;
  assign n14646 = n14645 ^ n14622;
  assign n14647 = ~n14641 & n14646;
  assign n14648 = n14618 & n14647;
  assign n14649 = ~n14640 & ~n14648;
  assign n14650 = ~n14404 & n14606;
  assign n14651 = n14405 & n14611;
  assign n14652 = ~n14614 & ~n14651;
  assign n14653 = ~n14628 & n14652;
  assign n14654 = ~n14650 & n14653;
  assign n14655 = n14402 & ~n14654;
  assign n14656 = n14405 & n14620;
  assign n14657 = n14606 & n14610;
  assign n14658 = ~n14656 & ~n14657;
  assign n14659 = ~n14607 & n14658;
  assign n14660 = n14609 & ~n14659;
  assign n14661 = ~n14651 & ~n14657;
  assign n14662 = ~n14612 & n14661;
  assign n14663 = n14627 & ~n14662;
  assign n14664 = ~n14660 & ~n14663;
  assign n14665 = ~n14655 & n14664;
  assign n14666 = n14606 & n14624;
  assign n14667 = n14611 & n14618;
  assign n14668 = ~n14666 & ~n14667;
  assign n14669 = n14668 ^ n14622;
  assign n14670 = n14668 ^ n14609;
  assign n14671 = n14670 ^ n14609;
  assign n14672 = n14610 & n14620;
  assign n14673 = ~n14607 & ~n14672;
  assign n14674 = ~n14614 & ~n14656;
  assign n14675 = n14673 & n14674;
  assign n14676 = n14675 ^ n14609;
  assign n14677 = n14671 & n14676;
  assign n14678 = n14677 ^ n14609;
  assign n14679 = ~n14669 & n14678;
  assign n14680 = n14679 ^ n14622;
  assign n14681 = n14665 & ~n14680;
  assign n14682 = n14649 & n14681;
  assign n14683 = n14638 & n14682;
  assign n14684 = n14631 & n14683;
  assign n14685 = n14617 & n14684;
  assign n14686 = n14685 ^ n13668;
  assign n14687 = n14686 ^ x106;
  assign n14688 = n13734 & ~n14182;
  assign n14689 = ~n13722 & ~n13735;
  assign n14690 = ~n13754 & ~n14689;
  assign n14691 = n13738 & ~n13754;
  assign n14692 = ~n13629 & n13714;
  assign n14693 = ~n14691 & ~n14692;
  assign n14694 = ~n13710 & ~n13762;
  assign n14695 = n13705 & ~n14694;
  assign n14696 = ~n13722 & ~n13751;
  assign n14697 = ~n13707 & n14696;
  assign n14698 = n13742 & n14697;
  assign n14699 = n13737 & ~n14698;
  assign n14700 = ~n14695 & ~n14699;
  assign n14701 = n14693 & n14700;
  assign n14702 = ~n14690 & n14701;
  assign n14703 = ~n14688 & n14702;
  assign n14704 = n13701 & n13709;
  assign n14705 = n13742 & ~n14704;
  assign n14706 = ~n13730 & n14705;
  assign n14707 = n14706 ^ n13729;
  assign n14708 = n14707 ^ n13729;
  assign n14709 = n13729 ^ n13628;
  assign n14710 = n14709 ^ n13729;
  assign n14711 = ~n14708 & n14710;
  assign n14712 = n14711 ^ n13729;
  assign n14713 = ~n13629 & n14712;
  assign n14714 = n14713 ^ n13729;
  assign n14715 = n14703 & ~n14714;
  assign n14716 = ~n13704 & n14715;
  assign n14717 = n14174 & n14716;
  assign n14718 = ~n13756 & n14717;
  assign n14719 = n14718 ^ n11724;
  assign n14720 = n14719 ^ x104;
  assign n14721 = ~n14540 & ~n14566;
  assign n14722 = n14564 & ~n14721;
  assign n14723 = ~n14541 & ~n14567;
  assign n14724 = n14536 & ~n14723;
  assign n14725 = ~n14722 & ~n14724;
  assign n14726 = ~n14537 & n14561;
  assign n14727 = ~n14545 & ~n14572;
  assign n14728 = ~n14588 & n14727;
  assign n14729 = n14441 & ~n14728;
  assign n14730 = ~n14726 & ~n14729;
  assign n14731 = n14572 ^ n14439;
  assign n14732 = n14731 ^ n14572;
  assign n14733 = n14572 ^ n14565;
  assign n14734 = n14733 ^ n14572;
  assign n14735 = n14732 & n14734;
  assign n14736 = n14735 ^ n14572;
  assign n14737 = n14440 & n14736;
  assign n14738 = n14737 ^ n14572;
  assign n14739 = n14730 & ~n14738;
  assign n14740 = n14550 & n14564;
  assign n14741 = ~n14541 & ~n14560;
  assign n14742 = n14527 & ~n14741;
  assign n14743 = ~n14532 & ~n14546;
  assign n14744 = ~n14576 & n14743;
  assign n14745 = ~n14588 & n14744;
  assign n14746 = n14536 & ~n14745;
  assign n14747 = ~n14550 & ~n14567;
  assign n14748 = n14721 & n14747;
  assign n14749 = n14441 & ~n14748;
  assign n14750 = ~n14525 & ~n14588;
  assign n14751 = n14533 & n14750;
  assign n14752 = n14564 & ~n14751;
  assign n14753 = n14548 & ~n14576;
  assign n14754 = n14527 & ~n14753;
  assign n14755 = ~n14752 & ~n14754;
  assign n14756 = ~n14749 & n14755;
  assign n14757 = ~n14746 & n14756;
  assign n14758 = ~n14742 & n14757;
  assign n14759 = ~n14740 & n14758;
  assign n14760 = n14739 & n14759;
  assign n14761 = ~n14526 & n14760;
  assign n14762 = n14725 & n14761;
  assign n14763 = n14762 ^ n11760;
  assign n14764 = n14763 ^ x66;
  assign n14765 = ~n14720 & ~n14764;
  assign n14766 = n12658 & n12666;
  assign n14767 = n14205 & ~n14766;
  assign n14768 = n11846 & n12651;
  assign n14769 = n12662 & n12671;
  assign n14770 = ~n14768 & ~n14769;
  assign n14771 = n12688 & ~n12691;
  assign n14772 = n11847 & ~n14771;
  assign n14773 = n12684 & ~n12687;
  assign n14774 = n12666 & ~n14773;
  assign n14775 = ~n14772 & ~n14774;
  assign n14776 = ~n11846 & n12697;
  assign n14777 = ~n12681 & n12704;
  assign n14778 = n12652 & ~n14777;
  assign n14779 = ~n14776 & ~n14778;
  assign n14780 = n14775 & n14779;
  assign n14781 = n14770 & n14780;
  assign n14782 = n12660 & n14781;
  assign n14783 = n12675 & n14782;
  assign n14784 = n14767 & n14783;
  assign n14785 = ~n12648 & n14784;
  assign n14786 = ~n14212 & n14785;
  assign n14787 = n14786 ^ n11415;
  assign n14788 = n14787 ^ x64;
  assign n14789 = n14263 ^ n13513;
  assign n14790 = n14789 ^ n14263;
  assign n14791 = n14263 ^ n13578;
  assign n14792 = n14791 ^ n14263;
  assign n14793 = n14790 & ~n14792;
  assign n14794 = n14793 ^ n14263;
  assign n14795 = ~n13571 & ~n14794;
  assign n14796 = n14795 ^ n14263;
  assign n14798 = ~n13567 & ~n13603;
  assign n14797 = ~n13573 & n14250;
  assign n14799 = n14798 ^ n14797;
  assign n14800 = n14799 ^ n14798;
  assign n14801 = n14798 ^ n13527;
  assign n14802 = n14801 ^ n14798;
  assign n14803 = ~n14800 & ~n14802;
  assign n14804 = n14803 ^ n14798;
  assign n14805 = ~n13560 & ~n14804;
  assign n14806 = n14805 ^ n14798;
  assign n14807 = n14796 & n14806;
  assign n14808 = n13563 & n13599;
  assign n14809 = n13589 & n13607;
  assign n14810 = n13578 & ~n14809;
  assign n14811 = n13568 & ~n13586;
  assign n14812 = n13578 & ~n14811;
  assign n14813 = n13585 & n14261;
  assign n14814 = n13563 & ~n14813;
  assign n14815 = ~n14812 & ~n14814;
  assign n14816 = ~n13584 & n13596;
  assign n14817 = n13561 & ~n14816;
  assign n14818 = ~n13587 & n13609;
  assign n14819 = ~n13583 & n14818;
  assign n14820 = n13571 & ~n14819;
  assign n14821 = ~n14817 & ~n14820;
  assign n14822 = n14815 & n14821;
  assign n14823 = n14246 & n14822;
  assign n14824 = ~n14810 & n14823;
  assign n14825 = ~n14808 & n14824;
  assign n14826 = n14807 & n14825;
  assign n14827 = n14826 ^ n11449;
  assign n14828 = n14827 ^ x90;
  assign n14829 = n14788 & ~n14828;
  assign n14830 = n13136 & n13177;
  assign n14831 = ~n13182 & n14145;
  assign n14832 = ~n13164 & n14831;
  assign n14833 = n12967 & ~n14832;
  assign n14834 = ~n14830 & ~n14833;
  assign n14835 = n13125 & ~n13188;
  assign n14836 = n13165 & n14155;
  assign n14837 = ~n13148 & n14836;
  assign n14838 = n13149 & ~n14837;
  assign n14839 = ~n13140 & n13154;
  assign n14840 = ~n13148 & n14839;
  assign n14841 = ~n13125 & n14840;
  assign n14842 = n13142 & ~n13153;
  assign n14843 = ~n13152 & n14842;
  assign n14844 = ~n13136 & n14843;
  assign n14845 = ~n14841 & ~n14844;
  assign n14846 = n13150 & n14845;
  assign n14847 = ~n14838 & ~n14846;
  assign n14848 = ~n14835 & n14847;
  assign n14849 = n14834 & n14848;
  assign n14850 = n13162 ^ n13140;
  assign n14851 = n14850 ^ n13162;
  assign n14852 = n13162 ^ n12966;
  assign n14853 = n14852 ^ n13162;
  assign n14854 = n14851 & n14853;
  assign n14855 = n14854 ^ n13162;
  assign n14856 = n12838 & n14855;
  assign n14857 = n14856 ^ n13162;
  assign n14858 = n14849 & ~n14857;
  assign n14859 = n13161 & n14858;
  assign n14860 = ~n13158 & n14859;
  assign n14861 = n14142 & n14860;
  assign n14862 = n14861 ^ n11693;
  assign n14863 = n14862 ^ x81;
  assign n14864 = ~n13935 & ~n13943;
  assign n14865 = n13894 & ~n14864;
  assign n14866 = n13887 & n13894;
  assign n14867 = n13813 ^ n13781;
  assign n14868 = n13886 & n13891;
  assign n14869 = ~n13926 & ~n14868;
  assign n14870 = n14867 & ~n14869;
  assign n14871 = n13897 & n14867;
  assign n14872 = n13939 & n14294;
  assign n14873 = n13894 & ~n14872;
  assign n14874 = ~n14871 & ~n14873;
  assign n14875 = n13814 & ~n14290;
  assign n14876 = n13925 & ~n13942;
  assign n14877 = n13939 & n14876;
  assign n14878 = n13911 & ~n14877;
  assign n14879 = n13814 & n13908;
  assign n14880 = ~n13892 & ~n13935;
  assign n14881 = n14280 & n14880;
  assign n14882 = n14294 & n14881;
  assign n14883 = ~n13943 & n14882;
  assign n14884 = n13889 & ~n14883;
  assign n14885 = ~n14879 & ~n14884;
  assign n14886 = ~n14878 & n14885;
  assign n14887 = ~n14875 & n14886;
  assign n14888 = n14874 & n14887;
  assign n14889 = ~n14870 & n14888;
  assign n14890 = ~n14866 & n14889;
  assign n14891 = n13907 & n14890;
  assign n14892 = ~n14865 & n14891;
  assign n14893 = ~n14293 & n14892;
  assign n14894 = ~n13888 & n14893;
  assign n14895 = n14894 ^ n11552;
  assign n14896 = n14895 ^ x107;
  assign n14897 = n14863 & n14896;
  assign n14898 = n14829 & n14897;
  assign n14899 = n14765 & n14898;
  assign n14900 = n14720 & n14764;
  assign n14901 = ~n14863 & n14896;
  assign n14902 = n14829 & n14901;
  assign n14903 = n14900 & n14902;
  assign n14904 = ~n14899 & ~n14903;
  assign n14905 = n14720 & ~n14764;
  assign n14906 = ~n14788 & n14828;
  assign n14907 = n14863 & ~n14896;
  assign n14908 = n14906 & n14907;
  assign n14909 = n14905 & n14908;
  assign n14910 = ~n14720 & n14764;
  assign n14911 = n14829 & n14907;
  assign n14912 = ~n14788 & ~n14828;
  assign n14913 = ~n14863 & ~n14896;
  assign n14914 = n14912 & n14913;
  assign n14915 = ~n14911 & ~n14914;
  assign n14916 = n14910 & ~n14915;
  assign n14917 = ~n14909 & ~n14916;
  assign n14918 = n14904 & n14917;
  assign n14919 = n14788 & n14828;
  assign n14920 = n14897 & n14919;
  assign n14921 = n14905 & n14920;
  assign n14922 = n14897 & n14912;
  assign n14923 = n14900 & n14922;
  assign n14924 = ~n14921 & ~n14923;
  assign n14925 = ~n14765 & ~n14900;
  assign n14926 = n14907 & n14912;
  assign n14927 = ~n14925 & n14926;
  assign n14928 = n14901 & n14912;
  assign n14929 = n14906 & n14913;
  assign n14930 = ~n14928 & ~n14929;
  assign n14931 = n14765 & ~n14930;
  assign n14932 = ~n14927 & ~n14931;
  assign n14933 = ~n14898 & ~n14902;
  assign n14934 = n14910 & ~n14933;
  assign n14935 = ~n14902 & ~n14926;
  assign n14936 = n14930 & n14935;
  assign n14937 = n14905 & ~n14936;
  assign n14938 = n14897 & n14906;
  assign n14939 = ~n14920 & ~n14938;
  assign n14940 = n14913 & n14919;
  assign n14941 = n14907 & n14919;
  assign n14942 = ~n14940 & ~n14941;
  assign n14943 = n14939 & n14942;
  assign n14944 = n14900 & ~n14943;
  assign n14945 = ~n14937 & ~n14944;
  assign n14948 = n14901 & n14919;
  assign n14949 = ~n14938 & ~n14948;
  assign n14950 = n14942 & n14949;
  assign n14946 = n14938 ^ n14906;
  assign n14947 = ~n14940 & ~n14946;
  assign n14951 = n14950 ^ n14947;
  assign n14952 = n14950 ^ n14764;
  assign n14953 = n14952 ^ n14950;
  assign n14954 = n14951 & n14953;
  assign n14955 = n14954 ^ n14950;
  assign n14956 = ~n14720 & ~n14955;
  assign n14957 = n14945 & ~n14956;
  assign n14958 = ~n14934 & n14957;
  assign n14959 = n14932 & n14958;
  assign n14960 = n14914 ^ n14764;
  assign n14961 = n14960 ^ n14914;
  assign n14962 = n14901 & n14906;
  assign n14963 = ~n14941 & ~n14962;
  assign n14964 = n14963 ^ n14914;
  assign n14965 = ~n14961 & ~n14964;
  assign n14966 = n14965 ^ n14914;
  assign n14967 = n14720 & n14966;
  assign n14968 = n14959 & ~n14967;
  assign n14969 = n14924 & n14968;
  assign n14970 = n14918 & n14969;
  assign n14971 = n14970 ^ n13699;
  assign n14972 = n14971 ^ x80;
  assign n14973 = n14687 & n14972;
  assign n14974 = n14399 & n14973;
  assign n14975 = n14006 & n14398;
  assign n14976 = n14973 & n14975;
  assign n14977 = ~n14687 & n14972;
  assign n14978 = n14399 & n14977;
  assign n14979 = ~n14976 & ~n14978;
  assign n14980 = ~n14106 & n14123;
  assign n14981 = ~n14097 & n14109;
  assign n14982 = ~n14980 & ~n14981;
  assign n14983 = n14009 & ~n14121;
  assign n14984 = n14099 & n14134;
  assign n14985 = ~n14983 & ~n14984;
  assign n14986 = n14982 & n14985;
  assign n14987 = n14986 ^ n11915;
  assign n14988 = n14987 ^ x102;
  assign n14989 = n14169 ^ x85;
  assign n14990 = ~n14988 & n14989;
  assign n14991 = ~n13381 & n13400;
  assign n14992 = n13343 & ~n14991;
  assign n14993 = ~n13376 & n14426;
  assign n14994 = n13384 & ~n14993;
  assign n14995 = ~n14992 & ~n14994;
  assign n14996 = ~n13388 & ~n13393;
  assign n14997 = ~n14406 & ~n14996;
  assign n14998 = ~n13381 & ~n13404;
  assign n14999 = ~n13377 & n14998;
  assign n15000 = n13371 & ~n14999;
  assign n15001 = ~n13373 & n13406;
  assign n15002 = ~n13355 & n15001;
  assign n15003 = n13384 & ~n15002;
  assign n15004 = ~n15000 & ~n15003;
  assign n15005 = ~n14997 & n15004;
  assign n15006 = n14995 & n15005;
  assign n15007 = ~n13363 & n15006;
  assign n15008 = n13380 & n15007;
  assign n15009 = n13370 & n15008;
  assign n15010 = n14409 & n15009;
  assign n15011 = n15010 ^ n11957;
  assign n15012 = n15011 ^ x75;
  assign n15013 = n13513 & n13560;
  assign n15014 = n13571 & ~n14250;
  assign n15015 = ~n15013 & ~n15014;
  assign n15016 = n13563 & n13577;
  assign n15017 = n13590 & n14263;
  assign n15018 = n13561 & ~n15017;
  assign n15019 = ~n13563 & n13597;
  assign n15020 = ~n13571 & n14816;
  assign n15021 = ~n15019 & ~n15020;
  assign n15022 = n15021 ^ n13527;
  assign n15023 = n15022 ^ n15021;
  assign n15024 = n13607 & ~n13608;
  assign n15025 = n13568 & n15024;
  assign n15026 = n15025 ^ n15021;
  assign n15027 = n15026 ^ n15021;
  assign n15028 = n15023 & ~n15027;
  assign n15029 = n15028 ^ n15021;
  assign n15030 = ~n13560 & n15029;
  assign n15031 = n15030 ^ n15021;
  assign n15032 = ~n15018 & ~n15031;
  assign n15033 = ~n15016 & n15032;
  assign n15034 = n15015 & n15033;
  assign n15035 = ~n14244 & n15034;
  assign n15036 = n13580 & n15035;
  assign n15037 = n14252 & n15036;
  assign n15038 = n13570 & n15037;
  assign n15039 = n15038 ^ n11985;
  assign n15040 = n15039 ^ x92;
  assign n15041 = n15012 & ~n15040;
  assign n15042 = n14990 & n15041;
  assign n15043 = n14988 & n14989;
  assign n15044 = ~n15012 & ~n15040;
  assign n15045 = n15043 & n15044;
  assign n15046 = ~n15042 & ~n15045;
  assign n15047 = n14241 ^ x125;
  assign n15048 = ~n14545 & ~n14576;
  assign n15049 = n14564 & ~n15048;
  assign n15050 = ~n14550 & ~n14565;
  assign n15051 = n14441 & ~n15050;
  assign n15052 = ~n15049 & ~n15051;
  assign n15053 = ~n14566 & ~n14572;
  assign n15054 = ~n14537 & ~n15053;
  assign n15055 = ~n14540 & n14548;
  assign n15056 = n14536 & ~n15055;
  assign n15057 = ~n14530 & n14589;
  assign n15058 = ~n14560 & n15057;
  assign n15059 = n14441 & ~n15058;
  assign n15060 = ~n15056 & ~n15059;
  assign n15061 = ~n15054 & n15060;
  assign n15062 = n14564 & ~n14750;
  assign n15063 = n14561 ^ n14440;
  assign n15064 = n14565 ^ n14439;
  assign n15065 = n15064 ^ n14565;
  assign n15066 = n14542 & ~n14567;
  assign n15067 = n15066 ^ n14565;
  assign n15068 = ~n15065 & ~n15067;
  assign n15069 = n15068 ^ n14565;
  assign n15070 = n15069 ^ n14561;
  assign n15071 = n15063 & n15070;
  assign n15072 = n15071 ^ n15068;
  assign n15073 = n15072 ^ n14565;
  assign n15074 = n15073 ^ n14440;
  assign n15075 = ~n14561 & n15074;
  assign n15076 = n15075 ^ n14561;
  assign n15077 = n15076 ^ n14440;
  assign n15078 = ~n15062 & ~n15077;
  assign n15079 = n15061 & n15078;
  assign n15080 = n15052 & n15079;
  assign n15081 = ~n14534 & n15080;
  assign n15082 = ~n14526 & n15081;
  assign n15083 = n14725 & n15082;
  assign n15084 = n15083 ^ n11902;
  assign n15085 = n15084 ^ x116;
  assign n15086 = ~n15047 & n15085;
  assign n15087 = ~n15046 & n15086;
  assign n15088 = n15047 & n15085;
  assign n15089 = ~n15012 & n15040;
  assign n15090 = n15043 & n15089;
  assign n15091 = n14990 & n15089;
  assign n15092 = n15041 & n15043;
  assign n15093 = ~n15091 & ~n15092;
  assign n15094 = ~n15090 & n15093;
  assign n15095 = n15088 & ~n15094;
  assign n15096 = n14988 & ~n14989;
  assign n15097 = n15044 & n15096;
  assign n15098 = n15012 & n15040;
  assign n15099 = n15096 & n15098;
  assign n15100 = ~n15042 & ~n15099;
  assign n15101 = ~n15097 & n15100;
  assign n15102 = n15088 & ~n15101;
  assign n15103 = n15089 & n15096;
  assign n15104 = ~n14988 & ~n14989;
  assign n15105 = n15041 & n15104;
  assign n15106 = ~n15103 & ~n15105;
  assign n15107 = n15098 & n15104;
  assign n15108 = ~n15097 & ~n15107;
  assign n15109 = n15106 & n15108;
  assign n15110 = ~n15091 & n15109;
  assign n15111 = n15086 & ~n15110;
  assign n15112 = ~n15102 & ~n15111;
  assign n15114 = n15043 & n15098;
  assign n15113 = n15047 & ~n15085;
  assign n15115 = n15114 ^ n15113;
  assign n15116 = n15113 ^ n15086;
  assign n15117 = n15116 ^ n15086;
  assign n15118 = ~n15045 & n15106;
  assign n15119 = n15093 & n15118;
  assign n15120 = n15119 ^ n15086;
  assign n15121 = n15117 & n15120;
  assign n15122 = n15121 ^ n15086;
  assign n15123 = n15115 & ~n15122;
  assign n15124 = n15123 ^ n15114;
  assign n15125 = n15112 & ~n15124;
  assign n15128 = n15041 & n15096;
  assign n15129 = n15044 & n15104;
  assign n15130 = ~n15128 & ~n15129;
  assign n15126 = n15100 & n15109;
  assign n15127 = n15093 & n15126;
  assign n15131 = n15130 ^ n15127;
  assign n15132 = n15131 ^ n15130;
  assign n15133 = n15130 ^ n15085;
  assign n15134 = n15133 ^ n15130;
  assign n15135 = n15132 & ~n15134;
  assign n15136 = n15135 ^ n15130;
  assign n15137 = ~n15047 & ~n15136;
  assign n15138 = n15137 ^ n15130;
  assign n15139 = n15125 & n15138;
  assign n15140 = ~n15095 & n15139;
  assign n15141 = ~n15087 & n15140;
  assign n15142 = n15141 ^ n13455;
  assign n15143 = n15142 ^ x121;
  assign n15144 = n14058 & n14093;
  assign n15145 = n14091 & ~n14093;
  assign n15146 = ~n15144 & ~n15145;
  assign n15147 = ~n14086 & n15146;
  assign n15148 = ~n14101 & n15147;
  assign n15149 = n14109 & ~n15148;
  assign n15150 = ~n14010 & n14094;
  assign n15151 = n14118 & ~n15150;
  assign n15152 = n14009 & ~n15151;
  assign n15153 = ~n15149 & ~n15152;
  assign n15154 = n14058 & n14081;
  assign n15155 = n14114 & ~n15154;
  assign n15156 = ~n14102 & n15155;
  assign n15157 = n15156 ^ n14008;
  assign n15158 = n15157 ^ n15156;
  assign n15159 = ~n14113 & ~n14117;
  assign n15160 = n15148 & n15159;
  assign n15161 = n15160 ^ n15156;
  assign n15162 = n15158 & ~n15161;
  assign n15163 = n15162 ^ n15156;
  assign n15164 = ~n14007 & ~n15163;
  assign n15165 = n15153 & ~n15164;
  assign n15166 = n14112 & n15165;
  assign n15167 = n15166 ^ n12496;
  assign n15168 = n15167 ^ x91;
  assign n15169 = n15011 ^ x109;
  assign n15170 = n15168 & n15169;
  assign n15171 = ~n12647 & n12700;
  assign n15172 = n12656 & ~n15171;
  assign n15173 = n12652 & n12665;
  assign n15174 = ~n12655 & n12704;
  assign n15175 = n11847 & ~n15174;
  assign n15176 = ~n15173 & ~n15175;
  assign n15177 = n12687 ^ n11382;
  assign n15178 = n15177 ^ n12687;
  assign n15179 = n12687 ^ n12677;
  assign n15180 = n15179 ^ n12687;
  assign n15181 = n15178 & n15180;
  assign n15182 = n15181 ^ n12687;
  assign n15183 = ~n11846 & n15182;
  assign n15184 = n15183 ^ n12687;
  assign n15185 = n15176 & ~n15184;
  assign n15186 = ~n15172 & n15185;
  assign n15187 = n12703 & n14229;
  assign n15188 = n15187 ^ n11846;
  assign n15189 = n15188 ^ n15187;
  assign n15190 = n12688 & n12699;
  assign n15191 = ~n12681 & n15190;
  assign n15192 = n15191 ^ n15187;
  assign n15193 = ~n15189 & n15192;
  assign n15194 = n15193 ^ n15187;
  assign n15195 = ~n11382 & ~n15194;
  assign n15196 = n15186 & ~n15195;
  assign n15197 = n12661 & n15196;
  assign n15198 = n14767 & n15197;
  assign n15199 = ~n14212 & n15198;
  assign n15200 = n15199 ^ n12862;
  assign n15201 = n15200 ^ x77;
  assign n15202 = n13737 & ~n14179;
  assign n15203 = n13705 & ~n13743;
  assign n15204 = ~n13718 & n14696;
  assign n15205 = ~n13730 & n15204;
  assign n15206 = n13734 & ~n15205;
  assign n15207 = ~n15203 & ~n15206;
  assign n15208 = n13737 & ~n13746;
  assign n15212 = ~n13700 & n13709;
  assign n15213 = ~n13756 & ~n15212;
  assign n15209 = ~n13714 & ~n13735;
  assign n15210 = ~n13738 & n15209;
  assign n15211 = ~n13729 & n15210;
  assign n15214 = n15213 ^ n15211;
  assign n15215 = n15213 ^ n13630;
  assign n15216 = n15213 & n15215;
  assign n15217 = n15216 ^ n15213;
  assign n15218 = n15214 & n15217;
  assign n15219 = n15218 ^ n15216;
  assign n15220 = n15219 ^ n15213;
  assign n15221 = n15220 ^ n13630;
  assign n15222 = ~n15208 & n15221;
  assign n15223 = n15222 ^ n15208;
  assign n15224 = n15207 & ~n15223;
  assign n15225 = n14174 & n15224;
  assign n15226 = ~n15202 & n15225;
  assign n15227 = n13740 ^ n13734;
  assign n15228 = n13740 ^ n13705;
  assign n15229 = n15228 ^ n13705;
  assign n15230 = n13705 ^ n13703;
  assign n15231 = n15229 & ~n15230;
  assign n15232 = n15231 ^ n13705;
  assign n15233 = ~n15227 & n15232;
  assign n15234 = n15233 ^ n13734;
  assign n15235 = n15226 & ~n15234;
  assign n15236 = ~n13712 & n15235;
  assign n15237 = n14177 & n15236;
  assign n15238 = ~n13704 & n15237;
  assign n15239 = n15238 ^ n12889;
  assign n15240 = n15239 ^ x126;
  assign n15241 = n15201 & n15240;
  assign n15242 = n13905 & n14867;
  assign n15243 = n13814 & n13943;
  assign n15244 = ~n15242 & ~n15243;
  assign n15245 = n13889 & n13923;
  assign n15246 = n14290 & n14869;
  assign n15247 = n13894 & ~n15246;
  assign n15248 = n13927 & n14305;
  assign n15249 = n14280 & n15248;
  assign n15250 = n13911 & ~n15249;
  assign n15251 = ~n15247 & ~n15250;
  assign n15252 = ~n15245 & n15251;
  assign n15253 = n15244 & n15252;
  assign n15254 = ~n13902 & n15253;
  assign n15255 = ~n13910 & n15254;
  assign n15256 = ~n14865 & n15255;
  assign n15257 = ~n14282 & n15256;
  assign n15258 = ~n14293 & n15257;
  assign n15259 = n15258 ^ n12578;
  assign n15260 = n15259 ^ x84;
  assign n15261 = n15084 ^ x78;
  assign n15262 = ~n15260 & n15261;
  assign n15263 = n15241 & n15262;
  assign n15264 = n15170 & n15263;
  assign n15265 = ~n15168 & ~n15169;
  assign n15266 = n15201 & ~n15240;
  assign n15267 = n15260 & n15261;
  assign n15268 = n15266 & n15267;
  assign n15269 = n15265 & n15268;
  assign n15270 = n15168 & ~n15169;
  assign n15271 = ~n15201 & n15240;
  assign n15272 = n15262 & n15271;
  assign n15273 = n15241 & n15267;
  assign n15274 = ~n15272 & ~n15273;
  assign n15275 = n15270 & ~n15274;
  assign n15276 = n15262 & n15266;
  assign n15277 = n15170 & n15276;
  assign n15278 = n15267 & n15271;
  assign n15279 = n15170 & n15278;
  assign n15280 = ~n15277 & ~n15279;
  assign n15281 = ~n15168 & n15169;
  assign n15282 = n15260 & ~n15261;
  assign n15283 = n15271 & n15282;
  assign n15284 = n15281 & n15283;
  assign n15285 = n15266 & n15282;
  assign n15286 = ~n15201 & ~n15240;
  assign n15287 = ~n15260 & ~n15261;
  assign n15288 = n15286 & n15287;
  assign n15289 = ~n15285 & ~n15288;
  assign n15290 = ~n15276 & n15289;
  assign n15291 = n15270 & ~n15290;
  assign n15292 = ~n15284 & ~n15291;
  assign n15293 = n15169 & n15288;
  assign n15294 = n15282 & n15286;
  assign n15295 = n15266 & n15287;
  assign n15296 = ~n15294 & ~n15295;
  assign n15297 = n15265 & ~n15296;
  assign n15298 = ~n15293 & ~n15297;
  assign n15299 = n15267 & n15286;
  assign n15300 = ~n15268 & ~n15299;
  assign n15301 = n15281 & ~n15300;
  assign n15302 = n15241 & n15282;
  assign n15303 = ~n15169 & n15302;
  assign n15304 = ~n15268 & n15296;
  assign n15305 = n15170 & ~n15304;
  assign n15306 = ~n15303 & ~n15305;
  assign n15307 = ~n15170 & ~n15265;
  assign n15308 = n15283 & ~n15307;
  assign n15309 = n15241 & n15287;
  assign n15310 = ~n15299 & ~n15309;
  assign n15311 = n15270 & ~n15310;
  assign n15312 = ~n15308 & ~n15311;
  assign n15313 = n15274 & ~n15276;
  assign n15314 = n15265 & ~n15313;
  assign n15315 = n15262 & n15286;
  assign n15316 = n15271 & n15287;
  assign n15317 = ~n15302 & ~n15316;
  assign n15318 = ~n15315 & n15317;
  assign n15319 = ~n15263 & n15318;
  assign n15320 = n15281 & ~n15319;
  assign n15321 = ~n15314 & ~n15320;
  assign n15322 = n15312 & n15321;
  assign n15323 = n15306 & n15322;
  assign n15324 = ~n15301 & n15323;
  assign n15325 = n15298 & n15324;
  assign n15326 = n15292 & n15325;
  assign n15327 = n15280 & n15326;
  assign n15328 = ~n15275 & n15327;
  assign n15329 = ~n15269 & n15328;
  assign n15330 = ~n15264 & n15329;
  assign n15331 = n15330 ^ n13237;
  assign n15332 = n15331 ^ x99;
  assign n15333 = ~n15143 & ~n15332;
  assign n15334 = ~n14979 & n15333;
  assign n15335 = ~n14687 & ~n14972;
  assign n15336 = n14399 & n15335;
  assign n15337 = n15333 & n15336;
  assign n15338 = n14687 & ~n14972;
  assign n15339 = n14399 & n15338;
  assign n15340 = n15143 & n15332;
  assign n15341 = n15339 & n15340;
  assign n15342 = ~n14006 & n14398;
  assign n15343 = n14973 & n15342;
  assign n15344 = ~n15143 & n15332;
  assign n15345 = n15343 & n15344;
  assign n15346 = ~n15341 & ~n15345;
  assign n15347 = ~n15337 & n15346;
  assign n15348 = ~n15334 & n15347;
  assign n15349 = n15336 & n15340;
  assign n15350 = n14975 & n14977;
  assign n15351 = ~n14006 & ~n14398;
  assign n15352 = n14973 & n15351;
  assign n15353 = ~n15350 & ~n15352;
  assign n15354 = n15340 & ~n15353;
  assign n15355 = ~n15349 & ~n15354;
  assign n15356 = n15344 & n15350;
  assign n15357 = n15335 & n15342;
  assign n15358 = n15143 & ~n15332;
  assign n15359 = n15357 & n15358;
  assign n15360 = ~n15356 & ~n15359;
  assign n15361 = n15340 & n15343;
  assign n15362 = n15333 & n15339;
  assign n15363 = ~n15361 & ~n15362;
  assign n15364 = n15332 ^ n15143;
  assign n15365 = n14977 & n15351;
  assign n15366 = n15338 & n15342;
  assign n15367 = ~n15365 & ~n15366;
  assign n15368 = ~n15364 & ~n15367;
  assign n15369 = n14975 & n15335;
  assign n15370 = n14977 & n15342;
  assign n15371 = n15338 & n15351;
  assign n15372 = ~n15366 & ~n15371;
  assign n15373 = ~n15370 & n15372;
  assign n15374 = ~n15369 & n15373;
  assign n15375 = n15344 & ~n15374;
  assign n15376 = n15335 & n15351;
  assign n15377 = n14975 & n15338;
  assign n15378 = n14979 & ~n15377;
  assign n15379 = ~n15370 & n15378;
  assign n15380 = ~n15376 & n15379;
  assign n15381 = ~n15352 & n15380;
  assign n15382 = n15358 & ~n15381;
  assign n15383 = ~n15375 & ~n15382;
  assign n15384 = ~n15368 & n15383;
  assign n15385 = n15363 & n15384;
  assign n15386 = n15376 ^ n15332;
  assign n15387 = n15386 ^ n15376;
  assign n15388 = n15376 ^ n15357;
  assign n15389 = ~n15387 & n15388;
  assign n15390 = n15389 ^ n15376;
  assign n15391 = ~n15143 & n15390;
  assign n15392 = n15385 & ~n15391;
  assign n15393 = n15360 & n15392;
  assign n15394 = n15355 & n15393;
  assign n15395 = n15348 & n15394;
  assign n15396 = ~n14974 & n15395;
  assign n15397 = n15396 ^ n14719;
  assign n15398 = n15397 ^ x65;
  assign n15399 = n13967 ^ n13962;
  assign n15400 = n13967 ^ n13624;
  assign n15401 = n15400 ^ n13967;
  assign n15402 = n15399 & n15401;
  assign n15403 = n15402 ^ n13967;
  assign n15404 = ~n13977 & ~n15403;
  assign n15405 = ~n13627 & n15404;
  assign n15406 = n13997 & ~n15405;
  assign n15407 = n13206 & n13959;
  assign n15408 = n13625 & n13962;
  assign n15409 = ~n13998 & ~n15408;
  assign n15410 = n13981 & n15409;
  assign n15411 = ~n15407 & n15410;
  assign n15412 = n13972 & n15411;
  assign n15413 = n13958 & ~n15412;
  assign n15414 = ~n15406 & ~n15413;
  assign n15415 = ~n13625 & ~n13961;
  assign n15416 = n13207 & ~n15415;
  assign n15417 = ~n15407 & ~n15416;
  assign n15418 = n13624 & n13962;
  assign n15419 = n13961 & n13967;
  assign n15420 = ~n15418 & ~n15419;
  assign n15421 = n15409 & n15420;
  assign n15422 = n15417 & n15421;
  assign n15423 = n15422 ^ n13957;
  assign n15424 = n15423 ^ n15422;
  assign n15425 = n13419 & n13967;
  assign n15426 = n15417 & ~n15425;
  assign n15427 = n13964 & n15426;
  assign n15428 = n15427 ^ n15422;
  assign n15429 = ~n15424 & ~n15428;
  assign n15430 = n15429 ^ n15422;
  assign n15431 = ~n13780 & n15430;
  assign n15432 = n15414 & ~n15431;
  assign n15433 = n15432 ^ n13012;
  assign n15434 = n15433 ^ x91;
  assign n15435 = n14609 & n14656;
  assign n15436 = ~n14614 & ~n14632;
  assign n15437 = ~n14625 & n15436;
  assign n15438 = n14402 & ~n15437;
  assign n15439 = ~n15435 & ~n15438;
  assign n15440 = n14613 & n14619;
  assign n15441 = n14627 & ~n14668;
  assign n15442 = ~n15440 & ~n15441;
  assign n15443 = n14606 & n14619;
  assign n15444 = ~n14657 & ~n14672;
  assign n15445 = n14402 & ~n15444;
  assign n15446 = ~n15443 & ~n15445;
  assign n15447 = n14609 & n14651;
  assign n15448 = n14618 & n14641;
  assign n15449 = ~n14639 & ~n15448;
  assign n15450 = n14661 & n14673;
  assign n15451 = n15449 & n15450;
  assign n15452 = n14622 & ~n15451;
  assign n15453 = n14653 & ~n14672;
  assign n15454 = ~n14609 & n15453;
  assign n15455 = n14654 & ~n14672;
  assign n15456 = ~n14639 & n15455;
  assign n15457 = n14404 & ~n14628;
  assign n15458 = n14609 & ~n15457;
  assign n15459 = ~n14627 & ~n15458;
  assign n15460 = ~n15456 & ~n15459;
  assign n15461 = ~n15454 & n15460;
  assign n15462 = ~n15452 & ~n15461;
  assign n15463 = ~n15447 & n15462;
  assign n15464 = n15446 & n15463;
  assign n15465 = n15442 & n15464;
  assign n15466 = n15439 & n15465;
  assign n15467 = n14638 & n15466;
  assign n15468 = n14617 & n15467;
  assign n15469 = n15468 ^ n13883;
  assign n15470 = n15469 ^ x77;
  assign n15471 = ~n15434 & ~n15470;
  assign n15472 = n14827 ^ x115;
  assign n15473 = n15259 ^ x72;
  assign n15474 = n15472 & ~n15473;
  assign n15475 = ~n13349 & n14425;
  assign n15476 = n13343 & ~n15475;
  assign n15477 = ~n13367 & n14998;
  assign n15478 = ~n13376 & n15477;
  assign n15479 = ~n13388 & n15478;
  assign n15480 = n13346 & ~n15479;
  assign n15481 = ~n15476 & ~n15480;
  assign n15482 = n13371 & n13397;
  assign n15483 = ~n13373 & ~n13398;
  assign n15484 = ~n14406 & ~n15483;
  assign n15485 = n13341 & n13355;
  assign n15486 = n13343 & ~n14998;
  assign n15487 = ~n15485 & ~n15486;
  assign n15488 = n13396 & ~n13404;
  assign n15489 = n13371 & ~n15488;
  assign n15490 = n13378 & n13403;
  assign n15491 = ~n13393 & n15490;
  assign n15492 = n13384 & ~n15491;
  assign n15493 = ~n15489 & ~n15492;
  assign n15494 = n15487 & n15493;
  assign n15495 = ~n15484 & n15494;
  assign n15496 = ~n15482 & n15495;
  assign n15497 = n15481 & n15496;
  assign n15498 = n14418 & n15497;
  assign n15499 = ~n13345 & n15498;
  assign n15500 = n15499 ^ n12556;
  assign n15501 = n15500 ^ x96;
  assign n15502 = ~n13133 & ~n13177;
  assign n15503 = ~n13152 & n15502;
  assign n15504 = n13125 & ~n15503;
  assign n15505 = n12967 & ~n14155;
  assign n15506 = ~n15504 & ~n15505;
  assign n15507 = n13150 & ~n13165;
  assign n15508 = n13171 & n13183;
  assign n15509 = n13154 & n15508;
  assign n15510 = n13149 & ~n15509;
  assign n15511 = ~n12838 & n13157;
  assign n15512 = ~n13123 & ~n13132;
  assign n15513 = n13136 & ~n15512;
  assign n15514 = ~n13178 & n13183;
  assign n15515 = ~n13132 & n15514;
  assign n15516 = n12967 & ~n15515;
  assign n15517 = ~n15513 & ~n15516;
  assign n15518 = ~n15511 & n15517;
  assign n15519 = ~n15510 & n15518;
  assign n15520 = ~n15507 & n15519;
  assign n15521 = n15506 & n15520;
  assign n15522 = ~n13163 & n15521;
  assign n15523 = ~n14857 & n15522;
  assign n15524 = ~n13158 & n15523;
  assign n15525 = n14142 & n15524;
  assign n15526 = n15525 ^ n12532;
  assign n15527 = n15526 ^ x122;
  assign n15528 = n15501 & ~n15527;
  assign n15529 = n15167 ^ x113;
  assign n15530 = n14763 ^ x82;
  assign n15531 = n15529 & ~n15530;
  assign n15532 = n15528 & n15531;
  assign n15533 = n15474 & n15532;
  assign n15534 = ~n15472 & n15473;
  assign n15535 = ~n15501 & n15527;
  assign n15536 = ~n15529 & n15530;
  assign n15537 = n15535 & n15536;
  assign n15538 = n15534 & n15537;
  assign n15539 = n15472 & n15473;
  assign n15540 = n15528 & n15536;
  assign n15541 = ~n15529 & ~n15530;
  assign n15542 = n15535 & n15541;
  assign n15543 = ~n15540 & ~n15542;
  assign n15544 = n15539 & ~n15543;
  assign n15545 = ~n15538 & ~n15544;
  assign n15546 = ~n15533 & n15545;
  assign n15547 = n15473 ^ n15472;
  assign n15548 = ~n15501 & ~n15527;
  assign n15549 = n15536 & n15548;
  assign n15550 = ~n15547 & n15549;
  assign n15551 = n15528 & n15541;
  assign n15552 = n15539 & n15551;
  assign n15553 = ~n15550 & ~n15552;
  assign n15554 = n15531 & n15535;
  assign n15555 = n15529 & n15530;
  assign n15556 = n15528 & n15555;
  assign n15557 = n15501 & n15527;
  assign n15558 = n15555 & n15557;
  assign n15559 = ~n15556 & ~n15558;
  assign n15560 = ~n15554 & n15559;
  assign n15561 = n15474 & ~n15560;
  assign n15562 = ~n15472 & ~n15473;
  assign n15563 = n15536 & n15557;
  assign n15564 = ~n15542 & ~n15563;
  assign n15565 = ~n15537 & n15564;
  assign n15566 = n15562 & ~n15565;
  assign n15567 = ~n15561 & ~n15566;
  assign n15568 = n15541 & n15548;
  assign n15569 = ~n15549 & ~n15551;
  assign n15570 = ~n15568 & n15569;
  assign n15571 = n15534 & ~n15570;
  assign n15572 = n15534 & n15554;
  assign n15573 = n15534 & n15558;
  assign n15574 = n15474 & n15563;
  assign n15575 = n15541 & n15557;
  assign n15576 = n15539 & n15575;
  assign n15577 = ~n15574 & ~n15576;
  assign n15578 = ~n15573 & n15577;
  assign n15579 = n15531 & n15548;
  assign n15580 = n15539 & n15579;
  assign n15581 = n15474 & n15568;
  assign n15582 = ~n15580 & ~n15581;
  assign n15583 = n15548 & n15555;
  assign n15584 = n15531 & n15557;
  assign n15585 = ~n15583 & ~n15584;
  assign n15586 = n15534 & ~n15585;
  assign n15587 = ~n15537 & ~n15575;
  assign n15588 = n15474 & ~n15587;
  assign n15589 = ~n15586 & ~n15588;
  assign n15590 = n15539 & ~n15559;
  assign n15591 = n15535 & n15555;
  assign n15592 = ~n15584 & ~n15591;
  assign n15593 = ~n15532 & ~n15556;
  assign n15594 = n15592 & n15593;
  assign n15595 = n15562 & ~n15594;
  assign n15596 = ~n15590 & ~n15595;
  assign n15597 = n15589 & n15596;
  assign n15598 = n15582 & n15597;
  assign n15599 = n15578 & n15598;
  assign n15600 = ~n15572 & n15599;
  assign n15601 = ~n15571 & n15600;
  assign n15602 = n15567 & n15601;
  assign n15603 = n15553 & n15602;
  assign n15604 = n15546 & n15603;
  assign n15605 = n15604 ^ n14522;
  assign n15606 = n15605 ^ x101;
  assign n15607 = n15085 ^ n15047;
  assign n15608 = n14990 & n15044;
  assign n15609 = n15089 & n15104;
  assign n15610 = ~n15107 & ~n15609;
  assign n15611 = ~n15608 & n15610;
  assign n15612 = n15611 ^ n15085;
  assign n15613 = n15612 ^ n15611;
  assign n15614 = ~n15128 & ~n15609;
  assign n15615 = ~n15103 & n15614;
  assign n15616 = n15615 ^ n15611;
  assign n15617 = ~n15613 & n15616;
  assign n15618 = n15617 ^ n15611;
  assign n15619 = n15607 & ~n15618;
  assign n15620 = ~n15097 & ~n15105;
  assign n15621 = n15610 & n15620;
  assign n15622 = ~n15047 & ~n15085;
  assign n15623 = ~n15621 & n15622;
  assign n15624 = n14990 & n15098;
  assign n15625 = ~n15090 & ~n15624;
  assign n15626 = ~n15092 & n15625;
  assign n15627 = ~n15129 & n15626;
  assign n15628 = n15118 & n15627;
  assign n15629 = n15088 & ~n15628;
  assign n15630 = ~n15623 & ~n15629;
  assign n15631 = ~n15086 & ~n15113;
  assign n15632 = n15624 ^ n14990;
  assign n15633 = ~n15086 & ~n15632;
  assign n15634 = ~n15092 & ~n15113;
  assign n15635 = ~n15633 & ~n15634;
  assign n15636 = ~n15114 & ~n15635;
  assign n15637 = ~n15631 & ~n15636;
  assign n15638 = n15630 & ~n15637;
  assign n15639 = ~n15087 & n15638;
  assign n15640 = ~n15608 & n15626;
  assign n15641 = n15640 ^ n15622;
  assign n15642 = n15641 ^ n15640;
  assign n15643 = n15640 ^ n15099;
  assign n15644 = ~n15642 & ~n15643;
  assign n15645 = n15644 ^ n15640;
  assign n15646 = n15639 & n15645;
  assign n15647 = ~n15619 & n15646;
  assign n15648 = n15647 ^ n14484;
  assign n15649 = n15648 ^ x116;
  assign n15650 = n15606 & ~n15649;
  assign n15651 = n13418 ^ x120;
  assign n15652 = n14862 ^ x65;
  assign n15653 = n15651 & n15652;
  assign n15654 = n14008 & ~n14112;
  assign n15655 = n15151 ^ n14008;
  assign n15656 = n15655 ^ n15151;
  assign n15657 = n14112 & n15148;
  assign n15658 = n15657 ^ n15151;
  assign n15659 = ~n15656 & ~n15658;
  assign n15660 = n15659 ^ n15151;
  assign n15661 = n14007 & ~n15660;
  assign n15662 = ~n15654 & ~n15661;
  assign n15663 = n14099 & ~n15156;
  assign n15664 = n14123 & ~n15160;
  assign n15665 = ~n15663 & ~n15664;
  assign n15666 = n15662 & n15665;
  assign n15667 = n15666 ^ n12734;
  assign n15668 = n15667 ^ x88;
  assign n15669 = n13956 ^ x106;
  assign n15670 = n15668 & n15669;
  assign n15671 = n14719 ^ x97;
  assign n15672 = n14527 & n14546;
  assign n15673 = ~n14572 & ~n14576;
  assign n15674 = n14547 & n15673;
  assign n15675 = n14441 & ~n15674;
  assign n15676 = ~n15672 & ~n15675;
  assign n15677 = ~n14530 & n14723;
  assign n15678 = n14564 & ~n15677;
  assign n15679 = ~n14527 & n14583;
  assign n15680 = n14562 & n14747;
  assign n15681 = ~n14536 & n15680;
  assign n15682 = ~n15679 & ~n15681;
  assign n15683 = ~n14537 & n15682;
  assign n15684 = ~n15678 & ~n15683;
  assign n15685 = n15676 & n15684;
  assign n15686 = n14588 ^ n14536;
  assign n15687 = n14588 ^ n14527;
  assign n15688 = n15687 ^ n14527;
  assign n15689 = n14527 ^ n14525;
  assign n15690 = ~n15688 & ~n15689;
  assign n15691 = n15690 ^ n14527;
  assign n15692 = n15686 & n15691;
  assign n15693 = n15692 ^ n14536;
  assign n15694 = n15685 & ~n15693;
  assign n15695 = n15052 & n15694;
  assign n15696 = n14582 & n15695;
  assign n15697 = ~n14534 & n15696;
  assign n15698 = n14725 & n15697;
  assign n15699 = n15698 ^ n12766;
  assign n15700 = n15699 ^ x123;
  assign n15701 = ~n15671 & n15700;
  assign n15702 = n15670 & n15701;
  assign n15703 = n15653 & n15702;
  assign n15704 = n15651 & ~n15652;
  assign n15705 = ~n15668 & n15669;
  assign n15706 = ~n15671 & ~n15700;
  assign n15707 = n15705 & n15706;
  assign n15708 = n15704 & n15707;
  assign n15709 = ~n15703 & ~n15708;
  assign n15710 = ~n15651 & ~n15652;
  assign n15711 = n15671 & ~n15700;
  assign n15712 = n15670 & n15711;
  assign n15713 = n15710 & n15712;
  assign n15714 = ~n15653 & ~n15710;
  assign n15715 = n15671 & n15700;
  assign n15716 = n15705 & n15715;
  assign n15717 = ~n15714 & n15716;
  assign n15718 = ~n15651 & n15652;
  assign n15719 = n15668 & ~n15669;
  assign n15720 = n15711 & n15719;
  assign n15721 = n15705 & n15711;
  assign n15722 = ~n15720 & ~n15721;
  assign n15723 = n15718 & ~n15722;
  assign n15724 = ~n15717 & ~n15723;
  assign n15725 = n15653 & n15712;
  assign n15726 = n15670 & n15715;
  assign n15727 = ~n15668 & ~n15669;
  assign n15728 = n15715 & n15727;
  assign n15729 = ~n15726 & ~n15728;
  assign n15730 = n15704 & ~n15729;
  assign n15731 = ~n15725 & ~n15730;
  assign n15732 = n15706 & n15719;
  assign n15733 = n15701 & n15727;
  assign n15734 = n15670 & n15706;
  assign n15735 = ~n15733 & ~n15734;
  assign n15736 = n15701 & n15719;
  assign n15737 = n15711 & n15727;
  assign n15738 = ~n15736 & ~n15737;
  assign n15739 = n15735 & n15738;
  assign n15740 = ~n15732 & n15739;
  assign n15741 = n15704 & ~n15740;
  assign n15742 = n15669 ^ n15668;
  assign n15743 = n15700 ^ n15669;
  assign n15744 = n15671 ^ n15669;
  assign n15745 = n15744 ^ n15669;
  assign n15746 = n15743 & n15745;
  assign n15747 = n15746 ^ n15669;
  assign n15748 = n15742 & n15747;
  assign n15749 = n15748 ^ n15700;
  assign n15750 = n15718 & n15749;
  assign n15751 = ~n15741 & ~n15750;
  assign n15752 = n15706 & n15727;
  assign n15753 = n15653 & n15752;
  assign n15754 = n15715 & n15719;
  assign n15755 = ~n15737 & ~n15754;
  assign n15756 = n15701 & n15705;
  assign n15757 = ~n15732 & ~n15756;
  assign n15758 = ~n15710 & n15757;
  assign n15759 = ~n15702 & ~n15707;
  assign n15760 = ~n15734 & n15759;
  assign n15761 = ~n15732 & n15760;
  assign n15762 = ~n15653 & n15761;
  assign n15763 = ~n15758 & ~n15762;
  assign n15764 = n15755 & ~n15763;
  assign n15765 = ~n15714 & n15764;
  assign n15766 = n15765 ^ n15714;
  assign n15767 = ~n15753 & n15766;
  assign n15768 = n15751 & n15767;
  assign n15769 = n15731 & n15768;
  assign n15770 = n15724 & n15769;
  assign n15771 = ~n15713 & n15770;
  assign n15772 = n15709 & n15771;
  assign n15773 = n15772 ^ n13812;
  assign n15774 = n15773 ^ x67;
  assign n15775 = ~n15273 & ~n15315;
  assign n15776 = n15281 & ~n15775;
  assign n15777 = n15272 & n15281;
  assign n15778 = ~n15283 & ~n15295;
  assign n15779 = n15270 & ~n15778;
  assign n15780 = ~n15777 & ~n15779;
  assign n15781 = n15263 & n15265;
  assign n15782 = n15169 & n15299;
  assign n15783 = ~n15781 & ~n15782;
  assign n15784 = n15278 & ~n15307;
  assign n15785 = n15270 & n15302;
  assign n15786 = ~n15784 & ~n15785;
  assign n15787 = ~n15169 & n15315;
  assign n15788 = ~n15268 & ~n15276;
  assign n15789 = n15270 & ~n15788;
  assign n15790 = ~n15287 & n15289;
  assign n15791 = n15170 & ~n15790;
  assign n15792 = ~n15789 & ~n15791;
  assign n15793 = ~n15285 & n15317;
  assign n15794 = ~n15309 & n15793;
  assign n15795 = n15281 & ~n15794;
  assign n15796 = ~n15294 & n15778;
  assign n15797 = ~n15316 & n15796;
  assign n15798 = n15265 & ~n15797;
  assign n15799 = ~n15795 & ~n15798;
  assign n15800 = n15792 & n15799;
  assign n15801 = ~n15275 & n15800;
  assign n15802 = ~n15787 & n15801;
  assign n15803 = n15786 & n15802;
  assign n15804 = n15783 & n15803;
  assign n15805 = n15780 & n15804;
  assign n15806 = ~n15776 & n15805;
  assign n15807 = ~n15269 & n15806;
  assign n15808 = ~n15264 & n15807;
  assign n15809 = n15808 ^ n12965;
  assign n15810 = n15809 ^ x78;
  assign n15811 = ~n15774 & n15810;
  assign n15812 = n15650 & n15811;
  assign n15813 = n15606 & n15649;
  assign n15814 = n15774 & n15810;
  assign n15815 = n15813 & n15814;
  assign n15816 = ~n15812 & ~n15815;
  assign n15817 = n15471 & ~n15816;
  assign n15818 = n15470 ^ n15434;
  assign n15819 = ~n15606 & n15649;
  assign n15820 = n15811 & n15819;
  assign n15821 = ~n15818 & n15820;
  assign n15822 = n15650 & n15814;
  assign n15823 = ~n15606 & ~n15649;
  assign n15824 = n15811 & n15823;
  assign n15825 = ~n15822 & ~n15824;
  assign n15826 = n15434 & ~n15825;
  assign n15827 = ~n15821 & ~n15826;
  assign n15828 = n15814 & n15819;
  assign n15829 = n15471 & n15828;
  assign n15830 = n15434 & ~n15470;
  assign n15831 = n15811 & n15813;
  assign n15832 = ~n15815 & ~n15831;
  assign n15833 = n15830 & ~n15832;
  assign n15834 = ~n15774 & ~n15810;
  assign n15835 = n15819 & n15834;
  assign n15836 = n15774 & ~n15810;
  assign n15837 = n15813 & n15836;
  assign n15838 = ~n15835 & ~n15837;
  assign n15839 = n15830 & ~n15838;
  assign n15840 = n15434 & n15470;
  assign n15841 = n15814 & n15823;
  assign n15842 = n15813 & n15834;
  assign n15843 = ~n15837 & ~n15842;
  assign n15844 = ~n15841 & n15843;
  assign n15845 = n15840 & ~n15844;
  assign n15846 = n15819 & n15836;
  assign n15847 = ~n15842 & ~n15846;
  assign n15848 = n15650 & n15836;
  assign n15849 = n15650 & n15834;
  assign n15850 = ~n15848 & ~n15849;
  assign n15851 = n15847 & n15850;
  assign n15852 = n15471 & ~n15851;
  assign n15853 = ~n15845 & ~n15852;
  assign n15864 = n15823 & n15836;
  assign n15865 = ~n15849 & ~n15864;
  assign n15854 = n15774 ^ n15649;
  assign n15855 = n15854 ^ n15649;
  assign n15856 = n15649 ^ n15606;
  assign n15857 = n15856 ^ n15774;
  assign n15858 = n15857 ^ n15649;
  assign n15859 = n15858 ^ n15649;
  assign n15860 = n15855 & n15859;
  assign n15861 = n15860 ^ n15649;
  assign n15862 = ~n15810 & n15861;
  assign n15863 = n15862 ^ n15857;
  assign n15866 = n15865 ^ n15863;
  assign n15867 = n15866 ^ n15865;
  assign n15868 = n15865 ^ n15470;
  assign n15869 = n15868 ^ n15865;
  assign n15870 = ~n15867 & n15869;
  assign n15871 = n15870 ^ n15865;
  assign n15872 = ~n15434 & ~n15871;
  assign n15873 = n15872 ^ n15865;
  assign n15874 = n15853 & n15873;
  assign n15875 = ~n15839 & n15874;
  assign n15876 = ~n15833 & n15875;
  assign n15877 = ~n15829 & n15876;
  assign n15878 = n15827 & n15877;
  assign n15879 = ~n15817 & n15878;
  assign n15880 = n15879 ^ n15699;
  assign n15881 = n15880 ^ x120;
  assign n15882 = ~n15398 & n15881;
  assign n15883 = ~n15607 & n15608;
  assign n15884 = ~n15090 & ~n15099;
  assign n15885 = n15086 & ~n15884;
  assign n15886 = n15088 & ~n15109;
  assign n15887 = ~n15885 & ~n15886;
  assign n15888 = n15113 & n15127;
  assign n15889 = n15106 & n15614;
  assign n15890 = ~n15047 & ~n15889;
  assign n15891 = n15093 & ~n15114;
  assign n15892 = n15622 & ~n15891;
  assign n15893 = ~n15890 & ~n15892;
  assign n15894 = ~n15888 & n15893;
  assign n15895 = n15887 & n15894;
  assign n15896 = ~n15095 & n15895;
  assign n15897 = ~n15883 & n15896;
  assign n15898 = ~n15087 & n15897;
  assign n15899 = n15898 ^ n12087;
  assign n15900 = n15899 ^ x105;
  assign n15901 = n15537 & ~n15547;
  assign n15902 = n15549 ^ n15473;
  assign n15903 = n15902 ^ n15549;
  assign n15904 = n15579 ^ n15549;
  assign n15905 = ~n15903 & n15904;
  assign n15906 = n15905 ^ n15549;
  assign n15907 = ~n15472 & n15906;
  assign n15908 = ~n15901 & ~n15907;
  assign n15909 = n15539 & n15554;
  assign n15910 = n15532 & n15534;
  assign n15911 = ~n15909 & ~n15910;
  assign n15912 = ~n15556 & ~n15583;
  assign n15913 = ~n15547 & ~n15912;
  assign n15914 = n15534 & ~n15559;
  assign n15915 = ~n15913 & ~n15914;
  assign n15916 = ~n15551 & ~n15584;
  assign n15917 = n15562 & ~n15916;
  assign n15918 = ~n15558 & ~n15579;
  assign n15919 = ~n15540 & ~n15568;
  assign n15920 = n15918 & n15919;
  assign n15921 = n15592 & n15920;
  assign n15922 = n15474 & ~n15921;
  assign n15923 = ~n15917 & ~n15922;
  assign n15924 = ~n15563 & ~n15575;
  assign n15925 = n15924 ^ n15473;
  assign n15926 = n15925 ^ n15924;
  assign n15927 = n15924 ^ n15532;
  assign n15928 = n15927 ^ n15924;
  assign n15929 = n15926 & n15928;
  assign n15930 = n15929 ^ n15924;
  assign n15931 = n15472 & ~n15930;
  assign n15932 = n15931 ^ n15924;
  assign n15933 = n15923 & n15932;
  assign n15934 = n15915 & n15933;
  assign n15935 = n15911 & n15934;
  assign n15936 = n15577 & n15935;
  assign n15937 = n15908 & n15936;
  assign n15938 = n15546 & n15937;
  assign n15939 = ~n15572 & n15938;
  assign n15940 = n15939 ^ n13120;
  assign n15941 = n15940 ^ x123;
  assign n15942 = n15900 & n15941;
  assign n15943 = n14402 & ~n14658;
  assign n15944 = n14637 & ~n15943;
  assign n15945 = n14402 & n14612;
  assign n15946 = n14627 & ~n14658;
  assign n15947 = ~n15945 & ~n15946;
  assign n15948 = n14401 ^ n14400;
  assign n15949 = ~n14632 & n15449;
  assign n15950 = n14673 & n15949;
  assign n15951 = n15950 ^ n14401;
  assign n15952 = n15951 ^ n15950;
  assign n15953 = ~n14625 & n15455;
  assign n15954 = n15953 ^ n15950;
  assign n15955 = n15952 & n15954;
  assign n15956 = n15955 ^ n15950;
  assign n15957 = ~n15948 & ~n15956;
  assign n15958 = n15947 & ~n15957;
  assign n15959 = n15442 & n15958;
  assign n15960 = n14628 ^ n14401;
  assign n15961 = n15960 ^ n14628;
  assign n15962 = n14613 & n14618;
  assign n15963 = n15962 ^ n14628;
  assign n15964 = n15961 & n15963;
  assign n15965 = n15964 ^ n14628;
  assign n15966 = n15948 & n15965;
  assign n15967 = n15959 & ~n15966;
  assign n15968 = n15944 & n15967;
  assign n15969 = n14631 & n15968;
  assign n15970 = n14617 & n15969;
  assign n15971 = n15970 ^ n14079;
  assign n15972 = n15971 ^ x82;
  assign n15973 = n14898 & n14900;
  assign n15974 = n14765 & ~n14935;
  assign n15975 = n14765 & ~n14963;
  assign n15976 = ~n14911 & ~n14928;
  assign n15977 = n14905 & ~n15976;
  assign n15978 = ~n15975 & ~n15977;
  assign n15979 = n14905 & n14940;
  assign n15980 = n14918 & ~n15979;
  assign n15981 = ~n14898 & ~n14928;
  assign n15982 = n14910 & ~n15981;
  assign n15983 = ~n14914 & ~n14922;
  assign n15984 = ~n14962 & n15983;
  assign n15985 = n14905 & ~n15984;
  assign n15986 = ~n15982 & ~n15985;
  assign n15987 = n14765 & n14948;
  assign n15988 = n14829 & n14913;
  assign n15989 = ~n14908 & ~n15988;
  assign n15990 = ~n14925 & ~n15989;
  assign n15991 = ~n14941 & n14949;
  assign n15992 = ~n14929 & n15991;
  assign n15993 = n14910 & ~n15992;
  assign n15994 = n14942 & ~n14962;
  assign n15995 = n14900 & ~n15994;
  assign n15996 = ~n15993 & ~n15995;
  assign n15997 = ~n15990 & n15996;
  assign n15998 = ~n15987 & n15997;
  assign n15999 = n15986 & n15998;
  assign n16000 = n15980 & n15999;
  assign n16001 = n15978 & n16000;
  assign n16002 = n14924 & n16001;
  assign n16003 = ~n15974 & n16002;
  assign n16004 = ~n15973 & n16003;
  assign n16005 = n16004 ^ n11845;
  assign n16006 = n16005 ^ x112;
  assign n16007 = n15972 & n16006;
  assign n16008 = n15718 & n15752;
  assign n16009 = n15718 & n15726;
  assign n16010 = n15704 & n15752;
  assign n16011 = ~n16009 & ~n16010;
  assign n16012 = ~n15712 & ~n15726;
  assign n16013 = n15653 & ~n16012;
  assign n16014 = ~n15734 & ~n15736;
  assign n16015 = n15704 & ~n16014;
  assign n16016 = ~n15732 & ~n15733;
  assign n16017 = ~n15737 & n16016;
  assign n16018 = n15653 & ~n16017;
  assign n16019 = ~n16015 & ~n16018;
  assign n16020 = ~n15720 & ~n15754;
  assign n16021 = ~n15707 & n16020;
  assign n16022 = n15735 & n16021;
  assign n16023 = n15718 & ~n16022;
  assign n16024 = ~n15721 & ~n15728;
  assign n16025 = ~n15714 & ~n16024;
  assign n16026 = ~n15651 & n15716;
  assign n16027 = ~n15728 & n16020;
  assign n16028 = ~n15716 & n16027;
  assign n16029 = n15704 & ~n16028;
  assign n16030 = ~n15736 & n15757;
  assign n16031 = ~n15702 & n16030;
  assign n16032 = n15710 & ~n16031;
  assign n16033 = ~n16029 & ~n16032;
  assign n16034 = ~n16026 & n16033;
  assign n16035 = ~n16025 & n16034;
  assign n16036 = ~n16023 & n16035;
  assign n16037 = n16019 & n16036;
  assign n16038 = ~n16013 & n16037;
  assign n16039 = n16011 & n16038;
  assign n16040 = ~n15713 & n16039;
  assign n16041 = ~n16008 & n16040;
  assign n16042 = n15709 & n16041;
  assign n16043 = n16042 ^ n12837;
  assign n16044 = n16043 ^ x64;
  assign n16045 = n15270 & n15278;
  assign n16046 = n15281 & n15302;
  assign n16047 = ~n16045 & ~n16046;
  assign n16048 = ~n15169 & n15309;
  assign n16049 = n15270 & ~n15304;
  assign n16050 = ~n16048 & ~n16049;
  assign n16051 = ~n15283 & ~n15316;
  assign n16052 = n15170 & ~n16051;
  assign n16053 = ~n15273 & ~n15276;
  assign n16054 = ~n15265 & n16053;
  assign n16055 = n15274 & ~n15277;
  assign n16056 = ~n15278 & n16055;
  assign n16057 = ~n16054 & ~n16056;
  assign n16058 = ~n15315 & ~n16057;
  assign n16059 = ~n15307 & ~n16058;
  assign n16060 = ~n16052 & ~n16059;
  assign n16061 = ~n15294 & ~n15309;
  assign n16062 = ~n15272 & n16061;
  assign n16063 = ~n15276 & n16062;
  assign n16064 = n16063 ^ n15285;
  assign n16065 = n15169 & ~n16064;
  assign n16066 = ~n15168 & n16065;
  assign n16067 = n16066 ^ n15285;
  assign n16068 = n16060 & ~n16067;
  assign n16069 = n16050 & n16068;
  assign n16070 = n16047 & n16069;
  assign n16071 = ~n15301 & n16070;
  assign n16072 = n15298 & n16071;
  assign n16073 = ~n15275 & n16072;
  assign n16074 = ~n15264 & n16073;
  assign n16075 = n16074 ^ n14056;
  assign n16076 = n16075 ^ x73;
  assign n16077 = ~n16044 & n16076;
  assign n16078 = n16007 & n16077;
  assign n16079 = n15942 & n16078;
  assign n16080 = ~n15900 & n15941;
  assign n16081 = ~n15972 & n16006;
  assign n16082 = n16077 & n16081;
  assign n16083 = n16044 & ~n16076;
  assign n16084 = n16007 & n16083;
  assign n16085 = ~n16082 & ~n16084;
  assign n16086 = n16080 & ~n16085;
  assign n16087 = ~n16079 & ~n16086;
  assign n16088 = n15900 & ~n15941;
  assign n16089 = n15972 & ~n16006;
  assign n16090 = ~n16044 & ~n16076;
  assign n16091 = n16089 & n16090;
  assign n16092 = ~n16078 & ~n16091;
  assign n16093 = n16007 & n16090;
  assign n16094 = ~n15972 & ~n16006;
  assign n16095 = n16077 & n16094;
  assign n16096 = n16044 & n16076;
  assign n16097 = n16007 & n16096;
  assign n16098 = ~n16095 & ~n16097;
  assign n16099 = ~n16093 & n16098;
  assign n16100 = ~n16006 & n16096;
  assign n16101 = n16081 & n16083;
  assign n16102 = ~n16100 & ~n16101;
  assign n16103 = n16099 & n16102;
  assign n16104 = n16092 & n16103;
  assign n16105 = n16088 & n16104;
  assign n16106 = ~n15900 & ~n15941;
  assign n16107 = n16044 & n16089;
  assign n16108 = n16090 & n16094;
  assign n16109 = ~n16107 & ~n16108;
  assign n16110 = n16103 & n16109;
  assign n16111 = n16106 & ~n16110;
  assign n16112 = ~n16105 & ~n16111;
  assign n16113 = ~n16095 & ~n16107;
  assign n16114 = ~n16101 & n16113;
  assign n16115 = n16092 & n16114;
  assign n16116 = n16080 & ~n16115;
  assign n16117 = n16006 & n16096;
  assign n16118 = ~n16077 & n16094;
  assign n16119 = ~n16117 & ~n16118;
  assign n16120 = ~n16084 & n16119;
  assign n16121 = ~n16091 & n16120;
  assign n16122 = n15942 & ~n16121;
  assign n16123 = ~n16116 & ~n16122;
  assign n16124 = n16112 & n16123;
  assign n16125 = n16087 & n16124;
  assign n16126 = n16125 ^ n15667;
  assign n16127 = n16126 ^ x121;
  assign n16128 = n15773 ^ x109;
  assign n16129 = n14171 & n14367;
  assign n16130 = n14332 & n14357;
  assign n16131 = ~n16129 & ~n16130;
  assign n16132 = ~n14357 & ~n14365;
  assign n16133 = n14171 & ~n16132;
  assign n16134 = n14351 ^ n14171;
  assign n16135 = n14351 ^ n14332;
  assign n16136 = n16135 ^ n14332;
  assign n16137 = n14371 ^ n14332;
  assign n16138 = ~n16136 & ~n16137;
  assign n16139 = n16138 ^ n14332;
  assign n16140 = n16134 & n16139;
  assign n16141 = n16140 ^ n14171;
  assign n16142 = n14170 ^ n14139;
  assign n16143 = n14346 ^ n14170;
  assign n16144 = n16143 ^ n14346;
  assign n16145 = n14386 ^ n14346;
  assign n16146 = ~n16144 & ~n16145;
  assign n16147 = n16146 ^ n14346;
  assign n16148 = ~n16142 & n16147;
  assign n16149 = ~n16141 & ~n16148;
  assign n16150 = ~n14335 & n14360;
  assign n16151 = n14341 & ~n16150;
  assign n16152 = ~n14330 & ~n14375;
  assign n16153 = ~n14352 & n16152;
  assign n16154 = n14332 & ~n16153;
  assign n16155 = ~n14337 & n14378;
  assign n16156 = n14341 & ~n16155;
  assign n16157 = n14338 & n14360;
  assign n16158 = ~n14346 & n16157;
  assign n16159 = n14342 & ~n16158;
  assign n16160 = ~n16156 & ~n16159;
  assign n16161 = ~n16154 & n16160;
  assign n16162 = ~n14352 & ~n14385;
  assign n16163 = n16162 ^ n14344;
  assign n16164 = n16163 ^ n14344;
  assign n16165 = n14344 ^ n14139;
  assign n16166 = n16165 ^ n14344;
  assign n16167 = ~n16164 & ~n16166;
  assign n16168 = n16167 ^ n14344;
  assign n16169 = n14170 & n16168;
  assign n16170 = n16169 ^ n14344;
  assign n16171 = n16161 & ~n16170;
  assign n16172 = ~n16151 & n16171;
  assign n16173 = n16149 & n16172;
  assign n16174 = ~n16133 & n16173;
  assign n16175 = n14340 & n16174;
  assign n16176 = n16131 & n16175;
  assign n16177 = n16176 ^ n13437;
  assign n16178 = n16177 ^ x100;
  assign n16179 = ~n16128 & ~n16178;
  assign n16180 = n13986 & ~n15405;
  assign n16181 = n13976 & ~n15412;
  assign n16182 = ~n16180 & ~n16181;
  assign n16183 = n13780 & ~n15430;
  assign n16184 = n16182 & ~n16183;
  assign n16185 = n16184 ^ n13822;
  assign n16186 = n16185 ^ x86;
  assign n16187 = ~n15307 & ~n16061;
  assign n16188 = ~n15263 & ~n15273;
  assign n16189 = n15270 & ~n16188;
  assign n16190 = n15274 & n15289;
  assign n16191 = n15170 & ~n16190;
  assign n16192 = ~n16189 & ~n16191;
  assign n16193 = ~n16187 & n16192;
  assign n16194 = n15281 & ~n15304;
  assign n16195 = ~n15299 & n15318;
  assign n16196 = ~n15272 & n16195;
  assign n16197 = n15265 & ~n16196;
  assign n16198 = ~n16194 & ~n16197;
  assign n16199 = n16193 & n16198;
  assign n16200 = n15780 & n16199;
  assign n16201 = n16047 & n16200;
  assign n16202 = ~n15776 & n16201;
  assign n16203 = n15292 & n16202;
  assign n16204 = n15280 & n16203;
  assign n16205 = ~n15269 & n16204;
  assign n16206 = n16205 ^ n13854;
  assign n16207 = n16206 ^ x76;
  assign n16208 = n16186 & n16207;
  assign n16209 = n15469 ^ x69;
  assign n16210 = n14900 & n14940;
  assign n16211 = ~n14908 & n14949;
  assign n16212 = n14915 & n16211;
  assign n16213 = n14963 & n16212;
  assign n16214 = ~n14902 & n16213;
  assign n16215 = n14905 & ~n16214;
  assign n16216 = ~n16210 & ~n16215;
  assign n16217 = n14942 & ~n14948;
  assign n16218 = ~n14908 & n16217;
  assign n16219 = n14910 & ~n16218;
  assign n16220 = n14765 & ~n15976;
  assign n16221 = ~n14920 & ~n14929;
  assign n16222 = ~n14925 & ~n16221;
  assign n16223 = ~n14926 & ~n14928;
  assign n16224 = ~n14910 & n16223;
  assign n16225 = ~n14898 & n15983;
  assign n16226 = ~n14900 & n16225;
  assign n16227 = ~n16224 & ~n16226;
  assign n16228 = ~n15988 & ~n16227;
  assign n16229 = n14764 & ~n16228;
  assign n16230 = ~n16222 & ~n16229;
  assign n16231 = ~n16220 & n16230;
  assign n16232 = ~n14923 & n16231;
  assign n16233 = ~n15974 & n16232;
  assign n16234 = ~n16219 & n16233;
  assign n16235 = n16216 & n16234;
  assign n16236 = ~n15975 & n16235;
  assign n16237 = ~n15973 & n16236;
  assign n16238 = n16237 ^ n13559;
  assign n16239 = n16238 ^ x126;
  assign n16240 = n16209 & n16239;
  assign n16241 = n16208 & n16240;
  assign n16242 = n16179 & n16241;
  assign n16243 = ~n16128 & n16178;
  assign n16247 = ~n16209 & ~n16239;
  assign n16248 = n16208 & n16247;
  assign n16244 = ~n16186 & ~n16207;
  assign n16245 = n16209 & ~n16239;
  assign n16246 = n16244 & n16245;
  assign n16249 = n16248 ^ n16246;
  assign n16250 = n16249 ^ n16248;
  assign n16251 = n16128 & ~n16178;
  assign n16252 = n16251 ^ n16248;
  assign n16253 = n16252 ^ n16248;
  assign n16254 = n16250 & ~n16253;
  assign n16255 = n16254 ^ n16248;
  assign n16256 = ~n16243 & n16255;
  assign n16257 = n16256 ^ n16248;
  assign n16258 = ~n16242 & ~n16257;
  assign n16259 = n16128 & n16178;
  assign n16260 = n16208 & n16245;
  assign n16261 = n16186 & ~n16207;
  assign n16262 = n16240 & n16261;
  assign n16263 = ~n16186 & n16207;
  assign n16264 = n16245 & n16263;
  assign n16265 = ~n16262 & ~n16264;
  assign n16266 = ~n16260 & n16265;
  assign n16267 = n16259 & ~n16266;
  assign n16268 = ~n16209 & n16239;
  assign n16269 = n16263 & n16268;
  assign n16270 = n16244 & n16268;
  assign n16271 = n16247 & n16261;
  assign n16272 = ~n16270 & ~n16271;
  assign n16273 = ~n16269 & n16272;
  assign n16274 = ~n16248 & n16273;
  assign n16275 = n16259 & ~n16274;
  assign n16276 = n16209 ^ n16186;
  assign n16277 = n16276 ^ n16239;
  assign n16278 = n16277 ^ n16209;
  assign n16279 = n16278 ^ n16207;
  assign n16280 = n16279 ^ n16239;
  assign n16281 = n16239 ^ n16209;
  assign n16282 = n16209 ^ n16207;
  assign n16283 = n16282 ^ n16209;
  assign n16284 = n16281 & n16283;
  assign n16285 = n16284 ^ n16209;
  assign n16286 = ~n16280 & n16285;
  assign n16287 = n16286 ^ n16277;
  assign n16288 = n16251 & ~n16287;
  assign n16289 = ~n16275 & ~n16288;
  assign n16290 = n16240 & n16244;
  assign n16291 = n16245 & n16261;
  assign n16292 = ~n16290 & ~n16291;
  assign n16293 = n16208 & n16268;
  assign n16294 = n16261 & n16268;
  assign n16295 = n16247 & n16263;
  assign n16296 = ~n16294 & ~n16295;
  assign n16297 = ~n16293 & n16296;
  assign n16298 = n16292 & n16297;
  assign n16299 = ~n16260 & n16298;
  assign n16300 = ~n16270 & n16299;
  assign n16301 = n16243 & ~n16300;
  assign n16302 = n16265 & ~n16294;
  assign n16303 = ~n16270 & n16302;
  assign n16304 = ~n16248 & n16303;
  assign n16305 = ~n16295 & n16304;
  assign n16306 = n16179 & ~n16305;
  assign n16307 = ~n16301 & ~n16306;
  assign n16308 = n16289 & n16307;
  assign n16309 = ~n16267 & n16308;
  assign n16310 = n16258 & n16309;
  assign n16311 = n16310 ^ n13956;
  assign n16312 = n16311 ^ x74;
  assign n16313 = ~n16127 & n16312;
  assign n16314 = n15882 & n16313;
  assign n16315 = n16127 & ~n16312;
  assign n16316 = n15882 & n16315;
  assign n16317 = ~n16314 & ~n16316;
  assign n16318 = n14397 ^ x115;
  assign n16319 = n15539 & n15563;
  assign n16320 = n15549 & n15562;
  assign n16321 = ~n16319 & ~n16320;
  assign n16322 = ~n15591 & n15919;
  assign n16323 = ~n15575 & n16322;
  assign n16324 = n15534 & ~n16323;
  assign n16325 = ~n15537 & n15543;
  assign n16326 = n15474 & ~n16325;
  assign n16327 = ~n15554 & ~n15556;
  assign n16328 = n15539 & ~n16327;
  assign n16329 = ~n15554 & ~n15558;
  assign n16330 = n15562 & ~n16329;
  assign n16331 = ~n15532 & ~n16330;
  assign n16332 = ~n15472 & ~n16331;
  assign n16333 = ~n16328 & ~n16332;
  assign n16334 = ~n16326 & n16333;
  assign n16335 = n15582 & n16334;
  assign n16336 = ~n16324 & n16335;
  assign n16337 = n16321 & n16336;
  assign n16338 = n15912 ^ n15551;
  assign n16339 = n16338 ^ n15551;
  assign n16340 = n15551 ^ n15473;
  assign n16341 = n16340 ^ n15551;
  assign n16342 = ~n16339 & ~n16341;
  assign n16343 = n16342 ^ n15551;
  assign n16344 = n15547 & n16343;
  assign n16345 = n16344 ^ n15551;
  assign n16346 = n16337 & ~n16345;
  assign n16347 = n15908 & n16346;
  assign n16348 = n15578 & n16347;
  assign n16349 = ~n15584 & n16348;
  assign n16350 = n16349 ^ n12643;
  assign n16351 = n16350 ^ x88;
  assign n16352 = ~n16318 & n16351;
  assign n16353 = n15735 & ~n15752;
  assign n16354 = n15653 & ~n16353;
  assign n16355 = ~n15714 & ~n15722;
  assign n16356 = ~n15734 & ~n15756;
  assign n16357 = n15718 & ~n16356;
  assign n16358 = ~n15702 & n15735;
  assign n16359 = n15710 & ~n16358;
  assign n16360 = ~n16357 & ~n16359;
  assign n16361 = ~n16355 & n16360;
  assign n16362 = ~n15754 & n15757;
  assign n16363 = ~n15712 & n16362;
  assign n16364 = n16363 ^ n15738;
  assign n16365 = n16364 ^ n15738;
  assign n16366 = n15738 ^ n15652;
  assign n16367 = n16366 ^ n15738;
  assign n16368 = ~n16365 & ~n16367;
  assign n16369 = n16368 ^ n15738;
  assign n16370 = n15651 & ~n16369;
  assign n16371 = n16370 ^ n15738;
  assign n16372 = n16361 & n16371;
  assign n16373 = n16011 & n16372;
  assign n16374 = n15731 & n16373;
  assign n16375 = n15724 & n16374;
  assign n16376 = ~n16354 & n16375;
  assign n16377 = ~n16008 & n16376;
  assign n16378 = n15709 & n16377;
  assign n16379 = n16378 ^ n13308;
  assign n16380 = n16379 ^ x113;
  assign n16381 = n14609 & n14628;
  assign n16382 = n14402 & ~n14668;
  assign n16383 = ~n16381 & ~n16382;
  assign n16384 = n14606 & n14618;
  assign n16385 = n14622 & n16384;
  assign n16386 = ~n14666 & n15450;
  assign n16387 = n14627 & ~n16386;
  assign n16394 = ~n14625 & ~n14639;
  assign n16388 = ~n14612 & ~n14622;
  assign n16389 = ~n14615 & ~n16388;
  assign n16390 = ~n14607 & n14615;
  assign n16391 = ~n14609 & n16390;
  assign n16392 = ~n14673 & ~n16391;
  assign n16393 = ~n16389 & ~n16392;
  assign n16395 = n16394 ^ n16393;
  assign n16396 = n16393 ^ n14623;
  assign n16397 = n16393 & ~n16396;
  assign n16398 = n16397 ^ n16393;
  assign n16399 = n16395 & n16398;
  assign n16400 = n16399 ^ n16397;
  assign n16401 = n16400 ^ n16393;
  assign n16402 = n16401 ^ n14623;
  assign n16403 = ~n16387 & ~n16402;
  assign n16404 = n16403 ^ n16387;
  assign n16405 = ~n16385 & ~n16404;
  assign n16406 = n16383 & n16405;
  assign n16407 = ~n15966 & n16406;
  assign n16408 = n14649 & n16407;
  assign n16409 = n15439 & n16408;
  assign n16410 = n15944 & n16409;
  assign n16411 = n16410 ^ n11381;
  assign n16412 = n16411 ^ x65;
  assign n16413 = n15086 & ~n15093;
  assign n16414 = n15103 & ~n15631;
  assign n16415 = ~n16413 & ~n16414;
  assign n16416 = n15092 & n15113;
  assign n16417 = ~n15099 & n15620;
  assign n16418 = n15622 & ~n16417;
  assign n16419 = ~n15607 & n15624;
  assign n16420 = n15042 & ~n15622;
  assign n16421 = ~n16419 & ~n16420;
  assign n16422 = ~n15045 & ~n15091;
  assign n16423 = ~n15114 & n16422;
  assign n16424 = n15622 & ~n16423;
  assign n16425 = ~n15609 & n16417;
  assign n16426 = n15088 & ~n16425;
  assign n16427 = ~n16424 & ~n16426;
  assign n16428 = n15047 & n15090;
  assign n16429 = n15130 & n15610;
  assign n16430 = ~n15631 & ~n16429;
  assign n16431 = ~n16428 & ~n16430;
  assign n16432 = n16427 & n16431;
  assign n16433 = n16421 & n16432;
  assign n16434 = ~n16418 & n16433;
  assign n16435 = ~n16416 & n16434;
  assign n16436 = n16415 & n16435;
  assign n16437 = ~n15883 & n16436;
  assign n16438 = n16437 ^ n13273;
  assign n16439 = n16438 ^ x120;
  assign n16440 = n15331 ^ x74;
  assign n16441 = ~n16439 & ~n16440;
  assign n16442 = n16412 & n16441;
  assign n16443 = n16380 & n16442;
  assign n16444 = n16352 & n16443;
  assign n16445 = ~n16318 & ~n16351;
  assign n16446 = n16380 & n16440;
  assign n16447 = n16412 & n16446;
  assign n16448 = ~n16439 & n16447;
  assign n16449 = ~n16412 & n16439;
  assign n16450 = n16440 & n16449;
  assign n16451 = ~n16380 & n16450;
  assign n16452 = ~n16448 & ~n16451;
  assign n16453 = n16445 & ~n16452;
  assign n16454 = ~n16444 & ~n16453;
  assign n16455 = n16318 & n16351;
  assign n16456 = n16412 & n16439;
  assign n16457 = ~n16440 & n16456;
  assign n16458 = n16380 & n16457;
  assign n16459 = n16455 & n16458;
  assign n16460 = ~n16380 & n16412;
  assign n16461 = ~n16439 & n16460;
  assign n16462 = n16440 & n16461;
  assign n16463 = n16352 & n16462;
  assign n16464 = ~n16459 & ~n16463;
  assign n16465 = n16445 & n16458;
  assign n16466 = n16441 & n16460;
  assign n16467 = n16445 & n16466;
  assign n16468 = n16446 & n16456;
  assign n16469 = n16468 ^ n16318;
  assign n16470 = n16469 ^ n16468;
  assign n16471 = n16439 & n16460;
  assign n16472 = ~n16440 & n16471;
  assign n16473 = n16472 ^ n16468;
  assign n16474 = n16470 & n16473;
  assign n16475 = n16474 ^ n16468;
  assign n16476 = n16351 & n16475;
  assign n16477 = ~n16467 & ~n16476;
  assign n16478 = n16318 & ~n16351;
  assign n16479 = ~n16412 & n16441;
  assign n16480 = ~n16380 & n16479;
  assign n16481 = ~n16448 & ~n16480;
  assign n16482 = ~n16458 & n16481;
  assign n16483 = n16478 & ~n16482;
  assign n16484 = ~n16412 & ~n16439;
  assign n16485 = n16446 & n16484;
  assign n16486 = n16352 & n16485;
  assign n16487 = n16443 & n16478;
  assign n16488 = ~n16486 & ~n16487;
  assign n16489 = ~n16462 & ~n16485;
  assign n16490 = n16452 & n16489;
  assign n16491 = n16455 & ~n16490;
  assign n16492 = n16439 ^ n16412;
  assign n16493 = n16440 ^ n16439;
  assign n16494 = ~n16492 & ~n16493;
  assign n16495 = n16494 ^ n16439;
  assign n16496 = ~n16380 & n16495;
  assign n16497 = n16352 & n16496;
  assign n16498 = ~n16491 & ~n16497;
  assign n16499 = n16446 & n16449;
  assign n16500 = ~n16462 & ~n16499;
  assign n16501 = n16445 & ~n16500;
  assign n16502 = ~n16445 & ~n16455;
  assign n16503 = n16380 & n16479;
  assign n16504 = ~n16440 & n16449;
  assign n16505 = n16380 & n16504;
  assign n16506 = ~n16503 & ~n16505;
  assign n16507 = ~n16502 & ~n16506;
  assign n16508 = n16440 & n16471;
  assign n16509 = ~n16499 & ~n16508;
  assign n16510 = n16440 & n16484;
  assign n16511 = ~n16380 & n16510;
  assign n16512 = ~n16380 & n16504;
  assign n16513 = ~n16511 & ~n16512;
  assign n16514 = n16509 & n16513;
  assign n16515 = n16478 & ~n16514;
  assign n16516 = ~n16507 & ~n16515;
  assign n16517 = ~n16501 & n16516;
  assign n16518 = n16498 & n16517;
  assign n16519 = n16488 & n16518;
  assign n16520 = ~n16483 & n16519;
  assign n16521 = n16477 & n16520;
  assign n16522 = ~n16465 & n16521;
  assign n16523 = n16464 & n16522;
  assign n16524 = n16454 & n16523;
  assign n16525 = n16524 ^ n13418;
  assign n16526 = n16525 ^ x88;
  assign n16527 = n16043 ^ x70;
  assign n16528 = n15809 ^ x84;
  assign n16529 = ~n16527 & n16528;
  assign n16530 = n15940 ^ x108;
  assign n16531 = ~n14337 & ~n14358;
  assign n16532 = n14171 & ~n16531;
  assign n16533 = ~n14170 & ~n14377;
  assign n16534 = n14332 & ~n14353;
  assign n16535 = n14335 & n16142;
  assign n16536 = n14332 & ~n14382;
  assign n16537 = ~n16535 & ~n16536;
  assign n16538 = ~n14330 & n14378;
  assign n16539 = n14171 & ~n16538;
  assign n16540 = ~n14344 & ~n14367;
  assign n16541 = ~n14342 & n16540;
  assign n16542 = ~n14365 & n14387;
  assign n16543 = ~n16541 & ~n16542;
  assign n16544 = n16531 & ~n16543;
  assign n16545 = ~n14343 & ~n16544;
  assign n16546 = ~n16539 & ~n16545;
  assign n16547 = n16537 & n16546;
  assign n16548 = n16131 & n16547;
  assign n16549 = ~n16534 & n16548;
  assign n16550 = ~n16533 & n16549;
  assign n16551 = n14386 ^ n14341;
  assign n16552 = n14386 ^ n14342;
  assign n16553 = n16552 ^ n14342;
  assign n16554 = ~n14346 & ~n14375;
  assign n16555 = n16554 ^ n14342;
  assign n16556 = n16553 & n16555;
  assign n16557 = n16556 ^ n14342;
  assign n16558 = ~n16551 & n16557;
  assign n16559 = n16558 ^ n14341;
  assign n16560 = n16550 & ~n16559;
  assign n16561 = ~n16532 & n16560;
  assign n16562 = n16561 ^ n13082;
  assign n16563 = n16562 ^ x102;
  assign n16564 = ~n16530 & ~n16563;
  assign n16565 = n15433 ^ x85;
  assign n16566 = ~n14720 & n15988;
  assign n16567 = n14764 & n14926;
  assign n16568 = ~n16566 & ~n16567;
  assign n16569 = ~n14929 & ~n14938;
  assign n16570 = n14905 & ~n16569;
  assign n16571 = n14905 & ~n14933;
  assign n16572 = ~n14962 & n16211;
  assign n16573 = n14910 & ~n16572;
  assign n16574 = ~n14900 & ~n14920;
  assign n16575 = ~n14765 & n16211;
  assign n16576 = ~n16574 & ~n16575;
  assign n16577 = ~n14940 & ~n16576;
  assign n16578 = ~n14925 & ~n16577;
  assign n16579 = ~n16573 & ~n16578;
  assign n16580 = ~n16571 & n16579;
  assign n16581 = n15978 & n16580;
  assign n16582 = ~n16570 & n16581;
  assign n16583 = n14928 ^ n14765;
  assign n16584 = n14922 ^ n14900;
  assign n16585 = n14928 ^ n14900;
  assign n16586 = n16585 ^ n14900;
  assign n16587 = ~n16584 & ~n16586;
  assign n16588 = n16587 ^ n14900;
  assign n16589 = n16583 & n16588;
  assign n16590 = n16589 ^ n14765;
  assign n16591 = n16582 & ~n16590;
  assign n16592 = n16568 & n16591;
  assign n16593 = n15980 & n16592;
  assign n16594 = ~n15973 & n16593;
  assign n16595 = n16594 ^ n13053;
  assign n16596 = n16595 ^ x83;
  assign n16597 = n16565 & ~n16596;
  assign n16598 = n16564 & n16597;
  assign n16599 = n16529 & n16598;
  assign n16600 = n16527 & n16528;
  assign n16601 = ~n16565 & ~n16596;
  assign n16602 = n16564 & n16601;
  assign n16603 = n16600 & n16602;
  assign n16604 = ~n16527 & ~n16528;
  assign n16605 = n16530 & n16563;
  assign n16606 = n16565 & n16596;
  assign n16607 = n16605 & n16606;
  assign n16608 = ~n16565 & n16596;
  assign n16609 = n16530 & ~n16563;
  assign n16610 = n16608 & n16609;
  assign n16611 = ~n16607 & ~n16610;
  assign n16612 = n16604 & ~n16611;
  assign n16613 = ~n16603 & ~n16612;
  assign n16614 = ~n16599 & n16613;
  assign n16615 = n16598 & n16600;
  assign n16616 = n16527 & ~n16528;
  assign n16617 = n16564 & n16606;
  assign n16618 = ~n16530 & n16563;
  assign n16619 = n16606 & n16618;
  assign n16620 = ~n16617 & ~n16619;
  assign n16621 = n16616 & ~n16620;
  assign n16622 = ~n16615 & ~n16621;
  assign n16623 = n16598 & n16604;
  assign n16624 = n16601 & n16618;
  assign n16625 = ~n16619 & ~n16624;
  assign n16626 = n16600 & ~n16625;
  assign n16627 = ~n16623 & ~n16626;
  assign n16628 = n16597 & n16605;
  assign n16629 = n16600 & n16628;
  assign n16630 = n16597 & n16609;
  assign n16631 = n16616 & n16630;
  assign n16632 = ~n16629 & ~n16631;
  assign n16633 = n16600 & n16630;
  assign n16634 = n16605 & n16608;
  assign n16635 = ~n16628 & ~n16634;
  assign n16636 = n16604 & ~n16635;
  assign n16637 = ~n16633 & ~n16636;
  assign n16638 = n16529 & n16602;
  assign n16639 = n16607 & n16616;
  assign n16640 = n16600 & n16617;
  assign n16641 = ~n16639 & ~n16640;
  assign n16642 = ~n16638 & n16641;
  assign n16643 = n16600 & n16610;
  assign n16644 = n16608 & n16618;
  assign n16645 = ~n16617 & ~n16644;
  assign n16646 = n16604 & ~n16645;
  assign n16647 = ~n16643 & ~n16646;
  assign n16648 = n16601 & n16609;
  assign n16649 = ~n16528 & n16648;
  assign n16650 = n16528 ^ n16527;
  assign n16651 = n16601 & n16605;
  assign n16652 = n16564 & n16608;
  assign n16653 = n16597 & n16618;
  assign n16654 = ~n16652 & ~n16653;
  assign n16655 = ~n16651 & n16654;
  assign n16656 = n16655 ^ n16528;
  assign n16657 = n16656 ^ n16655;
  assign n16658 = n16596 ^ n16565;
  assign n16659 = n16596 ^ n16563;
  assign n16660 = n16563 ^ n16530;
  assign n16661 = n16660 ^ n16563;
  assign n16662 = n16659 & n16661;
  assign n16663 = n16662 ^ n16563;
  assign n16664 = ~n16658 & n16663;
  assign n16665 = n16664 ^ n16563;
  assign n16666 = n16665 ^ n16655;
  assign n16667 = n16657 & ~n16666;
  assign n16668 = n16667 ^ n16655;
  assign n16669 = n16650 & ~n16668;
  assign n16670 = ~n16649 & ~n16669;
  assign n16671 = n16647 & n16670;
  assign n16672 = n16642 & n16671;
  assign n16673 = n16637 & n16672;
  assign n16674 = n16632 & n16673;
  assign n16675 = n16627 & n16674;
  assign n16676 = n16622 & n16675;
  assign n16677 = n16614 & n16676;
  assign n16678 = n16677 ^ n14862;
  assign n16679 = n16678 ^ x98;
  assign n16680 = ~n16526 & ~n16679;
  assign n16681 = ~n16317 & n16680;
  assign n16682 = ~n15398 & ~n15881;
  assign n16683 = ~n16127 & ~n16312;
  assign n16684 = n16682 & n16683;
  assign n16685 = n16526 & n16679;
  assign n16686 = n16684 & n16685;
  assign n16691 = n15882 & n16683;
  assign n16687 = n16127 & n16312;
  assign n16688 = n15882 & n16687;
  assign n16689 = n16315 & n16682;
  assign n16690 = ~n16688 & ~n16689;
  assign n16692 = n16691 ^ n16690;
  assign n16693 = n16692 ^ n16690;
  assign n16694 = n16690 ^ n16685;
  assign n16695 = n16694 ^ n16690;
  assign n16696 = n16693 & ~n16695;
  assign n16697 = n16696 ^ n16690;
  assign n16698 = ~n16680 & ~n16697;
  assign n16699 = n16698 ^ n16690;
  assign n16700 = ~n16686 & n16699;
  assign n16701 = n15398 & n15881;
  assign n16702 = n16315 & n16701;
  assign n16703 = n16526 & ~n16679;
  assign n16704 = n16702 & n16703;
  assign n16705 = n16313 & n16701;
  assign n16706 = ~n16680 & ~n16685;
  assign n16707 = n16705 & n16706;
  assign n16708 = ~n16704 & ~n16707;
  assign n16709 = n16313 & n16682;
  assign n16710 = n16706 & n16709;
  assign n16711 = n15398 & ~n15881;
  assign n16712 = n16683 & n16711;
  assign n16713 = n16712 ^ n16526;
  assign n16714 = n16713 ^ n16712;
  assign n16715 = n16712 ^ n16684;
  assign n16716 = ~n16714 & n16715;
  assign n16717 = n16716 ^ n16712;
  assign n16718 = n16679 & n16717;
  assign n16719 = ~n16710 & ~n16718;
  assign n16720 = n16682 & n16687;
  assign n16721 = ~n16526 & n16679;
  assign n16722 = n16720 & n16721;
  assign n16723 = n16683 & n16701;
  assign n16724 = n16687 & n16711;
  assign n16725 = ~n16723 & ~n16724;
  assign n16726 = n16315 & n16711;
  assign n16727 = ~n16688 & ~n16726;
  assign n16728 = n16317 & n16727;
  assign n16729 = n16725 & n16728;
  assign n16730 = n16685 & ~n16729;
  assign n16731 = ~n16722 & ~n16730;
  assign n16732 = n16687 & n16701;
  assign n16733 = ~n16726 & ~n16732;
  assign n16734 = ~n16724 & n16733;
  assign n16735 = ~n16680 & n16734;
  assign n16736 = n16313 & n16711;
  assign n16737 = n16721 & ~n16733;
  assign n16738 = ~n16712 & ~n16737;
  assign n16739 = ~n16736 & n16738;
  assign n16740 = n16725 & n16739;
  assign n16741 = ~n16735 & ~n16740;
  assign n16742 = n16741 ^ n16679;
  assign n16743 = n16742 ^ n16741;
  assign n16744 = n16733 & ~n16736;
  assign n16745 = ~n16689 & n16744;
  assign n16746 = n16745 ^ n16741;
  assign n16747 = n16746 ^ n16741;
  assign n16748 = ~n16743 & ~n16747;
  assign n16749 = n16748 ^ n16741;
  assign n16750 = n16526 & n16749;
  assign n16751 = n16750 ^ n16741;
  assign n16752 = n16731 & ~n16751;
  assign n16753 = n16719 & n16752;
  assign n16754 = n16708 & n16753;
  assign n16755 = n16700 & n16754;
  assign n16756 = ~n16681 & n16755;
  assign n16757 = n16756 ^ n16043;
  assign n16758 = n16757 ^ x101;
  assign n16759 = n15941 ^ n15900;
  assign n16760 = n16120 ^ n15941;
  assign n16761 = n16760 ^ n16120;
  assign n16762 = n16120 ^ n16110;
  assign n16763 = n16761 & ~n16762;
  assign n16764 = n16763 ^ n16120;
  assign n16765 = n16759 & ~n16764;
  assign n16766 = n16103 ^ n15941;
  assign n16767 = n16766 ^ n16103;
  assign n16768 = n16085 & n16114;
  assign n16769 = n16768 ^ n16103;
  assign n16770 = ~n16767 & n16769;
  assign n16771 = n16770 ^ n16103;
  assign n16772 = ~n16759 & ~n16771;
  assign n16773 = ~n16765 & ~n16772;
  assign n16774 = n16092 & n16773;
  assign n16775 = n16774 ^ n15167;
  assign n16776 = n16775 ^ x126;
  assign n16777 = n16478 & ~n16489;
  assign n16778 = n16455 & n16466;
  assign n16779 = n16352 & ~n16452;
  assign n16780 = ~n16778 & ~n16779;
  assign n16781 = ~n16777 & n16780;
  assign n16782 = n16455 & n16485;
  assign n16783 = ~n16472 & ~n16503;
  assign n16784 = n16318 & ~n16783;
  assign n16785 = ~n16782 & ~n16784;
  assign n16786 = ~n16480 & ~n16505;
  assign n16787 = n16509 & n16786;
  assign n16788 = n16352 & ~n16787;
  assign n16789 = ~n16468 & n16513;
  assign n16790 = ~n16502 & ~n16789;
  assign n16791 = ~n16788 & ~n16790;
  assign n16792 = n16499 ^ n16318;
  assign n16793 = n16792 ^ n16499;
  assign n16794 = ~n16466 & ~n16505;
  assign n16795 = ~n16443 & n16794;
  assign n16796 = n16795 ^ n16499;
  assign n16797 = ~n16793 & ~n16796;
  assign n16798 = n16797 ^ n16499;
  assign n16799 = ~n16351 & n16798;
  assign n16800 = n16791 & ~n16799;
  assign n16801 = n16785 & n16800;
  assign n16802 = ~n16483 & n16801;
  assign n16803 = n16781 & n16802;
  assign n16804 = n16464 & n16803;
  assign n16805 = n16454 & n16804;
  assign n16806 = n16805 ^ n15011;
  assign n16807 = n16806 ^ x77;
  assign n16808 = ~n16776 & n16807;
  assign n16809 = n15143 & n15343;
  assign n16810 = ~n15352 & ~n15370;
  assign n16811 = ~n15364 & ~n16810;
  assign n16812 = ~n16809 & ~n16811;
  assign n16813 = n15340 & n15376;
  assign n16814 = ~n14978 & ~n15377;
  assign n16815 = ~n14974 & n16814;
  assign n16816 = n15344 & ~n16815;
  assign n16817 = ~n16813 & ~n16816;
  assign n16818 = n16812 & n16817;
  assign n16819 = n15333 & ~n15372;
  assign n16820 = ~n15336 & ~n15365;
  assign n16821 = n15358 & ~n16820;
  assign n16822 = n15339 & n15358;
  assign n16823 = n15333 & n15350;
  assign n16824 = ~n16822 & ~n16823;
  assign n16825 = n15358 & ~n16815;
  assign n16826 = ~n14976 & ~n15369;
  assign n16827 = ~n15336 & n16826;
  assign n16828 = n15340 & ~n16827;
  assign n16829 = ~n15357 & ~n15371;
  assign n16830 = ~n15352 & n16829;
  assign n16831 = n15344 & ~n16830;
  assign n16832 = ~n16828 & ~n16831;
  assign n16833 = ~n16825 & n16832;
  assign n16834 = n15348 & n16833;
  assign n16835 = n16824 & n16834;
  assign n16836 = ~n16821 & n16835;
  assign n16837 = ~n16819 & n16836;
  assign n16838 = n16818 & n16837;
  assign n16839 = n15360 & n16838;
  assign n16840 = n16839 ^ n15239;
  assign n16841 = n16840 ^ x94;
  assign n16842 = n16005 ^ x104;
  assign n16843 = n16411 ^ x114;
  assign n16844 = n16842 & n16843;
  assign n16845 = n15899 ^ x90;
  assign n16846 = ~n14343 & n14367;
  assign n16847 = n14341 & ~n16153;
  assign n16848 = ~n16846 & ~n16847;
  assign n16849 = n16142 & ~n16554;
  assign n16850 = n14372 & n14382;
  assign n16851 = ~n14344 & n16850;
  assign n16852 = n14342 & ~n16851;
  assign n16853 = ~n14385 & n16157;
  assign n16854 = n14332 & ~n16853;
  assign n16855 = ~n16852 & ~n16854;
  assign n16856 = ~n16849 & n16855;
  assign n16857 = n16848 & n16856;
  assign n16858 = ~n16151 & n16857;
  assign n16859 = n16149 & n16858;
  assign n16860 = ~n16133 & n16859;
  assign n16861 = ~n16532 & n16860;
  assign n16862 = n16861 ^ n12457;
  assign n16863 = n16862 ^ x107;
  assign n16864 = n16845 & ~n16863;
  assign n16865 = n13986 & n14000;
  assign n16866 = ~n13627 & n16865;
  assign n16867 = ~n13974 & n13976;
  assign n16868 = ~n16866 & ~n16867;
  assign n16869 = n13995 & n13997;
  assign n16870 = ~n13957 & ~n13983;
  assign n16871 = ~n13627 & ~n16870;
  assign n16872 = n13780 & ~n16871;
  assign n16873 = ~n16869 & ~n16872;
  assign n16874 = n16868 & n16873;
  assign n16875 = n16874 ^ n12291;
  assign n16876 = n16875 ^ x72;
  assign n16877 = n16350 ^ x81;
  assign n16878 = n16876 & n16877;
  assign n16879 = n16864 & n16878;
  assign n16880 = n16844 & n16879;
  assign n16881 = n16842 & ~n16843;
  assign n16882 = ~n16845 & ~n16863;
  assign n16883 = ~n16876 & ~n16877;
  assign n16884 = n16882 & n16883;
  assign n16885 = n16881 & n16884;
  assign n16886 = ~n16880 & ~n16885;
  assign n16887 = ~n16876 & n16877;
  assign n16888 = n16864 & n16887;
  assign n16889 = ~n16842 & n16888;
  assign n16890 = ~n16842 & ~n16843;
  assign n16891 = n16845 & n16863;
  assign n16892 = n16878 & n16891;
  assign n16893 = ~n16845 & n16863;
  assign n16894 = n16887 & n16893;
  assign n16895 = ~n16892 & ~n16894;
  assign n16896 = n16890 & ~n16895;
  assign n16897 = ~n16889 & ~n16896;
  assign n16898 = n16876 & ~n16877;
  assign n16899 = n16893 & n16898;
  assign n16900 = ~n16892 & ~n16899;
  assign n16901 = n16844 & ~n16900;
  assign n16902 = n16883 & n16891;
  assign n16903 = n16864 & n16898;
  assign n16904 = n16883 & n16893;
  assign n16905 = ~n16903 & ~n16904;
  assign n16906 = ~n16902 & n16905;
  assign n16907 = n16881 & ~n16906;
  assign n16908 = ~n16901 & ~n16907;
  assign n16909 = ~n16842 & n16843;
  assign n16910 = n16891 & n16898;
  assign n16911 = n16878 & n16882;
  assign n16912 = n16887 & n16891;
  assign n16913 = ~n16911 & ~n16912;
  assign n16914 = ~n16910 & n16913;
  assign n16915 = n16909 & ~n16914;
  assign n16916 = n16876 ^ n16863;
  assign n16917 = n16916 ^ n16845;
  assign n16918 = n16877 & n16917;
  assign n16919 = n16881 & n16918;
  assign n16920 = ~n16884 & ~n16902;
  assign n16921 = n16905 & n16920;
  assign n16922 = n16844 & ~n16921;
  assign n16923 = ~n16919 & ~n16922;
  assign n16924 = n16882 & n16898;
  assign n16925 = n16920 & ~n16924;
  assign n16926 = n16909 & ~n16925;
  assign n16927 = n16882 & n16887;
  assign n16928 = n16864 & n16883;
  assign n16929 = ~n16910 & ~n16928;
  assign n16930 = ~n16904 & n16929;
  assign n16931 = ~n16927 & n16930;
  assign n16932 = ~n16904 & n16925;
  assign n16933 = ~n16890 & n16932;
  assign n16934 = ~n16931 & ~n16933;
  assign n16935 = ~n16926 & ~n16934;
  assign n16936 = n16923 & n16935;
  assign n16937 = ~n16915 & n16936;
  assign n16938 = n16908 & n16937;
  assign n16939 = n16897 & n16938;
  assign n16940 = n16886 & n16939;
  assign n16941 = n16843 ^ n16842;
  assign n16942 = n16879 ^ n16843;
  assign n16943 = n16942 ^ n16879;
  assign n16944 = n16927 ^ n16879;
  assign n16945 = n16943 & n16944;
  assign n16946 = n16945 ^ n16879;
  assign n16947 = ~n16941 & n16946;
  assign n16948 = n16940 & ~n16947;
  assign n16949 = n16948 ^ n15200;
  assign n16950 = n16949 ^ x108;
  assign n16951 = n16841 & ~n16950;
  assign n16952 = ~n16271 & ~n16293;
  assign n16953 = n16259 & ~n16952;
  assign n16954 = ~n16243 & ~n16251;
  assign n16955 = n16241 & ~n16954;
  assign n16956 = n16243 & ~n16292;
  assign n16957 = ~n16955 & ~n16956;
  assign n16958 = n16244 & n16247;
  assign n16959 = ~n16294 & ~n16958;
  assign n16960 = ~n16290 & n16959;
  assign n16961 = n16259 & ~n16960;
  assign n16962 = ~n16264 & n16274;
  assign n16963 = n16243 & ~n16962;
  assign n16964 = ~n16961 & ~n16963;
  assign n16965 = n16179 & ~n16287;
  assign n16966 = n16304 & ~n16958;
  assign n16967 = ~n16291 & n16966;
  assign n16968 = n16251 & ~n16967;
  assign n16969 = ~n16965 & ~n16968;
  assign n16970 = n16964 & n16969;
  assign n16971 = ~n16267 & n16970;
  assign n16972 = n16957 & n16971;
  assign n16973 = ~n16953 & n16972;
  assign n16974 = n16973 ^ n15259;
  assign n16975 = n16974 ^ x83;
  assign n16976 = n15823 & n15834;
  assign n16977 = n15830 & n16976;
  assign n16978 = ~n15434 & n15470;
  assign n16979 = ~n15828 & ~n15831;
  assign n16980 = n16978 & ~n16979;
  assign n16981 = ~n16977 & ~n16980;
  assign n16982 = ~n15470 & n15846;
  assign n16983 = ~n15835 & ~n15864;
  assign n16984 = n15471 & ~n16983;
  assign n16985 = ~n16982 & ~n16984;
  assign n16986 = ~n15818 & n15849;
  assign n16987 = n15838 & ~n15864;
  assign n16988 = n15840 & ~n16987;
  assign n16989 = ~n16986 & ~n16988;
  assign n16990 = ~n15815 & ~n15820;
  assign n16991 = n16978 & ~n16990;
  assign n16992 = ~n15831 & ~n15841;
  assign n16993 = ~n15820 & n16992;
  assign n16994 = ~n15822 & n16993;
  assign n16995 = n15830 & ~n16994;
  assign n16996 = ~n15824 & ~n15837;
  assign n16997 = ~n15812 & n16979;
  assign n16998 = n15840 & ~n16997;
  assign n16999 = n16996 & ~n16998;
  assign n17000 = ~n15818 & ~n16999;
  assign n17001 = ~n15848 & ~n16976;
  assign n17002 = n15841 & ~n16994;
  assign n17003 = n17001 & ~n17002;
  assign n17004 = ~n15842 & n17003;
  assign n17005 = n16978 & ~n17004;
  assign n17006 = ~n17000 & ~n17005;
  assign n17007 = ~n16995 & n17006;
  assign n17008 = ~n15817 & n17007;
  assign n17009 = ~n16991 & n17008;
  assign n17010 = n16989 & n17009;
  assign n17011 = n16985 & n17010;
  assign n17012 = n16981 & n17011;
  assign n17013 = ~n15839 & n17012;
  assign n17014 = n17013 ^ n15084;
  assign n17015 = n17014 ^ x109;
  assign n17016 = ~n16975 & n17015;
  assign n17017 = n16951 & n17016;
  assign n17018 = n16808 & n17017;
  assign n17019 = ~n16776 & ~n16807;
  assign n17020 = n16841 & n16950;
  assign n17021 = n16975 & n17015;
  assign n17022 = n17020 & n17021;
  assign n17023 = n17019 & n17022;
  assign n17024 = ~n17018 & ~n17023;
  assign n17025 = n17017 & n17019;
  assign n17026 = n16776 & ~n16807;
  assign n17027 = ~n16975 & ~n17015;
  assign n17028 = n17020 & n17027;
  assign n17029 = ~n16841 & ~n16950;
  assign n17030 = n16975 & ~n17015;
  assign n17031 = n17029 & n17030;
  assign n17032 = ~n17028 & ~n17031;
  assign n17033 = n17026 & ~n17032;
  assign n17034 = ~n17025 & ~n17033;
  assign n17035 = ~n16841 & n16950;
  assign n17036 = n17021 & n17035;
  assign n17037 = n16951 & n17021;
  assign n17038 = n17016 & n17029;
  assign n17039 = ~n17037 & ~n17038;
  assign n17040 = ~n17036 & n17039;
  assign n17041 = n16808 & ~n17040;
  assign n17042 = n16776 & n16807;
  assign n17043 = n17027 & n17035;
  assign n17044 = ~n17037 & ~n17043;
  assign n17045 = n17042 & ~n17044;
  assign n17046 = ~n17041 & ~n17045;
  assign n17047 = ~n16808 & ~n17026;
  assign n17048 = n17016 & n17035;
  assign n17049 = n17021 & n17029;
  assign n17050 = ~n17048 & ~n17049;
  assign n17051 = n17047 & ~n17050;
  assign n17052 = n17030 & n17035;
  assign n17053 = ~n17017 & ~n17052;
  assign n17054 = n17026 & ~n17053;
  assign n17055 = n17022 & n17026;
  assign n17056 = n17027 & n17029;
  assign n17057 = n17020 & n17030;
  assign n17058 = n16951 & n17027;
  assign n17059 = ~n17057 & ~n17058;
  assign n17060 = ~n17056 & n17059;
  assign n17061 = n17042 & ~n17060;
  assign n17062 = ~n17055 & ~n17061;
  assign n17063 = n17016 & n17020;
  assign n17064 = ~n17036 & ~n17038;
  assign n17065 = ~n17063 & n17064;
  assign n17066 = n17026 & ~n17065;
  assign n17067 = ~n17043 & ~n17057;
  assign n17068 = ~n17052 & ~n17056;
  assign n17069 = n17067 & n17068;
  assign n17070 = n16808 & ~n17069;
  assign n17071 = ~n17066 & ~n17070;
  assign n17072 = n17028 & n17042;
  assign n17073 = n16951 & n17030;
  assign n17074 = ~n17028 & ~n17073;
  assign n17075 = ~n17031 & n17074;
  assign n17076 = ~n17056 & n17075;
  assign n17077 = n17019 & ~n17076;
  assign n17078 = ~n17072 & ~n17077;
  assign n17079 = n17071 & n17078;
  assign n17080 = n17062 & n17079;
  assign n17081 = ~n17054 & n17080;
  assign n17082 = ~n17051 & n17081;
  assign n17083 = n17046 & n17082;
  assign n17084 = n17034 & n17083;
  assign n17085 = n17024 & n17084;
  assign n17086 = n17085 ^ n15809;
  assign n17087 = n17086 ^ x83;
  assign n17088 = n16758 & n17087;
  assign n17089 = n16083 & n16094;
  assign n17090 = n16098 & ~n17089;
  assign n17091 = n16076 & n16089;
  assign n17092 = ~n16093 & ~n17091;
  assign n17093 = n17090 & n17092;
  assign n17094 = n16080 & ~n17093;
  assign n17095 = n16076 ^ n15972;
  assign n17096 = n17095 ^ n15972;
  assign n17097 = n16076 ^ n16044;
  assign n17098 = n17097 ^ n15972;
  assign n17099 = n17098 ^ n15972;
  assign n17100 = n17096 & n17099;
  assign n17101 = n17100 ^ n15972;
  assign n17102 = ~n16006 & ~n17101;
  assign n17103 = n17102 ^ n17097;
  assign n17104 = n16088 & n17103;
  assign n17105 = ~n17094 & ~n17104;
  assign n17106 = n16081 & n16090;
  assign n17107 = ~n16091 & ~n17106;
  assign n17108 = n16081 & n16096;
  assign n17109 = ~n16108 & ~n17108;
  assign n17110 = n16113 & n17109;
  assign n17111 = n17107 & n17110;
  assign n17112 = n15942 & ~n17111;
  assign n17113 = ~n16082 & n17092;
  assign n17114 = n16102 & n17113;
  assign n17115 = n17107 & n17114;
  assign n17116 = n16106 & ~n17115;
  assign n17117 = ~n17112 & ~n17116;
  assign n17118 = n17105 & n17117;
  assign n17119 = n16087 & n17118;
  assign n17120 = n17119 ^ n14138;
  assign n17121 = n17120 ^ x75;
  assign n17122 = n16529 & n16644;
  assign n17123 = n16600 & n16634;
  assign n17124 = n16604 & n16630;
  assign n17125 = ~n17123 & ~n17124;
  assign n17126 = ~n17122 & n17125;
  assign n17127 = n16529 & ~n16654;
  assign n17128 = n16627 & ~n17127;
  assign n17129 = n16602 & n16616;
  assign n17130 = n16606 & n16609;
  assign n17131 = ~n16648 & ~n17130;
  assign n17132 = ~n16630 & ~n16634;
  assign n17133 = n17131 & n17132;
  assign n17134 = ~n16619 & n17133;
  assign n17135 = n16529 & ~n17134;
  assign n17136 = ~n16628 & ~n16651;
  assign n17137 = ~n17130 & n17136;
  assign n17138 = n16600 & ~n17137;
  assign n17139 = n17132 & n17136;
  assign n17140 = n16616 & ~n17139;
  assign n17141 = ~n16653 & n17131;
  assign n17142 = n16611 & n17141;
  assign n17143 = n16604 & ~n17142;
  assign n17144 = ~n17140 & ~n17143;
  assign n17145 = ~n17138 & n17144;
  assign n17146 = ~n17135 & n17145;
  assign n17147 = ~n17129 & n17146;
  assign n17148 = n16624 ^ n16527;
  assign n17149 = n17148 ^ n16624;
  assign n17150 = n16652 ^ n16624;
  assign n17151 = n17150 ^ n16624;
  assign n17152 = n17149 & n17151;
  assign n17153 = n17152 ^ n16624;
  assign n17154 = n16528 & n17153;
  assign n17155 = n17154 ^ n16624;
  assign n17156 = n17147 & ~n17155;
  assign n17157 = n17128 & n17156;
  assign n17158 = n17126 & n17157;
  assign n17159 = n16622 & n17158;
  assign n17160 = n17159 ^ n14169;
  assign n17161 = n17160 ^ x124;
  assign n17162 = n17121 & ~n17161;
  assign n17163 = n14005 ^ x75;
  assign n17164 = n16238 ^ x93;
  assign n17165 = ~n17163 & n17164;
  assign n17166 = n15142 ^ x68;
  assign n17167 = n15539 & n15583;
  assign n17168 = n15534 & ~n15592;
  assign n17169 = ~n17167 & ~n17168;
  assign n17170 = n15562 & ~n15593;
  assign n17171 = ~n15542 & n15924;
  assign n17172 = ~n15549 & n17171;
  assign n17173 = n15474 & ~n17172;
  assign n17174 = ~n15547 & ~n15918;
  assign n17175 = n15569 & ~n15579;
  assign n17176 = ~n15563 & n17175;
  assign n17177 = n15534 & ~n17176;
  assign n17178 = ~n17174 & ~n17177;
  assign n17179 = n15474 & ~n15594;
  assign n17180 = n15919 & n15924;
  assign n17181 = n15539 & ~n17180;
  assign n17182 = ~n15575 & n16325;
  assign n17183 = n15562 & ~n17182;
  assign n17184 = ~n17181 & ~n17183;
  assign n17185 = ~n17179 & n17184;
  assign n17186 = n17178 & n17185;
  assign n17187 = ~n17173 & n17186;
  assign n17188 = ~n17170 & n17187;
  assign n17189 = n17169 & n17188;
  assign n17190 = n15911 & n17189;
  assign n17191 = ~n15572 & n17190;
  assign n17192 = n17191 ^ n13510;
  assign n17193 = n17192 ^ x110;
  assign n17194 = n17166 & n17193;
  assign n17195 = n15738 & ~n15756;
  assign n17196 = n15653 & ~n17195;
  assign n17197 = ~n15756 & n16353;
  assign n17198 = n15729 & n17197;
  assign n17199 = n15722 & n17198;
  assign n17200 = n15704 & ~n17199;
  assign n17201 = ~n17196 & ~n17200;
  assign n17202 = n15718 & ~n15757;
  assign n17203 = ~n15737 & n15759;
  assign n17204 = n15710 & ~n17203;
  assign n17207 = ~n15721 & n15729;
  assign n17205 = ~n15716 & n15722;
  assign n17206 = ~n15702 & n17205;
  assign n17208 = n17207 ^ n17206;
  assign n17209 = n17207 ^ n15652;
  assign n17210 = n17209 ^ n17207;
  assign n17211 = n17208 & n17210;
  assign n17212 = n17211 ^ n17207;
  assign n17213 = ~n15651 & ~n17212;
  assign n17214 = ~n17204 & ~n17213;
  assign n17215 = ~n17202 & n17214;
  assign n17216 = n17201 & n17215;
  assign n17217 = ~n16013 & n17216;
  assign n17218 = ~n16354 & n17217;
  assign n17219 = ~n15713 & n17218;
  assign n17220 = ~n16008 & n17219;
  assign n17221 = ~n15733 & n17220;
  assign n17222 = n17221 ^ n13480;
  assign n17223 = n17222 ^ x124;
  assign n17224 = n16177 ^ x125;
  assign n17225 = n17223 & n17224;
  assign n17226 = n17194 & n17225;
  assign n17227 = ~n17166 & n17193;
  assign n17228 = ~n17223 & n17224;
  assign n17229 = n17227 & n17228;
  assign n17230 = ~n17226 & ~n17229;
  assign n17231 = n17165 & ~n17230;
  assign n17232 = ~n17166 & ~n17193;
  assign n17233 = n17228 & n17232;
  assign n17234 = ~n17163 & ~n17164;
  assign n17235 = n17233 & n17234;
  assign n17236 = n17223 & ~n17224;
  assign n17237 = n17232 & n17236;
  assign n17238 = n17163 & ~n17164;
  assign n17239 = n17237 & n17238;
  assign n17240 = ~n17235 & ~n17239;
  assign n17241 = ~n17231 & n17240;
  assign n17242 = ~n17223 & ~n17224;
  assign n17243 = n17227 & n17242;
  assign n17244 = n17163 & n17164;
  assign n17245 = n17243 & n17244;
  assign n17246 = n17232 & n17242;
  assign n17247 = n17166 & ~n17193;
  assign n17248 = n17236 & n17247;
  assign n17249 = ~n17246 & ~n17248;
  assign n17250 = n17244 & ~n17249;
  assign n17251 = ~n17245 & ~n17250;
  assign n17252 = n17225 & n17247;
  assign n17253 = n17238 & n17252;
  assign n17254 = n17228 & n17247;
  assign n17255 = n17165 & n17254;
  assign n17256 = n17225 & n17227;
  assign n17257 = n17244 & n17256;
  assign n17258 = ~n17255 & ~n17257;
  assign n17259 = ~n17253 & n17258;
  assign n17260 = n17229 & n17238;
  assign n17261 = n17165 & n17233;
  assign n17262 = n17194 & n17228;
  assign n17263 = n17244 & n17262;
  assign n17264 = n17193 ^ n17166;
  assign n17265 = n17225 & ~n17264;
  assign n17266 = n17238 & n17265;
  assign n17267 = ~n17263 & ~n17266;
  assign n17268 = ~n17261 & n17267;
  assign n17269 = ~n17260 & n17268;
  assign n17270 = n17194 & n17242;
  assign n17271 = n17194 & n17236;
  assign n17272 = ~n17270 & ~n17271;
  assign n17273 = ~n17233 & n17272;
  assign n17274 = n17238 & ~n17273;
  assign n17275 = n17227 & n17236;
  assign n17276 = ~n17248 & ~n17275;
  assign n17277 = ~n17243 & n17276;
  assign n17278 = ~n17271 & n17277;
  assign n17279 = n17165 & ~n17278;
  assign n17280 = ~n17274 & ~n17279;
  assign n17281 = ~n17237 & ~n17275;
  assign n17282 = ~n17254 & n17281;
  assign n17283 = n17244 & ~n17282;
  assign n17284 = n17242 & n17247;
  assign n17285 = ~n17237 & ~n17284;
  assign n17286 = ~n17243 & ~n17256;
  assign n17287 = ~n17252 & n17286;
  assign n17288 = ~n17270 & n17287;
  assign n17289 = ~n17262 & n17288;
  assign n17290 = n17285 & n17289;
  assign n17291 = n17234 & ~n17290;
  assign n17292 = ~n17283 & ~n17291;
  assign n17293 = n17280 & n17292;
  assign n17294 = n17269 & n17293;
  assign n17295 = n17259 & n17294;
  assign n17296 = n17251 & n17295;
  assign n17297 = n17241 & n17296;
  assign n17298 = n17297 ^ n14278;
  assign n17299 = n17298 ^ x125;
  assign n17300 = ~n16892 & ~n16911;
  assign n17301 = n16909 & ~n17300;
  assign n17302 = n16881 & ~n16895;
  assign n17303 = ~n16844 & ~n16890;
  assign n17304 = n16910 & ~n17303;
  assign n17305 = ~n17302 & ~n17304;
  assign n17306 = n16881 & n16899;
  assign n17307 = n16924 & ~n17303;
  assign n17308 = ~n17306 & ~n17307;
  assign n17309 = n16844 & ~n16920;
  assign n17310 = ~n16894 & ~n16899;
  assign n17311 = n16930 & n17310;
  assign n17312 = ~n16888 & n17311;
  assign n17313 = n16909 & ~n17312;
  assign n17314 = ~n16903 & ~n16928;
  assign n17315 = ~n16904 & n17314;
  assign n17316 = ~n16924 & n17315;
  assign n17317 = ~n16927 & n17316;
  assign n17318 = n16881 & ~n17317;
  assign n17319 = ~n17313 & ~n17318;
  assign n17320 = ~n17309 & n17319;
  assign n17321 = n16878 & n16893;
  assign n17322 = ~n16880 & ~n16927;
  assign n17323 = ~n16912 & n17322;
  assign n17324 = ~n17321 & n17323;
  assign n17325 = n17324 ^ n16890;
  assign n17326 = n17324 ^ n16844;
  assign n17327 = n17326 ^ n16844;
  assign n17328 = n17314 ^ n16844;
  assign n17329 = n17327 & n17328;
  assign n17330 = n17329 ^ n16844;
  assign n17331 = ~n17325 & n17330;
  assign n17332 = n17331 ^ n16890;
  assign n17333 = n17320 & ~n17332;
  assign n17334 = n17308 & n17333;
  assign n17335 = n17305 & n17334;
  assign n17336 = ~n17301 & n17335;
  assign n17337 = ~n16947 & n17336;
  assign n17338 = n17337 ^ n14241;
  assign n17339 = n17338 ^ x118;
  assign n17340 = ~n17299 & ~n17339;
  assign n17341 = ~n14974 & ~n15369;
  assign n17342 = n15358 & ~n17341;
  assign n17343 = n15372 & n16815;
  assign n17344 = ~n15343 & n17343;
  assign n17345 = n15333 & ~n17344;
  assign n17346 = ~n17342 & ~n17345;
  assign n17347 = n14976 & n15143;
  assign n17348 = ~n15343 & ~n15366;
  assign n17349 = ~n15352 & n17348;
  assign n17350 = n14979 & n17349;
  assign n17351 = ~n15350 & n17350;
  assign n17352 = ~n15339 & n17351;
  assign n17353 = n15344 & ~n17352;
  assign n17356 = ~n15370 & n16829;
  assign n17357 = ~n15365 & n17356;
  assign n17354 = n15367 & ~n15376;
  assign n17355 = ~n15357 & n17354;
  assign n17358 = n17357 ^ n17355;
  assign n17359 = n17357 ^ n15332;
  assign n17360 = n17359 ^ n17357;
  assign n17361 = n17358 & ~n17360;
  assign n17362 = n17361 ^ n17357;
  assign n17363 = n15143 & ~n17362;
  assign n17364 = ~n17353 & ~n17363;
  assign n17365 = ~n17347 & n17364;
  assign n17366 = n17346 & n17365;
  assign n17367 = ~n15391 & n17366;
  assign n17368 = n15355 & n17367;
  assign n17369 = n16824 & n17368;
  assign n17370 = n17369 ^ n14200;
  assign n17371 = n17370 ^ x85;
  assign n17372 = n16179 & ~n16272;
  assign n17373 = n16251 & n16290;
  assign n17374 = n16240 & n16263;
  assign n17375 = ~n16260 & ~n17374;
  assign n17376 = n16259 & ~n17375;
  assign n17377 = ~n17373 & ~n17376;
  assign n17378 = ~n17372 & n17377;
  assign n17379 = n16179 & n17374;
  assign n17380 = n16248 & n16251;
  assign n17381 = ~n17379 & ~n17380;
  assign n17382 = n16259 & n16291;
  assign n17383 = ~n16246 & n16297;
  assign n17384 = ~n16264 & n17383;
  assign n17385 = n16251 & ~n17384;
  assign n17386 = ~n17382 & ~n17385;
  assign n17387 = ~n16260 & ~n16262;
  assign n17388 = ~n16269 & ~n16295;
  assign n17389 = ~n16246 & n17388;
  assign n17390 = n17387 & n17389;
  assign n17391 = n16179 & ~n17390;
  assign n17392 = ~n16270 & ~n16958;
  assign n17393 = ~n16248 & n17392;
  assign n17394 = n17393 ^ n17389;
  assign n17395 = n16178 ^ n16128;
  assign n17396 = n17395 ^ n16128;
  assign n17397 = n17393 ^ n16128;
  assign n17398 = ~n17396 & n17397;
  assign n17399 = n17398 ^ n16128;
  assign n17400 = n17394 & n17399;
  assign n17401 = n17400 ^ n17389;
  assign n17402 = ~n16293 & n17401;
  assign n17403 = n17402 ^ n16262;
  assign n17404 = n17402 ^ n16178;
  assign n17405 = n17402 & n17404;
  assign n17406 = n17405 ^ n17402;
  assign n17407 = ~n17403 & n17406;
  assign n17408 = n17407 ^ n17405;
  assign n17409 = n17408 ^ n17402;
  assign n17410 = n17409 ^ n16178;
  assign n17411 = ~n17391 & n17410;
  assign n17412 = n17411 ^ n17391;
  assign n17413 = n17386 & ~n17412;
  assign n17414 = n17381 & n17413;
  assign n17415 = n17378 & n17414;
  assign n17416 = n16957 & n17415;
  assign n17417 = n17416 ^ n14327;
  assign n17418 = n17417 ^ x100;
  assign n17419 = n17371 & n17418;
  assign n17420 = n17340 & n17419;
  assign n17421 = n17162 & n17420;
  assign n17422 = ~n17121 & ~n17161;
  assign n17423 = ~n17299 & n17339;
  assign n17424 = n17419 & n17423;
  assign n17425 = n17422 & n17424;
  assign n17426 = n17121 & n17161;
  assign n17427 = n17299 & n17339;
  assign n17428 = n17419 & n17427;
  assign n17429 = n17299 & ~n17339;
  assign n17430 = ~n17371 & n17418;
  assign n17431 = n17429 & n17430;
  assign n17432 = ~n17428 & ~n17431;
  assign n17433 = n17426 & ~n17432;
  assign n17434 = ~n17425 & ~n17433;
  assign n17435 = ~n17421 & n17434;
  assign n17436 = ~n17422 & ~n17426;
  assign n17437 = n17423 & n17430;
  assign n17438 = ~n17371 & ~n17418;
  assign n17439 = n17340 & n17438;
  assign n17440 = ~n17437 & ~n17439;
  assign n17441 = ~n17436 & ~n17440;
  assign n17442 = n17371 & ~n17418;
  assign n17443 = n17429 & n17442;
  assign n17444 = n17162 & n17443;
  assign n17445 = n17419 & n17429;
  assign n17446 = n17427 & n17442;
  assign n17447 = ~n17445 & ~n17446;
  assign n17448 = n17422 & ~n17447;
  assign n17449 = ~n17444 & ~n17448;
  assign n17450 = ~n17441 & n17449;
  assign n17451 = n17427 & n17430;
  assign n17452 = n17427 & n17438;
  assign n17453 = ~n17443 & ~n17452;
  assign n17454 = ~n17451 & n17453;
  assign n17455 = ~n17121 & ~n17454;
  assign n17456 = n17340 & n17442;
  assign n17457 = n17423 & n17438;
  assign n17458 = n17447 & ~n17457;
  assign n17459 = ~n17456 & n17458;
  assign n17460 = n17426 & ~n17459;
  assign n17461 = ~n17455 & ~n17460;
  assign n17462 = n17339 ^ n17299;
  assign n17463 = n17371 ^ n17299;
  assign n17464 = n17463 ^ n17339;
  assign n17465 = n17463 ^ n17418;
  assign n17466 = ~n17464 & n17465;
  assign n17467 = n17466 ^ n17463;
  assign n17468 = ~n17462 & n17467;
  assign n17469 = n17468 ^ n17463;
  assign n17470 = n17162 & n17469;
  assign n17471 = ~n17121 & n17161;
  assign n17472 = n17423 & n17442;
  assign n17473 = ~n17439 & ~n17472;
  assign n17474 = ~n17437 & n17473;
  assign n17475 = ~n17445 & n17474;
  assign n17476 = ~n17456 & n17475;
  assign n17477 = n17471 & ~n17476;
  assign n17478 = ~n17470 & ~n17477;
  assign n17479 = n17461 & n17478;
  assign n17480 = n17450 & n17479;
  assign n17481 = n17435 & n17480;
  assign n17482 = n17481 ^ n16562;
  assign n17483 = n17482 ^ x70;
  assign n17484 = n15397 ^ x72;
  assign n17485 = n15471 & ~n16979;
  assign n17486 = n15434 & n15820;
  assign n17487 = n15828 & n15840;
  assign n17488 = ~n17486 & ~n17487;
  assign n17489 = ~n15812 & ~n15822;
  assign n17490 = ~n15818 & ~n17489;
  assign n17491 = n15816 & ~n15841;
  assign n17492 = n15830 & ~n17491;
  assign n17493 = ~n17490 & ~n17492;
  assign n17494 = n15838 & n15850;
  assign n17495 = n16978 & ~n17494;
  assign n17496 = ~n15824 & n16993;
  assign n17497 = n16978 & ~n17496;
  assign n17498 = n15865 & ~n16976;
  assign n17499 = ~n15846 & n17498;
  assign n17500 = n15840 & ~n17499;
  assign n17501 = ~n17497 & ~n17500;
  assign n17502 = n15824 ^ n15470;
  assign n17503 = n15847 & ~n15864;
  assign n17504 = n17503 ^ n15848;
  assign n17505 = n15848 ^ n15434;
  assign n17506 = n17505 ^ n15848;
  assign n17507 = ~n17504 & ~n17506;
  assign n17508 = n17507 ^ n15848;
  assign n17509 = n17508 ^ n15824;
  assign n17510 = n17502 & n17509;
  assign n17511 = n17510 ^ n17507;
  assign n17512 = n17511 ^ n15848;
  assign n17513 = n17512 ^ n15470;
  assign n17514 = ~n15824 & n17513;
  assign n17515 = n17514 ^ n15824;
  assign n17516 = n17515 ^ n15470;
  assign n17517 = n17501 & ~n17516;
  assign n17518 = ~n15839 & n17517;
  assign n17519 = ~n17495 & n17518;
  assign n17520 = n17493 & n17519;
  assign n17521 = n17488 & n17520;
  assign n17522 = ~n17485 & n17521;
  assign n17523 = n17522 ^ n14763;
  assign n17524 = n17523 ^ x99;
  assign n17525 = n17484 & n17524;
  assign n17526 = n16243 & ~n16265;
  assign n17527 = ~n16264 & ~n16291;
  assign n17528 = ~n16293 & n17527;
  assign n17529 = n16179 & ~n17528;
  assign n17530 = ~n17526 & ~n17529;
  assign n17531 = ~n16270 & ~n16295;
  assign n17532 = n16259 & ~n17531;
  assign n17533 = n16959 & n17388;
  assign n17534 = ~n16954 & ~n17533;
  assign n17535 = ~n17532 & ~n17534;
  assign n17536 = n17530 & n17535;
  assign n17537 = n17387 ^ n16290;
  assign n17538 = n17537 ^ n16290;
  assign n17539 = n16290 ^ n16128;
  assign n17540 = n17539 ^ n16290;
  assign n17541 = ~n17538 & n17540;
  assign n17542 = n17541 ^ n16290;
  assign n17543 = ~n16178 & n17542;
  assign n17544 = n17543 ^ n16290;
  assign n17545 = n17536 & ~n17544;
  assign n17546 = n17381 & n17545;
  assign n17547 = n16258 & n17546;
  assign n17548 = n17378 & n17547;
  assign n17549 = ~n16953 & n17548;
  assign n17550 = n17549 ^ n14895;
  assign n17551 = n17550 ^ x104;
  assign n17552 = n16890 & n16904;
  assign n17553 = n16909 & ~n16920;
  assign n17554 = ~n17552 & ~n17553;
  assign n17555 = ~n16884 & n16905;
  assign n17556 = n16844 & ~n17555;
  assign n17557 = n16925 & ~n16928;
  assign n17558 = ~n16879 & n17557;
  assign n17559 = ~n17321 & n17558;
  assign n17560 = n16881 & ~n17559;
  assign n17561 = ~n17556 & ~n17560;
  assign n17562 = ~n16927 & n17303;
  assign n17563 = n16842 & ~n16879;
  assign n17564 = ~n17322 & ~n17563;
  assign n17565 = n16913 & ~n17564;
  assign n17566 = ~n17562 & ~n17565;
  assign n17567 = ~n16888 & ~n17566;
  assign n17568 = n17567 ^ n16842;
  assign n17569 = n17567 ^ n16843;
  assign n17570 = n17569 ^ n16843;
  assign n17571 = ~n16899 & ~n16903;
  assign n17572 = n17571 ^ n16843;
  assign n17573 = n17570 & n17572;
  assign n17574 = n17573 ^ n16843;
  assign n17575 = n17568 & n17574;
  assign n17576 = n17575 ^ n16842;
  assign n17577 = n17561 & n17576;
  assign n17578 = n17554 & n17577;
  assign n17579 = n17305 & n17578;
  assign n17580 = ~n17301 & n17579;
  assign n17581 = n17580 ^ n14787;
  assign n17582 = n17581 ^ x97;
  assign n17583 = ~n17551 & ~n17582;
  assign n17584 = n17244 & n17270;
  assign n17585 = n17238 & ~n17276;
  assign n17586 = ~n17584 & ~n17585;
  assign n17587 = n17165 & n17246;
  assign n17588 = n17234 & ~n17285;
  assign n17589 = ~n17587 & ~n17588;
  assign n17590 = ~n17229 & ~n17252;
  assign n17591 = n17234 & ~n17590;
  assign n17592 = n17238 & n17246;
  assign n17593 = ~n17591 & ~n17592;
  assign n17594 = ~n17163 & ~n17272;
  assign n17595 = n17165 & ~n17287;
  assign n17596 = ~n17594 & ~n17595;
  assign n17597 = n17234 & n17265;
  assign n17598 = ~n17254 & ~n17271;
  assign n17599 = n17238 & ~n17598;
  assign n17600 = n17225 & n17232;
  assign n17601 = ~n17252 & ~n17600;
  assign n17602 = ~n17246 & n17601;
  assign n17603 = n17285 & n17602;
  assign n17604 = n17244 & ~n17603;
  assign n17605 = ~n17599 & ~n17604;
  assign n17606 = ~n17597 & n17605;
  assign n17607 = n17596 & n17606;
  assign n17608 = n17258 & n17607;
  assign n17609 = n17593 & n17608;
  assign n17610 = n17269 & n17609;
  assign n17611 = n17589 & n17610;
  assign n17612 = n17586 & n17611;
  assign n17613 = n17612 ^ n14827;
  assign n17614 = n17613 ^ x123;
  assign n17615 = n16678 ^ x114;
  assign n17616 = ~n17614 & ~n17615;
  assign n17617 = n17583 & n17616;
  assign n17618 = n17525 & n17617;
  assign n17619 = n17484 & ~n17524;
  assign n17620 = n17551 & n17582;
  assign n17621 = n17614 & ~n17615;
  assign n17622 = n17620 & n17621;
  assign n17623 = n17619 & n17622;
  assign n17624 = ~n17618 & ~n17623;
  assign n17625 = ~n17614 & n17615;
  assign n17626 = n17583 & n17625;
  assign n17627 = n17525 & n17626;
  assign n17628 = ~n17484 & ~n17524;
  assign n17629 = n17617 & n17628;
  assign n17630 = ~n17627 & ~n17629;
  assign n17631 = n17524 ^ n17484;
  assign n17632 = ~n17551 & n17582;
  assign n17633 = n17625 & n17632;
  assign n17634 = ~n17631 & n17633;
  assign n17635 = n17621 & n17632;
  assign n17636 = n17614 & n17615;
  assign n17637 = n17620 & n17636;
  assign n17638 = ~n17582 & n17636;
  assign n17639 = n17551 & n17638;
  assign n17640 = ~n17637 & ~n17639;
  assign n17641 = ~n17635 & n17640;
  assign n17642 = n17619 & ~n17641;
  assign n17643 = ~n17634 & ~n17642;
  assign n17644 = ~n17484 & n17524;
  assign n17645 = n17551 & ~n17582;
  assign n17646 = n17625 & n17645;
  assign n17647 = n17620 & n17625;
  assign n17648 = n17616 & n17645;
  assign n17649 = ~n17647 & ~n17648;
  assign n17650 = ~n17646 & n17649;
  assign n17651 = n17644 & ~n17650;
  assign n17652 = n17619 & n17626;
  assign n17653 = n17525 & n17639;
  assign n17654 = n17632 & n17636;
  assign n17655 = n17621 & n17645;
  assign n17656 = ~n17654 & ~n17655;
  assign n17657 = n17628 & ~n17656;
  assign n17658 = ~n17653 & ~n17657;
  assign n17659 = ~n17652 & n17658;
  assign n17660 = n17583 & n17621;
  assign n17661 = ~n17639 & ~n17660;
  assign n17662 = n17628 & ~n17661;
  assign n17663 = ~n17633 & ~n17648;
  assign n17664 = ~n17617 & n17663;
  assign n17665 = n17619 & ~n17664;
  assign n17666 = n17644 & n17654;
  assign n17667 = ~n17551 & n17638;
  assign n17668 = ~n17635 & ~n17667;
  assign n17669 = ~n17666 & n17668;
  assign n17670 = ~n17622 & n17669;
  assign n17671 = n17524 & ~n17670;
  assign n17672 = ~n17665 & ~n17671;
  assign n17673 = ~n17662 & n17672;
  assign n17674 = n17659 & n17673;
  assign n17675 = ~n17651 & n17674;
  assign n17676 = n17643 & n17675;
  assign n17679 = n17616 & n17620;
  assign n17677 = n17616 & n17632;
  assign n17678 = ~n17646 & ~n17677;
  assign n17680 = n17679 ^ n17678;
  assign n17681 = n17680 ^ n17679;
  assign n17682 = n17679 ^ n17484;
  assign n17683 = n17682 ^ n17679;
  assign n17684 = ~n17681 & ~n17683;
  assign n17685 = n17684 ^ n17679;
  assign n17686 = ~n17524 & n17685;
  assign n17687 = n17686 ^ n17679;
  assign n17688 = n17676 & ~n17687;
  assign n17689 = n17630 & n17688;
  assign n17690 = n17624 & n17689;
  assign n17691 = n17690 ^ n16595;
  assign n17692 = n17691 ^ x118;
  assign n17693 = ~n17483 & n17692;
  assign n17694 = ~n15365 & n17349;
  assign n17695 = ~n14974 & n17694;
  assign n17696 = n15333 & ~n17695;
  assign n17697 = ~n14974 & n15380;
  assign n17698 = ~n15336 & n17697;
  assign n17699 = n15344 & ~n17698;
  assign n17700 = ~n17696 & ~n17699;
  assign n17701 = ~n15364 & n15369;
  assign n17702 = ~n14978 & n15373;
  assign n17703 = n15340 & ~n17702;
  assign n17704 = ~n15357 & n17351;
  assign n17705 = n15358 & ~n17704;
  assign n17706 = ~n17703 & ~n17705;
  assign n17707 = ~n17701 & n17706;
  assign n17708 = n17700 & n17707;
  assign n17709 = ~n15354 & n17708;
  assign n17710 = n15347 & n17709;
  assign n17711 = n16824 & n17710;
  assign n17712 = n17711 ^ n13779;
  assign n17713 = n17712 ^ x107;
  assign n17714 = n16311 ^ x89;
  assign n17715 = ~n17713 & n17714;
  assign n17716 = n16909 & n17321;
  assign n17717 = n16881 & ~n17314;
  assign n17718 = ~n17716 & ~n17717;
  assign n17719 = n16895 & ~n16904;
  assign n17720 = n16844 & ~n17719;
  assign n17721 = ~n16902 & n17310;
  assign n17722 = n16890 & ~n17721;
  assign n17723 = ~n17720 & ~n17722;
  assign n17724 = n17718 & n17723;
  assign n17725 = ~n16842 & n16912;
  assign n17726 = ~n16888 & ~n16910;
  assign n17727 = ~n17303 & ~n17726;
  assign n17728 = ~n16894 & n16913;
  assign n17729 = ~n17321 & n17728;
  assign n17730 = n16881 & ~n17729;
  assign n17731 = ~n16884 & n17315;
  assign n17732 = n16909 & ~n17731;
  assign n17733 = ~n17730 & ~n17732;
  assign n17734 = ~n17727 & n17733;
  assign n17735 = ~n17725 & n17734;
  assign n17736 = n17724 & n17735;
  assign n17737 = n17308 & n17736;
  assign n17738 = n16886 & n17737;
  assign n17739 = ~n17301 & n17738;
  assign n17740 = ~n16947 & n17739;
  assign n17741 = n17740 ^ n12716;
  assign n17742 = n17741 ^ x113;
  assign n17743 = n16529 & n16651;
  assign n17744 = n17126 & ~n17743;
  assign n17745 = ~n16528 & n16610;
  assign n17746 = n16616 & ~n17136;
  assign n17747 = ~n17745 & ~n17746;
  assign n17748 = n16600 & ~n17141;
  assign n17749 = ~n16617 & ~n16648;
  assign n17750 = ~n16607 & n17749;
  assign n17751 = n16529 & ~n17750;
  assign n17752 = n16645 & ~n16648;
  assign n17753 = ~n16602 & n17752;
  assign n17754 = n16616 & ~n17753;
  assign n17755 = n16625 & ~n16652;
  assign n17756 = n16604 & ~n17755;
  assign n17757 = ~n17754 & ~n17756;
  assign n17758 = ~n17751 & n17757;
  assign n17759 = ~n17748 & n17758;
  assign n17760 = n17747 & n17759;
  assign n17761 = n16642 & n17760;
  assign n17762 = n16637 & n17761;
  assign n17763 = n17128 & n17762;
  assign n17764 = n17744 & n17763;
  assign n17765 = n17764 ^ n13205;
  assign n17766 = n17765 ^ x66;
  assign n17767 = n16525 ^ x96;
  assign n17768 = ~n17766 & ~n17767;
  assign n17769 = n17742 & n17768;
  assign n17770 = n17244 & n17265;
  assign n17771 = n17238 & n17262;
  assign n17772 = ~n17770 & ~n17771;
  assign n17773 = n17233 & n17244;
  assign n17774 = n17234 & ~n17276;
  assign n17775 = ~n17773 & ~n17774;
  assign n17776 = ~n17275 & ~n17284;
  assign n17777 = ~n17271 & n17776;
  assign n17778 = n17165 & ~n17777;
  assign n17779 = n17230 & n17285;
  assign n17780 = n17238 & ~n17779;
  assign n17783 = ~n17229 & n17601;
  assign n17781 = n17230 & ~n17262;
  assign n17782 = ~n17233 & n17781;
  assign n17784 = n17783 ^ n17782;
  assign n17785 = n17783 ^ n17164;
  assign n17786 = n17785 ^ n17783;
  assign n17787 = n17784 & ~n17786;
  assign n17788 = n17787 ^ n17783;
  assign n17789 = ~n17163 & ~n17788;
  assign n17790 = ~n17780 & ~n17789;
  assign n17791 = ~n17778 & n17790;
  assign n17792 = n17775 & n17791;
  assign n17793 = n17772 & n17792;
  assign n17794 = n17259 & n17793;
  assign n17795 = n17251 & n17794;
  assign n17796 = n17589 & n17795;
  assign n17797 = n17586 & n17796;
  assign n17798 = n17797 ^ n13622;
  assign n17799 = n17798 ^ x122;
  assign n17800 = ~n17742 & n17799;
  assign n17801 = n17800 ^ n17799;
  assign n17802 = n17766 & ~n17801;
  assign n17803 = n17802 ^ n17799;
  assign n17804 = n17803 ^ n17767;
  assign n17805 = n17804 ^ n17803;
  assign n17806 = n17799 ^ n17742;
  assign n17807 = n17806 ^ n17803;
  assign n17808 = n17805 & n17807;
  assign n17809 = n17808 ^ n17803;
  assign n17810 = ~n17769 & n17809;
  assign n17811 = n17715 & n17810;
  assign n17812 = n17713 & ~n17714;
  assign n17813 = ~n17767 & ~n17803;
  assign n17815 = n17766 ^ n17742;
  assign n17814 = ~n17766 & n17767;
  assign n17816 = n17815 ^ n17814;
  assign n17817 = n17815 ^ n17799;
  assign n17818 = n17817 ^ n17815;
  assign n17819 = ~n17816 & n17818;
  assign n17820 = n17819 ^ n17815;
  assign n17821 = ~n17813 & n17820;
  assign n17822 = n17812 & ~n17821;
  assign n17823 = ~n17811 & ~n17822;
  assign n17824 = n17713 & n17714;
  assign n17825 = n17767 ^ n17766;
  assign n17826 = n17825 ^ n17767;
  assign n17827 = n17815 ^ n17767;
  assign n17828 = n17827 ^ n17767;
  assign n17829 = n17828 ^ n17767;
  assign n17830 = ~n17826 & n17829;
  assign n17831 = n17830 ^ n17767;
  assign n17832 = n17799 & n17831;
  assign n17833 = n17832 ^ n17827;
  assign n17834 = n17824 & ~n17833;
  assign n17835 = ~n17713 & ~n17714;
  assign n17836 = n17825 ^ n17799;
  assign n17837 = n17836 ^ n17767;
  assign n17838 = n17806 ^ n17742;
  assign n17839 = n17767 ^ n17742;
  assign n17840 = n17839 ^ n17742;
  assign n17841 = n17838 & n17840;
  assign n17842 = n17841 ^ n17742;
  assign n17843 = n17837 & ~n17842;
  assign n17844 = n17843 ^ n17825;
  assign n17845 = n17835 & ~n17844;
  assign n17846 = ~n17834 & ~n17845;
  assign n17847 = n17823 & n17846;
  assign n17848 = n17847 ^ n15433;
  assign n17849 = n17848 ^ x116;
  assign n17850 = n17613 ^ x112;
  assign n17851 = n16974 ^ x105;
  assign n17852 = n17850 & n17851;
  assign n17853 = n16654 & n17136;
  assign n17854 = ~n16644 & n17853;
  assign n17855 = n16604 & ~n17854;
  assign n17856 = ~n16624 & n16645;
  assign n17857 = n17141 & n17856;
  assign n17858 = ~n16628 & n17857;
  assign n17859 = n16616 & ~n17858;
  assign n17860 = ~n17855 & ~n17859;
  assign n17861 = ~n16607 & ~n16619;
  assign n17862 = n16654 & n17861;
  assign n17863 = ~n16630 & n17862;
  assign n17864 = n16600 & ~n17863;
  assign n17865 = ~n16610 & n17131;
  assign n17866 = n17865 ^ n16620;
  assign n17867 = n16620 ^ n16529;
  assign n17868 = n16620 & n17867;
  assign n17869 = n17868 ^ n16620;
  assign n17870 = n17866 & n17869;
  assign n17871 = n17870 ^ n17868;
  assign n17872 = n17871 ^ n16620;
  assign n17873 = n17872 ^ n16529;
  assign n17874 = ~n17864 & n17873;
  assign n17875 = n17874 ^ n17864;
  assign n17876 = n17860 & ~n17875;
  assign n17877 = n16632 & n17876;
  assign n17878 = n17744 & n17877;
  assign n17879 = n16614 & n17878;
  assign n17880 = n17879 ^ n15526;
  assign n17881 = n17880 ^ x90;
  assign n17882 = n16445 & ~n16513;
  assign n17883 = ~n16451 & ~n16511;
  assign n17884 = ~n16443 & n17883;
  assign n17885 = ~n16458 & n17884;
  assign n17886 = n16478 & ~n17885;
  assign n17887 = ~n17882 & ~n17886;
  assign n17888 = n16318 & ~n16786;
  assign n17889 = n16513 & n16794;
  assign n17890 = ~n16462 & n17889;
  assign n17891 = n16352 & ~n17890;
  assign n17892 = ~n16455 & n16509;
  assign n17893 = ~n16468 & ~n16508;
  assign n17894 = ~n16445 & n17893;
  assign n17895 = ~n17892 & ~n17894;
  assign n17896 = ~n16448 & ~n17895;
  assign n17897 = ~n16485 & n17896;
  assign n17898 = ~n16502 & ~n17897;
  assign n17899 = ~n17891 & ~n17898;
  assign n17900 = ~n17888 & n17899;
  assign n17901 = n17887 & n17900;
  assign n17902 = n16477 & n17901;
  assign n17903 = n16781 & n17902;
  assign n17904 = ~n16465 & n17903;
  assign n17905 = n17904 ^ n15500;
  assign n17906 = n17905 ^ x64;
  assign n17907 = n17881 & n17906;
  assign n17908 = n16775 ^ x81;
  assign n17909 = n17523 ^ x115;
  assign n17910 = ~n17908 & n17909;
  assign n17911 = n17907 & n17910;
  assign n17912 = n17852 & n17911;
  assign n17913 = n17850 & ~n17851;
  assign n17914 = n17908 & ~n17909;
  assign n17915 = n17907 & n17914;
  assign n17916 = n17913 & n17915;
  assign n17917 = ~n17912 & ~n17916;
  assign n17918 = n17908 & n17909;
  assign n17919 = n17907 & n17918;
  assign n17920 = ~n17881 & n17906;
  assign n17921 = ~n17908 & ~n17909;
  assign n17922 = n17920 & n17921;
  assign n17923 = ~n17919 & ~n17922;
  assign n17924 = n17852 & ~n17923;
  assign n17925 = ~n17850 & ~n17851;
  assign n17926 = ~n17881 & ~n17906;
  assign n17927 = n17910 & n17926;
  assign n17928 = n17925 & n17927;
  assign n17929 = ~n17850 & n17851;
  assign n17930 = n17881 & ~n17906;
  assign n17931 = n17910 & n17930;
  assign n17932 = ~n17922 & ~n17931;
  assign n17933 = n17929 & ~n17932;
  assign n17934 = ~n17928 & ~n17933;
  assign n17935 = n17910 & n17920;
  assign n17936 = n17929 & n17935;
  assign n17937 = n17922 & n17925;
  assign n17938 = ~n17936 & ~n17937;
  assign n17939 = n17918 & n17930;
  assign n17940 = n17914 & n17926;
  assign n17941 = ~n17939 & ~n17940;
  assign n17942 = n17852 & ~n17941;
  assign n17943 = n17925 & n17935;
  assign n17944 = n17921 & n17926;
  assign n17945 = n17852 & n17944;
  assign n17946 = ~n17943 & ~n17945;
  assign n17947 = ~n17915 & ~n17927;
  assign n17948 = n17851 & ~n17947;
  assign n17949 = n17918 & n17920;
  assign n17950 = n17918 & n17926;
  assign n17951 = n17914 & n17920;
  assign n17952 = ~n17950 & ~n17951;
  assign n17953 = ~n17949 & n17952;
  assign n17954 = ~n17935 & n17953;
  assign n17955 = n17913 & ~n17954;
  assign n17956 = ~n17948 & ~n17955;
  assign n17957 = n17907 & n17921;
  assign n17958 = n17925 & n17957;
  assign n17959 = ~n17940 & ~n17949;
  assign n17960 = ~n17919 & n17959;
  assign n17961 = n17929 & ~n17960;
  assign n17963 = n17914 & n17930;
  assign n17966 = n17921 & n17930;
  assign n17967 = ~n17911 & ~n17966;
  assign n17968 = ~n17963 & n17967;
  assign n17962 = ~n17939 & ~n17951;
  assign n17964 = ~n17919 & ~n17963;
  assign n17965 = n17962 & n17964;
  assign n17969 = n17968 ^ n17965;
  assign n17970 = n17968 ^ n17850;
  assign n17971 = n17970 ^ n17968;
  assign n17972 = n17969 & ~n17971;
  assign n17973 = n17972 ^ n17968;
  assign n17974 = ~n17851 & ~n17973;
  assign n17975 = ~n17961 & ~n17974;
  assign n17976 = ~n17958 & n17975;
  assign n17977 = n17956 & n17976;
  assign n17978 = n17946 & n17977;
  assign n17979 = ~n17942 & n17978;
  assign n17980 = n17938 & n17979;
  assign n17981 = n17934 & n17980;
  assign n17982 = ~n17924 & n17981;
  assign n17983 = n17917 & n17982;
  assign n17984 = n17983 ^ n15940;
  assign n17985 = n17984 ^ x76;
  assign n17986 = ~n17849 & ~n17985;
  assign n17987 = n17693 & n17986;
  assign n17988 = n17088 & n17987;
  assign n17989 = n17849 & n17985;
  assign n17990 = n17483 & ~n17692;
  assign n17991 = n17989 & n17990;
  assign n17992 = n17991 ^ n16758;
  assign n17993 = n17992 ^ n17991;
  assign n17994 = n17849 & ~n17985;
  assign n17995 = n17990 & n17994;
  assign n17996 = n17995 ^ n17991;
  assign n17997 = n17993 & n17996;
  assign n17998 = n17997 ^ n17991;
  assign n17999 = n17087 & n17998;
  assign n18000 = ~n17988 & ~n17999;
  assign n18001 = ~n16758 & n17087;
  assign n18002 = n17693 & n17994;
  assign n18003 = n17483 & n17692;
  assign n18004 = ~n17849 & n17985;
  assign n18005 = n18003 & n18004;
  assign n18006 = ~n17483 & ~n17692;
  assign n18007 = n17989 & n18006;
  assign n18008 = ~n18005 & ~n18007;
  assign n18009 = ~n18002 & n18008;
  assign n18010 = n18001 & ~n18009;
  assign n18011 = ~n16758 & ~n17087;
  assign n18012 = n17990 & n18004;
  assign n18013 = n17693 & n17989;
  assign n18014 = n18004 & n18006;
  assign n18015 = ~n18013 & ~n18014;
  assign n18016 = ~n18012 & n18015;
  assign n18017 = n18011 & ~n18016;
  assign n18018 = ~n18010 & ~n18017;
  assign n18019 = n16758 & ~n17087;
  assign n18020 = n17693 & n18004;
  assign n18021 = ~n18007 & ~n18020;
  assign n18022 = n18019 & ~n18021;
  assign n18023 = n17986 & n17990;
  assign n18024 = n17994 & n18006;
  assign n18025 = ~n18023 & ~n18024;
  assign n18026 = n17088 & ~n18025;
  assign n18027 = n17986 & n18006;
  assign n18028 = ~n17995 & ~n18027;
  assign n18029 = n17994 & n18003;
  assign n18030 = ~n18023 & ~n18029;
  assign n18031 = n18028 & n18030;
  assign n18032 = n18001 & ~n18031;
  assign n18033 = n17989 & n18003;
  assign n18034 = ~n18014 & n18021;
  assign n18035 = ~n18033 & n18034;
  assign n18036 = n17088 & ~n18035;
  assign n18037 = ~n18032 & ~n18036;
  assign n18038 = n17986 & n18003;
  assign n18039 = ~n18024 & ~n18038;
  assign n18040 = ~n18002 & ~n18029;
  assign n18041 = n18039 & n18040;
  assign n18042 = n18011 & ~n18041;
  assign n18043 = ~n17987 & ~n18029;
  assign n18044 = ~n17995 & n18043;
  assign n18045 = ~n18012 & n18044;
  assign n18046 = n18019 & ~n18045;
  assign n18047 = ~n18042 & ~n18046;
  assign n18048 = n18037 & n18047;
  assign n18049 = ~n18026 & n18048;
  assign n18050 = ~n18022 & n18049;
  assign n18051 = n18018 & n18050;
  assign n18052 = ~n18005 & ~n18013;
  assign n18053 = n18052 ^ n17991;
  assign n18054 = n17993 & ~n18053;
  assign n18055 = n18054 ^ n17991;
  assign n18056 = ~n17087 & n18055;
  assign n18057 = n18051 & ~n18056;
  assign n18058 = n18000 & n18057;
  assign n18059 = n18058 ^ n16678;
  assign n18060 = n17742 & ~n17799;
  assign n18061 = n17814 & n18060;
  assign n18062 = n17767 & n17800;
  assign n18063 = n18060 ^ n17766;
  assign n18064 = n18063 ^ n17766;
  assign n18065 = n17768 ^ n17766;
  assign n18066 = ~n18064 & n18065;
  assign n18067 = n18066 ^ n17766;
  assign n18068 = ~n18062 & ~n18067;
  assign n18069 = n17835 & ~n18068;
  assign n18070 = ~n17742 & ~n17799;
  assign n18071 = n17767 & n18070;
  assign n18072 = n17742 & n17799;
  assign n18073 = ~n17767 & n18072;
  assign n18074 = n17766 & n17767;
  assign n18075 = ~n17768 & ~n18074;
  assign n18076 = ~n17742 & n18075;
  assign n18077 = ~n18073 & ~n18076;
  assign n18078 = ~n18071 & n18077;
  assign n18079 = n17715 & ~n18078;
  assign n18080 = ~n18069 & ~n18079;
  assign n18081 = n17800 & n18074;
  assign n18082 = ~n17766 & ~n17806;
  assign n18083 = ~n17799 & n18075;
  assign n18084 = ~n18082 & ~n18083;
  assign n18085 = ~n18081 & n18084;
  assign n18086 = n17824 & ~n18085;
  assign n18087 = ~n17799 & n18074;
  assign n18088 = n17800 & n18075;
  assign n18089 = ~n18087 & ~n18088;
  assign n18090 = n17742 & n18089;
  assign n18091 = n18089 ^ n18075;
  assign n18092 = ~n17766 & ~n17799;
  assign n18093 = n18092 ^ n18090;
  assign n18094 = n18091 & n18093;
  assign n18095 = n18094 ^ n18092;
  assign n18096 = n18090 & n18095;
  assign n18097 = n18096 ^ n18089;
  assign n18098 = n17812 & ~n18097;
  assign n18099 = ~n18086 & ~n18098;
  assign n18100 = n18080 & n18099;
  assign n18101 = ~n18061 & n18100;
  assign n18102 = n18101 ^ n14005;
  assign n18103 = n18102 ^ x110;
  assign n18104 = n17644 & n17655;
  assign n18105 = n17619 & ~n17649;
  assign n18106 = ~n18104 & ~n18105;
  assign n18107 = ~n17626 & ~n17679;
  assign n18108 = n17628 & ~n18107;
  assign n18109 = ~n17617 & ~n17647;
  assign n18110 = n17644 & ~n18109;
  assign n18111 = n17619 & ~n17656;
  assign n18112 = ~n18110 & ~n18111;
  assign n18113 = ~n17633 & ~n17679;
  assign n18114 = n17525 & ~n18113;
  assign n18115 = n17628 & ~n17663;
  assign n18116 = ~n18114 & ~n18115;
  assign n18118 = ~n17637 & ~n17660;
  assign n18117 = ~n17622 & ~n17638;
  assign n18119 = n18118 ^ n18117;
  assign n18120 = n18119 ^ n18118;
  assign n18121 = n18118 ^ n17524;
  assign n18122 = n18121 ^ n18118;
  assign n18123 = ~n18120 & n18122;
  assign n18124 = n18123 ^ n18118;
  assign n18125 = n17631 & ~n18124;
  assign n18126 = n18125 ^ n18118;
  assign n18127 = n18116 & n18126;
  assign n18128 = n17678 ^ n17484;
  assign n18129 = n18128 ^ n17678;
  assign n18130 = n17678 ^ n17668;
  assign n18131 = n18130 ^ n17678;
  assign n18132 = n18129 & ~n18131;
  assign n18133 = n18132 ^ n17678;
  assign n18134 = ~n17524 & ~n18133;
  assign n18135 = n18134 ^ n17678;
  assign n18136 = n18127 & n18135;
  assign n18137 = n18112 & n18136;
  assign n18138 = ~n18108 & n18137;
  assign n18139 = n18106 & n18138;
  assign n18140 = n17659 & n18139;
  assign n18141 = n17624 & n18140;
  assign n18142 = n18141 ^ n16238;
  assign n18143 = n18142 ^ x124;
  assign n18144 = n18103 & ~n18143;
  assign n18145 = n16080 & n17115;
  assign n18146 = n15942 & ~n17103;
  assign n18147 = ~n18145 & ~n18146;
  assign n18148 = n16085 & n17093;
  assign n18149 = n16106 & ~n18148;
  assign n18150 = ~n16078 & n17111;
  assign n18151 = n16088 & ~n18150;
  assign n18152 = ~n18149 & ~n18151;
  assign n18153 = n18147 & n18152;
  assign n18154 = n18153 ^ n14987;
  assign n18155 = n18154 ^ x70;
  assign n18156 = n17165 & n17252;
  assign n18157 = ~n17248 & ~n17256;
  assign n18158 = ~n17270 & n18157;
  assign n18159 = n17238 & ~n18158;
  assign n18160 = ~n18156 & ~n18159;
  assign n18161 = n17234 & n17254;
  assign n18162 = ~n17243 & n17777;
  assign n18163 = ~n17165 & n18162;
  assign n18164 = n17272 & n17285;
  assign n18165 = ~n17234 & n18164;
  assign n18166 = ~n18163 & ~n18165;
  assign n18167 = n18166 ^ n17164;
  assign n18168 = n18167 ^ n18166;
  assign n18169 = ~n17229 & n17776;
  assign n18170 = n18169 ^ n18166;
  assign n18171 = n18170 ^ n18166;
  assign n18172 = n18168 & ~n18171;
  assign n18173 = n18172 ^ n18166;
  assign n18174 = n17163 & n18173;
  assign n18175 = n18174 ^ n18166;
  assign n18176 = ~n18161 & ~n18175;
  assign n18177 = n18160 & n18176;
  assign n18178 = n17268 & n18177;
  assign n18179 = ~n17250 & n18178;
  assign n18180 = n17593 & n18179;
  assign n18181 = n17772 & n18180;
  assign n18182 = n17241 & n18181;
  assign n18183 = n18182 ^ n15039;
  assign n18184 = n18183 ^ x91;
  assign n18185 = ~n18155 & n18184;
  assign n18186 = n16806 ^ x110;
  assign n18187 = n17160 ^ x116;
  assign n18188 = ~n18186 & ~n18187;
  assign n18189 = n18185 & n18188;
  assign n18190 = n17338 ^ x93;
  assign n18191 = n17014 ^ x84;
  assign n18192 = ~n18190 & n18191;
  assign n18193 = n18189 & n18192;
  assign n18194 = ~n18186 & n18187;
  assign n18195 = ~n18155 & ~n18184;
  assign n18196 = n18194 & n18195;
  assign n18197 = n18192 & n18196;
  assign n18198 = n18186 & n18187;
  assign n18199 = n18155 & ~n18184;
  assign n18200 = n18198 & n18199;
  assign n18201 = n18185 & n18198;
  assign n18202 = ~n18200 & ~n18201;
  assign n18203 = n18192 & ~n18202;
  assign n18204 = n18186 & ~n18187;
  assign n18205 = n18195 & n18204;
  assign n18206 = n18190 & ~n18191;
  assign n18207 = n18205 & n18206;
  assign n18208 = n18155 & n18184;
  assign n18209 = n18204 & n18208;
  assign n18210 = n18188 & n18195;
  assign n18211 = ~n18209 & ~n18210;
  assign n18212 = n18192 & ~n18211;
  assign n18213 = ~n18190 & ~n18191;
  assign n18214 = n18185 & n18204;
  assign n18215 = n18194 & n18208;
  assign n18216 = ~n18200 & ~n18215;
  assign n18217 = n18199 & n18204;
  assign n18218 = n18195 & n18198;
  assign n18219 = ~n18189 & ~n18218;
  assign n18220 = ~n18217 & n18219;
  assign n18221 = n18211 & n18220;
  assign n18222 = n18216 & n18221;
  assign n18223 = ~n18214 & n18222;
  assign n18224 = n18213 & n18223;
  assign n18225 = ~n18212 & ~n18224;
  assign n18226 = n18188 & n18199;
  assign n18227 = ~n18196 & ~n18201;
  assign n18228 = n18219 & n18227;
  assign n18229 = ~n18226 & n18228;
  assign n18230 = n18206 & ~n18229;
  assign n18231 = n18191 ^ n18190;
  assign n18239 = ~n18215 & ~n18217;
  assign n18232 = n18184 ^ n18155;
  assign n18233 = n18186 ^ n18184;
  assign n18234 = n18233 ^ n18187;
  assign n18235 = n18234 ^ n18184;
  assign n18236 = ~n18232 & n18235;
  assign n18237 = ~n18187 & n18236;
  assign n18238 = n18237 ^ n18234;
  assign n18240 = n18239 ^ n18238;
  assign n18241 = n18240 ^ n18239;
  assign n18242 = n18239 ^ n18191;
  assign n18243 = n18242 ^ n18239;
  assign n18244 = ~n18241 & n18243;
  assign n18245 = n18244 ^ n18239;
  assign n18246 = ~n18231 & ~n18245;
  assign n18247 = n18246 ^ n18239;
  assign n18248 = ~n18230 & n18247;
  assign n18249 = n18225 & n18248;
  assign n18250 = ~n18207 & n18249;
  assign n18251 = ~n18203 & n18250;
  assign n18252 = ~n18197 & n18251;
  assign n18253 = ~n18193 & n18252;
  assign n18254 = n18253 ^ n15142;
  assign n18255 = n18254 ^ x67;
  assign n18256 = n17913 & n17935;
  assign n18257 = n17915 & n17929;
  assign n18258 = ~n18256 & ~n18257;
  assign n18259 = n17915 & n17925;
  assign n18260 = n17852 & n17963;
  assign n18261 = ~n18259 & ~n18260;
  assign n18262 = ~n17949 & n17964;
  assign n18263 = n17925 & ~n18262;
  assign n18264 = n17932 & ~n17944;
  assign n18265 = n17913 & ~n18264;
  assign n18266 = ~n18263 & ~n18265;
  assign n18267 = n17852 & n17949;
  assign n18268 = ~n17940 & n17952;
  assign n18269 = n17929 & ~n18268;
  assign n18270 = ~n17931 & ~n17957;
  assign n18271 = ~n17963 & n18270;
  assign n18272 = n17929 & ~n18271;
  assign n18273 = ~n17919 & n17952;
  assign n18274 = n17913 & ~n18273;
  assign n18275 = ~n18272 & ~n18274;
  assign n18276 = n17906 ^ n17881;
  assign n18277 = n17906 & ~n17909;
  assign n18278 = ~n18276 & n18277;
  assign n18279 = n18278 ^ n18276;
  assign n18280 = ~n17908 & ~n18279;
  assign n18281 = n17925 & n18280;
  assign n18282 = ~n17922 & ~n17966;
  assign n18283 = ~n17935 & n18282;
  assign n18284 = n17852 & ~n18283;
  assign n18285 = ~n18281 & ~n18284;
  assign n18286 = n18275 & n18285;
  assign n18287 = n17938 & n18286;
  assign n18288 = n17917 & n18287;
  assign n18289 = ~n18269 & n18288;
  assign n18290 = ~n18267 & n18289;
  assign n18291 = n18266 & n18290;
  assign n18292 = n18261 & n18291;
  assign n18293 = n18258 & n18292;
  assign n18294 = ~n17942 & n18293;
  assign n18295 = n18294 ^ n17192;
  assign n18296 = n18295 ^ x78;
  assign n18297 = ~n18255 & n18296;
  assign n18298 = n16688 & n16721;
  assign n18299 = ~n16314 & ~n16689;
  assign n18300 = n16685 & ~n18299;
  assign n18301 = ~n18298 & ~n18300;
  assign n18302 = ~n16709 & ~n16732;
  assign n18303 = n16680 & ~n18302;
  assign n18304 = ~n16316 & ~n16720;
  assign n18305 = n16703 & ~n18304;
  assign n18306 = ~n18303 & ~n18305;
  assign n18307 = ~n16702 & ~n16709;
  assign n18308 = n16721 & ~n18307;
  assign n18309 = ~n16684 & n18299;
  assign n18310 = n16703 & ~n18309;
  assign n18311 = ~n18308 & ~n18310;
  assign n18312 = ~n16691 & n16725;
  assign n18313 = n16680 & ~n18312;
  assign n18314 = ~n16723 & n16733;
  assign n18315 = n16685 & ~n18314;
  assign n18316 = ~n18313 & ~n18315;
  assign n18317 = n18311 & n18316;
  assign n18318 = ~n16706 & ~n18304;
  assign n18319 = ~n16685 & ~n16706;
  assign n18320 = n16736 & ~n18319;
  assign n18321 = ~n18318 & ~n18320;
  assign n18322 = n18317 & n18321;
  assign n18323 = n16708 & n18322;
  assign n18324 = n18306 & n18323;
  assign n18325 = n18301 & n18324;
  assign n18326 = ~n16737 & n18325;
  assign n18327 = ~n16689 & n18326;
  assign n18328 = n18327 ^ n17222;
  assign n18329 = n18328 ^ x92;
  assign n18330 = n17420 & ~n17436;
  assign n18331 = ~n17453 & n17471;
  assign n18332 = ~n18330 & ~n18331;
  assign n18333 = n17422 & n17457;
  assign n18334 = n17426 & n17472;
  assign n18335 = ~n18333 & ~n18334;
  assign n18336 = n17431 & ~n17436;
  assign n18337 = n17422 & n17472;
  assign n18338 = ~n18336 & ~n18337;
  assign n18339 = n17429 & n17438;
  assign n18340 = ~n17446 & ~n18339;
  assign n18341 = n17471 & ~n18340;
  assign n18342 = n17340 & n17430;
  assign n18343 = n17473 & ~n18342;
  assign n18344 = ~n17457 & n18343;
  assign n18345 = n17162 & ~n18344;
  assign n18346 = ~n18341 & ~n18345;
  assign n18347 = ~n17445 & n17453;
  assign n18348 = n17426 & ~n18347;
  assign n18349 = n17161 ^ n17121;
  assign n18352 = ~n17424 & ~n18342;
  assign n18353 = ~n17451 & n18352;
  assign n18354 = ~n17456 & n18353;
  assign n18350 = ~n17451 & ~n18339;
  assign n18351 = ~n17428 & n18350;
  assign n18355 = n18354 ^ n18351;
  assign n18356 = n18354 ^ n17161;
  assign n18357 = n18356 ^ n18354;
  assign n18358 = n18355 & ~n18357;
  assign n18359 = n18358 ^ n18354;
  assign n18360 = n18349 & ~n18359;
  assign n18361 = ~n18348 & ~n18360;
  assign n18362 = n18346 & n18361;
  assign n18363 = n18338 & n18362;
  assign n18364 = n18335 & n18363;
  assign n18365 = n18332 & n18364;
  assign n18366 = n17450 & n18365;
  assign n18367 = n18366 ^ n16177;
  assign n18368 = n18367 ^ x93;
  assign n18369 = n18329 & ~n18368;
  assign n18370 = n18297 & n18369;
  assign n18371 = ~n18329 & ~n18368;
  assign n18372 = n18255 & ~n18296;
  assign n18373 = n18371 & n18372;
  assign n18374 = ~n18370 & ~n18373;
  assign n18375 = n18144 & ~n18374;
  assign n18376 = n18103 & n18143;
  assign n18377 = n18297 & n18371;
  assign n18378 = n18255 & n18296;
  assign n18379 = n18369 & n18378;
  assign n18380 = ~n18377 & ~n18379;
  assign n18381 = n18376 & ~n18380;
  assign n18382 = ~n18375 & ~n18381;
  assign n18383 = ~n18103 & ~n18143;
  assign n18384 = ~n18329 & n18368;
  assign n18385 = n18297 & n18384;
  assign n18386 = n18383 & n18385;
  assign n18387 = n18329 & n18368;
  assign n18388 = n18378 & n18387;
  assign n18389 = n18383 & n18388;
  assign n18390 = n18296 ^ n18255;
  assign n18391 = n18387 & n18390;
  assign n18392 = n18144 & n18391;
  assign n18393 = ~n18389 & ~n18392;
  assign n18394 = ~n18386 & n18393;
  assign n18395 = ~n18103 & n18143;
  assign n18396 = n18385 & n18395;
  assign n18397 = n18371 & n18378;
  assign n18398 = ~n18370 & ~n18397;
  assign n18399 = ~n18373 & n18398;
  assign n18400 = n18383 & ~n18399;
  assign n18401 = n18378 & n18384;
  assign n18402 = n18395 & n18401;
  assign n18403 = ~n18255 & ~n18296;
  assign n18404 = n18387 & n18403;
  assign n18405 = n18372 & n18384;
  assign n18406 = ~n18404 & ~n18405;
  assign n18407 = n18376 & ~n18406;
  assign n18408 = ~n18402 & ~n18407;
  assign n18409 = n18144 & n18388;
  assign n18410 = n18371 & n18403;
  assign n18411 = n18376 & n18410;
  assign n18412 = ~n18409 & ~n18411;
  assign n18413 = n18144 & n18385;
  assign n18414 = n18383 & ~n18406;
  assign n18415 = ~n18413 & ~n18414;
  assign n18416 = ~n18103 & n18410;
  assign n18417 = n18369 & n18403;
  assign n18418 = n18143 & n18417;
  assign n18419 = ~n18416 & ~n18418;
  assign n18420 = ~n18370 & ~n18401;
  assign n18421 = n18376 & ~n18420;
  assign n18422 = n18384 & n18403;
  assign n18423 = n18372 & n18387;
  assign n18424 = ~n18422 & ~n18423;
  assign n18425 = ~n18379 & n18424;
  assign n18426 = n18395 & ~n18425;
  assign n18427 = ~n18421 & ~n18426;
  assign n18428 = n18419 & n18427;
  assign n18429 = n18415 & n18428;
  assign n18430 = n18369 & n18372;
  assign n18431 = n18430 ^ n18144;
  assign n18432 = n18422 ^ n18395;
  assign n18433 = n18430 ^ n18395;
  assign n18434 = n18433 ^ n18395;
  assign n18435 = ~n18432 & ~n18434;
  assign n18436 = n18435 ^ n18395;
  assign n18437 = n18431 & n18436;
  assign n18438 = n18437 ^ n18144;
  assign n18439 = n18429 & ~n18438;
  assign n18440 = n18412 & n18439;
  assign n18441 = n18408 & n18440;
  assign n18442 = ~n18400 & n18441;
  assign n18443 = ~n18396 & n18442;
  assign n18444 = n18394 & n18443;
  assign n18445 = n18382 & n18444;
  assign n18446 = n18445 ^ n17298;
  assign n18447 = n18446 ^ x75;
  assign n18448 = n17715 & n18085;
  assign n18449 = n17835 & n18097;
  assign n18450 = ~n18448 & ~n18449;
  assign n18451 = ~n18061 & n18068;
  assign n18452 = n18451 ^ n17714;
  assign n18453 = n18452 ^ n18451;
  assign n18454 = ~n17799 & n17814;
  assign n18455 = n17766 & n18070;
  assign n18456 = ~n18454 & ~n18455;
  assign n18457 = n18077 & n18456;
  assign n18458 = n18457 ^ n18451;
  assign n18459 = n18453 & n18458;
  assign n18460 = n18459 ^ n18451;
  assign n18461 = n17713 & ~n18460;
  assign n18462 = n18450 & ~n18461;
  assign n18463 = n18462 ^ n16875;
  assign n18464 = n18463 ^ x105;
  assign n18465 = ~n17940 & ~n17957;
  assign n18466 = ~n17927 & n18465;
  assign n18467 = ~n17935 & n18466;
  assign n18468 = n17852 & ~n18467;
  assign n18469 = ~n17950 & n17967;
  assign n18470 = ~n17949 & n18469;
  assign n18471 = n17929 & ~n18470;
  assign n18472 = n17959 & n18271;
  assign n18473 = n17925 & ~n18472;
  assign n18475 = ~n17906 & ~n17908;
  assign n18474 = n17881 & n17909;
  assign n18476 = n18475 ^ n18474;
  assign n18477 = n17913 & n18476;
  assign n18478 = ~n18473 & ~n18477;
  assign n18479 = ~n18471 & n18478;
  assign n18480 = ~n18468 & n18479;
  assign n18481 = n18261 & n18480;
  assign n18482 = n18258 & n18481;
  assign n18483 = n17934 & n18482;
  assign n18484 = ~n17951 & n18483;
  assign n18485 = ~n17924 & n18484;
  assign n18486 = n18485 ^ n16350;
  assign n18487 = n18486 ^ x114;
  assign n18488 = n18464 & n18487;
  assign n18489 = n18192 & n18205;
  assign n18490 = n18213 & n18215;
  assign n18491 = ~n18489 & ~n18490;
  assign n18492 = n18185 & n18194;
  assign n18493 = ~n18218 & ~n18492;
  assign n18494 = n18190 & n18191;
  assign n18495 = ~n18493 & n18494;
  assign n18496 = n18188 & n18208;
  assign n18497 = n18213 & n18496;
  assign n18498 = ~n18495 & ~n18497;
  assign n18499 = ~n18214 & ~n18496;
  assign n18500 = n18192 & ~n18499;
  assign n18501 = n18206 & n18223;
  assign n18502 = n18194 & n18199;
  assign n18503 = ~n18217 & ~n18502;
  assign n18504 = n18211 & n18503;
  assign n18505 = ~n18215 & n18504;
  assign n18506 = ~n18189 & n18505;
  assign n18507 = n18494 & ~n18506;
  assign n18508 = ~n18501 & ~n18507;
  assign n18509 = ~n18200 & ~n18492;
  assign n18510 = ~n18217 & n18509;
  assign n18511 = n18192 & ~n18510;
  assign n18512 = ~n18201 & ~n18502;
  assign n18513 = n18220 & n18512;
  assign n18514 = ~n18205 & n18513;
  assign n18515 = n18213 & ~n18514;
  assign n18516 = ~n18511 & ~n18515;
  assign n18517 = n18508 & n18516;
  assign n18518 = ~n18500 & n18517;
  assign n18519 = n18498 & n18518;
  assign n18520 = n18491 & n18519;
  assign n18521 = ~n18197 & n18520;
  assign n18522 = ~n18193 & n18521;
  assign n18523 = n18522 ^ n15899;
  assign n18524 = n18523 ^ x123;
  assign n18525 = ~n17436 & n17456;
  assign n18526 = n17299 & n17438;
  assign n18527 = n17422 & n18526;
  assign n18528 = ~n18525 & ~n18527;
  assign n18529 = ~n17432 & n17436;
  assign n18530 = ~n17437 & n18350;
  assign n18531 = n17426 & ~n18530;
  assign n18532 = ~n18529 & ~n18531;
  assign n18533 = n17440 & n18352;
  assign n18534 = n17471 & ~n18533;
  assign n18535 = ~n17446 & n17474;
  assign n18536 = n17162 & ~n18535;
  assign n18537 = ~n18534 & ~n18536;
  assign n18538 = n18532 & n18537;
  assign n18539 = n18528 & n18538;
  assign n18540 = n18335 & n18539;
  assign n18541 = n18332 & n18540;
  assign n18542 = n17449 & n18541;
  assign n18543 = n17435 & n18542;
  assign n18544 = n18543 ^ n16862;
  assign n18545 = n18544 ^ x104;
  assign n18546 = n18524 & ~n18545;
  assign n18547 = n18488 & n18546;
  assign n18548 = ~n18524 & ~n18545;
  assign n18549 = n18488 & n18548;
  assign n18550 = ~n18547 & ~n18549;
  assign n18551 = n17525 & n17677;
  assign n18552 = n17630 & ~n18551;
  assign n18553 = n17525 & ~n17656;
  assign n18554 = n17628 & n17667;
  assign n18555 = ~n17622 & ~n17646;
  assign n18556 = ~n17631 & ~n18555;
  assign n18557 = ~n18554 & ~n18556;
  assign n18558 = ~n18553 & n18557;
  assign n18559 = ~n17637 & n17663;
  assign n18560 = n17668 & n18559;
  assign n18561 = n17644 & ~n18560;
  assign n18562 = n17619 & n17661;
  assign n18563 = n17661 ^ n17632;
  assign n18564 = n18562 ^ n17621;
  assign n18565 = n18563 & n18564;
  assign n18566 = n18565 ^ n17621;
  assign n18567 = n18562 & n18566;
  assign n18568 = n18567 ^ n17619;
  assign n18569 = ~n18561 & ~n18568;
  assign n18570 = n18558 & n18569;
  assign n18571 = ~n18110 & n18570;
  assign n18572 = n18552 & n18571;
  assign n18573 = n17658 & n18572;
  assign n18574 = ~n18108 & n18573;
  assign n18575 = n18106 & n18574;
  assign n18576 = n17624 & n18575;
  assign n18577 = n18576 ^ n16005;
  assign n18578 = n18577 ^ x72;
  assign n18579 = n17298 ^ x68;
  assign n18580 = n17741 ^ x117;
  assign n18581 = ~n18579 & n18580;
  assign n18582 = n17120 ^ x69;
  assign n18583 = n15812 & n16978;
  assign n18584 = n15471 & n15848;
  assign n18585 = ~n18583 & ~n18584;
  assign n18586 = ~n15818 & ~n16983;
  assign n18587 = ~n15434 & n15841;
  assign n18588 = n15816 & n15825;
  assign n18589 = n15847 & n18588;
  assign n18590 = n15840 & ~n18589;
  assign n18591 = n15843 & n16983;
  assign n18592 = n16978 & ~n18591;
  assign n18593 = ~n18590 & ~n18592;
  assign n18594 = n16979 ^ n15830;
  assign n18595 = n16979 ^ n15471;
  assign n18596 = n18595 ^ n15471;
  assign n18597 = n15850 & n16996;
  assign n18598 = ~n15820 & n18597;
  assign n18599 = n18598 ^ n15471;
  assign n18600 = n18596 & n18599;
  assign n18601 = n18600 ^ n15471;
  assign n18602 = ~n18594 & n18601;
  assign n18603 = n18602 ^ n15830;
  assign n18604 = n18593 & ~n18603;
  assign n18605 = ~n15817 & n18604;
  assign n18606 = ~n18587 & n18605;
  assign n18607 = ~n18586 & n18606;
  assign n18608 = n18585 & n18607;
  assign n18609 = n16981 & n18608;
  assign n18610 = n18609 ^ n14604;
  assign n18611 = n18610 ^ x86;
  assign n18612 = n18582 & n18611;
  assign n18613 = n17712 ^ x92;
  assign n18614 = n16445 & ~n16783;
  assign n18615 = n16455 & ~n16794;
  assign n18616 = ~n18614 & ~n18615;
  assign n18617 = ~n16502 & n16512;
  assign n18618 = ~n16508 & ~n16511;
  assign n18619 = n16352 & ~n18618;
  assign n18620 = ~n18617 & ~n18619;
  assign n18621 = ~n16466 & ~n16479;
  assign n18622 = n16478 & ~n18621;
  assign n18623 = ~n16468 & ~n16485;
  assign n18624 = n16445 & ~n18623;
  assign n18625 = ~n16505 & ~n16512;
  assign n18626 = ~n16458 & n18625;
  assign n18627 = n16352 & ~n18626;
  assign n18628 = ~n18624 & ~n18627;
  assign n18629 = ~n16451 & ~n16462;
  assign n18630 = n18629 ^ n16489;
  assign n18631 = n18629 ^ n16478;
  assign n18632 = n18631 ^ n16478;
  assign n18633 = n16478 ^ n16455;
  assign n18634 = n18632 & ~n18633;
  assign n18635 = n18634 ^ n16478;
  assign n18636 = n18630 & n18635;
  assign n18637 = n18636 ^ n16489;
  assign n18638 = n16509 & n18637;
  assign n18639 = n16318 & ~n18638;
  assign n18640 = n18628 & ~n18639;
  assign n18641 = n16454 & n18640;
  assign n18642 = ~n18622 & n18641;
  assign n18643 = n18620 & n18642;
  assign n18644 = n18616 & n18643;
  assign n18645 = n16488 & n18644;
  assign n18646 = ~n16465 & n18645;
  assign n18647 = n16464 & n18646;
  assign n18648 = n18647 ^ n14437;
  assign n18649 = n18648 ^ x67;
  assign n18650 = ~n18613 & ~n18649;
  assign n18651 = n18612 & n18650;
  assign n18652 = n18581 & n18651;
  assign n18653 = ~n18582 & ~n18611;
  assign n18654 = ~n18613 & n18649;
  assign n18655 = n18653 & n18654;
  assign n18656 = n18581 & n18655;
  assign n18657 = n18579 & n18580;
  assign n18658 = n18613 & ~n18649;
  assign n18659 = n18653 & n18658;
  assign n18660 = n18657 & n18659;
  assign n18661 = ~n18656 & ~n18660;
  assign n18662 = n18579 & ~n18580;
  assign n18663 = n18651 & n18662;
  assign n18664 = n18613 & n18649;
  assign n18665 = n18612 & n18664;
  assign n18666 = n18653 & n18664;
  assign n18667 = ~n18665 & ~n18666;
  assign n18668 = n18657 & ~n18667;
  assign n18669 = ~n18663 & ~n18668;
  assign n18670 = ~n18582 & n18611;
  assign n18671 = n18658 & n18670;
  assign n18672 = n18581 & n18671;
  assign n18673 = n18650 & n18653;
  assign n18674 = n18612 & n18654;
  assign n18675 = n18650 & n18670;
  assign n18676 = ~n18674 & ~n18675;
  assign n18677 = ~n18673 & n18676;
  assign n18678 = n18662 & ~n18677;
  assign n18679 = n18654 ^ n18650;
  assign n18680 = ~n18611 & n18679;
  assign n18681 = ~n18582 & n18680;
  assign n18682 = n18681 ^ n18650;
  assign n18683 = n18657 & n18682;
  assign n18684 = ~n18579 & ~n18580;
  assign n18685 = n18582 & ~n18611;
  assign n18686 = n18654 & n18685;
  assign n18687 = n18664 & n18685;
  assign n18688 = ~n18659 & ~n18687;
  assign n18689 = n18654 & n18670;
  assign n18690 = n18650 & n18685;
  assign n18691 = ~n18689 & ~n18690;
  assign n18692 = n18612 & n18658;
  assign n18693 = ~n18671 & ~n18692;
  assign n18694 = n18691 & n18693;
  assign n18695 = n18688 & n18694;
  assign n18696 = ~n18686 & n18695;
  assign n18697 = n18684 & ~n18696;
  assign n18698 = ~n18581 & ~n18662;
  assign n18699 = n18664 & n18670;
  assign n18700 = n18658 & n18685;
  assign n18701 = ~n18699 & ~n18700;
  assign n18702 = ~n18666 & ~n18687;
  assign n18703 = ~n18662 & n18702;
  assign n18704 = ~n18686 & ~n18692;
  assign n18705 = ~n18581 & n18704;
  assign n18706 = ~n18703 & ~n18705;
  assign n18707 = n18701 & ~n18706;
  assign n18708 = ~n18698 & ~n18707;
  assign n18709 = ~n18697 & ~n18708;
  assign n18710 = ~n18683 & n18709;
  assign n18711 = ~n18678 & n18710;
  assign n18712 = ~n18672 & n18711;
  assign n18713 = n18700 ^ n18674;
  assign n18714 = n18713 ^ n18674;
  assign n18715 = n18674 ^ n18580;
  assign n18716 = n18715 ^ n18674;
  assign n18717 = n18714 & n18716;
  assign n18718 = n18717 ^ n18674;
  assign n18719 = n18579 & n18718;
  assign n18720 = n18719 ^ n18674;
  assign n18721 = n18712 & ~n18720;
  assign n18722 = n18669 & n18721;
  assign n18723 = n18661 & n18722;
  assign n18724 = ~n18652 & n18723;
  assign n18725 = n18724 ^ n16411;
  assign n18726 = n18725 ^ x82;
  assign n18727 = ~n18578 & n18726;
  assign n18728 = ~n18550 & n18727;
  assign n18729 = ~n18464 & n18487;
  assign n18730 = n18524 & n18729;
  assign n18731 = ~n18545 & n18730;
  assign n18732 = ~n18549 & ~n18731;
  assign n18733 = n18578 & ~n18726;
  assign n18734 = ~n18732 & n18733;
  assign n18735 = ~n18728 & ~n18734;
  assign n18736 = n18524 & n18545;
  assign n18737 = n18488 & n18736;
  assign n18738 = n18545 & n18730;
  assign n18739 = ~n18737 & ~n18738;
  assign n18740 = ~n18727 & ~n18733;
  assign n18741 = ~n18739 & ~n18740;
  assign n18742 = n18548 & n18729;
  assign n18743 = ~n18524 & n18545;
  assign n18744 = n18729 & n18743;
  assign n18745 = ~n18547 & ~n18744;
  assign n18746 = ~n18742 & n18745;
  assign n18747 = ~n18731 & n18746;
  assign n18748 = ~n18578 & ~n18726;
  assign n18749 = ~n18747 & n18748;
  assign n18750 = ~n18464 & ~n18487;
  assign n18751 = n18546 & n18750;
  assign n18752 = n18733 & n18751;
  assign n18753 = n18464 & ~n18487;
  assign n18754 = n18548 & n18753;
  assign n18755 = n18748 & n18754;
  assign n18756 = n18733 & n18754;
  assign n18757 = ~n18755 & ~n18756;
  assign n18758 = n18743 & n18753;
  assign n18759 = n18736 & n18753;
  assign n18760 = n18736 & n18750;
  assign n18761 = ~n18759 & ~n18760;
  assign n18762 = ~n18758 & n18761;
  assign n18763 = n18748 & ~n18762;
  assign n18764 = n18578 & n18726;
  assign n18765 = n18548 & n18750;
  assign n18766 = n18746 & n18762;
  assign n18767 = ~n18549 & n18766;
  assign n18768 = ~n18765 & n18767;
  assign n18769 = n18764 & ~n18768;
  assign n18770 = ~n18763 & ~n18769;
  assign n18771 = n18743 & n18750;
  assign n18775 = n18488 & n18743;
  assign n18772 = n18546 & n18753;
  assign n18773 = ~n18751 & ~n18765;
  assign n18774 = ~n18772 & n18773;
  assign n18776 = n18775 ^ n18774;
  assign n18777 = n18733 ^ n18727;
  assign n18778 = n18774 ^ n18727;
  assign n18779 = n18778 ^ n18727;
  assign n18780 = ~n18777 & n18779;
  assign n18781 = n18780 ^ n18727;
  assign n18782 = ~n18776 & n18781;
  assign n18783 = n18782 ^ n18775;
  assign n18784 = ~n18771 & ~n18783;
  assign n18785 = ~n18740 & ~n18784;
  assign n18786 = n18770 & ~n18785;
  assign n18787 = n18757 & n18786;
  assign n18788 = ~n18752 & n18787;
  assign n18789 = ~n18749 & n18788;
  assign n18790 = ~n18741 & n18789;
  assign n18791 = n18735 & n18790;
  assign n18792 = n18791 ^ n17741;
  assign n18793 = n18792 ^ x93;
  assign n18794 = n18447 & n18793;
  assign n18795 = ~n16706 & n16736;
  assign n18796 = ~n16684 & ~n16723;
  assign n18797 = n16680 & ~n18796;
  assign n18798 = ~n16691 & n16727;
  assign n18799 = n16685 & ~n18798;
  assign n18800 = ~n18797 & ~n18799;
  assign n18801 = ~n18795 & n18800;
  assign n18802 = n16314 & n16721;
  assign n18803 = n16127 ^ n15398;
  assign n18804 = n18803 ^ n16312;
  assign n18805 = n18804 ^ n15881;
  assign n18806 = n16312 ^ n15398;
  assign n18807 = n15881 ^ n15398;
  assign n18808 = n18806 & ~n18807;
  assign n18809 = n18808 ^ n15398;
  assign n18810 = n18805 & n18809;
  assign n18811 = n16706 & n18810;
  assign n18812 = ~n18802 & ~n18811;
  assign n18813 = n16680 & n16726;
  assign n18814 = n16702 & ~n18319;
  assign n18815 = ~n18813 & ~n18814;
  assign n18816 = n18812 & n18815;
  assign n18817 = n16700 & n18816;
  assign n18818 = n18306 & n18817;
  assign n18819 = n18301 & n18818;
  assign n18820 = n18801 & n18819;
  assign n18821 = n18820 ^ n15773;
  assign n18822 = n18821 ^ x102;
  assign n18823 = n17086 ^ x109;
  assign n18824 = ~n18822 & n18823;
  assign n18825 = ~n17850 & n17927;
  assign n18826 = n17851 & ~n18270;
  assign n18827 = ~n18825 & ~n18826;
  assign n18828 = n17929 & n17966;
  assign n18829 = ~n17919 & ~n17927;
  assign n18830 = n18283 & n18829;
  assign n18831 = n17959 & n18830;
  assign n18832 = n17913 & ~n18831;
  assign n18833 = ~n18828 & ~n18832;
  assign n18834 = ~n17929 & ~n17949;
  assign n18835 = n17959 & n17962;
  assign n18836 = ~n18834 & ~n18835;
  assign n18837 = n17851 & n18836;
  assign n18839 = ~n17931 & ~n17944;
  assign n18838 = ~n17915 & n18273;
  assign n18840 = n18839 ^ n18838;
  assign n18841 = n18839 ^ n17925;
  assign n18842 = n18839 & n18841;
  assign n18843 = n18842 ^ n18839;
  assign n18844 = n18840 & n18843;
  assign n18845 = n18844 ^ n18842;
  assign n18846 = n18845 ^ n18839;
  assign n18847 = n18846 ^ n17925;
  assign n18848 = ~n18837 & n18847;
  assign n18849 = n18848 ^ n18837;
  assign n18850 = n18833 & ~n18849;
  assign n18851 = n18827 & n18850;
  assign n18852 = ~n18260 & n18851;
  assign n18853 = n17946 & n18852;
  assign n18854 = ~n17924 & n18853;
  assign n18855 = n17917 & n18854;
  assign n18856 = n18855 ^ n15605;
  assign n18857 = n18856 ^ x69;
  assign n18858 = n18198 & n18208;
  assign n18859 = n18213 & n18858;
  assign n18860 = ~n18207 & ~n18859;
  assign n18861 = n18494 & n18858;
  assign n18862 = n18192 & n18218;
  assign n18863 = ~n18861 & ~n18862;
  assign n18864 = n18216 & n18512;
  assign n18865 = n18206 & ~n18864;
  assign n18866 = n18493 & n18504;
  assign n18867 = n18213 & ~n18866;
  assign n18868 = ~n18865 & ~n18867;
  assign n18869 = n18196 & n18494;
  assign n18870 = ~n18494 & ~n18496;
  assign n18871 = ~n18217 & ~n18226;
  assign n18872 = ~n18206 & n18871;
  assign n18873 = ~n18870 & ~n18872;
  assign n18874 = ~n18214 & ~n18873;
  assign n18875 = ~n18189 & n18874;
  assign n18876 = n18875 ^ n18191;
  assign n18877 = n18876 ^ n18875;
  assign n18878 = ~n18209 & ~n18502;
  assign n18879 = n18878 ^ n18875;
  assign n18880 = n18879 ^ n18875;
  assign n18881 = n18877 & ~n18880;
  assign n18882 = n18881 ^ n18875;
  assign n18883 = ~n18190 & ~n18882;
  assign n18884 = n18883 ^ n18875;
  assign n18885 = ~n18869 & n18884;
  assign n18886 = n18868 & n18885;
  assign n18887 = ~n18500 & n18886;
  assign n18888 = n18498 & n18887;
  assign n18889 = n18863 & n18888;
  assign n18890 = ~n18203 & n18889;
  assign n18891 = n18860 & n18890;
  assign n18892 = ~n18197 & n18891;
  assign n18893 = n18892 ^ n15648;
  assign n18894 = n18893 ^ x84;
  assign n18895 = n18857 & n18894;
  assign n18896 = n18824 & n18895;
  assign n18897 = n17848 ^ x126;
  assign n18898 = n18684 & n18700;
  assign n18899 = n18662 & ~n18667;
  assign n18900 = ~n18655 & n18691;
  assign n18901 = n18657 & ~n18900;
  assign n18902 = ~n18899 & ~n18901;
  assign n18903 = ~n18580 & n18659;
  assign n18904 = ~n18579 & n18692;
  assign n18905 = ~n18903 & ~n18904;
  assign n18906 = n18666 & n18684;
  assign n18907 = n18657 & n18686;
  assign n18908 = n18662 & n18686;
  assign n18909 = n18657 & n18671;
  assign n18910 = ~n18908 & ~n18909;
  assign n18911 = ~n18665 & ~n18699;
  assign n18912 = ~n18687 & n18911;
  assign n18913 = n18581 & ~n18912;
  assign n18914 = ~n18673 & ~n18689;
  assign n18915 = ~n18700 & n18914;
  assign n18916 = n18662 & ~n18915;
  assign n18917 = ~n18913 & ~n18916;
  assign n18918 = n18657 & n18692;
  assign n18920 = ~n18673 & ~n18690;
  assign n18921 = ~n18671 & n18920;
  assign n18919 = n18677 & ~n18686;
  assign n18922 = n18921 ^ n18919;
  assign n18923 = n18921 ^ n18580;
  assign n18924 = n18923 ^ n18921;
  assign n18925 = n18922 & ~n18924;
  assign n18926 = n18925 ^ n18921;
  assign n18927 = ~n18579 & ~n18926;
  assign n18928 = ~n18918 & ~n18927;
  assign n18929 = n18917 & n18928;
  assign n18930 = n18669 & n18929;
  assign n18931 = ~n18652 & n18930;
  assign n18932 = n18910 & n18931;
  assign n18933 = ~n18907 & n18932;
  assign n18934 = ~n18906 & n18933;
  assign n18935 = n18905 & n18934;
  assign n18936 = n18902 & n18935;
  assign n18937 = ~n18898 & n18936;
  assign n18938 = n18937 ^ n15469;
  assign n18939 = n18938 ^ x108;
  assign n18940 = n18897 & n18939;
  assign n18941 = n18896 & n18940;
  assign n18942 = ~n18857 & ~n18894;
  assign n18943 = n18824 & n18942;
  assign n18944 = n18897 & ~n18939;
  assign n18945 = n18943 & n18944;
  assign n18946 = ~n18941 & ~n18945;
  assign n18947 = ~n18857 & n18894;
  assign n18948 = n18824 & n18947;
  assign n18949 = n18944 & n18948;
  assign n18950 = ~n18822 & ~n18823;
  assign n18951 = n18947 & n18950;
  assign n18952 = n18944 & n18951;
  assign n18953 = ~n18897 & n18939;
  assign n18954 = n18857 & ~n18894;
  assign n18955 = n18824 & n18954;
  assign n18956 = n18822 & n18823;
  assign n18957 = n18942 & n18956;
  assign n18958 = ~n18955 & ~n18957;
  assign n18959 = n18953 & ~n18958;
  assign n18960 = ~n18952 & ~n18959;
  assign n18961 = ~n18897 & ~n18939;
  assign n18962 = n18954 & n18956;
  assign n18963 = ~n18896 & ~n18962;
  assign n18964 = n18961 & ~n18963;
  assign n18965 = n18950 & n18954;
  assign n18966 = n18822 & ~n18823;
  assign n18967 = n18954 & n18966;
  assign n18968 = n18947 & n18966;
  assign n18969 = n18942 & n18950;
  assign n18970 = ~n18968 & ~n18969;
  assign n18971 = ~n18967 & n18970;
  assign n18972 = ~n18965 & n18971;
  assign n18973 = n18953 & ~n18972;
  assign n18974 = n18896 & n18953;
  assign n18975 = ~n18940 & ~n18961;
  assign n18976 = ~n18970 & ~n18975;
  assign n18977 = ~n18974 & ~n18976;
  assign n18984 = n18895 & n18966;
  assign n18985 = n18958 & ~n18984;
  assign n18978 = n18942 & n18966;
  assign n18979 = n18895 & n18956;
  assign n18980 = ~n18948 & ~n18979;
  assign n18981 = ~n18962 & ~n18965;
  assign n18982 = n18980 & n18981;
  assign n18983 = ~n18978 & n18982;
  assign n18986 = n18985 ^ n18983;
  assign n18987 = n18986 ^ n18985;
  assign n18988 = n18985 ^ n18897;
  assign n18989 = n18988 ^ n18985;
  assign n18990 = ~n18987 & n18989;
  assign n18991 = n18990 ^ n18985;
  assign n18992 = n18939 & ~n18991;
  assign n18993 = n18992 ^ n18985;
  assign n18994 = n18977 & n18993;
  assign n18995 = ~n18973 & n18994;
  assign n18998 = n18947 & n18956;
  assign n18996 = n18895 & n18950;
  assign n18997 = ~n18967 & ~n18996;
  assign n18999 = n18998 ^ n18997;
  assign n19000 = n18999 ^ n18998;
  assign n19001 = n18998 ^ n18939;
  assign n19002 = n19001 ^ n18998;
  assign n19003 = ~n19000 & ~n19002;
  assign n19004 = n19003 ^ n18998;
  assign n19005 = n18897 & n19004;
  assign n19006 = n19005 ^ n18998;
  assign n19007 = n18995 & ~n19006;
  assign n19008 = ~n18964 & n19007;
  assign n19009 = n18960 & n19008;
  assign n19010 = ~n18949 & n19009;
  assign n19011 = n18946 & n19010;
  assign n19012 = n19011 ^ n18610;
  assign n19013 = n19012 ^ x125;
  assign n19014 = n17984 ^ x120;
  assign n19096 = n18523 ^ x73;
  assign n19015 = n18577 ^ x80;
  assign n19016 = n16757 ^ x97;
  assign n19017 = ~n18579 & n18699;
  assign n19018 = n18657 & ~n18676;
  assign n19019 = ~n19017 & ~n19018;
  assign n19020 = ~n18666 & ~n18700;
  assign n19021 = ~n18692 & n19020;
  assign n19022 = n18581 & ~n19021;
  assign n19023 = n18693 & n18920;
  assign n19024 = ~n18674 & n19023;
  assign n19025 = n18662 & ~n19024;
  assign n19026 = ~n18688 & n18698;
  assign n19027 = ~n18686 & n18914;
  assign n19028 = n18581 & ~n19027;
  assign n19029 = ~n18655 & n18676;
  assign n19030 = ~n18671 & n19029;
  assign n19031 = n18684 & ~n19030;
  assign n19032 = ~n19028 & ~n19031;
  assign n19033 = ~n19026 & n19032;
  assign n19034 = ~n18652 & n19033;
  assign n19035 = ~n19025 & n19034;
  assign n19036 = ~n19022 & n19035;
  assign n19037 = n19019 & n19036;
  assign n19038 = n18902 & n19037;
  assign n19039 = ~n18898 & n19038;
  assign n19040 = n18910 & n19039;
  assign n19041 = n19040 ^ n15971;
  assign n19042 = n19041 ^ x115;
  assign n19043 = n19016 & n19042;
  assign n19044 = n19015 & n19043;
  assign n19045 = n16808 & n17022;
  assign n19046 = ~n16807 & ~n17064;
  assign n19047 = n17026 & ~n17067;
  assign n19048 = ~n19046 & ~n19047;
  assign n19049 = n17017 & n17047;
  assign n19050 = ~n17031 & ~n17048;
  assign n19051 = ~n17036 & n19050;
  assign n19052 = n17042 & ~n19051;
  assign n19053 = ~n19049 & ~n19052;
  assign n19054 = ~n17049 & n17074;
  assign n19055 = ~n16807 & ~n19054;
  assign n19056 = ~n17052 & ~n17058;
  assign n19057 = ~n17043 & ~n17073;
  assign n19058 = n19056 & n19057;
  assign n19059 = n17039 & n19058;
  assign n19060 = n16808 & ~n19059;
  assign n19061 = ~n19055 & ~n19060;
  assign n19062 = n19053 & n19061;
  assign n19063 = n17067 ^ n17063;
  assign n19064 = n19063 ^ n17063;
  assign n19065 = n17063 ^ n16776;
  assign n19066 = n19065 ^ n17063;
  assign n19067 = ~n19064 & ~n19066;
  assign n19068 = n19067 ^ n17063;
  assign n19069 = ~n16807 & n19068;
  assign n19070 = n19069 ^ n17063;
  assign n19071 = n19062 & ~n19070;
  assign n19072 = n19048 & n19071;
  assign n19073 = n17062 & n19072;
  assign n19074 = ~n19045 & n19073;
  assign n19075 = n19074 ^ n16075;
  assign n19076 = n19075 ^ x106;
  assign n19077 = n19044 & n19076;
  assign n19078 = ~n19015 & ~n19042;
  assign n19079 = n19016 & n19078;
  assign n19080 = n19076 & n19079;
  assign n19081 = ~n19077 & ~n19080;
  assign n19082 = ~n19076 & n19078;
  assign n19083 = n19015 & ~n19042;
  assign n19084 = n19016 & n19083;
  assign n19085 = n19076 & n19084;
  assign n19086 = ~n19082 & ~n19085;
  assign n19089 = ~n19015 & ~n19016;
  assign n19087 = ~n19016 & n19042;
  assign n19088 = n19015 & n19087;
  assign n19090 = n19089 ^ n19088;
  assign n19091 = n19076 & n19090;
  assign n19092 = n19091 ^ n19089;
  assign n19093 = n19086 & ~n19092;
  assign n19094 = n19081 & n19093;
  assign n19095 = ~n19044 & n19094;
  assign n19097 = n19096 ^ n19095;
  assign n19098 = n19097 ^ n19095;
  assign n19099 = ~n19016 & n19083;
  assign n19100 = ~n19076 & n19099;
  assign n19101 = ~n19076 & n19088;
  assign n19102 = ~n19015 & n19087;
  assign n19103 = n19076 & n19102;
  assign n19104 = n19086 & ~n19103;
  assign n19105 = ~n19101 & n19104;
  assign n19106 = n19081 & n19105;
  assign n19107 = ~n19100 & n19106;
  assign n19108 = n19107 ^ n19095;
  assign n19109 = n19098 & ~n19108;
  assign n19110 = n19109 ^ n19095;
  assign n19111 = ~n19014 & ~n19110;
  assign n19112 = ~n19015 & n19043;
  assign n19113 = ~n19076 & n19112;
  assign n19114 = ~n19085 & ~n19113;
  assign n19115 = ~n19100 & n19114;
  assign n19116 = ~n19082 & ~n19103;
  assign n19117 = n19099 ^ n19044;
  assign n19118 = n19076 & n19117;
  assign n19119 = n19118 ^ n19044;
  assign n19120 = n19116 & ~n19119;
  assign n19121 = n19115 & n19120;
  assign n19122 = n19121 ^ n19096;
  assign n19123 = n19122 ^ n19121;
  assign n19124 = n19042 ^ n19015;
  assign n19125 = n19124 ^ n19015;
  assign n19126 = n19016 ^ n19015;
  assign n19127 = n19126 ^ n19042;
  assign n19128 = n19127 ^ n19015;
  assign n19129 = n19128 ^ n19015;
  assign n19130 = ~n19125 & n19129;
  assign n19131 = n19130 ^ n19015;
  assign n19132 = n19076 & n19131;
  assign n19133 = n19132 ^ n19127;
  assign n19134 = n19133 ^ n19121;
  assign n19135 = n19123 & n19134;
  assign n19136 = n19135 ^ n19121;
  assign n19137 = n19014 & ~n19136;
  assign n19138 = ~n19111 & ~n19137;
  assign n19139 = n19138 ^ n17120;
  assign n19140 = n19139 ^ x108;
  assign n19141 = n18102 ^ x65;
  assign n19142 = n17420 & n17471;
  assign n19143 = n17426 & n18526;
  assign n19144 = ~n19142 & ~n19143;
  assign n19145 = n17422 & ~n17453;
  assign n19146 = ~n17428 & ~n17445;
  assign n19147 = ~n17436 & ~n19146;
  assign n19148 = n17447 & n18350;
  assign n19149 = n17162 & ~n19148;
  assign n19150 = ~n17420 & ~n18342;
  assign n19151 = ~n17422 & n19150;
  assign n19152 = ~n17431 & ~n17456;
  assign n19153 = ~n17426 & n19152;
  assign n19154 = ~n19151 & ~n19153;
  assign n19155 = ~n17437 & ~n19154;
  assign n19156 = ~n17457 & n19155;
  assign n19157 = n19156 ^ n17436;
  assign n19158 = n19157 ^ n19156;
  assign n19159 = ~n17443 & n18350;
  assign n19160 = n17471 & ~n19159;
  assign n19161 = ~n17424 & ~n19160;
  assign n19162 = n17473 & n19161;
  assign n19163 = ~n17431 & n19162;
  assign n19164 = n19163 ^ n19156;
  assign n19165 = n19158 & n19164;
  assign n19166 = n19165 ^ n19156;
  assign n19167 = ~n19149 & n19166;
  assign n19168 = ~n19147 & n19167;
  assign n19169 = ~n19145 & n19168;
  assign n19170 = n19144 & n19169;
  assign n19171 = n19170 ^ n14397;
  assign n19172 = n19171 ^ x99;
  assign n19173 = n19141 & ~n19172;
  assign n19174 = n17525 & n17647;
  assign n19175 = ~n17633 & ~n17637;
  assign n19176 = n17628 & ~n19175;
  assign n19177 = ~n19174 & ~n19176;
  assign n19178 = ~n17631 & n17679;
  assign n19179 = ~n17622 & ~n17660;
  assign n19180 = n17619 & ~n19179;
  assign n19181 = ~n19178 & ~n19180;
  assign n19182 = ~n17626 & ~n17648;
  assign n19183 = n17644 & ~n19182;
  assign n19184 = ~n17639 & ~n17655;
  assign n19185 = n17668 & n19184;
  assign n19186 = n17628 & ~n19185;
  assign n19187 = n17640 & ~n17654;
  assign n19188 = ~n17622 & n19187;
  assign n19189 = n17644 & ~n19188;
  assign n19190 = n18107 & n19175;
  assign n19191 = n17619 & ~n19190;
  assign n19192 = ~n17635 & n17661;
  assign n19193 = ~n17655 & n19192;
  assign n19194 = n17525 & ~n19193;
  assign n19195 = ~n19191 & ~n19194;
  assign n19196 = ~n19189 & n19195;
  assign n19197 = ~n19186 & n19196;
  assign n19198 = ~n19183 & n19197;
  assign n19199 = n19181 & n19198;
  assign n19200 = n19177 & n19199;
  assign n19201 = n18552 & n19200;
  assign n19202 = n18112 & n19201;
  assign n19203 = n19202 ^ n14971;
  assign n19204 = n19203 ^ x113;
  assign n19205 = n18673 & n18684;
  assign n19206 = ~n18651 & n18911;
  assign n19207 = ~n18686 & n19206;
  assign n19208 = n18657 & ~n19207;
  assign n19209 = ~n19205 & ~n19208;
  assign n19210 = ~n18579 & n18690;
  assign n19211 = ~n18689 & ~n18692;
  assign n19212 = n18581 & ~n19211;
  assign n19213 = ~n18665 & n18693;
  assign n19214 = n18684 & ~n19213;
  assign n19215 = n18688 & n18701;
  assign n19216 = n18581 & ~n19215;
  assign n19217 = ~n19214 & ~n19216;
  assign n19218 = n18691 & n19021;
  assign n19219 = ~n18675 & n19218;
  assign n19220 = ~n18687 & n19219;
  assign n19221 = n19220 ^ n18581;
  assign n19222 = n19221 ^ n19220;
  assign n19223 = ~n18655 & ~n18674;
  assign n19224 = n19223 ^ n19220;
  assign n19225 = n19224 ^ n19220;
  assign n19226 = ~n19222 & ~n19225;
  assign n19227 = n19226 ^ n19220;
  assign n19228 = ~n18662 & ~n19227;
  assign n19229 = n19228 ^ n19220;
  assign n19230 = n19217 & n19229;
  assign n19231 = ~n18898 & n19230;
  assign n19232 = ~n19212 & n19231;
  assign n19233 = ~n19210 & n19232;
  assign n19234 = n19209 & n19233;
  assign n19235 = n18661 & n19234;
  assign n19236 = n18910 & n19235;
  assign n19237 = n19236 ^ n14686;
  assign n19238 = n19237 ^ x74;
  assign n19239 = ~n19204 & ~n19238;
  assign n19240 = n19173 & n19239;
  assign n19241 = n18254 ^ x89;
  assign n19242 = n17026 & n17063;
  assign n19243 = n17042 & n17049;
  assign n19244 = ~n19242 & ~n19243;
  assign n19245 = n17037 & ~n17047;
  assign n19246 = ~n17052 & n17075;
  assign n19247 = n17019 & ~n19246;
  assign n19248 = ~n19245 & ~n19247;
  assign n19249 = n17022 & n17042;
  assign n19250 = n17026 & ~n19056;
  assign n19251 = ~n19249 & ~n19250;
  assign n19252 = n17047 & n17063;
  assign n19253 = n17048 ^ n16807;
  assign n19255 = ~n17056 & n19056;
  assign n19256 = ~n17031 & n19255;
  assign n19254 = ~n17058 & n17075;
  assign n19257 = n19256 ^ n19254;
  assign n19258 = n19256 ^ n16776;
  assign n19259 = n19258 ^ n19256;
  assign n19260 = n19257 & n19259;
  assign n19261 = n19260 ^ n19256;
  assign n19262 = n19261 ^ n17048;
  assign n19263 = ~n19253 & ~n19262;
  assign n19264 = n19263 ^ n19260;
  assign n19265 = n19264 ^ n19256;
  assign n19266 = n19265 ^ n16807;
  assign n19267 = ~n17048 & n19266;
  assign n19268 = n19267 ^ n17048;
  assign n19269 = n19268 ^ n16807;
  assign n19270 = ~n19252 & n19269;
  assign n19271 = n19251 & n19270;
  assign n19272 = n19248 & n19271;
  assign n19273 = n19244 & n19272;
  assign n19274 = n19048 & n19273;
  assign n19275 = ~n19045 & n19274;
  assign n19276 = n17024 & n19275;
  assign n19277 = n19276 ^ n15331;
  assign n19278 = n19277 ^ x96;
  assign n19279 = n19241 & ~n19278;
  assign n19280 = n19240 & n19279;
  assign n19281 = ~n19141 & n19172;
  assign n19282 = n19239 & n19281;
  assign n19283 = ~n19241 & ~n19278;
  assign n19284 = n19282 & n19283;
  assign n19285 = ~n19241 & n19278;
  assign n19286 = n19204 & ~n19238;
  assign n19287 = n19173 & n19286;
  assign n19288 = n19141 & n19172;
  assign n19289 = n19239 & n19288;
  assign n19290 = ~n19287 & ~n19289;
  assign n19291 = n19285 & ~n19290;
  assign n19292 = ~n19284 & ~n19291;
  assign n19293 = n19241 & n19278;
  assign n19294 = ~n19204 & n19238;
  assign n19295 = n19288 & n19294;
  assign n19296 = ~n19240 & ~n19295;
  assign n19297 = n19293 & ~n19296;
  assign n19298 = n19204 & n19238;
  assign n19299 = n19288 & n19298;
  assign n19300 = n19173 & n19298;
  assign n19301 = n19286 & n19288;
  assign n19302 = ~n19300 & ~n19301;
  assign n19303 = ~n19299 & n19302;
  assign n19304 = n19279 & ~n19303;
  assign n19305 = ~n19141 & ~n19172;
  assign n19306 = n19298 & n19305;
  assign n19307 = n19281 & n19286;
  assign n19308 = n19286 & n19305;
  assign n19309 = ~n19307 & ~n19308;
  assign n19310 = n19173 & n19294;
  assign n19311 = ~n19287 & ~n19310;
  assign n19312 = ~n19299 & n19311;
  assign n19313 = n19309 & n19312;
  assign n19314 = ~n19306 & n19313;
  assign n19315 = ~n19295 & n19314;
  assign n19316 = n19283 & ~n19315;
  assign n19317 = ~n19304 & ~n19316;
  assign n19318 = n19239 & n19305;
  assign n19319 = n19281 & n19298;
  assign n19320 = ~n19308 & ~n19319;
  assign n19321 = ~n19318 & n19320;
  assign n19322 = ~n19300 & n19321;
  assign n19323 = ~n19299 & n19322;
  assign n19324 = ~n19282 & n19323;
  assign n19325 = n19293 & ~n19324;
  assign n19326 = n19281 & n19294;
  assign n19327 = ~n19282 & n19309;
  assign n19328 = ~n19326 & n19327;
  assign n19329 = n19279 & ~n19328;
  assign n19330 = n19204 ^ n19172;
  assign n19331 = n19330 ^ n19172;
  assign n19332 = n19331 ^ n19238;
  assign n19333 = n19172 ^ n19141;
  assign n19334 = n19238 ^ n19141;
  assign n19335 = n19334 ^ n19141;
  assign n19336 = ~n19333 & ~n19335;
  assign n19337 = n19336 ^ n19141;
  assign n19338 = ~n19332 & n19337;
  assign n19339 = n19338 ^ n19330;
  assign n19340 = n19285 & ~n19339;
  assign n19341 = ~n19329 & ~n19340;
  assign n19342 = ~n19325 & n19341;
  assign n19343 = n19317 & n19342;
  assign n19344 = ~n19297 & n19343;
  assign n19345 = n19292 & n19344;
  assign n19346 = ~n19280 & n19345;
  assign n19347 = n19346 ^ n17712;
  assign n19348 = n19347 ^ x68;
  assign n19349 = n19140 & n19348;
  assign n19350 = n18486 ^ x121;
  assign n19351 = n19171 ^ x112;
  assign n19352 = n19350 & n19351;
  assign n19353 = ~n16316 & ~n16732;
  assign n19354 = ~n16705 & n19353;
  assign n19355 = n16703 & ~n19354;
  assign n19356 = ~n16705 & n18304;
  assign n19357 = n16685 & ~n19356;
  assign n19358 = ~n19355 & ~n19357;
  assign n19359 = n16680 & n16720;
  assign n19360 = ~n16702 & ~n16732;
  assign n19361 = ~n16526 & ~n19360;
  assign n19362 = n16725 & n18299;
  assign n19363 = n16706 & ~n19362;
  assign n19364 = ~n19361 & ~n19363;
  assign n19365 = ~n19359 & n19364;
  assign n19366 = n19358 & n19365;
  assign n19367 = n16719 & n19366;
  assign n19368 = ~n16681 & n19367;
  assign n19369 = n18801 & n19368;
  assign n19370 = n19369 ^ n16379;
  assign n19371 = n19370 ^ x81;
  assign n19372 = n18213 & ~n18227;
  assign n19373 = ~n18209 & ~n18226;
  assign n19374 = ~n18496 & n19373;
  assign n19375 = n18231 & ~n19374;
  assign n19376 = ~n19372 & ~n19375;
  assign n19377 = ~n18210 & ~n18214;
  assign n19378 = ~n18496 & n19377;
  assign n19379 = ~n18217 & n19378;
  assign n19380 = n18494 & ~n19379;
  assign n19381 = n18192 & ~n18216;
  assign n19382 = ~n18502 & n18509;
  assign n19383 = n18494 & ~n19382;
  assign n19384 = ~n19381 & ~n19383;
  assign n19385 = ~n18200 & n18493;
  assign n19386 = ~n18189 & n19385;
  assign n19387 = n19386 ^ n18190;
  assign n19388 = n19387 ^ n19386;
  assign n19389 = n18503 & n19377;
  assign n19390 = n19389 ^ n19386;
  assign n19391 = ~n19388 & n19390;
  assign n19392 = n19391 ^ n19386;
  assign n19393 = ~n18191 & ~n19392;
  assign n19394 = n19384 & ~n19393;
  assign n19395 = n18863 & n19394;
  assign n19396 = ~n18193 & n19395;
  assign n19397 = ~n19380 & n19396;
  assign n19398 = n19376 & n19397;
  assign n19399 = n18491 & n19398;
  assign n19400 = n18860 & n19399;
  assign n19401 = n19400 ^ n16438;
  assign n19402 = n19401 ^ x88;
  assign n19403 = ~n19371 & ~n19402;
  assign n19404 = n19277 ^ x107;
  assign n19405 = n18725 ^ x98;
  assign n19406 = ~n19404 & n19405;
  assign n19407 = n19403 & n19406;
  assign n19408 = n19352 & n19407;
  assign n19409 = n19350 & ~n19351;
  assign n19410 = n19371 & n19402;
  assign n19411 = n19404 & ~n19405;
  assign n19412 = n19410 & n19411;
  assign n19413 = n19409 & n19412;
  assign n19414 = ~n19350 & n19351;
  assign n19415 = ~n19371 & n19402;
  assign n19416 = ~n19404 & ~n19405;
  assign n19417 = n19415 & n19416;
  assign n19418 = n19406 & n19410;
  assign n19419 = ~n19417 & ~n19418;
  assign n19420 = n19414 & ~n19419;
  assign n19421 = ~n19413 & ~n19420;
  assign n19422 = ~n19408 & n19421;
  assign n19423 = n19371 & ~n19402;
  assign n19424 = n19406 & n19423;
  assign n19425 = n19409 & n19424;
  assign n19426 = n19404 & n19405;
  assign n19427 = n19415 & n19426;
  assign n19428 = n19352 & n19427;
  assign n19429 = n19409 & n19417;
  assign n19430 = ~n19428 & ~n19429;
  assign n19431 = ~n19425 & n19430;
  assign n19432 = ~n19350 & ~n19351;
  assign n19433 = ~n19352 & ~n19432;
  assign n19434 = n19403 & n19416;
  assign n19435 = ~n19424 & ~n19434;
  assign n19436 = ~n19433 & ~n19435;
  assign n19437 = ~n19352 & ~n19414;
  assign n19438 = n19403 & n19426;
  assign n19439 = n19411 & n19423;
  assign n19440 = ~n19438 & ~n19439;
  assign n19441 = ~n19412 & n19440;
  assign n19442 = ~n19437 & ~n19441;
  assign n19443 = ~n19436 & ~n19442;
  assign n19444 = n19410 & n19416;
  assign n19445 = n19414 & n19444;
  assign n19446 = n19410 & n19426;
  assign n19447 = ~n19434 & ~n19446;
  assign n19448 = ~n19439 & n19447;
  assign n19449 = ~n19427 & n19448;
  assign n19450 = n19409 & ~n19449;
  assign n19451 = ~n19445 & ~n19450;
  assign n19452 = n19443 & n19451;
  assign n19453 = n19406 & n19415;
  assign n19454 = n19453 ^ n19432;
  assign n19455 = n19453 ^ n19414;
  assign n19456 = n19455 ^ n19414;
  assign n19457 = n19416 & n19423;
  assign n19458 = n19403 & n19411;
  assign n19459 = ~n19457 & ~n19458;
  assign n19460 = ~n19427 & n19459;
  assign n19461 = n19460 ^ n19414;
  assign n19462 = ~n19456 & n19461;
  assign n19463 = n19462 ^ n19414;
  assign n19464 = n19454 & n19463;
  assign n19465 = n19464 ^ n19432;
  assign n19466 = n19452 & ~n19465;
  assign n19467 = n19423 & n19426;
  assign n19468 = n19467 ^ n19350;
  assign n19469 = n19468 ^ n19467;
  assign n19470 = n19467 ^ n19444;
  assign n19471 = n19469 & n19470;
  assign n19472 = n19471 ^ n19467;
  assign n19473 = n19351 & n19472;
  assign n19474 = n19466 & ~n19473;
  assign n19475 = n19407 ^ n19350;
  assign n19476 = n19475 ^ n19407;
  assign n19477 = n19411 & n19415;
  assign n19478 = ~n19467 & ~n19477;
  assign n19479 = n19478 ^ n19407;
  assign n19480 = ~n19476 & ~n19479;
  assign n19481 = n19480 ^ n19407;
  assign n19482 = ~n19351 & n19481;
  assign n19483 = n19474 & ~n19482;
  assign n19484 = n19431 & n19483;
  assign n19485 = n19422 & n19484;
  assign n19486 = n19485 ^ n18648;
  assign n19487 = n19486 ^ x110;
  assign n19488 = n19349 & ~n19487;
  assign n19489 = ~n19013 & n19488;
  assign n19490 = n18794 & n19489;
  assign n19491 = ~n18447 & ~n18793;
  assign n19492 = ~n19140 & n19487;
  assign n19493 = n19348 & n19492;
  assign n19494 = ~n19013 & n19493;
  assign n19495 = n19013 & n19488;
  assign n19496 = ~n19494 & ~n19495;
  assign n19497 = n19491 & ~n19496;
  assign n19498 = ~n19490 & ~n19497;
  assign n19499 = n18794 & n19495;
  assign n19500 = ~n18447 & n18793;
  assign n19501 = ~n19013 & ~n19348;
  assign n19502 = n19140 & n19501;
  assign n19503 = n19487 & n19502;
  assign n19504 = n19500 & n19503;
  assign n19505 = ~n19499 & ~n19504;
  assign n19506 = n19013 & ~n19348;
  assign n19507 = n19492 & n19506;
  assign n19508 = ~n19140 & ~n19487;
  assign n19509 = n19348 & n19508;
  assign n19510 = ~n19013 & n19509;
  assign n19511 = ~n19507 & ~n19510;
  assign n19512 = n19491 & ~n19511;
  assign n19513 = n19140 & n19506;
  assign n19514 = n19487 & n19513;
  assign n19515 = n19501 & n19508;
  assign n19516 = n19506 & n19508;
  assign n19517 = ~n19515 & ~n19516;
  assign n19518 = ~n19514 & n19517;
  assign n19519 = ~n19494 & n19518;
  assign n19520 = n18794 & ~n19519;
  assign n19521 = ~n19512 & ~n19520;
  assign n19522 = n18447 & ~n18793;
  assign n19523 = n19349 & n19487;
  assign n19524 = ~n19013 & n19523;
  assign n19525 = n19013 & n19493;
  assign n19526 = ~n19524 & ~n19525;
  assign n19527 = n19013 & n19509;
  assign n19528 = ~n19495 & ~n19527;
  assign n19529 = n19526 & n19528;
  assign n19530 = n19522 & ~n19529;
  assign n19531 = n19013 & n19523;
  assign n19532 = n19491 & n19531;
  assign n19533 = n19507 & n19522;
  assign n19534 = ~n19532 & ~n19533;
  assign n19535 = ~n19487 & n19502;
  assign n19536 = n19522 & n19535;
  assign n19537 = ~n19489 & ~n19510;
  assign n19538 = n19500 & ~n19537;
  assign n19539 = ~n19536 & ~n19538;
  assign n19540 = n19491 & n19525;
  assign n19541 = n18793 ^ n18447;
  assign n19542 = ~n19487 & n19513;
  assign n19543 = ~n19515 & ~n19542;
  assign n19544 = n19543 ^ n18793;
  assign n19545 = n19544 ^ n19543;
  assign n19546 = ~n19527 & ~n19531;
  assign n19547 = n19546 ^ n19543;
  assign n19548 = n19545 & n19547;
  assign n19549 = n19548 ^ n19543;
  assign n19550 = n19541 & ~n19549;
  assign n19551 = ~n19540 & ~n19550;
  assign n19552 = n19539 & n19551;
  assign n19553 = n19534 & n19552;
  assign n19554 = ~n19530 & n19553;
  assign n19555 = n19521 & n19554;
  assign n19556 = n19492 & n19501;
  assign n19557 = ~n19542 & ~n19556;
  assign n19558 = ~n19514 & n19557;
  assign n19559 = n19558 ^ n19502;
  assign n19560 = n19559 ^ n19558;
  assign n19561 = n19558 ^ n19522;
  assign n19562 = n19561 ^ n19558;
  assign n19563 = n19560 & ~n19562;
  assign n19564 = n19563 ^ n19558;
  assign n19565 = ~n19500 & ~n19564;
  assign n19566 = n19565 ^ n19558;
  assign n19567 = n19555 & n19566;
  assign n19568 = n19505 & n19567;
  assign n19569 = n19498 & n19568;
  assign n19570 = n19569 ^ n18725;
  assign n19571 = n18059 ^ x74;
  assign n19572 = n19352 & n19457;
  assign n19573 = ~n19434 & ~n19453;
  assign n19574 = n19352 & ~n19573;
  assign n19575 = n19407 & n19432;
  assign n19576 = n19409 & n19418;
  assign n19577 = n19414 & n19477;
  assign n19578 = ~n19576 & ~n19577;
  assign n19579 = ~n19575 & n19578;
  assign n19580 = ~n19412 & n19478;
  assign n19581 = ~n19433 & ~n19580;
  assign n19582 = n19440 & n19447;
  assign n19583 = ~n19424 & n19582;
  assign n19584 = n19414 & ~n19583;
  assign n19585 = ~n19581 & ~n19584;
  assign n19586 = n19460 & ~n19467;
  assign n19587 = n19409 & ~n19586;
  assign n19588 = ~n19438 & n19573;
  assign n19589 = ~n19444 & n19588;
  assign n19590 = n19432 & ~n19589;
  assign n19591 = ~n19587 & ~n19590;
  assign n19592 = n19585 & n19591;
  assign n19593 = n19579 & n19592;
  assign n19594 = ~n19574 & n19593;
  assign n19595 = n19431 & n19594;
  assign n19596 = ~n19572 & n19595;
  assign n19597 = n19422 & n19596;
  assign n19598 = n19597 ^ n16525;
  assign n19599 = n19598 ^ x64;
  assign n19600 = ~n19571 & ~n19599;
  assign n19601 = n18821 ^ x77;
  assign n19602 = n18367 ^ x68;
  assign n19603 = n19601 & n19602;
  assign n19604 = ~n17810 & n17824;
  assign n19605 = n17812 & n17844;
  assign n19606 = ~n19604 & ~n19605;
  assign n19607 = n17833 ^ n17714;
  assign n19608 = n19607 ^ n17833;
  assign n19609 = n17833 ^ n17821;
  assign n19610 = ~n19608 & n19609;
  assign n19611 = n19610 ^ n17833;
  assign n19612 = ~n17713 & ~n19611;
  assign n19613 = n19606 & ~n19612;
  assign n19614 = n19613 ^ n16185;
  assign n19615 = n19614 ^ x117;
  assign n19616 = n18142 ^ x94;
  assign n19617 = n19615 & ~n19616;
  assign n19618 = n17042 & n17063;
  assign n19619 = n17019 & ~n17039;
  assign n19620 = ~n19618 & ~n19619;
  assign n19621 = n17050 & n17059;
  assign n19622 = ~n17036 & n19621;
  assign n19623 = n19622 ^ n17064;
  assign n19624 = n19623 ^ n17064;
  assign n19625 = n17064 ^ n16776;
  assign n19626 = n19625 ^ n17064;
  assign n19627 = ~n19624 & n19626;
  assign n19628 = n19627 ^ n17064;
  assign n19629 = ~n16807 & ~n19628;
  assign n19630 = n19629 ^ n17064;
  assign n19631 = n19620 & n19630;
  assign n19632 = n17068 ^ n17059;
  assign n19633 = n17068 ^ n17019;
  assign n19634 = n19633 ^ n17019;
  assign n19635 = n17042 ^ n17019;
  assign n19636 = n19634 & ~n19635;
  assign n19637 = n19636 ^ n17019;
  assign n19638 = n19632 & n19637;
  assign n19639 = n19638 ^ n17059;
  assign n19640 = n19057 & n19639;
  assign n19641 = n19640 ^ n19246;
  assign n19642 = n19641 ^ n19246;
  assign n19643 = n19246 ^ n17026;
  assign n19644 = n19643 ^ n19246;
  assign n19645 = ~n19642 & ~n19644;
  assign n19646 = n19645 ^ n19246;
  assign n19647 = ~n16808 & ~n19646;
  assign n19648 = n19647 ^ n19246;
  assign n19649 = n19631 & n19648;
  assign n19650 = n19244 & n19649;
  assign n19651 = n17034 & n19650;
  assign n19652 = ~n19045 & n19651;
  assign n19653 = n17024 & n19652;
  assign n19654 = n19653 ^ n16206;
  assign n19655 = n19654 ^ x75;
  assign n19656 = n18938 ^ x100;
  assign n19657 = n19655 & n19656;
  assign n19658 = n19617 & n19657;
  assign n19659 = n19603 & n19658;
  assign n19660 = ~n19615 & n19616;
  assign n19661 = ~n19655 & n19656;
  assign n19662 = n19660 & n19661;
  assign n19663 = ~n19615 & ~n19616;
  assign n19664 = n19657 & n19663;
  assign n19665 = ~n19662 & ~n19664;
  assign n19666 = n19603 & ~n19665;
  assign n19667 = ~n19659 & ~n19666;
  assign n19668 = ~n19601 & ~n19602;
  assign n19669 = n19655 & ~n19656;
  assign n19670 = n19663 & n19669;
  assign n19671 = n19615 & n19616;
  assign n19672 = ~n19655 & ~n19656;
  assign n19673 = n19671 & n19672;
  assign n19674 = ~n19670 & ~n19673;
  assign n19675 = n19668 & ~n19674;
  assign n19676 = n19601 & ~n19602;
  assign n19677 = n19669 & n19671;
  assign n19678 = n19661 & n19671;
  assign n19679 = ~n19658 & ~n19678;
  assign n19680 = ~n19670 & n19679;
  assign n19681 = n19660 & n19669;
  assign n19682 = n19663 & n19672;
  assign n19683 = ~n19673 & ~n19682;
  assign n19684 = ~n19681 & n19683;
  assign n19685 = n19680 & n19684;
  assign n19686 = ~n19677 & n19685;
  assign n19687 = ~n19662 & n19686;
  assign n19688 = n19676 & n19687;
  assign n19689 = ~n19675 & ~n19688;
  assign n19690 = n19617 & n19661;
  assign n19691 = n19603 & n19690;
  assign n19692 = ~n19601 & n19602;
  assign n19693 = ~n19664 & ~n19678;
  assign n19694 = n19661 & n19663;
  assign n19695 = ~n19673 & ~n19694;
  assign n19696 = n19693 & n19695;
  assign n19697 = ~n19681 & n19696;
  assign n19698 = n19692 & ~n19697;
  assign n19699 = ~n19691 & ~n19698;
  assign n19700 = ~n19668 & ~n19692;
  assign n19701 = n19617 & n19669;
  assign n19702 = n19660 & n19672;
  assign n19703 = ~n19701 & ~n19702;
  assign n19704 = ~n19700 & ~n19703;
  assign n19705 = ~n19603 & ~n19670;
  assign n19706 = ~n19677 & ~n19682;
  assign n19707 = n19674 & n19706;
  assign n19708 = ~n19705 & ~n19707;
  assign n19709 = n19708 ^ n19601;
  assign n19710 = n19709 ^ n19708;
  assign n19711 = n19657 & n19660;
  assign n19712 = ~n19658 & ~n19711;
  assign n19713 = ~n19690 & n19712;
  assign n19714 = ~n19662 & n19713;
  assign n19715 = n19714 ^ n19708;
  assign n19716 = n19715 ^ n19708;
  assign n19717 = ~n19710 & ~n19716;
  assign n19718 = n19717 ^ n19708;
  assign n19719 = ~n19602 & n19718;
  assign n19720 = n19719 ^ n19708;
  assign n19721 = ~n19704 & ~n19720;
  assign n19722 = n19699 & n19721;
  assign n19723 = n19689 & n19722;
  assign n19724 = n19667 & n19723;
  assign n19725 = n19724 ^ n16311;
  assign n19726 = n19725 ^ x115;
  assign n19727 = ~n18968 & ~n18996;
  assign n19728 = n18940 & ~n19727;
  assign n19729 = n18953 & n18984;
  assign n19730 = n18951 & n18953;
  assign n19731 = ~n18964 & ~n19730;
  assign n19732 = n18971 & ~n18996;
  assign n19733 = n18944 & ~n19732;
  assign n19734 = n18940 & n18967;
  assign n19735 = ~n18955 & ~n18979;
  assign n19736 = ~n18940 & n19735;
  assign n19737 = ~n18962 & n19736;
  assign n19738 = ~n18943 & ~n18998;
  assign n19739 = n18980 & n19738;
  assign n19740 = ~n18944 & n19739;
  assign n19741 = ~n19737 & ~n19740;
  assign n19742 = n18897 & n19741;
  assign n19743 = n18970 & n18980;
  assign n19744 = n18958 & n19743;
  assign n19745 = n18953 & ~n19744;
  assign n19746 = n18965 ^ n18961;
  assign n19747 = n18961 ^ n18940;
  assign n19748 = n19747 ^ n18940;
  assign n19749 = n18823 & n18942;
  assign n19750 = ~n18978 & ~n19749;
  assign n19751 = ~n18984 & n19750;
  assign n19752 = ~n18996 & n19751;
  assign n19753 = n19752 ^ n18940;
  assign n19754 = n19748 & n19753;
  assign n19755 = n19754 ^ n18940;
  assign n19756 = n19746 & ~n19755;
  assign n19757 = n19756 ^ n18965;
  assign n19758 = ~n19745 & ~n19757;
  assign n19759 = ~n19742 & n19758;
  assign n19760 = ~n19734 & n19759;
  assign n19761 = ~n19733 & n19760;
  assign n19762 = n19731 & n19761;
  assign n19763 = ~n19729 & n19762;
  assign n19764 = ~n19728 & n19763;
  assign n19765 = ~n18949 & n19764;
  assign n19766 = n19765 ^ n15880;
  assign n19767 = n19766 ^ x96;
  assign n19768 = n19726 & n19767;
  assign n19769 = n19014 & ~n19096;
  assign n19770 = ~n19016 & n19078;
  assign n19771 = ~n19113 & ~n19770;
  assign n19772 = n19076 & n19088;
  assign n19773 = ~n19119 & ~n19772;
  assign n19774 = n19771 & n19773;
  assign n19775 = n19769 & ~n19774;
  assign n19776 = ~n19014 & ~n19096;
  assign n19777 = n19076 & n19112;
  assign n19778 = ~n19092 & n19115;
  assign n19779 = ~n19770 & n19778;
  assign n19780 = ~n19777 & n19779;
  assign n19781 = n19776 & ~n19780;
  assign n19782 = ~n19775 & ~n19781;
  assign n19783 = ~n19076 & n19084;
  assign n19784 = ~n19080 & ~n19783;
  assign n19785 = n19014 & ~n19784;
  assign n19786 = ~n19014 & n19096;
  assign n19787 = n19778 & n19784;
  assign n19788 = n19786 & n19787;
  assign n19789 = n19014 & n19096;
  assign n19790 = n19076 & n19099;
  assign n19791 = ~n19102 & ~n19790;
  assign n19792 = ~n19101 & n19791;
  assign n19793 = ~n19777 & n19792;
  assign n19794 = ~n19100 & n19793;
  assign n19795 = n19789 & ~n19794;
  assign n19796 = ~n19788 & ~n19795;
  assign n19797 = ~n19785 & n19796;
  assign n19798 = n19782 & n19797;
  assign n19799 = n19798 ^ n16126;
  assign n19800 = n19799 ^ x97;
  assign n19801 = n19285 & n19299;
  assign n19802 = n19279 & n19326;
  assign n19803 = ~n19801 & ~n19802;
  assign n19804 = n19294 & n19305;
  assign n19805 = n19279 & n19804;
  assign n19806 = ~n19284 & ~n19805;
  assign n19807 = n19278 ^ n19241;
  assign n19808 = n19306 & ~n19807;
  assign n19809 = n19293 & ~n19327;
  assign n19810 = ~n19808 & ~n19809;
  assign n19811 = n19279 & ~n19320;
  assign n19812 = ~n19295 & ~n19307;
  assign n19813 = n19285 & ~n19812;
  assign n19814 = ~n19240 & n19302;
  assign n19815 = ~n19326 & n19814;
  assign n19816 = ~n19310 & n19815;
  assign n19817 = n19283 & ~n19816;
  assign n19818 = ~n19289 & n19302;
  assign n19819 = n19279 & ~n19818;
  assign n19820 = ~n19319 & ~n19804;
  assign n19821 = ~n19318 & n19820;
  assign n19822 = ~n19282 & n19821;
  assign n19823 = n19285 & ~n19822;
  assign n19824 = ~n19287 & ~n19293;
  assign n19825 = ~n19240 & n19312;
  assign n19826 = ~n19824 & ~n19825;
  assign n19827 = ~n19823 & ~n19826;
  assign n19828 = ~n19819 & n19827;
  assign n19829 = ~n19817 & n19828;
  assign n19830 = ~n19813 & n19829;
  assign n19831 = ~n19811 & n19830;
  assign n19832 = n19810 & n19831;
  assign n19833 = n19806 & n19832;
  assign n19834 = n19803 & n19833;
  assign n19835 = n19834 ^ n15397;
  assign n19836 = n19835 ^ x106;
  assign n19837 = n19800 & ~n19836;
  assign n19838 = n19768 & n19837;
  assign n19839 = n19600 & n19838;
  assign n19840 = n19571 & n19599;
  assign n19841 = ~n19726 & n19767;
  assign n19842 = ~n19800 & ~n19836;
  assign n19843 = n19841 & n19842;
  assign n19844 = n19840 & n19843;
  assign n19845 = ~n19571 & n19599;
  assign n19846 = ~n19726 & ~n19767;
  assign n19847 = n19842 & n19846;
  assign n19848 = n19845 & n19847;
  assign n19849 = ~n19844 & ~n19848;
  assign n19850 = ~n19839 & n19849;
  assign n19851 = n19571 & ~n19599;
  assign n19852 = n19800 & n19836;
  assign n19853 = n19768 & n19852;
  assign n19854 = n19846 & n19852;
  assign n19855 = ~n19853 & ~n19854;
  assign n19856 = n19851 & ~n19855;
  assign n19857 = n19845 & n19854;
  assign n19858 = ~n19800 & n19836;
  assign n19859 = n19846 & n19858;
  assign n19860 = n19726 & ~n19767;
  assign n19861 = n19852 & n19860;
  assign n19862 = ~n19859 & ~n19861;
  assign n19863 = n19840 & ~n19862;
  assign n19864 = ~n19857 & ~n19863;
  assign n19865 = n19838 & n19840;
  assign n19866 = n19837 & n19846;
  assign n19867 = ~n19600 & ~n19840;
  assign n19868 = n19866 & ~n19867;
  assign n19869 = ~n19865 & ~n19868;
  assign n19870 = ~n19843 & ~n19847;
  assign n19871 = n19851 & ~n19870;
  assign n19872 = n19841 & n19858;
  assign n19873 = n19845 & n19872;
  assign n19874 = n19599 ^ n19571;
  assign n19875 = n19837 & n19860;
  assign n19876 = n19842 & n19860;
  assign n19877 = ~n19875 & ~n19876;
  assign n19878 = n19874 & ~n19877;
  assign n19879 = ~n19873 & ~n19878;
  assign n19880 = n19858 & n19860;
  assign n19881 = ~n19872 & ~n19880;
  assign n19882 = ~n19867 & ~n19881;
  assign n19883 = n19837 & n19841;
  assign n19884 = ~n19571 & n19883;
  assign n19885 = n19768 & n19858;
  assign n19886 = n19768 & n19842;
  assign n19887 = ~n19861 & ~n19886;
  assign n19888 = ~n19885 & n19887;
  assign n19889 = n19600 & ~n19888;
  assign n19890 = ~n19884 & ~n19889;
  assign n19891 = n19841 & n19852;
  assign n19892 = ~n19885 & ~n19891;
  assign n19893 = n19892 ^ n19853;
  assign n19894 = n19893 ^ n19853;
  assign n19895 = n19853 ^ n19600;
  assign n19896 = n19895 ^ n19853;
  assign n19897 = ~n19894 & ~n19896;
  assign n19898 = n19897 ^ n19853;
  assign n19899 = ~n19840 & n19898;
  assign n19900 = n19899 ^ n19853;
  assign n19901 = n19890 & ~n19900;
  assign n19902 = ~n19882 & n19901;
  assign n19903 = n19879 & n19902;
  assign n19904 = ~n19871 & n19903;
  assign n19905 = n19869 & n19904;
  assign n19906 = n19864 & n19905;
  assign n19907 = ~n19856 & n19906;
  assign n19908 = n19850 & n19907;
  assign n19909 = n19908 ^ n16757;
  assign n19910 = ~n18732 & n18764;
  assign n19911 = n18764 & n18771;
  assign n19912 = ~n18737 & ~n18744;
  assign n19913 = n18748 & ~n19912;
  assign n19914 = ~n19911 & ~n19913;
  assign n19915 = ~n18732 & n18748;
  assign n19916 = ~n18765 & ~n18775;
  assign n19917 = n18761 & n19916;
  assign n19918 = ~n18754 & n19917;
  assign n19919 = n18764 & ~n19918;
  assign n19920 = ~n18758 & ~n18772;
  assign n19921 = ~n18771 & n19920;
  assign n19922 = n18733 & ~n19921;
  assign n19923 = n18524 ^ n18464;
  assign n19924 = n19923 ^ n18545;
  assign n19925 = n18487 & ~n19924;
  assign n19926 = ~n18740 & n19925;
  assign n19927 = n18761 & ~n18771;
  assign n19928 = ~n18751 & n19927;
  assign n19929 = n19928 ^ n18726;
  assign n19930 = n19929 ^ n19928;
  assign n19931 = ~n18759 & n18773;
  assign n19932 = ~n18754 & n19931;
  assign n19933 = n19932 ^ n19928;
  assign n19934 = ~n19930 & n19933;
  assign n19935 = n19934 ^ n19928;
  assign n19936 = ~n18578 & ~n19935;
  assign n19937 = ~n19926 & ~n19936;
  assign n19938 = ~n19922 & n19937;
  assign n19939 = ~n19919 & n19938;
  assign n19940 = ~n19915 & n19939;
  assign n19941 = n19914 & n19940;
  assign n19942 = ~n18752 & n19941;
  assign n19943 = ~n19910 & n19942;
  assign n19944 = n19943 ^ n17338;
  assign n19945 = n19838 & n19851;
  assign n19946 = ~n19853 & ~n19872;
  assign n19947 = n19845 & ~n19946;
  assign n19948 = ~n19945 & ~n19947;
  assign n19949 = n19600 & ~n19862;
  assign n19950 = n19840 & n19847;
  assign n19951 = n19883 ^ n19599;
  assign n19952 = n19951 ^ n19883;
  assign n19953 = n19883 ^ n19866;
  assign n19954 = n19952 & n19953;
  assign n19955 = n19954 ^ n19883;
  assign n19956 = n19874 & n19955;
  assign n19957 = ~n19950 & ~n19956;
  assign n19958 = ~n19867 & ~n19892;
  assign n19959 = ~n19876 & n19881;
  assign n19960 = n19851 & ~n19959;
  assign n19961 = ~n19958 & ~n19960;
  assign n19962 = n19843 & n19867;
  assign n19963 = ~n19859 & ~n19883;
  assign n19964 = n19845 & ~n19963;
  assign n19965 = ~n19962 & ~n19964;
  assign n19966 = n19877 ^ n19599;
  assign n19967 = n19966 ^ n19877;
  assign n19968 = n19886 ^ n19877;
  assign n19969 = n19968 ^ n19877;
  assign n19970 = n19967 & n19969;
  assign n19971 = n19970 ^ n19877;
  assign n19972 = n19571 & ~n19971;
  assign n19973 = n19972 ^ n19877;
  assign n19974 = n19965 & n19973;
  assign n19975 = n19961 & n19974;
  assign n19976 = n19957 & n19975;
  assign n19977 = ~n19839 & n19976;
  assign n19978 = ~n19863 & n19977;
  assign n19979 = ~n19949 & n19978;
  assign n19980 = n19869 & n19979;
  assign n19981 = n19948 & n19980;
  assign n19982 = ~n19856 & n19981;
  assign n19983 = n19982 ^ n18821;
  assign n19984 = n19677 & n19692;
  assign n19985 = n19617 & n19672;
  assign n19986 = ~n19681 & ~n19985;
  assign n19987 = n19603 & ~n19986;
  assign n19988 = ~n19984 & ~n19987;
  assign n19989 = n19692 & n19711;
  assign n19990 = ~n19680 & n19692;
  assign n19991 = n19602 & n19682;
  assign n19992 = n19668 & n19687;
  assign n19993 = ~n19991 & ~n19992;
  assign n19994 = ~n19676 & ~n19692;
  assign n19995 = ~n19695 & ~n19994;
  assign n19996 = ~n19678 & ~n19702;
  assign n19997 = n19996 ^ n19602;
  assign n19998 = n19997 ^ n19996;
  assign n19999 = ~n19702 & ~n19985;
  assign n20000 = ~n19662 & n19999;
  assign n20001 = n19712 & n20000;
  assign n20002 = ~n19670 & n20001;
  assign n20003 = n20002 ^ n19996;
  assign n20004 = ~n19998 & n20003;
  assign n20005 = n20004 ^ n19996;
  assign n20006 = n19601 & ~n20005;
  assign n20007 = ~n19995 & ~n20006;
  assign n20008 = n19993 & n20007;
  assign n20009 = ~n19990 & n20008;
  assign n20010 = ~n19989 & n20009;
  assign n20011 = n19988 & n20010;
  assign n20012 = n19667 & n20011;
  assign n20013 = n20012 ^ n16974;
  assign n20014 = n19944 ^ x69;
  assign n20015 = ~n18939 & n18978;
  assign n20016 = ~n18948 & n19732;
  assign n20017 = n18961 & ~n20016;
  assign n20018 = ~n18967 & ~n18969;
  assign n20019 = ~n18998 & n19736;
  assign n20020 = ~n18948 & n18958;
  assign n20021 = ~n18944 & n20020;
  assign n20022 = ~n20019 & ~n20021;
  assign n20023 = n20018 & ~n20022;
  assign n20024 = n20023 ^ n18939;
  assign n20025 = n20024 ^ n20023;
  assign n20026 = n18981 & n19738;
  assign n20027 = n20026 ^ n20023;
  assign n20028 = n20027 ^ n20023;
  assign n20029 = n20025 & ~n20028;
  assign n20030 = n20029 ^ n20023;
  assign n20031 = ~n18897 & ~n20030;
  assign n20032 = n20031 ^ n20023;
  assign n20033 = ~n20017 & n20032;
  assign n20034 = ~n20015 & n20033;
  assign n20035 = n19731 & n20034;
  assign n20036 = n18960 & n20035;
  assign n20037 = ~n19729 & n20036;
  assign n20038 = ~n19728 & n20037;
  assign n20039 = n18946 & n20038;
  assign n20040 = n20039 ^ n17014;
  assign n20041 = n20040 ^ x91;
  assign n20042 = ~n20014 & n20041;
  assign n20043 = n18388 & n18395;
  assign n20044 = n18383 & n18422;
  assign n20045 = ~n20043 & ~n20044;
  assign n20046 = n18144 & ~n18380;
  assign n20047 = n20045 & ~n20046;
  assign n20048 = ~n18397 & ~n18430;
  assign n20049 = ~n18103 & ~n20048;
  assign n20050 = ~n18374 & n18395;
  assign n20051 = ~n20049 & ~n20050;
  assign n20052 = ~n18397 & ~n18417;
  assign n20053 = n18376 & ~n20052;
  assign n20054 = n18144 & ~n18406;
  assign n20055 = ~n20053 & ~n20054;
  assign n20056 = ~n18396 & ~n18405;
  assign n20057 = ~n18391 & n20056;
  assign n20058 = ~n18422 & n20057;
  assign n20059 = ~n18385 & n18424;
  assign n20060 = ~n18376 & n20059;
  assign n20061 = ~n20058 & ~n20060;
  assign n20062 = n20061 ^ n18103;
  assign n20063 = n20062 ^ n20061;
  assign n20064 = ~n18401 & ~n18417;
  assign n20065 = ~n18410 & n20064;
  assign n20066 = n20065 ^ n20061;
  assign n20067 = n20066 ^ n20061;
  assign n20068 = ~n20063 & ~n20067;
  assign n20069 = n20068 ^ n20061;
  assign n20070 = ~n18143 & n20069;
  assign n20071 = n20070 ^ n20061;
  assign n20072 = n20055 & ~n20071;
  assign n20073 = n20051 & n20072;
  assign n20074 = n20047 & n20073;
  assign n20075 = n18394 & n20074;
  assign n20076 = n18382 & n20075;
  assign n20077 = n20076 ^ n18183;
  assign n20078 = n20077 ^ x67;
  assign n20079 = n17991 & n18019;
  assign n20080 = n17088 & ~n18039;
  assign n20081 = ~n20079 & ~n20080;
  assign n20082 = n18011 & ~n18034;
  assign n20083 = ~n18012 & ~n18033;
  assign n20084 = n18028 & n20083;
  assign n20085 = ~n18024 & n20084;
  assign n20086 = n18019 & ~n20085;
  assign n20087 = ~n20082 & ~n20086;
  assign n20088 = ~n18020 & n20083;
  assign n20089 = ~n17991 & n20088;
  assign n20090 = ~n18002 & n20089;
  assign n20091 = n17088 & ~n20090;
  assign n20092 = ~n18027 & n18030;
  assign n20093 = ~n18002 & n20092;
  assign n20094 = n18011 & ~n20093;
  assign n20095 = n17692 ^ n17483;
  assign n20096 = n20095 ^ n17849;
  assign n20097 = ~n17985 & ~n20096;
  assign n20098 = n18035 & ~n20097;
  assign n20099 = n18001 & ~n20098;
  assign n20100 = ~n20094 & ~n20099;
  assign n20101 = ~n20091 & n20100;
  assign n20102 = n20087 & n20101;
  assign n20103 = ~n18056 & n20102;
  assign n20104 = n20081 & n20103;
  assign n20105 = ~n17988 & n20104;
  assign n20106 = n20105 ^ n17160;
  assign n20107 = n20106 ^ x92;
  assign n20108 = ~n20078 & n20107;
  assign n20109 = ~n19121 & n19776;
  assign n20110 = ~n19133 & n19786;
  assign n20111 = ~n20109 & ~n20110;
  assign n20112 = n19095 & n19769;
  assign n20113 = ~n19107 & n19789;
  assign n20114 = ~n20112 & ~n20113;
  assign n20115 = n20111 & n20114;
  assign n20116 = n20115 ^ n18154;
  assign n20117 = n20116 ^ x109;
  assign n20118 = ~n19424 & ~n19444;
  assign n20119 = n19432 & ~n20118;
  assign n20120 = n19412 & n19414;
  assign n20121 = n19409 & ~n19478;
  assign n20122 = ~n20120 & ~n20121;
  assign n20123 = ~n20119 & n20122;
  assign n20124 = n19417 & n19432;
  assign n20125 = n19409 & ~n19441;
  assign n20126 = ~n20124 & ~n20125;
  assign n20127 = ~n19446 & ~n19458;
  assign n20128 = ~n19433 & ~n20127;
  assign n20129 = n19352 & ~n20118;
  assign n20130 = ~n19418 & ~n19427;
  assign n20131 = n19588 & n20130;
  assign n20132 = ~n19457 & n20131;
  assign n20133 = n19414 & ~n20132;
  assign n20134 = ~n20129 & ~n20133;
  assign n20135 = ~n20128 & n20134;
  assign n20136 = n20126 & n20135;
  assign n20137 = ~n19482 & n20136;
  assign n20138 = n19430 & n20137;
  assign n20139 = n19579 & n20138;
  assign n20140 = ~n19574 & n20139;
  assign n20141 = n20123 & n20140;
  assign n20142 = ~n19572 & n20141;
  assign n20143 = n20142 ^ n16806;
  assign n20144 = n20143 ^ x86;
  assign n20145 = ~n20117 & n20144;
  assign n20146 = n20108 & n20145;
  assign n20147 = n20117 & ~n20144;
  assign n20148 = n20108 & n20147;
  assign n20149 = ~n20146 & ~n20148;
  assign n20150 = n20042 & ~n20149;
  assign n20151 = n20014 & n20041;
  assign n20152 = n20078 & n20107;
  assign n20153 = ~n20117 & ~n20144;
  assign n20154 = n20152 & n20153;
  assign n20155 = n20117 & n20144;
  assign n20156 = n20108 & n20155;
  assign n20157 = n20147 & n20152;
  assign n20158 = ~n20156 & ~n20157;
  assign n20159 = ~n20154 & n20158;
  assign n20160 = n20151 & ~n20159;
  assign n20161 = n20014 & ~n20041;
  assign n20162 = ~n20148 & ~n20156;
  assign n20163 = n20161 & ~n20162;
  assign n20164 = n20078 & ~n20107;
  assign n20165 = n20155 & n20164;
  assign n20166 = ~n20078 & ~n20107;
  assign n20167 = n20147 & n20166;
  assign n20168 = ~n20165 & ~n20167;
  assign n20169 = ~n20146 & n20168;
  assign n20170 = n20151 & ~n20169;
  assign n20171 = ~n20163 & ~n20170;
  assign n20172 = n20152 & n20155;
  assign n20173 = ~n20154 & ~n20172;
  assign n20174 = n20145 & n20166;
  assign n20175 = n20147 & n20164;
  assign n20176 = ~n20174 & ~n20175;
  assign n20177 = n20173 & n20176;
  assign n20178 = n20177 ^ n20042;
  assign n20179 = n20177 ^ n20161;
  assign n20180 = n20179 ^ n20161;
  assign n20181 = n20145 & n20164;
  assign n20182 = ~n20167 & ~n20181;
  assign n20183 = n20182 ^ n20161;
  assign n20184 = n20180 & n20183;
  assign n20185 = n20184 ^ n20161;
  assign n20186 = ~n20178 & n20185;
  assign n20187 = n20186 ^ n20042;
  assign n20188 = n20171 & ~n20187;
  assign n20189 = n20155 & n20166;
  assign n20190 = n20153 & n20166;
  assign n20191 = ~n20189 & ~n20190;
  assign n20192 = ~n20151 & ~n20161;
  assign n20193 = ~n20191 & ~n20192;
  assign n20194 = ~n20014 & ~n20041;
  assign n20195 = n20144 ^ n20107;
  assign n20196 = n20117 ^ n20107;
  assign n20197 = n20196 ^ n20107;
  assign n20198 = n20195 & n20197;
  assign n20199 = n20198 ^ n20107;
  assign n20200 = n20107 ^ n20078;
  assign n20201 = n20200 ^ n20144;
  assign n20202 = n20201 ^ n20107;
  assign n20203 = n20202 ^ n20117;
  assign n20204 = n20203 ^ n20144;
  assign n20205 = ~n20199 & ~n20204;
  assign n20206 = n20205 ^ n20201;
  assign n20207 = n20194 & n20206;
  assign n20208 = ~n20193 & ~n20207;
  assign n20209 = n20188 & n20208;
  assign n20210 = ~n20160 & n20209;
  assign n20211 = ~n20150 & n20210;
  assign n20212 = n20211 ^ n18254;
  assign n20213 = n19657 & n19671;
  assign n20214 = ~n19694 & ~n20213;
  assign n20215 = n19713 & n20214;
  assign n20216 = n19684 & n20215;
  assign n20217 = n19668 & ~n20216;
  assign n20218 = ~n19990 & ~n20217;
  assign n20219 = n19676 & ~n19693;
  assign n20220 = ~n19677 & n20000;
  assign n20221 = ~n19994 & ~n20220;
  assign n20222 = ~n19701 & ~n20213;
  assign n20223 = ~n19690 & n20222;
  assign n20224 = n19684 & n20223;
  assign n20225 = n19693 & n20224;
  assign n20226 = n19603 & ~n20225;
  assign n20227 = ~n20221 & ~n20226;
  assign n20228 = ~n20219 & n20227;
  assign n20229 = n20218 & n20228;
  assign n20230 = n19701 ^ n19676;
  assign n20231 = n19701 ^ n19692;
  assign n20232 = n20231 ^ n19692;
  assign n20233 = n19692 ^ n19670;
  assign n20234 = ~n20232 & ~n20233;
  assign n20235 = n20234 ^ n19692;
  assign n20236 = n20230 & n20235;
  assign n20237 = n20236 ^ n19676;
  assign n20238 = n20229 & ~n20237;
  assign n20239 = n20238 ^ n17550;
  assign n20240 = n20151 & n20174;
  assign n20241 = n20108 & n20153;
  assign n20242 = n20194 & n20241;
  assign n20243 = ~n20240 & ~n20242;
  assign n20244 = n20173 & ~n20174;
  assign n20245 = n20194 & ~n20244;
  assign n20246 = n20145 & n20152;
  assign n20247 = n20151 & n20246;
  assign n20248 = n20194 & n20246;
  assign n20249 = ~n20042 & ~n20161;
  assign n20250 = n20175 & ~n20249;
  assign n20251 = ~n20154 & ~n20156;
  assign n20252 = ~n20146 & n20251;
  assign n20253 = n20042 & ~n20252;
  assign n20254 = ~n20250 & ~n20253;
  assign n20255 = n20148 & n20194;
  assign n20256 = n20146 & ~n20192;
  assign n20257 = ~n20255 & ~n20256;
  assign n20258 = ~n20158 & n20161;
  assign n20259 = n20153 & n20164;
  assign n20260 = ~n20241 & ~n20259;
  assign n20261 = ~n20157 & n20260;
  assign n20262 = n20151 & ~n20261;
  assign n20263 = ~n20258 & ~n20262;
  assign n20264 = n20257 & n20263;
  assign n20265 = n20254 & n20264;
  assign n20266 = ~n20189 & ~n20259;
  assign n20267 = ~n20181 & ~n20190;
  assign n20268 = n20266 & n20267;
  assign n20269 = n20268 ^ n20249;
  assign n20270 = n20269 ^ n20268;
  assign n20271 = n20268 ^ n20168;
  assign n20272 = n20270 & n20271;
  assign n20273 = n20272 ^ n20268;
  assign n20274 = n20265 & n20273;
  assign n20275 = ~n20248 & n20274;
  assign n20276 = ~n20247 & n20275;
  assign n20277 = ~n20245 & n20276;
  assign n20278 = n20243 & n20277;
  assign n20279 = n20278 ^ n19401;
  assign n20280 = ~n18405 & n18424;
  assign n20281 = n18144 & ~n20280;
  assign n20282 = ~n18379 & n18398;
  assign n20283 = n18383 & ~n20282;
  assign n20284 = ~n20281 & ~n20283;
  assign n20285 = ~n18103 & n18417;
  assign n20286 = ~n18377 & n20048;
  assign n20287 = n18395 & ~n20286;
  assign n20288 = ~n20285 & ~n20287;
  assign n20289 = ~n18373 & n18380;
  assign n20290 = n18376 & ~n20289;
  assign n20291 = ~n18385 & ~n18404;
  assign n20292 = ~n18391 & n20291;
  assign n20293 = n18376 & ~n20292;
  assign n20294 = ~n18385 & n20280;
  assign n20295 = n18383 & ~n20294;
  assign n20296 = ~n20293 & ~n20295;
  assign n20297 = n18143 ^ n18103;
  assign n20298 = n18296 & n18387;
  assign n20299 = ~n18401 & ~n20298;
  assign n20300 = ~n18422 & n20299;
  assign n20301 = n20300 ^ n18143;
  assign n20302 = n20301 ^ n20300;
  assign n20303 = ~n18417 & n20282;
  assign n20304 = n20303 ^ n20300;
  assign n20305 = ~n20302 & n20304;
  assign n20306 = n20305 ^ n20300;
  assign n20307 = n20297 & ~n20306;
  assign n20308 = n20296 & ~n20307;
  assign n20309 = ~n20290 & n20308;
  assign n20310 = n20288 & n20309;
  assign n20311 = n20284 & n20310;
  assign n20312 = n18412 & n20311;
  assign n20313 = n20312 ^ n17798;
  assign n20314 = ~n19774 & n19776;
  assign n20315 = n19769 & n19780;
  assign n20316 = ~n20314 & ~n20315;
  assign n20317 = ~n19778 & n19789;
  assign n20318 = n19786 & ~n19794;
  assign n20319 = ~n20317 & ~n20318;
  assign n20320 = n20316 & n20319;
  assign n20321 = n19784 & n20320;
  assign n20322 = n20321 ^ n16775;
  assign n20323 = n20322 ^ x102;
  assign n20324 = n20143 ^ x116;
  assign n20325 = n20323 & n20324;
  assign n20327 = n18732 & n18739;
  assign n20328 = n18727 & ~n20327;
  assign n20329 = ~n18547 & ~n18751;
  assign n20330 = n18748 & ~n20329;
  assign n20331 = ~n20328 & ~n20330;
  assign n20332 = ~n18730 & n19916;
  assign n20333 = n18733 & ~n20332;
  assign n20334 = ~n18760 & n19920;
  assign n20335 = ~n18754 & n20334;
  assign n20336 = n18764 & ~n20335;
  assign n20337 = ~n18751 & ~n18754;
  assign n20338 = n18727 & ~n20337;
  assign n20339 = n18764 & ~n19912;
  assign n20340 = n18748 & ~n19921;
  assign n20341 = ~n20339 & ~n20340;
  assign n20342 = ~n18759 & ~n18775;
  assign n20343 = n18727 & ~n20342;
  assign n20344 = n18733 & ~n20334;
  assign n20345 = ~n20343 & ~n20344;
  assign n20346 = n20341 & n20345;
  assign n20347 = ~n20338 & n20346;
  assign n20348 = n18757 & n20347;
  assign n20349 = ~n19910 & n20348;
  assign n20350 = ~n20336 & n20349;
  assign n20351 = ~n20333 & n20350;
  assign n20352 = n20331 & n20351;
  assign n20353 = ~n19913 & n20352;
  assign n20354 = n20353 ^ n16949;
  assign n20355 = n20354 ^ x84;
  assign n20326 = n20013 ^ x126;
  assign n20356 = n20355 ^ n20326;
  assign n20357 = n19290 & ~n19300;
  assign n20358 = n19279 & ~n20357;
  assign n20359 = n19283 & ~n19323;
  assign n20360 = ~n20358 & ~n20359;
  assign n20361 = ~n19306 & ~n19310;
  assign n20362 = ~n19307 & n20361;
  assign n20363 = ~n19293 & n20362;
  assign n20364 = n19279 & ~n20361;
  assign n20365 = n19820 & ~n20364;
  assign n20366 = n19309 & n20365;
  assign n20367 = ~n20363 & ~n20366;
  assign n20368 = n19241 & n20367;
  assign n20372 = ~n19301 & ~n19310;
  assign n20369 = ~n19318 & ~n19326;
  assign n20370 = n19309 & n20369;
  assign n20371 = ~n19300 & n20370;
  assign n20373 = n20372 ^ n20371;
  assign n20374 = n20373 ^ n20372;
  assign n20375 = n20372 ^ n19278;
  assign n20376 = n20375 ^ n20372;
  assign n20377 = ~n20374 & n20376;
  assign n20378 = n20377 ^ n20372;
  assign n20379 = n19807 & ~n20378;
  assign n20380 = n20379 ^ n20372;
  assign n20381 = ~n20368 & n20380;
  assign n20382 = n20360 & n20381;
  assign n20383 = ~n19297 & n20382;
  assign n20384 = n19292 & n20383;
  assign n20385 = ~n19280 & n20384;
  assign n20386 = n19803 & n20385;
  assign n20387 = n20386 ^ n16840;
  assign n20388 = n20387 ^ x70;
  assign n20389 = n20040 ^ x85;
  assign n20390 = ~n20388 & ~n20389;
  assign n20391 = ~n20356 & n20390;
  assign n20392 = n20325 & n20391;
  assign n20393 = ~n20323 & ~n20324;
  assign n20394 = n20326 & ~n20355;
  assign n20395 = n20388 & n20389;
  assign n20396 = n20394 & n20395;
  assign n20397 = n20393 & n20396;
  assign n20398 = ~n20326 & n20355;
  assign n20399 = n20395 & n20398;
  assign n20400 = n20325 & n20399;
  assign n20401 = ~n20397 & ~n20400;
  assign n20402 = n20323 & ~n20324;
  assign n20403 = n20396 & n20402;
  assign n20404 = ~n20388 & n20389;
  assign n20405 = n20398 & n20404;
  assign n20406 = n20326 & n20355;
  assign n20407 = n20395 & n20406;
  assign n20408 = ~n20405 & ~n20407;
  assign n20409 = n20325 & ~n20408;
  assign n20410 = ~n20403 & ~n20409;
  assign n20411 = ~n20323 & n20324;
  assign n20412 = n20324 & ~n20411;
  assign n20413 = n20388 & ~n20389;
  assign n20414 = n20398 & n20413;
  assign n20415 = n20390 & n20394;
  assign n20416 = ~n20414 & ~n20415;
  assign n20417 = ~n20412 & ~n20416;
  assign n20418 = ~n20326 & ~n20355;
  assign n20419 = n20390 & n20411;
  assign n20420 = n20411 ^ n20388;
  assign n20421 = n20420 ^ n20411;
  assign n20422 = ~n20325 & ~n20393;
  assign n20423 = n20422 ^ n20411;
  assign n20424 = ~n20421 & ~n20423;
  assign n20425 = n20424 ^ n20411;
  assign n20426 = n20389 & n20425;
  assign n20427 = ~n20419 & ~n20426;
  assign n20428 = n20418 & ~n20427;
  assign n20429 = ~n20417 & ~n20428;
  assign n20430 = n20404 & n20406;
  assign n20431 = n20430 ^ n20411;
  assign n20432 = n20406 & n20413;
  assign n20433 = ~n20405 & ~n20432;
  assign n20434 = n20433 ^ n20402;
  assign n20435 = n20430 ^ n20402;
  assign n20436 = n20435 ^ n20402;
  assign n20437 = n20434 & ~n20436;
  assign n20438 = n20437 ^ n20402;
  assign n20439 = n20431 & n20438;
  assign n20440 = n20439 ^ n20411;
  assign n20441 = n20429 & ~n20440;
  assign n20445 = n20355 & n20390;
  assign n20442 = n20413 & n20418;
  assign n20443 = n20394 & n20413;
  assign n20444 = ~n20442 & ~n20443;
  assign n20446 = n20445 ^ n20444;
  assign n20447 = n20446 ^ n20445;
  assign n20448 = n20445 ^ n20323;
  assign n20449 = n20448 ^ n20445;
  assign n20450 = ~n20447 & n20449;
  assign n20451 = n20450 ^ n20445;
  assign n20452 = n20324 & n20451;
  assign n20453 = n20452 ^ n20445;
  assign n20454 = n20441 & ~n20453;
  assign n20456 = ~n20356 & n20395;
  assign n20455 = n20394 & n20404;
  assign n20457 = n20456 ^ n20455;
  assign n20458 = n20457 ^ n20456;
  assign n20459 = n20456 ^ n20323;
  assign n20460 = n20459 ^ n20456;
  assign n20461 = n20458 & ~n20460;
  assign n20462 = n20461 ^ n20456;
  assign n20463 = n20324 & n20462;
  assign n20464 = n20463 ^ n20456;
  assign n20465 = n20454 & ~n20464;
  assign n20466 = n20410 & n20465;
  assign n20467 = n20401 & n20466;
  assign n20468 = ~n20392 & n20467;
  assign n20469 = n20468 ^ n19075;
  assign n20470 = n19241 & n19306;
  assign n20471 = n19293 & n19319;
  assign n20472 = ~n20470 & ~n20471;
  assign n20473 = ~n19807 & ~n20369;
  assign n20474 = ~n19301 & n19824;
  assign n20475 = ~n19295 & n20474;
  assign n20476 = ~n19308 & n20372;
  assign n20477 = ~n19299 & n20476;
  assign n20478 = ~n19279 & n20477;
  assign n20479 = ~n20475 & ~n20478;
  assign n20480 = n19241 & n20479;
  assign n20481 = ~n19299 & n20357;
  assign n20482 = n19283 & ~n20481;
  assign n20483 = n19327 & n19814;
  assign n20484 = ~n19804 & n20483;
  assign n20485 = n19285 & ~n20484;
  assign n20486 = ~n20482 & ~n20485;
  assign n20487 = ~n20480 & n20486;
  assign n20488 = ~n19280 & n20487;
  assign n20489 = ~n20473 & n20488;
  assign n20490 = n20472 & n20489;
  assign n20491 = n19282 ^ n19241;
  assign n20492 = n20491 ^ n19282;
  assign n20493 = n19307 ^ n19282;
  assign n20494 = ~n20492 & n20493;
  assign n20495 = n20494 ^ n19282;
  assign n20496 = ~n19278 & n20495;
  assign n20497 = n20490 & ~n20496;
  assign n20498 = n19806 & n20497;
  assign n20499 = n19803 & n20498;
  assign n20500 = n20499 ^ n17370;
  assign n20501 = ~n18373 & ~n18377;
  assign n20502 = n18143 & ~n20501;
  assign n20503 = ~n18410 & n20291;
  assign n20504 = n18395 & ~n20503;
  assign n20505 = ~n20502 & ~n20504;
  assign n20506 = n18144 & ~n20064;
  assign n20507 = ~n18391 & ~n18430;
  assign n20508 = n18383 & ~n20507;
  assign n20509 = n18398 & ~n20298;
  assign n20510 = n18376 & ~n20509;
  assign n20511 = ~n20508 & ~n20510;
  assign n20512 = ~n20506 & n20511;
  assign n20513 = n20505 & n20512;
  assign n20514 = ~n18438 & n20513;
  assign n20515 = n20047 & n20514;
  assign n20516 = n18393 & n20515;
  assign n20517 = n18408 & n20516;
  assign n20518 = ~n18400 & n20517;
  assign n20519 = n20518 ^ n17613;
  assign n20520 = n20519 ^ x88;
  assign n20521 = n20013 ^ x81;
  assign n20522 = n20520 & n20521;
  assign n20523 = n17087 ^ n16758;
  assign n20524 = ~n20083 & ~n20523;
  assign n20525 = ~n18014 & n18040;
  assign n20526 = ~n18005 & n20525;
  assign n20527 = n17088 & ~n20526;
  assign n20528 = ~n20524 & ~n20527;
  assign n20529 = ~n18013 & n18021;
  assign n20530 = n18001 & ~n20529;
  assign n20531 = n18008 & n18015;
  assign n20532 = ~n17987 & n20531;
  assign n20533 = n18039 & n20532;
  assign n20534 = n18019 & ~n20533;
  assign n20535 = ~n20530 & ~n20534;
  assign n20536 = ~n17991 & ~n18007;
  assign n20537 = n18011 & ~n20536;
  assign n20538 = n18011 ^ n18001;
  assign n20541 = n17483 & n17986;
  assign n20542 = ~n18024 & ~n20541;
  assign n20543 = ~n18002 & n20542;
  assign n20539 = ~n18024 & ~n18027;
  assign n20540 = n18043 & n20539;
  assign n20544 = n20543 ^ n20540;
  assign n20545 = n20543 ^ n18011;
  assign n20546 = n20545 ^ n20543;
  assign n20547 = ~n20544 & n20546;
  assign n20548 = n20547 ^ n20543;
  assign n20549 = n20538 & n20548;
  assign n20550 = n20549 ^ n18001;
  assign n20551 = ~n20537 & ~n20550;
  assign n20552 = n20535 & n20551;
  assign n20553 = n20528 & n20552;
  assign n20554 = ~n20079 & n20553;
  assign n20555 = n18000 & n20554;
  assign n20556 = n20555 ^ n17880;
  assign n20557 = n20556 ^ x66;
  assign n20558 = ~n19414 & ~n19432;
  assign n20559 = ~n19447 & ~n20558;
  assign n20560 = n20118 & n20127;
  assign n20561 = ~n19407 & n20560;
  assign n20562 = n19409 & ~n20561;
  assign n20563 = ~n20559 & ~n20562;
  assign n20564 = n19352 & ~n20130;
  assign n20565 = ~n19407 & ~n19427;
  assign n20566 = n19414 & ~n20565;
  assign n20567 = ~n19439 & ~n19458;
  assign n20568 = ~n19432 & n20567;
  assign n20569 = ~n19427 & n19440;
  assign n20570 = ~n19352 & n20569;
  assign n20571 = ~n20568 & ~n20570;
  assign n20572 = ~n19477 & ~n20571;
  assign n20573 = ~n19433 & ~n20572;
  assign n20574 = ~n20566 & ~n20573;
  assign n20575 = ~n20564 & n20574;
  assign n20576 = n20563 & n20575;
  assign n20577 = ~n19473 & n20576;
  assign n20578 = n20123 & n20577;
  assign n20579 = ~n19572 & n20578;
  assign n20580 = n19422 & n20579;
  assign n20581 = n20580 ^ n17905;
  assign n20582 = n20581 ^ x105;
  assign n20583 = n20557 & n20582;
  assign n20584 = n20322 ^ x122;
  assign n20585 = ~n18962 & ~n18998;
  assign n20586 = n18944 & ~n20585;
  assign n20587 = ~n18975 & n18979;
  assign n20588 = ~n20586 & ~n20587;
  assign n20589 = n18896 & ~n18939;
  assign n20590 = ~n18996 & n20018;
  assign n20591 = n18953 & ~n20590;
  assign n20592 = ~n18958 & n18961;
  assign n20593 = ~n18955 & n19738;
  assign n20594 = ~n18948 & n20593;
  assign n20595 = n18953 & ~n20594;
  assign n20596 = ~n20592 & ~n20595;
  assign n20597 = n18940 & n19749;
  assign n20598 = ~n18984 & n20018;
  assign n20599 = n18944 & ~n20598;
  assign n20600 = ~n20597 & ~n20599;
  assign n20601 = ~n18951 & ~n18961;
  assign n20602 = ~n18965 & ~n18968;
  assign n20603 = ~n18948 & n20602;
  assign n20604 = ~n18940 & n20603;
  assign n20605 = ~n20601 & ~n20604;
  assign n20606 = ~n18978 & ~n20605;
  assign n20607 = ~n18975 & ~n20606;
  assign n20608 = n20600 & ~n20607;
  assign n20609 = n20596 & n20608;
  assign n20610 = ~n18949 & n20609;
  assign n20611 = ~n19728 & n20610;
  assign n20612 = ~n20591 & n20611;
  assign n20613 = ~n20589 & n20612;
  assign n20614 = n20588 & n20613;
  assign n20615 = ~n19729 & n20614;
  assign n20616 = n18946 & n20615;
  assign n20617 = n20616 ^ n17523;
  assign n20618 = n20617 ^ x120;
  assign n20619 = ~n20584 & ~n20618;
  assign n20620 = n20583 & n20619;
  assign n20621 = n20584 & n20618;
  assign n20622 = n20583 & n20621;
  assign n20623 = ~n20557 & ~n20582;
  assign n20624 = n20584 & ~n20618;
  assign n20625 = n20623 & n20624;
  assign n20626 = ~n20622 & ~n20625;
  assign n20627 = ~n20620 & n20626;
  assign n20628 = n20522 & ~n20627;
  assign n20629 = n20520 & ~n20521;
  assign n20630 = n20620 & n20629;
  assign n20631 = ~n20557 & n20582;
  assign n20632 = n20621 & n20631;
  assign n20633 = n20624 & n20631;
  assign n20634 = ~n20632 & ~n20633;
  assign n20635 = ~n20521 & ~n20634;
  assign n20636 = ~n20630 & ~n20635;
  assign n20637 = ~n20628 & n20636;
  assign n20638 = ~n20584 & n20618;
  assign n20639 = n20583 & n20638;
  assign n20640 = n20629 & n20639;
  assign n20641 = ~n20520 & n20521;
  assign n20642 = n20557 & ~n20582;
  assign n20643 = n20624 & n20642;
  assign n20644 = ~n20622 & ~n20643;
  assign n20645 = n20641 & ~n20644;
  assign n20646 = ~n20640 & ~n20645;
  assign n20647 = n20638 & n20642;
  assign n20648 = ~n20521 & n20647;
  assign n20649 = n20583 & n20624;
  assign n20650 = ~n20520 & n20649;
  assign n20651 = ~n20648 & ~n20650;
  assign n20652 = n20621 & n20623;
  assign n20653 = n20641 & n20652;
  assign n20654 = ~n20520 & ~n20521;
  assign n20655 = n20621 & n20642;
  assign n20656 = n20619 & n20642;
  assign n20657 = n20623 & n20638;
  assign n20658 = ~n20639 & ~n20657;
  assign n20659 = ~n20656 & n20658;
  assign n20660 = ~n20655 & n20659;
  assign n20661 = n20654 & ~n20660;
  assign n20662 = ~n20653 & ~n20661;
  assign n20663 = n20651 & n20662;
  assign n20664 = n20522 & n20632;
  assign n20665 = n20619 & n20623;
  assign n20666 = n20644 & ~n20665;
  assign n20667 = n20629 & ~n20666;
  assign n20668 = n20619 & n20631;
  assign n20669 = n20631 & n20638;
  assign n20670 = ~n20656 & ~n20669;
  assign n20671 = ~n20657 & n20670;
  assign n20672 = ~n20641 & n20671;
  assign n20673 = ~n20584 & n20623;
  assign n20674 = n20522 & ~n20670;
  assign n20675 = ~n20673 & ~n20674;
  assign n20676 = ~n20647 & n20675;
  assign n20677 = ~n20672 & ~n20676;
  assign n20678 = ~n20668 & ~n20677;
  assign n20679 = n20521 & ~n20678;
  assign n20680 = ~n20667 & ~n20679;
  assign n20681 = ~n20664 & n20680;
  assign n20682 = n20663 & n20681;
  assign n20683 = n20646 & n20682;
  assign n20684 = n20637 & n20683;
  assign n20685 = n20684 ^ n18856;
  assign n20686 = ~n20643 & ~n20652;
  assign n20687 = n20522 & ~n20686;
  assign n20688 = n20641 & ~n20658;
  assign n20689 = ~n20649 & ~n20655;
  assign n20690 = n20629 & ~n20689;
  assign n20691 = ~n20688 & ~n20690;
  assign n20692 = n20641 & n20655;
  assign n20693 = n20629 & n20656;
  assign n20694 = ~n20692 & ~n20693;
  assign n20695 = n20629 & ~n20658;
  assign n20696 = ~n20665 & ~n20669;
  assign n20697 = n20522 & ~n20696;
  assign n20698 = ~n20695 & ~n20697;
  assign n20699 = n20627 & n20670;
  assign n20700 = n20654 & ~n20699;
  assign n20701 = ~n20643 & ~n20668;
  assign n20702 = ~n20625 & n20701;
  assign n20703 = ~n20633 & n20702;
  assign n20704 = ~n20649 & n20703;
  assign n20705 = n20641 & ~n20704;
  assign n20706 = ~n20700 & ~n20705;
  assign n20707 = n20698 & n20706;
  assign n20708 = n20521 ^ n20520;
  assign n20709 = n20639 ^ n20521;
  assign n20710 = n20709 ^ n20639;
  assign n20711 = n20647 ^ n20639;
  assign n20712 = ~n20710 & n20711;
  assign n20713 = n20712 ^ n20639;
  assign n20714 = ~n20708 & n20713;
  assign n20715 = n20707 & ~n20714;
  assign n20716 = n20694 & n20715;
  assign n20717 = n20691 & n20716;
  assign n20718 = ~n20687 & n20717;
  assign n20719 = n20637 & n20718;
  assign n20720 = n20719 ^ n18295;
  assign n20721 = n18731 & n18748;
  assign n20722 = ~n18738 & ~n18742;
  assign n20723 = n19920 & n20722;
  assign n20724 = ~n18759 & n20723;
  assign n20725 = n18764 & ~n20724;
  assign n20726 = ~n20721 & ~n20725;
  assign n20727 = ~n18578 & n18775;
  assign n20728 = n18739 & ~n18758;
  assign n20729 = n18733 & ~n20728;
  assign n20730 = ~n18740 & ~n18745;
  assign n20731 = n18727 & n18737;
  assign n20732 = n18760 ^ n18578;
  assign n20733 = n18760 ^ n18726;
  assign n20734 = n20733 ^ n18726;
  assign n20735 = n18748 & ~n19920;
  assign n20736 = ~n18765 & ~n20735;
  assign n20737 = n20736 ^ n18726;
  assign n20738 = ~n20734 & ~n20737;
  assign n20739 = n20738 ^ n18726;
  assign n20740 = ~n20732 & ~n20739;
  assign n20741 = n20740 ^ n18578;
  assign n20742 = ~n20731 & n20741;
  assign n20743 = ~n20730 & n20742;
  assign n20744 = ~n20729 & n20743;
  assign n20745 = ~n20727 & n20744;
  assign n20746 = n20726 & n20745;
  assign n20747 = ~n18756 & n20746;
  assign n20748 = n19914 & n20747;
  assign n20749 = ~n20338 & n20748;
  assign n20750 = ~n18752 & n20749;
  assign n20751 = ~n19910 & n20750;
  assign n20752 = n20751 ^ n17581;
  assign n20753 = ~n19867 & n19875;
  assign n20754 = ~n19854 & ~n19885;
  assign n20755 = ~n19880 & n20754;
  assign n20756 = n19963 & n20755;
  assign n20757 = ~n19843 & n20756;
  assign n20758 = n19600 & ~n20757;
  assign n20759 = ~n20753 & ~n20758;
  assign n20760 = n19887 & ~n19891;
  assign n20761 = ~n19876 & n20760;
  assign n20762 = n19845 & ~n20761;
  assign n20763 = ~n19861 & n20755;
  assign n20764 = n19840 & ~n20763;
  assign n20765 = ~n19847 & ~n19886;
  assign n20766 = ~n19875 & n20765;
  assign n20767 = ~n19859 & n20766;
  assign n20768 = ~n19880 & n20767;
  assign n20769 = n19851 & ~n20768;
  assign n20770 = ~n20764 & ~n20769;
  assign n20771 = ~n20762 & n20770;
  assign n20772 = n20759 & n20771;
  assign n20773 = ~n19947 & n20772;
  assign n20774 = ~n19865 & n20773;
  assign n20775 = n19957 & n20774;
  assign n20776 = ~n19856 & n20775;
  assign n20777 = n19850 & n20776;
  assign n20778 = n20777 ^ n19370;
  assign n20779 = n18019 & n20097;
  assign n20780 = n18012 & ~n20523;
  assign n20781 = ~n18030 & ~n20523;
  assign n20782 = n17088 & ~n18015;
  assign n20783 = ~n20781 & ~n20782;
  assign n20784 = n18011 & ~n20532;
  assign n20785 = ~n18005 & n18021;
  assign n20786 = n18019 & ~n20785;
  assign n20787 = n20089 & n20539;
  assign n20788 = n18040 & n20787;
  assign n20789 = n18001 & ~n20788;
  assign n20790 = ~n20786 & ~n20789;
  assign n20791 = ~n20784 & n20790;
  assign n20792 = n20783 & n20791;
  assign n20793 = n20081 & n20792;
  assign n20794 = ~n20780 & n20793;
  assign n20795 = ~n20779 & n20794;
  assign n20796 = ~n17988 & n20795;
  assign n20797 = n20796 ^ n17765;
  assign n20798 = n18794 & ~n19526;
  assign n20799 = n19500 & ~n19528;
  assign n20800 = ~n20798 & ~n20799;
  assign n20801 = n19494 & n19500;
  assign n20802 = n18794 & n19510;
  assign n20803 = ~n20801 & ~n20802;
  assign n20804 = ~n19489 & ~n19525;
  assign n20805 = n19491 & ~n20804;
  assign n20806 = ~n19503 & n19557;
  assign n20807 = n19522 & ~n20806;
  assign n20808 = ~n18794 & ~n19504;
  assign n20809 = ~n19516 & ~n19542;
  assign n20810 = ~n19503 & ~n19514;
  assign n20811 = n20809 & n20810;
  assign n20812 = ~n20808 & ~n20811;
  assign n20813 = ~n20807 & ~n20812;
  assign n20814 = ~n19500 & ~n19522;
  assign n20815 = ~n19509 & ~n19515;
  assign n20816 = ~n19531 & n20815;
  assign n20817 = ~n19507 & n20816;
  assign n20818 = ~n20814 & ~n20817;
  assign n20819 = n19140 ^ n19013;
  assign n20820 = n20819 ^ n19487;
  assign n20821 = ~n19348 & n20820;
  assign n20822 = n19491 & n20821;
  assign n20823 = ~n20818 & ~n20822;
  assign n20824 = n20813 & n20823;
  assign n20825 = ~n20805 & n20824;
  assign n20826 = n20803 & n20825;
  assign n20827 = n20800 & n20826;
  assign n20828 = n19498 & n20827;
  assign n20829 = n20828 ^ n19041;
  assign n20830 = n19690 & n19692;
  assign n20831 = n19681 & ~n19994;
  assign n20832 = ~n20830 & ~n20831;
  assign n20833 = n19676 & n19702;
  assign n20835 = n19616 ^ n19615;
  assign n20836 = n20835 ^ n19655;
  assign n20837 = n20836 ^ n19656;
  assign n20834 = n19616 & n19669;
  assign n20838 = n20837 ^ n20834;
  assign n20839 = n19668 & ~n20838;
  assign n20840 = n19674 & n20214;
  assign n20841 = n19603 & ~n20840;
  assign n20842 = ~n19662 & ~n19694;
  assign n20843 = ~n19676 & n20842;
  assign n20844 = ~n19692 & n19713;
  assign n20845 = ~n20843 & ~n20844;
  assign n20846 = ~n19678 & ~n20845;
  assign n20847 = ~n19994 & ~n20846;
  assign n20848 = ~n20841 & ~n20847;
  assign n20849 = ~n20839 & n20848;
  assign n20850 = ~n20833 & n20849;
  assign n20851 = n20832 & n20850;
  assign n20852 = ~n19666 & n20851;
  assign n20853 = ~n19989 & n20852;
  assign n20854 = ~n20237 & n20853;
  assign n20855 = n19988 & n20854;
  assign n20856 = n20855 ^ n17417;
  assign n20857 = ~n20148 & n20158;
  assign n20858 = n20151 & ~n20857;
  assign n20859 = ~n20158 & n20194;
  assign n20860 = ~n20165 & n20266;
  assign n20861 = ~n20175 & n20860;
  assign n20862 = n20161 & ~n20861;
  assign n20863 = ~n20859 & ~n20862;
  assign n20864 = ~n20156 & ~n20172;
  assign n20865 = n20042 & ~n20864;
  assign n20866 = n20165 ^ n20041;
  assign n20868 = ~n20175 & ~n20190;
  assign n20867 = ~n20181 & n20260;
  assign n20869 = n20868 ^ n20867;
  assign n20870 = n20868 ^ n20014;
  assign n20871 = n20870 ^ n20868;
  assign n20872 = n20869 & ~n20871;
  assign n20873 = n20872 ^ n20868;
  assign n20874 = n20873 ^ n20165;
  assign n20875 = ~n20866 & ~n20874;
  assign n20876 = n20875 ^ n20872;
  assign n20877 = n20876 ^ n20868;
  assign n20878 = n20877 ^ n20041;
  assign n20879 = ~n20165 & n20878;
  assign n20880 = n20879 ^ n20165;
  assign n20881 = n20880 ^ n20041;
  assign n20882 = ~n20865 & n20881;
  assign n20883 = n20863 & n20882;
  assign n20884 = ~n20248 & n20883;
  assign n20885 = n20243 & n20884;
  assign n20886 = ~n20858 & n20885;
  assign n20887 = ~n20174 & ~n20259;
  assign n20888 = n20182 & n20887;
  assign n20889 = n20888 ^ n20014;
  assign n20890 = n20889 ^ n20888;
  assign n20891 = n20173 & ~n20241;
  assign n20892 = ~n20146 & n20891;
  assign n20893 = n20892 ^ n20888;
  assign n20894 = n20890 & n20893;
  assign n20895 = n20894 ^ n20888;
  assign n20896 = ~n20041 & ~n20895;
  assign n20897 = n20886 & ~n20896;
  assign n20898 = ~n20247 & n20897;
  assign n20899 = ~n20150 & n20898;
  assign n20900 = n20899 ^ n18893;
  assign n20901 = ~n19875 & ~n19880;
  assign n20902 = n19845 & ~n20901;
  assign n20903 = ~n19866 & n20755;
  assign n20904 = n19851 & ~n20903;
  assign n20905 = ~n20902 & ~n20904;
  assign n20906 = n19853 & ~n19867;
  assign n20907 = ~n19883 & n20766;
  assign n20908 = n19840 & ~n20907;
  assign n20909 = ~n20906 & ~n20908;
  assign n20910 = n20905 & n20909;
  assign n20911 = n19959 ^ n19886;
  assign n20912 = n20911 ^ n19886;
  assign n20913 = n19886 ^ n19599;
  assign n20914 = n20913 ^ n19886;
  assign n20915 = ~n20912 & ~n20914;
  assign n20916 = n20915 ^ n19886;
  assign n20917 = ~n19874 & n20916;
  assign n20918 = n20917 ^ n19886;
  assign n20919 = n20910 & ~n20918;
  assign n20920 = ~n19871 & n20919;
  assign n20921 = ~n19949 & n20920;
  assign n20922 = n19864 & n20921;
  assign n20923 = n19948 & n20922;
  assign n20924 = n19850 & n20923;
  assign n20925 = ~n19843 & n20924;
  assign n20926 = n20925 ^ n18328;
  assign n20927 = n20325 & n20396;
  assign n20928 = n20391 & n20402;
  assign n20929 = n20404 & n20418;
  assign n20930 = ~n20430 & ~n20929;
  assign n20931 = n20411 & ~n20930;
  assign n20932 = ~n20928 & ~n20931;
  assign n20933 = n20390 & n20398;
  assign n20934 = ~n20443 & ~n20933;
  assign n20935 = ~n20415 & n20934;
  assign n20936 = ~n20432 & n20935;
  assign n20937 = n20393 & ~n20936;
  assign n20938 = n20398 & n20426;
  assign n20939 = ~n20937 & ~n20938;
  assign n20940 = ~n20422 & n20430;
  assign n20941 = n20390 & n20418;
  assign n20942 = ~n20432 & n20444;
  assign n20943 = ~n20325 & n20942;
  assign n20944 = ~n20411 & n20935;
  assign n20945 = ~n20943 & ~n20944;
  assign n20946 = ~n20941 & ~n20945;
  assign n20947 = n20946 ^ n20323;
  assign n20948 = n20947 ^ n20946;
  assign n20949 = ~n20414 & ~n20455;
  assign n20950 = ~n20432 & n20949;
  assign n20951 = ~n20405 & n20950;
  assign n20952 = n20951 ^ n20946;
  assign n20953 = n20952 ^ n20946;
  assign n20954 = n20948 & ~n20953;
  assign n20955 = n20954 ^ n20946;
  assign n20956 = ~n20324 & ~n20955;
  assign n20957 = n20956 ^ n20946;
  assign n20958 = ~n20940 & n20957;
  assign n20959 = n20939 & n20958;
  assign n20960 = ~n20400 & n20959;
  assign n20961 = ~n20464 & n20960;
  assign n20962 = n20932 & n20961;
  assign n20963 = ~n20927 & n20962;
  assign n20964 = n20963 ^ n19277;
  assign n20965 = n19835 ^ x113;
  assign n20966 = n20617 ^ x104;
  assign n20967 = ~n20965 & ~n20966;
  assign n20968 = n18059 ^ x90;
  assign n20969 = n20239 ^ x80;
  assign n20970 = n20968 & ~n20969;
  assign n20971 = n20519 ^ x99;
  assign n20972 = n20752 ^ x73;
  assign n20973 = n20971 & n20972;
  assign n20974 = n20970 & n20973;
  assign n20975 = ~n20968 & n20969;
  assign n20976 = n20971 & ~n20972;
  assign n20977 = n20975 & n20976;
  assign n20978 = ~n20974 & ~n20977;
  assign n20979 = n20967 & ~n20978;
  assign n20980 = ~n20965 & n20966;
  assign n20981 = n20968 & n20969;
  assign n20982 = ~n20971 & n20972;
  assign n20983 = n20981 & n20982;
  assign n20984 = n20970 & n20982;
  assign n20985 = ~n20968 & ~n20969;
  assign n20986 = ~n20971 & ~n20972;
  assign n20987 = n20985 & n20986;
  assign n20988 = ~n20984 & ~n20987;
  assign n20989 = ~n20983 & n20988;
  assign n20990 = n20980 & ~n20989;
  assign n20991 = n20973 & n20975;
  assign n20992 = ~n20974 & ~n20991;
  assign n20993 = n20980 & ~n20992;
  assign n20994 = n20965 & ~n20966;
  assign n20995 = ~n20988 & n20994;
  assign n20996 = ~n20993 & ~n20995;
  assign n20997 = n20965 & n20966;
  assign n20998 = n20981 & n20986;
  assign n20999 = n20997 & n20998;
  assign n21000 = n20973 & n20981;
  assign n21001 = n20973 & n20985;
  assign n21002 = n20970 & n20976;
  assign n21003 = ~n21001 & ~n21002;
  assign n21004 = ~n20977 & n21003;
  assign n21005 = ~n20998 & n21004;
  assign n21006 = ~n21000 & n21005;
  assign n21007 = n20994 & ~n21006;
  assign n21008 = n20975 & n20986;
  assign n21009 = n20976 & n20981;
  assign n21010 = ~n21008 & ~n21009;
  assign n21011 = n20980 & ~n21010;
  assign n21012 = n20978 & ~n20983;
  assign n21013 = n20997 & ~n21012;
  assign n21014 = ~n20967 & ~n20997;
  assign n21015 = n20975 & n20982;
  assign n21016 = n20982 & n20985;
  assign n21017 = n20970 & n20986;
  assign n21018 = ~n20983 & ~n21017;
  assign n21019 = n20967 & ~n21018;
  assign n21020 = ~n21002 & ~n21019;
  assign n21021 = ~n21016 & n21020;
  assign n21022 = ~n21015 & n21021;
  assign n21023 = ~n21014 & ~n21022;
  assign n21024 = ~n21013 & ~n21023;
  assign n21025 = ~n21011 & n21024;
  assign n21026 = ~n21007 & n21025;
  assign n21027 = ~n20999 & n21026;
  assign n21028 = n20966 ^ n20965;
  assign n21029 = n21001 ^ n20966;
  assign n21030 = n21029 ^ n21001;
  assign n21031 = n21001 ^ n20991;
  assign n21032 = ~n21030 & n21031;
  assign n21033 = n21032 ^ n21001;
  assign n21034 = ~n21028 & n21033;
  assign n21035 = n21027 & ~n21034;
  assign n21036 = n20976 & n20985;
  assign n21037 = n21036 ^ n20966;
  assign n21038 = n21037 ^ n21036;
  assign n21039 = n21036 ^ n21008;
  assign n21040 = ~n21038 & n21039;
  assign n21041 = n21040 ^ n21036;
  assign n21042 = n21028 & n21041;
  assign n21043 = n21035 & ~n21042;
  assign n21044 = n20996 & n21043;
  assign n21045 = ~n20990 & n21044;
  assign n21046 = ~n20979 & n21045;
  assign n21047 = n21046 ^ n18577;
  assign n21048 = n20411 & n20456;
  assign n21049 = n20393 & ~n20930;
  assign n21050 = ~n21048 & ~n21049;
  assign n21051 = n20325 & n20414;
  assign n21052 = n20402 & ~n20934;
  assign n21053 = ~n21051 & ~n21052;
  assign n21054 = n20325 & n20455;
  assign n21055 = n20393 & n20399;
  assign n21056 = ~n21054 & ~n21055;
  assign n21057 = ~n20430 & n20433;
  assign n21058 = ~n20456 & n21057;
  assign n21059 = n20402 & ~n21058;
  assign n21060 = n20390 & n20406;
  assign n21061 = ~n20442 & n20950;
  assign n21062 = ~n21060 & n21061;
  assign n21063 = n20411 & ~n21062;
  assign n21064 = ~n21059 & ~n21063;
  assign n21065 = ~n20393 & ~n20398;
  assign n21066 = ~n20935 & ~n21065;
  assign n21067 = ~n20442 & ~n21066;
  assign n21068 = n21067 ^ n20422;
  assign n21069 = n21068 ^ n21067;
  assign n21070 = n21067 ^ n20929;
  assign n21071 = n21069 & ~n21070;
  assign n21072 = n21071 ^ n21067;
  assign n21073 = n21064 & n21072;
  assign n21074 = n21056 & n21073;
  assign n21075 = n21053 & n21074;
  assign n21076 = n20401 & n21075;
  assign n21077 = n21050 & n21076;
  assign n21078 = ~n20927 & n21077;
  assign n21079 = ~n20392 & n21078;
  assign n21080 = n21079 ^ n17086;
  assign n21081 = n19139 ^ x118;
  assign n21082 = n20106 ^ x100;
  assign n21083 = ~n21081 & n21082;
  assign n21084 = n18446 ^ x101;
  assign n21085 = n19944 ^ x94;
  assign n21086 = ~n21084 & n21085;
  assign n21087 = n20500 ^ x124;
  assign n21088 = n20856 ^ x76;
  assign n21089 = n21087 & ~n21088;
  assign n21090 = n21086 & n21089;
  assign n21091 = n21083 & n21090;
  assign n21092 = n21081 & ~n21082;
  assign n21093 = n21084 & ~n21085;
  assign n21094 = ~n21087 & n21088;
  assign n21095 = n21093 & n21094;
  assign n21096 = n21084 & n21085;
  assign n21097 = ~n21087 & ~n21088;
  assign n21098 = n21096 & n21097;
  assign n21099 = ~n21095 & ~n21098;
  assign n21100 = n21099 ^ n21083;
  assign n21101 = n21100 ^ n21099;
  assign n21102 = n21089 & n21093;
  assign n21103 = n21102 ^ n21099;
  assign n21104 = n21103 ^ n21099;
  assign n21105 = ~n21101 & n21104;
  assign n21106 = n21105 ^ n21099;
  assign n21107 = ~n21092 & ~n21106;
  assign n21108 = n21107 ^ n21099;
  assign n21109 = ~n21091 & n21108;
  assign n21110 = ~n21081 & ~n21082;
  assign n21111 = n21087 & n21088;
  assign n21112 = n21096 & n21111;
  assign n21113 = n21110 & n21112;
  assign n21114 = ~n21083 & ~n21092;
  assign n21115 = n21093 & n21097;
  assign n21116 = n21114 & n21115;
  assign n21117 = ~n21113 & ~n21116;
  assign n21118 = n21081 & n21082;
  assign n21119 = n21093 & n21111;
  assign n21120 = n21094 & n21096;
  assign n21121 = ~n21119 & ~n21120;
  assign n21122 = n21118 & ~n21121;
  assign n21123 = n21088 ^ n21087;
  assign n21125 = n21123 ^ n21088;
  assign n21126 = n21084 & ~n21125;
  assign n21124 = ~n21085 & ~n21123;
  assign n21127 = n21126 ^ n21124;
  assign n21128 = ~n21112 & ~n21127;
  assign n21129 = n21083 & ~n21128;
  assign n21130 = ~n21122 & ~n21129;
  assign n21131 = n21089 & n21096;
  assign n21132 = ~n21119 & ~n21131;
  assign n21133 = n21092 & ~n21132;
  assign n21134 = ~n21084 & ~n21085;
  assign n21135 = n21097 & n21134;
  assign n21136 = n21086 & n21094;
  assign n21137 = n21086 & n21111;
  assign n21138 = n21094 & n21134;
  assign n21139 = ~n21137 & ~n21138;
  assign n21140 = n21092 & ~n21139;
  assign n21141 = ~n21136 & ~n21140;
  assign n21142 = ~n21135 & n21141;
  assign n21143 = ~n21110 & n21142;
  assign n21144 = ~n21082 & ~n21143;
  assign n21145 = ~n21118 & ~n21144;
  assign n21146 = n21086 & n21097;
  assign n21147 = ~n21138 & ~n21146;
  assign n21148 = n21089 & n21134;
  assign n21149 = n21139 & ~n21148;
  assign n21150 = ~n21092 & n21141;
  assign n21151 = n21144 & ~n21150;
  assign n21152 = n21149 & ~n21151;
  assign n21153 = n21147 & n21152;
  assign n21154 = ~n21145 & ~n21153;
  assign n21155 = ~n21133 & ~n21154;
  assign n21156 = n21130 & n21155;
  assign n21157 = n21117 & n21156;
  assign n21158 = n21109 & n21157;
  assign n21159 = n21158 ^ n18367;
  assign n21160 = n21110 & n21120;
  assign n21161 = n21110 & n21119;
  assign n21162 = n21114 & n21131;
  assign n21163 = ~n21161 & ~n21162;
  assign n21164 = ~n21095 & ~n21120;
  assign n21165 = n21118 & ~n21164;
  assign n21166 = n21090 & n21092;
  assign n21167 = n21099 & ~n21119;
  assign n21168 = n21083 & ~n21167;
  assign n21169 = ~n21166 & ~n21168;
  assign n21170 = ~n21115 & n21169;
  assign n21171 = ~n21114 & ~n21170;
  assign n21172 = n21111 & n21134;
  assign n21173 = ~n21146 & ~n21172;
  assign n21174 = n21141 & n21173;
  assign n21175 = ~n21115 & n21174;
  assign n21176 = ~n21118 & n21175;
  assign n21177 = ~n21114 & ~n21140;
  assign n21178 = n21143 & ~n21148;
  assign n21179 = ~n21146 & n21178;
  assign n21180 = ~n21177 & ~n21179;
  assign n21181 = ~n21176 & n21180;
  assign n21182 = ~n21171 & ~n21181;
  assign n21183 = ~n21165 & n21182;
  assign n21184 = n21163 & n21183;
  assign n21185 = n21082 ^ n21081;
  assign n21186 = n21149 ^ n21082;
  assign n21187 = n21186 ^ n21149;
  assign n21188 = ~n21102 & ~n21112;
  assign n21189 = n21188 ^ n21149;
  assign n21190 = ~n21187 & n21189;
  assign n21191 = n21190 ^ n21149;
  assign n21192 = n21185 & ~n21191;
  assign n21193 = n21184 & ~n21192;
  assign n21194 = n21109 & n21193;
  assign n21195 = ~n21160 & n21194;
  assign n21196 = n21195 ^ n19171;
  assign n21197 = n20175 & n20249;
  assign n21198 = n20182 & ~n20241;
  assign n21199 = n20151 & ~n21198;
  assign n21200 = ~n20156 & n20266;
  assign n21201 = n20194 & ~n21200;
  assign n21202 = ~n21199 & ~n21201;
  assign n21203 = ~n21197 & n21202;
  assign n21204 = n20161 & n20206;
  assign n21205 = n20176 & n20860;
  assign n21206 = ~n20157 & n21205;
  assign n21207 = n20042 & ~n21206;
  assign n21208 = ~n21204 & ~n21207;
  assign n21209 = n21203 & n21208;
  assign n21210 = ~n20245 & n21209;
  assign n21211 = ~n20160 & n21210;
  assign n21212 = ~n20150 & n21211;
  assign n21213 = n20243 & n21212;
  assign n21214 = n21213 ^ n18523;
  assign n21215 = n19347 ^ x112;
  assign n21216 = n19725 ^ x65;
  assign n21217 = ~n21215 & n21216;
  assign n21218 = n20313 ^ x98;
  assign n21219 = n19598 ^ x72;
  assign n21220 = n21218 & n21219;
  assign n21221 = n18792 ^ x89;
  assign n21222 = n21220 & n21221;
  assign n21223 = n20797 ^ x107;
  assign n21224 = ~n21219 & ~n21223;
  assign n21225 = ~n21218 & ~n21221;
  assign n21226 = ~n21224 & n21225;
  assign n21227 = ~n21218 & n21221;
  assign n21228 = n21227 ^ n21218;
  assign n21229 = ~n21223 & n21228;
  assign n21230 = n21229 ^ n21218;
  assign n21231 = ~n21219 & n21230;
  assign n21232 = ~n21226 & ~n21231;
  assign n21233 = ~n21222 & n21232;
  assign n21234 = n21217 & n21233;
  assign n21235 = ~n21215 & ~n21216;
  assign n21237 = n21219 & n21227;
  assign n21236 = ~n21219 & n21225;
  assign n21238 = n21237 ^ n21236;
  assign n21239 = n21223 & n21238;
  assign n21240 = n21239 ^ n21237;
  assign n21241 = ~n21221 & ~n21223;
  assign n21242 = n21219 ^ n21218;
  assign n21243 = n21242 ^ n21218;
  assign n21244 = n21225 ^ n21218;
  assign n21245 = n21243 & ~n21244;
  assign n21246 = n21245 ^ n21218;
  assign n21247 = ~n21241 & n21246;
  assign n21248 = n21247 ^ n21219;
  assign n21249 = ~n21240 & ~n21248;
  assign n21250 = n21235 & ~n21249;
  assign n21251 = ~n21234 & ~n21250;
  assign n21252 = n21221 ^ n21219;
  assign n21253 = n21223 ^ n21219;
  assign n21254 = n21253 ^ n21221;
  assign n21255 = n21254 ^ n21219;
  assign n21256 = n21255 ^ n21219;
  assign n21257 = ~n21252 & n21256;
  assign n21258 = n21257 ^ n21219;
  assign n21259 = ~n21218 & n21258;
  assign n21260 = n21259 ^ n21254;
  assign n21261 = n21260 ^ n21216;
  assign n21262 = n21261 ^ n21260;
  assign n21263 = n21218 & n21241;
  assign n21265 = n21219 & n21223;
  assign n21264 = n21221 & n21223;
  assign n21266 = n21265 ^ n21264;
  assign n21267 = n21218 & n21266;
  assign n21268 = n21267 ^ n21265;
  assign n21269 = ~n21231 & ~n21268;
  assign n21270 = ~n21263 & n21269;
  assign n21271 = n21270 ^ n21260;
  assign n21272 = ~n21262 & n21271;
  assign n21273 = n21272 ^ n21260;
  assign n21274 = n21215 & ~n21273;
  assign n21275 = n21251 & ~n21274;
  assign n21276 = n21275 ^ n17848;
  assign n21277 = ~n20978 & n20994;
  assign n21278 = ~n20999 & ~n21277;
  assign n21279 = ~n21001 & ~n21016;
  assign n21280 = n20997 & ~n21279;
  assign n21281 = ~n20998 & ~n21016;
  assign n21282 = ~n20983 & n21281;
  assign n21283 = n21003 & n21282;
  assign n21284 = ~n20987 & n21283;
  assign n21285 = n20980 & ~n21284;
  assign n21286 = ~n21280 & ~n21285;
  assign n21287 = ~n20984 & ~n21015;
  assign n21288 = n20967 & ~n21287;
  assign n21289 = ~n21000 & ~n21036;
  assign n21290 = ~n21017 & n21289;
  assign n21291 = ~n21014 & ~n21290;
  assign n21292 = ~n20991 & ~n21002;
  assign n21293 = ~n21009 & n21292;
  assign n21294 = ~n21015 & n21293;
  assign n21295 = n20994 & ~n21294;
  assign n21296 = ~n21291 & ~n21295;
  assign n21297 = ~n21288 & n21296;
  assign n21298 = n21286 & n21297;
  assign n21299 = n21008 ^ n20997;
  assign n21300 = n21008 ^ n20983;
  assign n21301 = n21300 ^ n20983;
  assign n21302 = n20983 ^ n20967;
  assign n21303 = n21301 & ~n21302;
  assign n21304 = n21303 ^ n20983;
  assign n21305 = n21299 & ~n21304;
  assign n21306 = n21305 ^ n20997;
  assign n21307 = n21298 & ~n21306;
  assign n21308 = n20996 & n21307;
  assign n21309 = n21278 & n21308;
  assign n21310 = ~n20979 & n21309;
  assign n21311 = n21310 ^ n18142;
  assign n21312 = n19491 & n19527;
  assign n21313 = ~n19495 & ~n19524;
  assign n21314 = n19500 & ~n21313;
  assign n21315 = ~n21312 & ~n21314;
  assign n21316 = n19531 & n20814;
  assign n21317 = ~n19507 & n20810;
  assign n21318 = n19522 & ~n21317;
  assign n21319 = ~n19507 & n20809;
  assign n21320 = n19500 & ~n21319;
  assign n21321 = ~n19494 & ~n19524;
  assign n21322 = ~n19509 & n21321;
  assign n21323 = n19522 & ~n21322;
  assign n21324 = ~n21320 & ~n21323;
  assign n21325 = n18794 & n19525;
  assign n21326 = ~n19489 & n19557;
  assign n21327 = ~n19507 & n21326;
  assign n21328 = ~n18794 & n21327;
  assign n21329 = ~n19515 & n19558;
  assign n21330 = ~n19491 & n21329;
  assign n21331 = ~n21328 & ~n21330;
  assign n21332 = n20814 & n21331;
  assign n21333 = ~n21325 & ~n21332;
  assign n21334 = n21324 & n21333;
  assign n21335 = n19505 & n21334;
  assign n21336 = ~n21318 & n21335;
  assign n21337 = ~n21316 & n21336;
  assign n21338 = n21315 & n21337;
  assign n21339 = n19539 & n21338;
  assign n21340 = n19498 & n21339;
  assign n21341 = n21340 ^ n19237;
  assign n21342 = n21092 & n21148;
  assign n21343 = n21090 & n21110;
  assign n21344 = n21083 & ~n21121;
  assign n21345 = ~n21343 & ~n21344;
  assign n21346 = ~n21342 & n21345;
  assign n21347 = ~n21115 & ~n21131;
  assign n21348 = n21083 & ~n21347;
  assign n21349 = n21081 & n21146;
  assign n21350 = ~n21090 & ~n21135;
  assign n21351 = n21147 & n21350;
  assign n21352 = n21083 & ~n21351;
  assign n21353 = ~n21112 & n21347;
  assign n21354 = ~n21119 & n21353;
  assign n21355 = n21092 & ~n21354;
  assign n21356 = ~n21352 & ~n21355;
  assign n21357 = ~n21095 & n21188;
  assign n21358 = ~n21118 & n21357;
  assign n21359 = ~n21110 & n21347;
  assign n21360 = n21099 & n21359;
  assign n21361 = ~n21358 & ~n21360;
  assign n21362 = ~n21148 & ~n21361;
  assign n21363 = ~n21172 & n21362;
  assign n21364 = n21114 & ~n21363;
  assign n21365 = n21356 & ~n21364;
  assign n21366 = ~n21160 & n21365;
  assign n21367 = ~n21349 & n21366;
  assign n21368 = ~n21348 & n21367;
  assign n21369 = n21137 ^ n21082;
  assign n21370 = n21369 ^ n21137;
  assign n21371 = n21137 ^ n21136;
  assign n21372 = ~n21370 & n21371;
  assign n21373 = n21372 ^ n21137;
  assign n21374 = ~n21185 & n21373;
  assign n21375 = n21368 & ~n21374;
  assign n21376 = n21346 & n21375;
  assign n21377 = ~n21140 & n21376;
  assign n21378 = n21377 ^ n18544;
  assign n21379 = ~n21081 & n21098;
  assign n21380 = n21083 & n21102;
  assign n21381 = ~n21379 & ~n21380;
  assign n21382 = n21114 & ~n21147;
  assign n21383 = ~n21137 & n21350;
  assign n21384 = n21092 & ~n21383;
  assign n21385 = ~n21136 & ~n21172;
  assign n21386 = n21118 & ~n21385;
  assign n21387 = ~n21095 & n21121;
  assign n21388 = ~n21115 & n21387;
  assign n21389 = n21092 & ~n21388;
  assign n21390 = n21139 & n21173;
  assign n21391 = n21083 & ~n21390;
  assign n21392 = ~n21389 & ~n21391;
  assign n21393 = ~n21386 & n21392;
  assign n21394 = n21347 ^ n21119;
  assign n21395 = n21347 ^ n21110;
  assign n21396 = n21395 ^ n21110;
  assign n21397 = n21118 ^ n21110;
  assign n21398 = ~n21396 & ~n21397;
  assign n21399 = n21398 ^ n21110;
  assign n21400 = ~n21394 & ~n21399;
  assign n21401 = n21400 ^ n21119;
  assign n21402 = n21188 & ~n21401;
  assign n21403 = n21114 & ~n21402;
  assign n21404 = n21393 & ~n21403;
  assign n21405 = ~n21160 & n21404;
  assign n21406 = ~n21384 & n21405;
  assign n21407 = ~n21382 & n21406;
  assign n21408 = n21381 & n21407;
  assign n21409 = n21346 & n21408;
  assign n21410 = n21409 ^ n17482;
  assign n21411 = ~n20399 & n20408;
  assign n21412 = n20402 & ~n21411;
  assign n21413 = n20395 & n20418;
  assign n21414 = ~n20415 & ~n21413;
  assign n21415 = ~n20422 & ~n21414;
  assign n21416 = ~n21412 & ~n21415;
  assign n21417 = n20411 & ~n20936;
  assign n21418 = n20393 & ~n21061;
  assign n21419 = ~n21417 & ~n21418;
  assign n21420 = n21416 & n21419;
  assign n21421 = n21053 & n21420;
  assign n21422 = n20410 & n21421;
  assign n21423 = n20932 & n21422;
  assign n21424 = n21050 & n21423;
  assign n21425 = ~n20927 & n21424;
  assign n21426 = ~n20392 & n21425;
  assign n21427 = n21426 ^ n19654;
  assign n21428 = n20967 & n21001;
  assign n21429 = n20980 & ~n21004;
  assign n21430 = n21018 & ~n21036;
  assign n21431 = ~n21008 & n21430;
  assign n21432 = n20967 & ~n21431;
  assign n21433 = ~n21015 & ~n21017;
  assign n21434 = n21289 & n21433;
  assign n21435 = ~n21002 & n21434;
  assign n21436 = n20994 & ~n21435;
  assign n21437 = ~n21432 & ~n21436;
  assign n21438 = n20997 & n21000;
  assign n21439 = ~n20974 & ~n21009;
  assign n21440 = ~n21014 & ~n21439;
  assign n21441 = n20989 & ~n21015;
  assign n21442 = n20980 & ~n21441;
  assign n21443 = ~n20997 & ~n21442;
  assign n21444 = ~n20990 & n21433;
  assign n21445 = ~n20987 & n21444;
  assign n21446 = ~n21443 & ~n21445;
  assign n21447 = ~n21440 & ~n21446;
  assign n21448 = ~n21438 & n21447;
  assign n21449 = n21437 & n21448;
  assign n21450 = n21278 & n21449;
  assign n21451 = ~n21429 & n21450;
  assign n21452 = ~n21428 & n21451;
  assign n21453 = ~n21034 & n21452;
  assign n21454 = ~n21042 & n21453;
  assign n21455 = n21454 ^ n19203;
  assign n21456 = n21215 & n21216;
  assign n21457 = n21220 & ~n21221;
  assign n21458 = n21223 & n21457;
  assign n21459 = ~n21224 & ~n21265;
  assign n21460 = n21221 & ~n21459;
  assign n21461 = ~n21222 & ~n21460;
  assign n21462 = ~n21236 & n21461;
  assign n21463 = ~n21458 & n21462;
  assign n21464 = n21456 & ~n21463;
  assign n21465 = n21215 & ~n21216;
  assign n21466 = ~n21220 & n21264;
  assign n21467 = ~n21240 & ~n21458;
  assign n21468 = ~n21466 & n21467;
  assign n21469 = ~n21263 & n21468;
  assign n21470 = n21465 & ~n21469;
  assign n21471 = ~n21464 & ~n21470;
  assign n21472 = n21220 & ~n21223;
  assign n21473 = n21459 ^ n21221;
  assign n21474 = n21473 ^ n21221;
  assign n21475 = n21227 ^ n21221;
  assign n21476 = ~n21474 & ~n21475;
  assign n21477 = n21476 ^ n21221;
  assign n21478 = ~n21472 & n21477;
  assign n21479 = ~n21458 & n21478;
  assign n21480 = n21479 ^ n21216;
  assign n21481 = n21480 ^ n21479;
  assign n21482 = n21225 & n21265;
  assign n21483 = ~n21224 & ~n21264;
  assign n21484 = n21218 & ~n21483;
  assign n21485 = ~n21482 & ~n21484;
  assign n21486 = n21467 & n21485;
  assign n21487 = n21486 ^ n21479;
  assign n21488 = n21481 & n21487;
  assign n21489 = n21488 ^ n21479;
  assign n21490 = ~n21215 & n21489;
  assign n21491 = n21471 & ~n21490;
  assign n21492 = n21491 ^ n18463;
  assign n21493 = n20997 & ~n21433;
  assign n21494 = ~n21016 & ~n21017;
  assign n21495 = n20988 & n21494;
  assign n21496 = n20980 & ~n21495;
  assign n21497 = ~n21493 & ~n21496;
  assign n21498 = n20967 & ~n21282;
  assign n21499 = ~n20977 & n21293;
  assign n21500 = n20980 & ~n21499;
  assign n21501 = ~n20997 & ~n21000;
  assign n21502 = ~n20967 & n21293;
  assign n21503 = ~n21501 & ~n21502;
  assign n21504 = ~n21001 & ~n21503;
  assign n21505 = ~n21014 & ~n21504;
  assign n21506 = ~n21500 & ~n21505;
  assign n21509 = ~n21008 & n21287;
  assign n21510 = ~n20983 & n21509;
  assign n21507 = n21003 & ~n21009;
  assign n21508 = ~n21036 & n21507;
  assign n21511 = n21510 ^ n21508;
  assign n21512 = n21510 ^ n20994;
  assign n21513 = n21510 & n21512;
  assign n21514 = n21513 ^ n21510;
  assign n21515 = n21511 & n21514;
  assign n21516 = n21515 ^ n21513;
  assign n21517 = n21516 ^ n21510;
  assign n21518 = n21517 ^ n20994;
  assign n21519 = n21506 & n21518;
  assign n21520 = n21519 ^ n21506;
  assign n21521 = ~n21498 & n21520;
  assign n21522 = n21497 & n21521;
  assign n21523 = ~n21306 & n21522;
  assign n21524 = ~n20979 & n21523;
  assign n21525 = n21524 ^ n17691;
  assign n21526 = n21217 & ~n21260;
  assign n21527 = n21235 & ~n21270;
  assign n21528 = ~n21526 & ~n21527;
  assign n21529 = n21249 & n21465;
  assign n21530 = ~n21233 & n21456;
  assign n21531 = ~n21529 & ~n21530;
  assign n21532 = n21528 & n21531;
  assign n21533 = n21532 ^ n19614;
  assign n21534 = n21465 & ~n21479;
  assign n21535 = n21217 & ~n21462;
  assign n21536 = ~n21534 & ~n21535;
  assign n21537 = n21223 & n21236;
  assign n21538 = ~n21219 & n21264;
  assign n21539 = ~n21237 & ~n21538;
  assign n21540 = ~n21263 & n21539;
  assign n21541 = n21235 & ~n21540;
  assign n21542 = ~n21537 & ~n21541;
  assign n21543 = n21456 & ~n21486;
  assign n21544 = n21542 & ~n21543;
  assign n21545 = n21536 & n21544;
  assign n21546 = ~n21458 & n21545;
  assign n21547 = n21546 ^ n18102;
  assign n21548 = n20633 & n20641;
  assign n21549 = n20629 & ~n20696;
  assign n21550 = ~n21548 & ~n21549;
  assign n21551 = n20522 & n20620;
  assign n21552 = n20625 & n20654;
  assign n21553 = ~n21551 & ~n21552;
  assign n21554 = n20522 & n20647;
  assign n21555 = n20654 & n20668;
  assign n21556 = ~n21554 & ~n21555;
  assign n21557 = ~n20520 & n20657;
  assign n21558 = ~n20639 & ~n20652;
  assign n21559 = ~n20632 & n21558;
  assign n21560 = ~n20647 & n21559;
  assign n21561 = n20629 & ~n21560;
  assign n21562 = ~n20633 & n20644;
  assign n21563 = n20654 & ~n21562;
  assign n21564 = ~n21561 & ~n21563;
  assign n21565 = ~n21557 & n21564;
  assign n21566 = ~n20622 & n20696;
  assign n21567 = ~n20620 & n21566;
  assign n21568 = n20641 & ~n21567;
  assign n21569 = ~n20632 & n20702;
  assign n21570 = n20522 & ~n21569;
  assign n21571 = ~n21568 & ~n21570;
  assign n21572 = n21565 & n21571;
  assign n21573 = n21556 & n21572;
  assign n21574 = ~n20714 & n21573;
  assign n21575 = n20694 & n21574;
  assign n21576 = n21553 & n21575;
  assign n21577 = n21550 & n21576;
  assign n21578 = ~n20649 & n21577;
  assign n21579 = n21578 ^ n18486;
  assign n21580 = n20632 & n20641;
  assign n21581 = ~n20649 & n21559;
  assign n21582 = n20654 & ~n21581;
  assign n21583 = ~n21580 & ~n21582;
  assign n21584 = n20522 & ~n20634;
  assign n21586 = ~n20620 & ~n20647;
  assign n21585 = n20626 & ~n20633;
  assign n21587 = n21586 ^ n21585;
  assign n21588 = n21587 ^ n21586;
  assign n21589 = n21586 ^ n20521;
  assign n21590 = n21589 ^ n21586;
  assign n21591 = ~n21588 & ~n21590;
  assign n21592 = n21591 ^ n21586;
  assign n21593 = n20520 & ~n21592;
  assign n21594 = n21593 ^ n21586;
  assign n21595 = ~n21584 & n21594;
  assign n21596 = n21583 & n21595;
  assign n21597 = n21556 & n21596;
  assign n21598 = n21553 & n21597;
  assign n21599 = n21550 & n21598;
  assign n21600 = n20646 & n21599;
  assign n21601 = n20691 & n21600;
  assign n21602 = ~n20687 & n21601;
  assign n21603 = ~n20674 & n21602;
  assign n21604 = n21603 ^ n17984;
  assign n21605 = n19522 & ~n19558;
  assign n21606 = n18794 & ~n19528;
  assign n21607 = ~n21605 & ~n21606;
  assign n21608 = n19500 & ~n20804;
  assign n21609 = ~n19489 & n21321;
  assign n21610 = n19491 & ~n21609;
  assign n21611 = n19517 & n20810;
  assign n21612 = n19500 & ~n21611;
  assign n21613 = n19526 & n19537;
  assign n21614 = n19522 & ~n21613;
  assign n21615 = ~n21612 & ~n21614;
  assign n21616 = ~n19535 & n20809;
  assign n21617 = ~n19510 & n21616;
  assign n21618 = ~n18794 & n21617;
  assign n21619 = ~n19491 & ~n20821;
  assign n21620 = n20814 & ~n21619;
  assign n21621 = ~n21618 & n21620;
  assign n21622 = n21615 & ~n21621;
  assign n21623 = ~n21610 & n21622;
  assign n21624 = ~n21608 & n21623;
  assign n21625 = n21607 & n21624;
  assign n21626 = n20800 & n21625;
  assign n21627 = n19534 & n21626;
  assign n21628 = n21627 ^ n18938;
  assign y0 = n18059;
  assign y1 = n19570;
  assign y2 = n18792;
  assign y3 = n19909;
  assign y4 = n19944;
  assign y5 = n19983;
  assign y6 = n20013;
  assign y7 = n20212;
  assign y8 = n20239;
  assign y9 = n20279;
  assign y10 = n20313;
  assign y11 = n20469;
  assign y12 = n20500;
  assign y13 = n20685;
  assign y14 = n20387;
  assign y15 = n20720;
  assign y16 = n20752;
  assign y17 = n20778;
  assign y18 = n20797;
  assign y19 = n20829;
  assign y20 = n20856;
  assign y21 = n20900;
  assign y22 = n20354;
  assign y23 = n20926;
  assign y24 = n20519;
  assign y25 = n20964;
  assign y26 = n19598;
  assign y27 = n21047;
  assign y28 = n18446;
  assign y29 = n21080;
  assign y30 = n20040;
  assign y31 = n21159;
  assign y32 = n20617;
  assign y33 = n21196;
  assign y34 = n19725;
  assign y35 = n21214;
  assign y36 = n19139;
  assign y37 = n21276;
  assign y38 = n20143;
  assign y39 = n21311;
  assign y40 = n20556;
  assign y41 = n21341;
  assign y42 = n19766;
  assign y43 = n21378;
  assign y44 = n19012;
  assign y45 = n21410;
  assign y46 = n20077;
  assign y47 = n21427;
  assign y48 = n20581;
  assign y49 = n21455;
  assign y50 = n19799;
  assign y51 = n21492;
  assign y52 = n19486;
  assign y53 = n21525;
  assign y54 = n20116;
  assign y55 = n21533;
  assign y56 = n20322;
  assign y57 = n21547;
  assign y58 = n19835;
  assign y59 = n21579;
  assign y60 = n19347;
  assign y61 = n21604;
  assign y62 = n20106;
  assign y63 = n21628;
endmodule
