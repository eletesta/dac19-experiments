module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831, x832, x833, x834, x835, x836, x837, x838, x839, x840, x841, x842, x843, x844, x845, x846, x847, x848, x849, x850, x851, x852, x853, x854, x855, x856, x857, x858, x859, x860, x861, x862, x863, x864, x865, x866, x867, x868, x869, x870, x871, x872, x873, x874, x875, x876, x877, x878, x879, x880, x881, x882, x883, x884, x885, x886, x887, x888, x889, x890, x891, x892, x893, x894, x895, x896, x897, x898, x899, x900, x901, x902, x903, x904, x905, x906, x907, x908, x909, x910, x911, x912, x913, x914, x915, x916, x917, x918, x919, x920, x921, x922, x923, x924, x925, x926, x927, x928, x929, x930, x931, x932, x933, x934, x935, x936, x937, x938, x939, x940, x941, x942, x943, x944, x945, x946, x947, x948, x949, x950, x951, x952, x953, x954, x955, x956, x957, x958, x959, x960, x961, x962, x963, x964, x965, x966, x967, x968, x969, x970, x971, x972, x973, x974, x975, x976, x977, x978, x979, x980, x981, x982, x983, x984, x985, x986, x987, x988, x989, x990, x991, x992, x993, x994, x995, x996, x997, x998, x999, x1000, x1001, x1002, x1003, x1004, x1005, x1006, x1007, x1008, x1009, x1010, x1011, x1012, x1013, x1014, x1015, x1016, x1017, x1018, x1019, x1020, x1021, x1022, x1023, x1024, x1025, x1026, x1027, x1028, x1029, x1030, x1031, x1032, x1033, x1034, x1035, x1036, x1037, x1038, x1039, x1040, x1041, x1042, x1043, x1044, x1045, x1046, x1047, x1048, x1049, x1050, x1051, x1052, x1053, x1054, x1055, x1056, x1057, x1058, x1059, x1060, x1061, x1062, x1063, x1064, x1065, x1066, x1067, x1068, x1069, x1070, x1071, x1072, x1073, x1074, x1075, x1076, x1077, x1078, x1079, x1080, x1081, x1082, x1083, x1084, x1085, x1086, x1087, x1088, x1089, x1090, x1091, x1092, x1093, x1094, x1095, x1096, x1097, x1098, x1099, x1100, x1101, x1102, x1103, x1104, x1105, x1106, x1107, x1108, x1109, x1110, x1111, x1112, x1113, x1114, x1115, x1116, x1117, x1118, x1119, x1120, x1121, x1122, x1123, x1124, x1125, x1126, x1127, x1128, x1129, x1130, x1131, x1132, x1133, x1134, x1135, x1136, x1137, x1138, x1139, x1140, x1141, x1142, x1143, x1144, x1145, x1146, x1147, x1148, x1149, x1150, x1151, x1152, x1153, x1154, x1155, x1156, x1157, x1158, x1159, x1160, x1161, x1162, x1163, x1164, x1165, x1166, x1167, x1168, x1169, x1170, x1171, x1172, x1173, x1174, x1175, x1176, x1177, x1178, x1179, x1180, x1181, x1182, x1183, x1184, x1185, x1186, x1187, x1188, x1189, x1190, x1191, x1192, x1193, x1194, x1195, x1196, x1197, x1198, x1199, x1200, x1201, x1202, x1203, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141, y142, y143, y144, y145, y146, y147, y148, y149, y150, y151, y152, y153, y154, y155, y156, y157, y158, y159, y160, y161, y162, y163, y164, y165, y166, y167, y168, y169, y170, y171, y172, y173, y174, y175, y176, y177, y178, y179, y180, y181, y182, y183, y184, y185, y186, y187, y188, y189, y190, y191, y192, y193, y194, y195, y196, y197, y198, y199, y200, y201, y202, y203, y204, y205, y206, y207, y208, y209, y210, y211, y212, y213, y214, y215, y216, y217, y218, y219, y220, y221, y222, y223, y224, y225, y226, y227, y228, y229, y230, y231, y232, y233, y234, y235, y236, y237, y238, y239, y240, y241, y242, y243, y244, y245, y246, y247, y248, y249, y250, y251, y252, y253, y254, y255, y256, y257, y258, y259, y260, y261, y262, y263, y264, y265, y266, y267, y268, y269, y270, y271, y272, y273, y274, y275, y276, y277, y278, y279, y280, y281, y282, y283, y284, y285, y286, y287, y288, y289, y290, y291, y292, y293, y294, y295, y296, y297, y298, y299, y300, y301, y302, y303, y304, y305, y306, y307, y308, y309, y310, y311, y312, y313, y314, y315, y316, y317, y318, y319, y320, y321, y322, y323, y324, y325, y326, y327, y328, y329, y330, y331, y332, y333, y334, y335, y336, y337, y338, y339, y340, y341, y342, y343, y344, y345, y346, y347, y348, y349, y350, y351, y352, y353, y354, y355, y356, y357, y358, y359, y360, y361, y362, y363, y364, y365, y366, y367, y368, y369, y370, y371, y372, y373, y374, y375, y376, y377, y378, y379, y380, y381, y382, y383, y384, y385, y386, y387, y388, y389, y390, y391, y392, y393, y394, y395, y396, y397, y398, y399, y400, y401, y402, y403, y404, y405, y406, y407, y408, y409, y410, y411, y412, y413, y414, y415, y416, y417, y418, y419, y420, y421, y422, y423, y424, y425, y426, y427, y428, y429, y430, y431, y432, y433, y434, y435, y436, y437, y438, y439, y440, y441, y442, y443, y444, y445, y446, y447, y448, y449, y450, y451, y452, y453, y454, y455, y456, y457, y458, y459, y460, y461, y462, y463, y464, y465, y466, y467, y468, y469, y470, y471, y472, y473, y474, y475, y476, y477, y478, y479, y480, y481, y482, y483, y484, y485, y486, y487, y488, y489, y490, y491, y492, y493, y494, y495, y496, y497, y498, y499, y500, y501, y502, y503, y504, y505, y506, y507, y508, y509, y510, y511, y512, y513, y514, y515, y516, y517, y518, y519, y520, y521, y522, y523, y524, y525, y526, y527, y528, y529, y530, y531, y532, y533, y534, y535, y536, y537, y538, y539, y540, y541, y542, y543, y544, y545, y546, y547, y548, y549, y550, y551, y552, y553, y554, y555, y556, y557, y558, y559, y560, y561, y562, y563, y564, y565, y566, y567, y568, y569, y570, y571, y572, y573, y574, y575, y576, y577, y578, y579, y580, y581, y582, y583, y584, y585, y586, y587, y588, y589, y590, y591, y592, y593, y594, y595, y596, y597, y598, y599, y600, y601, y602, y603, y604, y605, y606, y607, y608, y609, y610, y611, y612, y613, y614, y615, y616, y617, y618, y619, y620, y621, y622, y623, y624, y625, y626, y627, y628, y629, y630, y631, y632, y633, y634, y635, y636, y637, y638, y639, y640, y641, y642, y643, y644, y645, y646, y647, y648, y649, y650, y651, y652, y653, y654, y655, y656, y657, y658, y659, y660, y661, y662, y663, y664, y665, y666, y667, y668, y669, y670, y671, y672, y673, y674, y675, y676, y677, y678, y679, y680, y681, y682, y683, y684, y685, y686, y687, y688, y689, y690, y691, y692, y693, y694, y695, y696, y697, y698, y699, y700, y701, y702, y703, y704, y705, y706, y707, y708, y709, y710, y711, y712, y713, y714, y715, y716, y717, y718, y719, y720, y721, y722, y723, y724, y725, y726, y727, y728, y729, y730, y731, y732, y733, y734, y735, y736, y737, y738, y739, y740, y741, y742, y743, y744, y745, y746, y747, y748, y749, y750, y751, y752, y753, y754, y755, y756, y757, y758, y759, y760, y761, y762, y763, y764, y765, y766, y767, y768, y769, y770, y771, y772, y773, y774, y775, y776, y777, y778, y779, y780, y781, y782, y783, y784, y785, y786, y787, y788, y789, y790, y791, y792, y793, y794, y795, y796, y797, y798, y799, y800, y801, y802, y803, y804, y805, y806, y807, y808, y809, y810, y811, y812, y813, y814, y815, y816, y817, y818, y819, y820, y821, y822, y823, y824, y825, y826, y827, y828, y829, y830, y831, y832, y833, y834, y835, y836, y837, y838, y839, y840, y841, y842, y843, y844, y845, y846, y847, y848, y849, y850, y851, y852, y853, y854, y855, y856, y857, y858, y859, y860, y861, y862, y863, y864, y865, y866, y867, y868, y869, y870, y871, y872, y873, y874, y875, y876, y877, y878, y879, y880, y881, y882, y883, y884, y885, y886, y887, y888, y889, y890, y891, y892, y893, y894, y895, y896, y897, y898, y899, y900, y901, y902, y903, y904, y905, y906, y907, y908, y909, y910, y911, y912, y913, y914, y915, y916, y917, y918, y919, y920, y921, y922, y923, y924, y925, y926, y927, y928, y929, y930, y931, y932, y933, y934, y935, y936, y937, y938, y939, y940, y941, y942, y943, y944, y945, y946, y947, y948, y949, y950, y951, y952, y953, y954, y955, y956, y957, y958, y959, y960, y961, y962, y963, y964, y965, y966, y967, y968, y969, y970, y971, y972, y973, y974, y975, y976, y977, y978, y979, y980, y981, y982, y983, y984, y985, y986, y987, y988, y989, y990, y991, y992, y993, y994, y995, y996, y997, y998, y999, y1000, y1001, y1002, y1003, y1004, y1005, y1006, y1007, y1008, y1009, y1010, y1011, y1012, y1013, y1014, y1015, y1016, y1017, y1018, y1019, y1020, y1021, y1022, y1023, y1024, y1025, y1026, y1027, y1028, y1029, y1030, y1031, y1032, y1033, y1034, y1035, y1036, y1037, y1038, y1039, y1040, y1041, y1042, y1043, y1044, y1045, y1046, y1047, y1048, y1049, y1050, y1051, y1052, y1053, y1054, y1055, y1056, y1057, y1058, y1059, y1060, y1061, y1062, y1063, y1064, y1065, y1066, y1067, y1068, y1069, y1070, y1071, y1072, y1073, y1074, y1075, y1076, y1077, y1078, y1079, y1080, y1081, y1082, y1083, y1084, y1085, y1086, y1087, y1088, y1089, y1090, y1091, y1092, y1093, y1094, y1095, y1096, y1097, y1098, y1099, y1100, y1101, y1102, y1103, y1104, y1105, y1106, y1107, y1108, y1109, y1110, y1111, y1112, y1113, y1114, y1115, y1116, y1117, y1118, y1119, y1120, y1121, y1122, y1123, y1124, y1125, y1126, y1127, y1128, y1129, y1130, y1131, y1132, y1133, y1134, y1135, y1136, y1137, y1138, y1139, y1140, y1141, y1142, y1143, y1144, y1145, y1146, y1147, y1148, y1149, y1150, y1151, y1152, y1153, y1154, y1155, y1156, y1157, y1158, y1159, y1160, y1161, y1162, y1163, y1164, y1165, y1166, y1167, y1168, y1169, y1170, y1171, y1172, y1173, y1174, y1175, y1176, y1177, y1178, y1179, y1180, y1181, y1182, y1183, y1184, y1185, y1186, y1187, y1188, y1189, y1190, y1191, y1192, y1193, y1194, y1195, y1196, y1197, y1198, y1199, y1200, y1201, y1202, y1203, y1204, y1205, y1206, y1207, y1208, y1209, y1210, y1211, y1212, y1213, y1214, y1215, y1216, y1217, y1218, y1219, y1220, y1221, y1222, y1223, y1224, y1225, y1226, y1227, y1228, y1229, y1230);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831, x832, x833, x834, x835, x836, x837, x838, x839, x840, x841, x842, x843, x844, x845, x846, x847, x848, x849, x850, x851, x852, x853, x854, x855, x856, x857, x858, x859, x860, x861, x862, x863, x864, x865, x866, x867, x868, x869, x870, x871, x872, x873, x874, x875, x876, x877, x878, x879, x880, x881, x882, x883, x884, x885, x886, x887, x888, x889, x890, x891, x892, x893, x894, x895, x896, x897, x898, x899, x900, x901, x902, x903, x904, x905, x906, x907, x908, x909, x910, x911, x912, x913, x914, x915, x916, x917, x918, x919, x920, x921, x922, x923, x924, x925, x926, x927, x928, x929, x930, x931, x932, x933, x934, x935, x936, x937, x938, x939, x940, x941, x942, x943, x944, x945, x946, x947, x948, x949, x950, x951, x952, x953, x954, x955, x956, x957, x958, x959, x960, x961, x962, x963, x964, x965, x966, x967, x968, x969, x970, x971, x972, x973, x974, x975, x976, x977, x978, x979, x980, x981, x982, x983, x984, x985, x986, x987, x988, x989, x990, x991, x992, x993, x994, x995, x996, x997, x998, x999, x1000, x1001, x1002, x1003, x1004, x1005, x1006, x1007, x1008, x1009, x1010, x1011, x1012, x1013, x1014, x1015, x1016, x1017, x1018, x1019, x1020, x1021, x1022, x1023, x1024, x1025, x1026, x1027, x1028, x1029, x1030, x1031, x1032, x1033, x1034, x1035, x1036, x1037, x1038, x1039, x1040, x1041, x1042, x1043, x1044, x1045, x1046, x1047, x1048, x1049, x1050, x1051, x1052, x1053, x1054, x1055, x1056, x1057, x1058, x1059, x1060, x1061, x1062, x1063, x1064, x1065, x1066, x1067, x1068, x1069, x1070, x1071, x1072, x1073, x1074, x1075, x1076, x1077, x1078, x1079, x1080, x1081, x1082, x1083, x1084, x1085, x1086, x1087, x1088, x1089, x1090, x1091, x1092, x1093, x1094, x1095, x1096, x1097, x1098, x1099, x1100, x1101, x1102, x1103, x1104, x1105, x1106, x1107, x1108, x1109, x1110, x1111, x1112, x1113, x1114, x1115, x1116, x1117, x1118, x1119, x1120, x1121, x1122, x1123, x1124, x1125, x1126, x1127, x1128, x1129, x1130, x1131, x1132, x1133, x1134, x1135, x1136, x1137, x1138, x1139, x1140, x1141, x1142, x1143, x1144, x1145, x1146, x1147, x1148, x1149, x1150, x1151, x1152, x1153, x1154, x1155, x1156, x1157, x1158, x1159, x1160, x1161, x1162, x1163, x1164, x1165, x1166, x1167, x1168, x1169, x1170, x1171, x1172, x1173, x1174, x1175, x1176, x1177, x1178, x1179, x1180, x1181, x1182, x1183, x1184, x1185, x1186, x1187, x1188, x1189, x1190, x1191, x1192, x1193, x1194, x1195, x1196, x1197, x1198, x1199, x1200, x1201, x1202, x1203;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141, y142, y143, y144, y145, y146, y147, y148, y149, y150, y151, y152, y153, y154, y155, y156, y157, y158, y159, y160, y161, y162, y163, y164, y165, y166, y167, y168, y169, y170, y171, y172, y173, y174, y175, y176, y177, y178, y179, y180, y181, y182, y183, y184, y185, y186, y187, y188, y189, y190, y191, y192, y193, y194, y195, y196, y197, y198, y199, y200, y201, y202, y203, y204, y205, y206, y207, y208, y209, y210, y211, y212, y213, y214, y215, y216, y217, y218, y219, y220, y221, y222, y223, y224, y225, y226, y227, y228, y229, y230, y231, y232, y233, y234, y235, y236, y237, y238, y239, y240, y241, y242, y243, y244, y245, y246, y247, y248, y249, y250, y251, y252, y253, y254, y255, y256, y257, y258, y259, y260, y261, y262, y263, y264, y265, y266, y267, y268, y269, y270, y271, y272, y273, y274, y275, y276, y277, y278, y279, y280, y281, y282, y283, y284, y285, y286, y287, y288, y289, y290, y291, y292, y293, y294, y295, y296, y297, y298, y299, y300, y301, y302, y303, y304, y305, y306, y307, y308, y309, y310, y311, y312, y313, y314, y315, y316, y317, y318, y319, y320, y321, y322, y323, y324, y325, y326, y327, y328, y329, y330, y331, y332, y333, y334, y335, y336, y337, y338, y339, y340, y341, y342, y343, y344, y345, y346, y347, y348, y349, y350, y351, y352, y353, y354, y355, y356, y357, y358, y359, y360, y361, y362, y363, y364, y365, y366, y367, y368, y369, y370, y371, y372, y373, y374, y375, y376, y377, y378, y379, y380, y381, y382, y383, y384, y385, y386, y387, y388, y389, y390, y391, y392, y393, y394, y395, y396, y397, y398, y399, y400, y401, y402, y403, y404, y405, y406, y407, y408, y409, y410, y411, y412, y413, y414, y415, y416, y417, y418, y419, y420, y421, y422, y423, y424, y425, y426, y427, y428, y429, y430, y431, y432, y433, y434, y435, y436, y437, y438, y439, y440, y441, y442, y443, y444, y445, y446, y447, y448, y449, y450, y451, y452, y453, y454, y455, y456, y457, y458, y459, y460, y461, y462, y463, y464, y465, y466, y467, y468, y469, y470, y471, y472, y473, y474, y475, y476, y477, y478, y479, y480, y481, y482, y483, y484, y485, y486, y487, y488, y489, y490, y491, y492, y493, y494, y495, y496, y497, y498, y499, y500, y501, y502, y503, y504, y505, y506, y507, y508, y509, y510, y511, y512, y513, y514, y515, y516, y517, y518, y519, y520, y521, y522, y523, y524, y525, y526, y527, y528, y529, y530, y531, y532, y533, y534, y535, y536, y537, y538, y539, y540, y541, y542, y543, y544, y545, y546, y547, y548, y549, y550, y551, y552, y553, y554, y555, y556, y557, y558, y559, y560, y561, y562, y563, y564, y565, y566, y567, y568, y569, y570, y571, y572, y573, y574, y575, y576, y577, y578, y579, y580, y581, y582, y583, y584, y585, y586, y587, y588, y589, y590, y591, y592, y593, y594, y595, y596, y597, y598, y599, y600, y601, y602, y603, y604, y605, y606, y607, y608, y609, y610, y611, y612, y613, y614, y615, y616, y617, y618, y619, y620, y621, y622, y623, y624, y625, y626, y627, y628, y629, y630, y631, y632, y633, y634, y635, y636, y637, y638, y639, y640, y641, y642, y643, y644, y645, y646, y647, y648, y649, y650, y651, y652, y653, y654, y655, y656, y657, y658, y659, y660, y661, y662, y663, y664, y665, y666, y667, y668, y669, y670, y671, y672, y673, y674, y675, y676, y677, y678, y679, y680, y681, y682, y683, y684, y685, y686, y687, y688, y689, y690, y691, y692, y693, y694, y695, y696, y697, y698, y699, y700, y701, y702, y703, y704, y705, y706, y707, y708, y709, y710, y711, y712, y713, y714, y715, y716, y717, y718, y719, y720, y721, y722, y723, y724, y725, y726, y727, y728, y729, y730, y731, y732, y733, y734, y735, y736, y737, y738, y739, y740, y741, y742, y743, y744, y745, y746, y747, y748, y749, y750, y751, y752, y753, y754, y755, y756, y757, y758, y759, y760, y761, y762, y763, y764, y765, y766, y767, y768, y769, y770, y771, y772, y773, y774, y775, y776, y777, y778, y779, y780, y781, y782, y783, y784, y785, y786, y787, y788, y789, y790, y791, y792, y793, y794, y795, y796, y797, y798, y799, y800, y801, y802, y803, y804, y805, y806, y807, y808, y809, y810, y811, y812, y813, y814, y815, y816, y817, y818, y819, y820, y821, y822, y823, y824, y825, y826, y827, y828, y829, y830, y831, y832, y833, y834, y835, y836, y837, y838, y839, y840, y841, y842, y843, y844, y845, y846, y847, y848, y849, y850, y851, y852, y853, y854, y855, y856, y857, y858, y859, y860, y861, y862, y863, y864, y865, y866, y867, y868, y869, y870, y871, y872, y873, y874, y875, y876, y877, y878, y879, y880, y881, y882, y883, y884, y885, y886, y887, y888, y889, y890, y891, y892, y893, y894, y895, y896, y897, y898, y899, y900, y901, y902, y903, y904, y905, y906, y907, y908, y909, y910, y911, y912, y913, y914, y915, y916, y917, y918, y919, y920, y921, y922, y923, y924, y925, y926, y927, y928, y929, y930, y931, y932, y933, y934, y935, y936, y937, y938, y939, y940, y941, y942, y943, y944, y945, y946, y947, y948, y949, y950, y951, y952, y953, y954, y955, y956, y957, y958, y959, y960, y961, y962, y963, y964, y965, y966, y967, y968, y969, y970, y971, y972, y973, y974, y975, y976, y977, y978, y979, y980, y981, y982, y983, y984, y985, y986, y987, y988, y989, y990, y991, y992, y993, y994, y995, y996, y997, y998, y999, y1000, y1001, y1002, y1003, y1004, y1005, y1006, y1007, y1008, y1009, y1010, y1011, y1012, y1013, y1014, y1015, y1016, y1017, y1018, y1019, y1020, y1021, y1022, y1023, y1024, y1025, y1026, y1027, y1028, y1029, y1030, y1031, y1032, y1033, y1034, y1035, y1036, y1037, y1038, y1039, y1040, y1041, y1042, y1043, y1044, y1045, y1046, y1047, y1048, y1049, y1050, y1051, y1052, y1053, y1054, y1055, y1056, y1057, y1058, y1059, y1060, y1061, y1062, y1063, y1064, y1065, y1066, y1067, y1068, y1069, y1070, y1071, y1072, y1073, y1074, y1075, y1076, y1077, y1078, y1079, y1080, y1081, y1082, y1083, y1084, y1085, y1086, y1087, y1088, y1089, y1090, y1091, y1092, y1093, y1094, y1095, y1096, y1097, y1098, y1099, y1100, y1101, y1102, y1103, y1104, y1105, y1106, y1107, y1108, y1109, y1110, y1111, y1112, y1113, y1114, y1115, y1116, y1117, y1118, y1119, y1120, y1121, y1122, y1123, y1124, y1125, y1126, y1127, y1128, y1129, y1130, y1131, y1132, y1133, y1134, y1135, y1136, y1137, y1138, y1139, y1140, y1141, y1142, y1143, y1144, y1145, y1146, y1147, y1148, y1149, y1150, y1151, y1152, y1153, y1154, y1155, y1156, y1157, y1158, y1159, y1160, y1161, y1162, y1163, y1164, y1165, y1166, y1167, y1168, y1169, y1170, y1171, y1172, y1173, y1174, y1175, y1176, y1177, y1178, y1179, y1180, y1181, y1182, y1183, y1184, y1185, y1186, y1187, y1188, y1189, y1190, y1191, y1192, y1193, y1194, y1195, y1196, y1197, y1198, y1199, y1200, y1201, y1202, y1203, y1204, y1205, y1206, y1207, y1208, y1209, y1210, y1211, y1212, y1213, y1214, y1215, y1216, y1217, y1218, y1219, y1220, y1221, y1222, y1223, y1224, y1225, y1226, y1227, y1228, y1229, y1230;
  wire n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909;
  assign n1205 = x32 & ~x95;
  assign n1206 = ~x85 & ~x106;
  assign n1207 = ~x76 & n1206;
  assign n1208 = ~x48 & ~x61;
  assign n1209 = n1207 & n1208;
  assign n1210 = ~x104 & n1209;
  assign n1211 = ~x89 & n1210;
  assign n1212 = ~x49 & n1211;
  assign n1213 = ~x45 & n1212;
  assign n1214 = ~x69 & ~x83;
  assign n1215 = ~x103 & n1214;
  assign n1216 = ~x82 & ~x111;
  assign n1217 = ~x36 & n1216;
  assign n1218 = ~x66 & n1217;
  assign n1219 = n1215 & n1218;
  assign n1220 = n1213 & n1219;
  assign n1221 = ~x73 & n1220;
  assign n1222 = ~x88 & ~x98;
  assign n1223 = ~x102 & ~x107;
  assign n1224 = n1222 & n1223;
  assign n1225 = ~x64 & ~x65;
  assign n1226 = ~x63 & n1225;
  assign n1227 = n1224 & n1226;
  assign n1228 = ~x81 & n1227;
  assign n1229 = n1221 & n1228;
  assign n1230 = ~x67 & ~x68;
  assign n1231 = ~x71 & ~x84;
  assign n1232 = n1230 & n1231;
  assign n1233 = n1229 & n1232;
  assign n1234 = ~x91 & ~x109;
  assign n1235 = ~x46 & ~x47;
  assign n1236 = n1234 & n1235;
  assign n1237 = ~x77 & ~x86;
  assign n1238 = ~x50 & ~x110;
  assign n1239 = n1237 & n1238;
  assign n1240 = n1236 & n1239;
  assign n1241 = ~x53 & ~x60;
  assign n1242 = ~x58 & n1241;
  assign n1243 = ~x97 & ~x108;
  assign n1244 = ~x94 & n1243;
  assign n1245 = n1242 & n1244;
  assign n1246 = n1240 & n1245;
  assign n1247 = n1233 & n1246;
  assign n1248 = ~x72 & ~x96;
  assign n1249 = ~x51 & ~x70;
  assign n1250 = n1248 & n1249;
  assign n1251 = ~x35 & ~x93;
  assign n1252 = ~x90 & n1251;
  assign n1253 = n1250 & n1252;
  assign n1254 = n1247 & n1253;
  assign n1255 = ~x40 & n1254;
  assign n1256 = n1205 & n1255;
  assign n1257 = x210 ^ x198;
  assign n1258 = x299 & n1257;
  assign n1259 = n1258 ^ x198;
  assign n1260 = ~x841 & ~n1259;
  assign n1261 = x225 & ~n1260;
  assign n1262 = n1256 & n1261;
  assign n1263 = n1247 & n1252;
  assign n1264 = ~x32 & ~x95;
  assign n1265 = ~x40 & n1264;
  assign n1266 = x51 & x70;
  assign n1267 = x72 & x96;
  assign n1268 = ~n1266 & ~n1267;
  assign n1269 = n1265 & n1268;
  assign n1270 = ~n1248 & ~n1249;
  assign n1271 = n1269 & ~n1270;
  assign n1272 = n1263 & n1271;
  assign n1273 = x96 & n1272;
  assign n1274 = x95 & ~x479;
  assign n1275 = ~n1273 & ~n1274;
  assign n1276 = n1250 & n1265;
  assign n1282 = ~x73 & ~x84;
  assign n1283 = ~x68 & n1282;
  assign n1284 = ~x66 & n1283;
  assign n1285 = n1213 & n1284;
  assign n1286 = n1215 & n1285;
  assign n1287 = ~x36 & ~x67;
  assign n1288 = x82 & x111;
  assign n1289 = n1287 & ~n1288;
  assign n1290 = x36 & x67;
  assign n1291 = n1216 & ~n1290;
  assign n1292 = ~n1289 & ~n1291;
  assign n1293 = n1286 & ~n1292;
  assign n1294 = n1216 & n1287;
  assign n1295 = n1215 & n1294;
  assign n1296 = ~n1293 & ~n1295;
  assign n1297 = x104 & ~n1209;
  assign n1298 = ~x49 & ~n1297;
  assign n1299 = ~n1211 & ~n1298;
  assign n1300 = x89 & ~n1210;
  assign n1301 = ~x45 & ~n1300;
  assign n1302 = ~n1299 & n1301;
  assign n1303 = ~n1212 & ~n1302;
  assign n1304 = x76 & ~n1206;
  assign n1305 = x85 & x106;
  assign n1306 = n1208 & ~n1305;
  assign n1307 = ~n1304 & n1306;
  assign n1308 = x61 ^ x48;
  assign n1309 = n1207 & n1308;
  assign n1310 = ~n1307 & ~n1309;
  assign n1311 = n1284 & ~n1310;
  assign n1312 = ~n1303 & n1311;
  assign n1313 = x68 & ~n1282;
  assign n1314 = ~n1284 & ~n1313;
  assign n1315 = x73 & x84;
  assign n1316 = ~x66 & ~n1315;
  assign n1317 = ~n1283 & ~n1316;
  assign n1318 = n1314 & ~n1317;
  assign n1319 = n1213 & n1318;
  assign n1320 = ~n1312 & ~n1319;
  assign n1321 = ~n1296 & ~n1320;
  assign n1322 = n1285 & n1294;
  assign n1323 = x83 ^ x69;
  assign n1324 = x103 ^ x83;
  assign n1325 = n1323 & ~n1324;
  assign n1326 = n1325 ^ x69;
  assign n1327 = n1322 & ~n1326;
  assign n1328 = ~n1321 & ~n1327;
  assign n1329 = n1229 & n1322;
  assign n1330 = ~x71 & ~x81;
  assign n1331 = n1227 & n1330;
  assign n1332 = ~n1329 & ~n1331;
  assign n1333 = ~n1328 & ~n1332;
  assign n1334 = n1221 & n1232;
  assign n1335 = ~x102 & n1232;
  assign n1336 = ~x81 & n1222;
  assign n1337 = n1335 & n1336;
  assign n1338 = x107 ^ x102;
  assign n1339 = x98 ^ x88;
  assign n1340 = ~n1338 & ~n1339;
  assign n1341 = ~n1222 & ~n1223;
  assign n1342 = ~n1340 & ~n1341;
  assign n1343 = n1342 ^ n1224;
  assign n1344 = ~x81 & n1343;
  assign n1345 = n1344 ^ n1224;
  assign n1346 = n1337 & ~n1345;
  assign n1347 = x64 & x65;
  assign n1348 = n1346 & ~n1347;
  assign n1349 = n1225 & n1345;
  assign n1350 = ~n1348 & ~n1349;
  assign n1351 = ~x63 & ~n1350;
  assign n1352 = n1225 & n1346;
  assign n1353 = ~n1351 & ~n1352;
  assign n1354 = n1334 & ~n1353;
  assign n1355 = ~n1333 & ~n1354;
  assign n1356 = ~x50 & n1241;
  assign n1357 = ~x77 & n1356;
  assign n1358 = n1243 & n1357;
  assign n1359 = ~x86 & ~x94;
  assign n1360 = n1358 & n1359;
  assign n1361 = ~n1355 & n1360;
  assign n1362 = n1357 ^ n1243;
  assign n1363 = x97 & x108;
  assign n1364 = n1359 & ~n1363;
  assign n1365 = n1364 ^ n1243;
  assign n1366 = n1362 & ~n1365;
  assign n1367 = n1366 ^ n1357;
  assign n1368 = n1233 & n1367;
  assign n1369 = ~n1361 & ~n1368;
  assign n1370 = x53 & x60;
  assign n1371 = ~x77 & ~n1370;
  assign n1372 = ~n1356 & ~n1371;
  assign n1373 = x50 & ~n1241;
  assign n1374 = ~x46 & ~x109;
  assign n1375 = ~n1373 & n1374;
  assign n1376 = ~n1372 & n1375;
  assign n1377 = ~n1369 & n1376;
  assign n1378 = x86 & x94;
  assign n1379 = n1377 & ~n1378;
  assign n1380 = n1233 & n1360;
  assign n1381 = n1379 & ~n1380;
  assign n1382 = ~x46 & ~n1234;
  assign n1383 = n1380 & n1382;
  assign n1384 = ~x58 & ~x90;
  assign n1385 = ~x47 & ~x110;
  assign n1386 = n1384 & n1385;
  assign n1387 = ~n1383 & n1386;
  assign n1388 = ~n1381 & n1387;
  assign n1389 = n1376 & n1380;
  assign n1390 = ~x91 & ~x93;
  assign n1391 = n1386 & n1390;
  assign n1392 = ~n1389 & ~n1391;
  assign n1393 = x91 ^ x47;
  assign n1394 = ~n1384 & n1393;
  assign n1395 = n1251 & ~n1394;
  assign n1396 = x91 & ~n1385;
  assign n1397 = n1395 & ~n1396;
  assign n1398 = ~x47 & n1384;
  assign n1399 = x58 & x90;
  assign n1400 = ~x110 & ~n1399;
  assign n1401 = ~n1398 & ~n1400;
  assign n1402 = n1397 & ~n1401;
  assign n1403 = ~n1392 & n1402;
  assign n1404 = ~n1388 & n1403;
  assign n1405 = ~x90 & n1247;
  assign n1406 = x93 ^ x35;
  assign n1407 = n1405 & n1406;
  assign n1408 = ~n1404 & ~n1407;
  assign n1409 = n1276 & ~n1408;
  assign n1410 = ~n1272 & ~n1409;
  assign n1277 = x40 ^ x32;
  assign n1278 = n1277 ^ x95;
  assign n1279 = x40 & x95;
  assign n1280 = n1278 & n1279;
  assign n1281 = n1280 ^ n1278;
  assign n1411 = n1410 ^ n1281;
  assign n1412 = n1254 & ~n1411;
  assign n1413 = n1412 ^ n1410;
  assign n1414 = ~n1276 & n1413;
  assign n1415 = x97 & n1391;
  assign n1416 = n1377 & n1415;
  assign n1417 = n1276 & n1391;
  assign n1418 = ~x35 & n1417;
  assign n1419 = n1416 & n1418;
  assign n1420 = ~n1273 & ~n1419;
  assign n1421 = x1091 & x1093;
  assign n1422 = ~x833 & x957;
  assign n1423 = n1421 & n1422;
  assign n1424 = ~x1091 & x1093;
  assign n1425 = ~n1423 & ~n1424;
  assign n1426 = x950 & x1092;
  assign n1427 = x829 & n1426;
  assign n1428 = n1425 & n1427;
  assign n1429 = ~x841 & n1428;
  assign n1430 = n1247 & n1429;
  assign n1431 = x1093 & n1428;
  assign n1432 = ~x46 & ~x94;
  assign n1433 = x97 ^ x36;
  assign n1434 = n1432 & n1433;
  assign n1435 = n1431 & n1434;
  assign n1436 = ~n1430 & ~n1435;
  assign n1437 = ~n1420 & ~n1436;
  assign n1438 = ~x174 & ~x189;
  assign n1439 = ~x144 & n1438;
  assign n1440 = ~x142 & ~x299;
  assign n1441 = ~n1439 & n1440;
  assign n1442 = ~x152 & ~x166;
  assign n1443 = ~x161 & n1442;
  assign n1444 = ~x146 & x299;
  assign n1445 = ~n1443 & n1444;
  assign n1446 = ~n1441 & ~n1445;
  assign n1447 = ~n1259 & n1446;
  assign n1448 = n1437 & n1447;
  assign n1449 = ~x35 & n1241;
  assign n1450 = ~x97 & ~n1449;
  assign n1451 = ~x137 & ~n1450;
  assign n1452 = ~n1448 & n1451;
  assign n1453 = n1385 & n1389;
  assign n1454 = ~x109 & ~x110;
  assign n1455 = ~n1235 & ~n1454;
  assign n1456 = n1380 & ~n1455;
  assign n1457 = ~n1453 & n1456;
  assign n1458 = n1384 & ~n1457;
  assign n1459 = n1403 & ~n1458;
  assign n1460 = ~x40 & ~x51;
  assign n1461 = n1248 & n1460;
  assign n1462 = n1251 & n1461;
  assign n1463 = ~x93 & x225;
  assign n1464 = x35 & ~n1463;
  assign n1465 = ~n1462 & ~n1464;
  assign n1466 = n1405 & n1465;
  assign n1467 = ~x95 & ~n1466;
  assign n1468 = ~n1459 & n1467;
  assign n1469 = ~n1404 & n1468;
  assign n1470 = ~n1452 & ~n1469;
  assign n1471 = ~n1414 & n1470;
  assign n1472 = n1471 ^ x234;
  assign n1473 = n1275 & n1472;
  assign n1474 = n1473 ^ x234;
  assign n1475 = ~n1262 & ~n1474;
  assign n1476 = ~x228 & ~n1413;
  assign n1477 = x105 & x228;
  assign n1478 = ~n1476 & ~n1477;
  assign n1479 = ~x216 & ~x221;
  assign n1480 = ~x215 & x299;
  assign n1481 = n1479 & n1480;
  assign n1482 = ~n1478 & n1481;
  assign n1483 = ~x223 & ~x224;
  assign n1484 = ~x222 & n1483;
  assign n1485 = ~x299 & n1484;
  assign n1486 = ~n1482 & ~n1485;
  assign n1487 = n1475 & ~n1486;
  assign n1488 = ~x215 & n1479;
  assign n1489 = ~n1478 & n1488;
  assign n1490 = ~x216 & x833;
  assign n1491 = ~x929 & n1490;
  assign n1492 = ~x221 & x265;
  assign n1493 = ~n1491 & ~n1492;
  assign n1494 = ~x215 & ~n1493;
  assign n1495 = x221 & ~n1490;
  assign n1496 = ~x215 & ~n1495;
  assign n1497 = ~x1144 & ~n1496;
  assign n1498 = ~n1494 & ~n1497;
  assign n1499 = ~x332 & ~n1498;
  assign n1500 = ~n1488 & ~n1499;
  assign n1501 = x299 & ~n1500;
  assign n1502 = x153 & ~n1477;
  assign n1503 = ~x332 & n1502;
  assign n1504 = n1488 & ~n1503;
  assign n1505 = n1501 & ~n1504;
  assign n1506 = ~n1489 & n1505;
  assign n1507 = ~n1487 & ~n1506;
  assign n1508 = ~x75 & ~x100;
  assign n1509 = ~x74 & n1508;
  assign n1510 = ~x38 & ~x54;
  assign n1511 = n1509 & n1510;
  assign n1512 = ~x87 & ~x92;
  assign n1513 = ~x39 & n1512;
  assign n1514 = n1511 & n1513;
  assign n1515 = ~x56 & ~x62;
  assign n1516 = ~x55 & n1515;
  assign n1517 = ~x57 & ~x59;
  assign n1518 = n1516 & n1517;
  assign n1519 = n1514 & n1518;
  assign n1520 = ~n1507 & n1519;
  assign n1521 = n1254 & n1265;
  assign n1522 = n1514 & n1521;
  assign n1523 = n1517 & n1522;
  assign n1524 = x57 & ~x59;
  assign n1525 = n1515 & n1524;
  assign n1526 = n1522 & n1525;
  assign n1527 = ~x55 & n1526;
  assign n1528 = n1518 & n1521;
  assign n1529 = ~x74 & ~x92;
  assign n1530 = ~x54 & n1529;
  assign n1531 = ~x87 & n1508;
  assign n1532 = n1530 & n1531;
  assign n1533 = x38 & ~x39;
  assign n1534 = n1532 & n1533;
  assign n1535 = n1528 & n1534;
  assign n1536 = ~x39 & ~x87;
  assign n1537 = ~x38 & n1536;
  assign n1538 = ~x92 & n1508;
  assign n1539 = n1537 & n1538;
  assign n1540 = ~x74 & n1539;
  assign n1541 = ~x57 & n1515;
  assign n1542 = x54 & x59;
  assign n1543 = n1541 & ~n1542;
  assign n1544 = ~x54 & ~x59;
  assign n1545 = n1544 ^ x55;
  assign n1546 = n1543 & ~n1545;
  assign n1547 = n1540 & n1546;
  assign n1548 = n1521 & n1547;
  assign n1549 = ~n1535 & ~n1548;
  assign n1550 = ~n1527 & n1549;
  assign n1551 = n1528 & n1537;
  assign n1552 = ~x54 & ~x75;
  assign n1553 = x92 ^ x74;
  assign n1554 = n1552 & n1553;
  assign n1555 = x75 ^ x54;
  assign n1556 = n1529 & n1555;
  assign n1557 = ~n1554 & ~n1556;
  assign n1558 = n1551 & ~n1557;
  assign n1559 = ~x100 & n1558;
  assign n1560 = n1550 & ~n1559;
  assign n1561 = x62 ^ x56;
  assign n1562 = ~x55 & n1561;
  assign n1563 = n1523 & n1562;
  assign n1564 = x92 ^ x87;
  assign n1565 = x100 ^ x39;
  assign n1566 = ~n1564 & ~n1565;
  assign n1567 = ~x39 & ~x100;
  assign n1568 = ~n1512 & ~n1567;
  assign n1569 = ~n1566 & ~n1568;
  assign n1570 = ~x74 & ~x75;
  assign n1571 = n1510 & n1570;
  assign n1572 = n1569 & n1571;
  assign n1573 = n1528 & n1572;
  assign n1574 = ~n1563 & ~n1573;
  assign n1575 = n1560 & n1574;
  assign n1576 = n1523 & ~n1575;
  assign n1577 = ~x228 & n1576;
  assign n1578 = n1488 & n1577;
  assign n1579 = n1488 & ~n1502;
  assign n1580 = ~n1578 & ~n1579;
  assign n1581 = x234 & n1274;
  assign n1582 = n1477 & ~n1581;
  assign n1583 = ~n1576 & n1582;
  assign n1584 = ~n1563 & ~n1583;
  assign n1585 = ~n1580 & n1584;
  assign n1586 = ~x105 & x228;
  assign n1587 = ~x137 & ~n1586;
  assign n1588 = n1488 & ~n1587;
  assign n1589 = ~x228 & n1517;
  assign n1590 = n1502 & ~n1589;
  assign n1591 = n1588 & ~n1590;
  assign n1592 = ~n1575 & n1591;
  assign n1593 = ~n1500 & ~n1518;
  assign n1594 = ~n1592 & n1593;
  assign n1595 = ~n1585 & n1594;
  assign n1596 = n1511 & n1564;
  assign n1597 = ~x39 & x252;
  assign n1598 = ~n1596 & n1597;
  assign n1599 = ~x146 & ~n1443;
  assign n1600 = n1598 & ~n1599;
  assign n1601 = ~x228 & n1572;
  assign n1602 = ~n1600 & n1601;
  assign n1603 = n1521 & n1602;
  assign n1604 = n1488 & n1603;
  assign n1605 = n1477 & n1481;
  assign n1606 = ~n1485 & ~n1605;
  assign n1607 = ~x332 & ~n1581;
  assign n1608 = ~n1606 & n1607;
  assign n1609 = ~n1604 & ~n1608;
  assign n1610 = ~x210 & ~n1599;
  assign n1611 = ~x137 & ~x332;
  assign n1612 = ~n1610 & n1611;
  assign n1613 = n1501 & n1612;
  assign n1614 = n1485 & n1611;
  assign n1615 = ~x142 & ~n1439;
  assign n1616 = ~x198 & ~n1615;
  assign n1617 = n1614 & ~n1616;
  assign n1618 = x100 ^ x75;
  assign n1619 = n1530 & n1618;
  assign n1620 = ~n1617 & n1619;
  assign n1621 = x137 & n1508;
  assign n1622 = ~n1557 & n1621;
  assign n1623 = ~n1620 & ~n1622;
  assign n1624 = ~n1613 & ~n1623;
  assign n1625 = n1521 & n1624;
  assign n1626 = n1537 & n1625;
  assign n1627 = ~n1609 & ~n1626;
  assign n1628 = n1505 & ~n1604;
  assign n1629 = ~n1627 & ~n1628;
  assign n1630 = ~n1505 & n1532;
  assign n1631 = ~n1596 & ~n1630;
  assign n1632 = ~x39 & ~n1631;
  assign n1633 = n1510 & n1529;
  assign n1634 = n1531 & n1633;
  assign n1635 = ~n1632 & ~n1634;
  assign n1636 = x153 & n1586;
  assign n1637 = n1588 & ~n1636;
  assign n1638 = ~x332 & ~n1637;
  assign n1639 = n1501 & n1638;
  assign n1640 = ~n1614 & ~n1639;
  assign n1641 = ~n1635 & n1640;
  assign n1642 = n1521 & n1641;
  assign n1643 = ~n1514 & n1518;
  assign n1644 = ~n1642 & n1643;
  assign n1645 = ~n1629 & n1644;
  assign n1646 = ~x224 & x833;
  assign n1647 = x222 & ~n1646;
  assign n1648 = ~x223 & ~n1647;
  assign n1649 = x1144 & ~n1648;
  assign n1650 = x929 & n1646;
  assign n1651 = x224 & x265;
  assign n1652 = ~x222 & ~n1651;
  assign n1653 = ~n1650 & ~n1652;
  assign n1654 = ~x223 & ~n1653;
  assign n1655 = ~n1649 & ~n1654;
  assign n1656 = ~x299 & n1518;
  assign n1657 = n1655 & n1656;
  assign n1658 = ~n1645 & ~n1657;
  assign n1659 = ~n1595 & n1658;
  assign n1660 = ~n1520 & n1659;
  assign n1661 = ~x332 & ~n1660;
  assign n1662 = ~n1413 & n1519;
  assign n1663 = ~n1576 & ~n1662;
  assign n1664 = ~x228 & ~n1663;
  assign n1665 = n1518 & n1603;
  assign n1666 = ~n1664 & ~n1665;
  assign n1667 = n1488 & ~n1666;
  assign n1668 = ~n1656 & ~n1667;
  assign n1669 = ~n1477 & n1488;
  assign n1670 = ~x154 & n1669;
  assign n1671 = ~x215 & x221;
  assign n1672 = n1490 & n1671;
  assign n1673 = x939 & n1672;
  assign n1674 = x216 & ~x221;
  assign n1675 = ~x215 & n1674;
  assign n1676 = x276 & n1675;
  assign n1677 = ~n1673 & ~n1676;
  assign n1678 = ~n1670 & n1677;
  assign n1679 = x1146 & ~n1496;
  assign n1680 = n1678 & ~n1679;
  assign n1681 = n1477 & n1488;
  assign n1682 = n1274 & n1681;
  assign n1683 = x239 & n1682;
  assign n1684 = n1680 & ~n1683;
  assign n1685 = n1668 & ~n1684;
  assign n1686 = n1488 & n1514;
  assign n1687 = x299 & n1686;
  assign n1688 = ~n1275 & n1687;
  assign n1689 = n1476 & n1688;
  assign n1690 = ~n1274 & ~n1514;
  assign n1691 = ~n1275 & ~n1690;
  assign n1692 = ~n1606 & n1691;
  assign n1693 = ~n1689 & ~n1692;
  assign n1694 = x239 & ~n1693;
  assign n1695 = ~x299 & ~n1648;
  assign n1696 = x1146 & n1695;
  assign n1697 = ~x223 & ~x299;
  assign n1698 = x222 & n1697;
  assign n1699 = n1646 & n1698;
  assign n1700 = x939 & n1699;
  assign n1701 = x224 & n1697;
  assign n1702 = ~x222 & n1701;
  assign n1703 = x276 & n1702;
  assign n1704 = ~n1700 & ~n1703;
  assign n1705 = ~n1696 & n1704;
  assign n1706 = ~n1694 & n1705;
  assign n1707 = n1518 & ~n1706;
  assign n1708 = ~n1685 & ~n1707;
  assign n1709 = x274 & n1675;
  assign n1710 = ~x151 & n1669;
  assign n1711 = n1710 ^ n1488;
  assign n1712 = ~n1709 & ~n1711;
  assign n1713 = ~x927 & n1672;
  assign n1714 = n1712 & ~n1713;
  assign n1715 = ~x1145 & ~n1496;
  assign n1716 = n1714 & ~n1715;
  assign n1717 = x235 & n1682;
  assign n1718 = ~n1716 & ~n1717;
  assign n1719 = n1668 & ~n1718;
  assign n1720 = x235 & ~n1693;
  assign n1721 = x1145 & n1695;
  assign n1722 = ~x274 & n1702;
  assign n1723 = x927 & n1699;
  assign n1724 = ~n1722 & ~n1723;
  assign n1725 = ~n1721 & n1724;
  assign n1726 = ~n1720 & n1725;
  assign n1727 = n1518 & ~n1726;
  assign n1728 = ~n1719 & ~n1727;
  assign n1729 = x284 & n1275;
  assign n1730 = n1729 ^ x146;
  assign n1731 = ~n1478 & ~n1730;
  assign n1732 = n1731 ^ x146;
  assign n1733 = n1686 & n1732;
  assign n1734 = ~n1274 & n1681;
  assign n1735 = ~x284 & n1734;
  assign n1736 = ~x264 & n1675;
  assign n1737 = x944 & n1672;
  assign n1738 = ~n1736 & ~n1737;
  assign n1739 = ~n1735 & n1738;
  assign n1740 = x146 & n1669;
  assign n1741 = x1143 & ~n1496;
  assign n1742 = ~n1740 & ~n1741;
  assign n1743 = n1739 & n1742;
  assign n1744 = ~n1604 & ~n1743;
  assign n1745 = x299 & ~n1744;
  assign n1746 = ~n1477 & ~n1603;
  assign n1747 = x284 & ~n1274;
  assign n1748 = n1488 & ~n1747;
  assign n1749 = ~n1586 & n1748;
  assign n1750 = ~n1746 & n1749;
  assign n1751 = n1745 & ~n1750;
  assign n1752 = ~n1687 & ~n1751;
  assign n1753 = ~n1733 & ~n1752;
  assign n1754 = ~x238 & ~n1693;
  assign n1755 = x284 & n1485;
  assign n1756 = ~n1691 & n1755;
  assign n1757 = x264 & n1702;
  assign n1758 = n1518 & ~n1757;
  assign n1759 = ~x944 & n1699;
  assign n1760 = n1758 & ~n1759;
  assign n1761 = ~x1143 & n1695;
  assign n1762 = n1760 & ~n1761;
  assign n1763 = ~n1756 & n1762;
  assign n1764 = ~n1754 & n1763;
  assign n1765 = ~n1753 & n1764;
  assign n1766 = x228 & x238;
  assign n1767 = ~n1578 & ~n1766;
  assign n1768 = n1749 & ~n1767;
  assign n1769 = ~n1578 & ~n1743;
  assign n1770 = ~n1768 & ~n1769;
  assign n1771 = ~n1518 & ~n1770;
  assign n1772 = ~n1765 & ~n1771;
  assign n1773 = ~n1477 & ~n1577;
  assign n1774 = ~n1665 & n1773;
  assign n1775 = ~x262 & ~n1774;
  assign n1776 = ~x172 & n1773;
  assign n1777 = n1274 & n1477;
  assign n1778 = ~n1776 & ~n1777;
  assign n1779 = ~n1775 & n1778;
  assign n1780 = n1488 & ~n1779;
  assign n1781 = ~x1142 & ~n1490;
  assign n1782 = x221 & ~n1781;
  assign n1783 = ~x932 & n1490;
  assign n1784 = n1782 & ~n1783;
  assign n1785 = ~x277 & n1674;
  assign n1786 = ~n1784 & ~n1785;
  assign n1787 = n1786 ^ x1142;
  assign n1788 = ~x215 & ~n1787;
  assign n1789 = n1788 ^ x1142;
  assign n1790 = ~n1780 & ~n1789;
  assign n1791 = x262 & n1518;
  assign n1792 = n1604 & n1791;
  assign n1793 = ~x249 & n1274;
  assign n1794 = n1681 & n1793;
  assign n1795 = ~n1656 & ~n1794;
  assign n1796 = ~n1792 & n1795;
  assign n1797 = ~n1790 & n1796;
  assign n1798 = x262 & ~n1691;
  assign n1799 = n1485 & ~n1793;
  assign n1800 = ~n1798 & n1799;
  assign n1801 = x1142 & n1695;
  assign n1802 = ~x277 & n1702;
  assign n1803 = x932 & n1699;
  assign n1804 = ~n1802 & ~n1803;
  assign n1805 = ~n1801 & n1804;
  assign n1806 = ~n1800 & n1805;
  assign n1807 = n1518 & ~n1806;
  assign n1808 = ~n1797 & ~n1807;
  assign n1809 = ~x249 & ~n1275;
  assign n1810 = n1485 & n1809;
  assign n1811 = n1480 & n1786;
  assign n1812 = ~n1810 & ~n1811;
  assign n1813 = n1519 & ~n1812;
  assign n1814 = ~n1808 & ~n1813;
  assign n1815 = x172 & n1478;
  assign n1816 = n1481 & n1813;
  assign n1817 = ~n1815 & n1816;
  assign n1818 = x262 ^ x249;
  assign n1819 = n1275 & ~n1818;
  assign n1820 = n1819 ^ x249;
  assign n1821 = ~n1478 & ~n1820;
  assign n1822 = n1817 & ~n1821;
  assign n1823 = ~n1814 & ~n1822;
  assign n1824 = x171 & n1669;
  assign n1825 = x861 & ~n1274;
  assign n1826 = n1681 & ~n1825;
  assign n1827 = ~n1824 & ~n1826;
  assign n1828 = ~x935 & n1672;
  assign n1829 = x270 & n1675;
  assign n1830 = ~n1828 & ~n1829;
  assign n1831 = ~x1141 & ~n1496;
  assign n1832 = n1830 & ~n1831;
  assign n1833 = n1827 & n1832;
  assign n1834 = ~n1489 & ~n1833;
  assign n1835 = n1514 & ~n1834;
  assign n1836 = x299 & ~n1835;
  assign n1837 = ~n1273 & n1825;
  assign n1838 = ~n1486 & ~n1837;
  assign n1839 = ~n1836 & ~n1838;
  assign n1840 = n1833 ^ x861;
  assign n1841 = ~n1604 & n1840;
  assign n1842 = n1841 ^ x861;
  assign n1843 = x299 & ~n1842;
  assign n1844 = ~x299 & ~n1825;
  assign n1845 = ~n1514 & ~n1844;
  assign n1846 = ~n1843 & n1845;
  assign n1847 = ~n1839 & ~n1846;
  assign n1848 = ~x1141 & n1695;
  assign n1849 = ~x935 & n1699;
  assign n1850 = x270 & n1702;
  assign n1851 = ~n1849 & ~n1850;
  assign n1852 = ~n1848 & n1851;
  assign n1853 = ~n1847 & n1852;
  assign n1854 = x241 & ~n1693;
  assign n1855 = n1518 & ~n1854;
  assign n1856 = ~n1853 & n1855;
  assign n1857 = ~n1578 & n1833;
  assign n1858 = ~n1518 & ~n1682;
  assign n1859 = ~x241 & ~n1518;
  assign n1860 = ~n1858 & ~n1859;
  assign n1861 = ~n1857 & ~n1860;
  assign n1862 = x861 & n1578;
  assign n1863 = n1861 & ~n1862;
  assign n1864 = ~n1856 & ~n1863;
  assign n1865 = n1476 & n1514;
  assign n1866 = n1746 & ~n1865;
  assign n1867 = x869 & ~n1866;
  assign n1868 = n1488 & ~n1867;
  assign n1869 = ~x170 & n1866;
  assign n1870 = n1868 & ~n1869;
  assign n1871 = x1140 & ~n1496;
  assign n1872 = x921 & n1490;
  assign n1873 = x216 & x282;
  assign n1874 = ~x221 & ~n1873;
  assign n1875 = ~n1872 & ~n1874;
  assign n1876 = ~x215 & ~n1875;
  assign n1877 = ~n1871 & ~n1876;
  assign n1878 = x299 & ~n1877;
  assign n1879 = ~n1870 & n1878;
  assign n1880 = x1140 & n1695;
  assign n1881 = x869 & ~n1274;
  assign n1882 = n1485 & n1881;
  assign n1883 = ~n1880 & ~n1882;
  assign n1884 = x921 & n1699;
  assign n1885 = ~x282 & n1702;
  assign n1886 = ~n1884 & ~n1885;
  assign n1887 = n1883 & n1886;
  assign n1888 = ~n1879 & n1887;
  assign n1889 = n1518 & n1693;
  assign n1890 = ~n1888 & n1889;
  assign n1891 = x248 & ~n1858;
  assign n1892 = ~n1889 & n1891;
  assign n1893 = ~n1578 & ~n1734;
  assign n1894 = x869 & ~n1893;
  assign n1895 = ~x170 & n1669;
  assign n1896 = n1895 ^ n1488;
  assign n1897 = ~n1877 & ~n1896;
  assign n1898 = ~n1578 & n1897;
  assign n1899 = ~n1894 & ~n1898;
  assign n1900 = ~n1518 & ~n1899;
  assign n1901 = ~n1892 & ~n1900;
  assign n1902 = ~n1890 & n1901;
  assign n1903 = ~x148 & n1478;
  assign n1904 = n1687 & ~n1903;
  assign n1905 = x862 ^ x247;
  assign n1906 = n1275 & n1905;
  assign n1907 = n1906 ^ x247;
  assign n1908 = ~n1478 & n1907;
  assign n1909 = n1904 & ~n1908;
  assign n1910 = ~n1691 & n1905;
  assign n1911 = n1910 ^ x247;
  assign n1912 = n1485 & ~n1911;
  assign n1913 = x148 & n1669;
  assign n1914 = ~x920 & n1672;
  assign n1915 = ~n1913 & ~n1914;
  assign n1916 = ~x1139 & ~n1496;
  assign n1917 = x281 & n1675;
  assign n1918 = ~n1916 & ~n1917;
  assign n1919 = n1915 & n1918;
  assign n1920 = ~x862 & n1734;
  assign n1921 = ~x247 & n1682;
  assign n1922 = ~n1920 & ~n1921;
  assign n1923 = n1919 & n1922;
  assign n1924 = ~n1686 & ~n1923;
  assign n1925 = n1924 ^ x862;
  assign n1926 = ~n1604 & ~n1925;
  assign n1927 = n1926 ^ x862;
  assign n1928 = x299 & ~n1927;
  assign n1929 = x281 & n1702;
  assign n1930 = n1518 & ~n1929;
  assign n1931 = ~x920 & n1699;
  assign n1932 = n1930 & ~n1931;
  assign n1933 = ~x1139 & n1695;
  assign n1934 = n1932 & ~n1933;
  assign n1935 = ~n1928 & n1934;
  assign n1936 = ~n1912 & n1935;
  assign n1937 = ~n1909 & n1936;
  assign n1938 = ~n1578 & ~n1923;
  assign n1939 = ~n1518 & ~n1938;
  assign n1940 = ~x862 & n1578;
  assign n1941 = n1939 & ~n1940;
  assign n1942 = ~n1937 & ~n1941;
  assign n1943 = x877 ^ x246;
  assign n1944 = n1275 & n1943;
  assign n1945 = n1944 ^ x246;
  assign n1946 = n1945 ^ x169;
  assign n1947 = ~n1478 & ~n1946;
  assign n1948 = n1947 ^ x169;
  assign n1949 = n1514 & ~n1948;
  assign n1950 = x877 & ~n1274;
  assign n1951 = n1950 ^ x169;
  assign n1952 = ~n1746 & ~n1951;
  assign n1953 = n1952 ^ x169;
  assign n1954 = n1488 & n1953;
  assign n1955 = ~n1686 & ~n1954;
  assign n1956 = ~n1949 & ~n1955;
  assign n1957 = ~x1138 & ~n1496;
  assign n1958 = x269 & n1675;
  assign n1959 = ~x940 & n1672;
  assign n1960 = ~n1958 & ~n1959;
  assign n1961 = ~n1957 & n1960;
  assign n1962 = x299 & n1961;
  assign n1963 = ~n1956 & n1962;
  assign n1964 = x1138 & n1695;
  assign n1965 = ~x269 & n1702;
  assign n1966 = x877 & n1485;
  assign n1967 = ~n1965 & ~n1966;
  assign n1968 = ~n1964 & n1967;
  assign n1969 = x940 & n1699;
  assign n1970 = n1968 & ~n1969;
  assign n1971 = n1970 ^ x246;
  assign n1972 = ~n1692 & ~n1971;
  assign n1973 = n1972 ^ x246;
  assign n1974 = n1518 & ~n1973;
  assign n1975 = ~n1963 & n1974;
  assign n1976 = ~n1773 & n1950;
  assign n1977 = n1488 & ~n1976;
  assign n1978 = ~x169 & n1773;
  assign n1979 = n1977 & ~n1978;
  assign n1980 = n1961 & ~n1979;
  assign n1981 = x246 & n1682;
  assign n1982 = ~n1518 & ~n1981;
  assign n1983 = ~n1980 & n1982;
  assign n1984 = ~n1975 & ~n1983;
  assign n1985 = x878 ^ x240;
  assign n1986 = n1275 & n1985;
  assign n1987 = n1986 ^ x240;
  assign n1988 = ~n1478 & ~n1987;
  assign n1989 = x168 & ~n1477;
  assign n1990 = ~n1476 & n1989;
  assign n1991 = ~n1514 & ~n1692;
  assign n1992 = n1481 & ~n1991;
  assign n1993 = ~n1990 & n1992;
  assign n1994 = ~n1988 & n1993;
  assign n1995 = x878 & ~n1274;
  assign n1996 = n1477 & ~n1995;
  assign n1997 = n1488 & ~n1989;
  assign n1998 = ~n1996 & n1997;
  assign n1999 = ~x280 & n1675;
  assign n2000 = ~n1998 & ~n1999;
  assign n2001 = ~n1604 & ~n2000;
  assign n2002 = x1137 & ~n1496;
  assign n2003 = x933 & n1672;
  assign n2004 = ~n2002 & ~n2003;
  assign n2005 = x299 & n2004;
  assign n2006 = ~n2001 & n2005;
  assign n2007 = x878 & n1604;
  assign n2008 = n2006 & ~n2007;
  assign n2009 = n1514 & n1692;
  assign n2010 = ~n2008 & ~n2009;
  assign n2011 = ~n1687 & n2010;
  assign n2012 = ~n1994 & ~n2011;
  assign n2013 = ~x1137 & n1695;
  assign n2014 = n1485 & ~n1995;
  assign n2015 = x280 & n1702;
  assign n2016 = ~n2014 & ~n2015;
  assign n2017 = ~n2013 & n2016;
  assign n2018 = ~x933 & n1699;
  assign n2019 = n2017 & ~n2018;
  assign n2020 = ~n2012 & n2019;
  assign n2021 = x240 & n1485;
  assign n2022 = n1691 & n2021;
  assign n2023 = n1518 & ~n2022;
  assign n2024 = ~n2020 & n2023;
  assign n2025 = x240 & n1682;
  assign n2026 = n2004 & ~n2025;
  assign n2027 = n2000 & n2026;
  assign n2028 = ~n1578 & ~n2027;
  assign n2029 = ~n1518 & ~n2028;
  assign n2030 = x878 & n1578;
  assign n2031 = n2029 & ~n2030;
  assign n2032 = ~n2024 & ~n2031;
  assign n2033 = n1478 & n1518;
  assign n2034 = x875 & ~n1274;
  assign n2035 = n2034 ^ x166;
  assign n2036 = ~n1746 & n2035;
  assign n2037 = n2036 ^ x166;
  assign n2038 = n2033 & ~n2037;
  assign n2039 = n1488 & ~n2038;
  assign n2040 = ~x875 & ~n1274;
  assign n2041 = n2040 ^ x166;
  assign n2042 = ~n1773 & ~n2041;
  assign n2043 = n2042 ^ x166;
  assign n2044 = ~n1519 & ~n2043;
  assign n2045 = ~n2033 & n2044;
  assign n2046 = ~n1519 & n2037;
  assign n2047 = x875 ^ x245;
  assign n2048 = n1275 & n2047;
  assign n2049 = n2048 ^ x245;
  assign n2050 = ~n2046 & ~n2049;
  assign n2051 = ~n1478 & n2050;
  assign n2052 = ~n2045 & ~n2051;
  assign n2053 = n2039 & n2052;
  assign n2054 = x1136 & ~n1496;
  assign n2055 = x928 & n1672;
  assign n2056 = x266 & n1675;
  assign n2057 = ~n2055 & ~n2056;
  assign n2058 = ~n2054 & n2057;
  assign n2059 = ~n1656 & n2058;
  assign n2060 = ~n2053 & n2059;
  assign n2061 = x245 & n1691;
  assign n2062 = n1485 & n1518;
  assign n2063 = ~n2061 & n2062;
  assign n2064 = x875 & ~n1691;
  assign n2065 = n2063 & ~n2064;
  assign n2066 = ~x1136 & n1695;
  assign n2067 = ~x266 & n1702;
  assign n2068 = ~x928 & n1699;
  assign n2069 = ~n2067 & ~n2068;
  assign n2070 = ~n2066 & n2069;
  assign n2071 = n1518 & ~n2070;
  assign n2072 = ~n2065 & ~n2071;
  assign n2073 = ~n2060 & n2072;
  assign n2074 = ~x161 & n1866;
  assign n2075 = n1488 & ~n2074;
  assign n2076 = x879 & ~n1691;
  assign n2077 = ~n1866 & ~n2076;
  assign n2078 = n2075 & ~n2077;
  assign n2079 = x244 & ~n1693;
  assign n2080 = n1481 & ~n1746;
  assign n2081 = ~n1485 & ~n2080;
  assign n2082 = n2076 & ~n2081;
  assign n2083 = x279 & n1702;
  assign n2084 = n1518 & ~n2083;
  assign n2085 = x938 & n1699;
  assign n2086 = n2084 & ~n2085;
  assign n2087 = x1135 & n1695;
  assign n2088 = n2086 & ~n2087;
  assign n2089 = ~n2082 & n2088;
  assign n2090 = ~n2079 & n2089;
  assign n2091 = ~n2078 & n2090;
  assign n2092 = x879 ^ x244;
  assign n2093 = ~n1274 & n2092;
  assign n2094 = n2093 ^ x244;
  assign n2095 = n2094 ^ x161;
  assign n2096 = ~n1773 & n2095;
  assign n2097 = n2096 ^ x161;
  assign n2098 = n1488 & n2097;
  assign n2099 = ~n1518 & ~n2098;
  assign n2100 = ~n2091 & ~n2099;
  assign n2101 = x1135 & ~n1496;
  assign n2102 = x938 & n1672;
  assign n2103 = x279 & n1675;
  assign n2104 = ~n2102 & ~n2103;
  assign n2105 = ~n2101 & n2104;
  assign n2106 = ~n2100 & n2105;
  assign n2107 = ~x299 & n2090;
  assign n2108 = ~n2106 & ~n2107;
  assign n2109 = x152 & n1866;
  assign n2110 = n1488 & ~n2109;
  assign n2111 = x846 ^ x242;
  assign n2112 = ~n1691 & n2111;
  assign n2113 = n2112 ^ x242;
  assign n2114 = ~n1866 & n2113;
  assign n2115 = n2110 & ~n2114;
  assign n2116 = n1485 & ~n2113;
  assign n2117 = ~x930 & n1699;
  assign n2118 = ~x278 & n1702;
  assign n2119 = ~n2117 & ~n2118;
  assign n2120 = n1518 & n2119;
  assign n2121 = ~n2116 & n2120;
  assign n2122 = ~n2115 & n2121;
  assign n2123 = ~n1274 & n2111;
  assign n2124 = n2123 ^ x242;
  assign n2125 = ~n1773 & n2124;
  assign n2126 = n1488 & ~n2125;
  assign n2127 = x152 & n1773;
  assign n2128 = n2126 & ~n2127;
  assign n2129 = ~n1518 & ~n2128;
  assign n2130 = ~n2122 & ~n2129;
  assign n2131 = ~x278 & n1675;
  assign n2132 = ~x930 & n1672;
  assign n2133 = ~n2131 & ~n2132;
  assign n2134 = ~n2130 & n2133;
  assign n2135 = ~x299 & n2121;
  assign n2136 = ~n2134 & ~n2135;
  assign n2137 = n1695 ^ n1496;
  assign n2138 = n1656 & ~n2137;
  assign n2139 = n2138 ^ n1496;
  assign n2140 = ~x1134 & ~n2139;
  assign n2141 = ~n2136 & ~n2140;
  assign n2142 = n1233 & n1244;
  assign n2143 = n1403 & ~n2142;
  assign n2144 = n1379 & n2143;
  assign n2145 = x93 & x841;
  assign n2146 = n1407 & ~n2145;
  assign n2147 = n1461 & ~n2146;
  assign n2148 = ~n1459 & n2147;
  assign n2149 = ~n2144 & n2148;
  assign n2150 = ~n1414 & ~n2149;
  assign n2151 = ~n1255 & ~n2150;
  assign n2152 = n1255 & ~n1260;
  assign n2153 = x32 & ~n2152;
  assign n2154 = ~x70 & ~x95;
  assign n2155 = n1241 & n2154;
  assign n2156 = ~n2153 & n2155;
  assign n2157 = x32 & ~n2156;
  assign n2158 = n1519 & ~n1521;
  assign n2159 = ~n2157 & n2158;
  assign n2160 = ~n2151 & n2159;
  assign n2161 = ~x332 & ~x468;
  assign n2162 = x299 & n2161;
  assign n2170 = ~x614 & ~x616;
  assign n2171 = ~x642 & n2170;
  assign n2172 = x603 & n2171;
  assign n2173 = ~x661 & ~x662;
  assign n2174 = ~x681 & n2173;
  assign n2175 = x680 & n2174;
  assign n2176 = ~n2172 & ~n2175;
  assign n2163 = ~x969 & ~x971;
  assign n2164 = ~x974 & ~x977;
  assign n2165 = n2163 & n2164;
  assign n2166 = ~x587 & ~x602;
  assign n2167 = ~x961 & ~x967;
  assign n2168 = n2166 & n2167;
  assign n2169 = n2165 & n2168;
  assign n2177 = n2176 ^ n2169;
  assign n2178 = n2161 & n2177;
  assign n2179 = n2178 ^ n2176;
  assign n2180 = ~n2162 & n2179;
  assign n2181 = x824 & n1426;
  assign n2182 = ~n1423 & n2181;
  assign n2183 = ~n1428 & ~n2182;
  assign n2184 = ~n2180 & ~n2183;
  assign n2185 = ~x979 & ~x984;
  assign n2186 = ~x287 & n2185;
  assign n2187 = ~x252 & ~x1001;
  assign n2188 = x835 & ~n2187;
  assign n2189 = n2186 & n2188;
  assign n2190 = n2184 & n2189;
  assign n2191 = ~n1480 & ~n1697;
  assign n2192 = n2190 & n2191;
  assign n2193 = ~x970 & ~x972;
  assign n2194 = ~x975 & ~x978;
  assign n2195 = n2193 & n2194;
  assign n2196 = ~x907 & ~x947;
  assign n2197 = ~x960 & ~x963;
  assign n2198 = n2196 & n2197;
  assign n2199 = n2195 & n2198;
  assign n2200 = n2161 & n2199;
  assign n2201 = x299 & n2200;
  assign n2202 = n2192 & ~n2201;
  assign n2203 = x39 & n2202;
  assign n2204 = ~x41 & ~x101;
  assign n2205 = ~x99 & n2204;
  assign n2206 = ~x113 & n2205;
  assign n2207 = ~x43 & ~x44;
  assign n2208 = ~x42 & ~x114;
  assign n2209 = n2207 & n2208;
  assign n2210 = ~x115 & ~x116;
  assign n2211 = n2209 & n2210;
  assign n2212 = n2206 & n2211;
  assign n2213 = ~x52 & n2212;
  assign n2214 = ~x129 & x250;
  assign n2215 = x683 & ~n2214;
  assign n2216 = ~n2213 & n2215;
  assign n2217 = ~n1446 & ~n2216;
  assign n2218 = ~x250 & ~n1446;
  assign n2219 = ~x1093 & n2181;
  assign n2220 = ~x1093 & n1427;
  assign n2221 = ~n2219 & ~n2220;
  assign n2222 = n2218 & ~n2221;
  assign n2223 = ~x252 & n1446;
  assign n2224 = ~n2222 & ~n2223;
  assign n2225 = ~n2217 & n2224;
  assign n2226 = x100 & ~n2225;
  assign n2227 = ~x87 & x100;
  assign n2228 = ~n1537 & ~n2227;
  assign n2229 = ~x74 & ~n2228;
  assign n2230 = ~n2226 & n2229;
  assign n2231 = x224 & n1698;
  assign n2232 = ~n2179 & n2231;
  assign n2233 = ~n2161 & n2176;
  assign n2234 = ~n2200 & ~n2233;
  assign n2235 = x299 & n1671;
  assign n2236 = x216 & n2235;
  assign n2237 = n2234 & n2236;
  assign n2238 = ~n2232 & ~n2237;
  assign n2239 = n1431 & n2189;
  assign n2240 = ~n2238 & n2239;
  assign n2241 = x39 & n2240;
  assign n2242 = ~n2230 & ~n2241;
  assign n2243 = ~n2203 & n2242;
  assign n2244 = ~n1575 & n2243;
  assign n2245 = ~n1527 & ~n1563;
  assign n2246 = ~n2244 & n2245;
  assign n2247 = ~n2160 & n2246;
  assign n2248 = n1276 & n1519;
  assign n2249 = n1459 & n2248;
  assign n2250 = ~n1662 & ~n2249;
  assign n2251 = x67 & ~n1214;
  assign n2252 = n1217 & ~n2251;
  assign n2253 = ~x67 & ~n1323;
  assign n2254 = n2252 & ~n2253;
  assign n2255 = n1285 & n2254;
  assign n2256 = ~x85 & n1330;
  assign n2257 = ~n1319 & n2256;
  assign n2258 = ~n2255 & n2257;
  assign n2259 = ~x82 & n2258;
  assign n2260 = ~n2142 & n2259;
  assign n2261 = ~x58 & n1385;
  assign n2262 = ~n2260 & n2261;
  assign n2263 = n2147 & n2262;
  assign n2264 = x103 & ~x314;
  assign n2265 = ~x109 & ~n2264;
  assign n2266 = ~n2263 & n2265;
  assign n2267 = ~n2250 & ~n2266;
  assign n2268 = ~x72 & ~n2267;
  assign n2269 = ~n1410 & n1519;
  assign n2270 = n1256 & n1260;
  assign n2271 = n1225 & n1337;
  assign n2272 = n1246 & n2271;
  assign n2273 = n1220 & n2272;
  assign n2274 = ~x73 & n1253;
  assign n2275 = n2273 & n2274;
  assign n2276 = ~x32 & n1274;
  assign n2277 = n2275 & n2276;
  assign n2278 = n1250 & n1264;
  assign n2279 = ~x58 & x841;
  assign n2280 = x90 ^ x58;
  assign n2281 = ~n2279 & n2280;
  assign n2282 = n2278 & n2281;
  assign n2283 = ~n2277 & ~n2282;
  assign n2284 = ~n2270 & n2283;
  assign n2285 = ~n1265 & n2284;
  assign n2286 = n1250 & n1519;
  assign n2287 = n1403 & n2286;
  assign n2288 = ~n2285 & n2287;
  assign n2289 = ~n2269 & ~n2288;
  assign n2290 = ~n2268 & ~n2289;
  assign n2291 = x158 & x159;
  assign n2292 = x197 & n2291;
  assign n2293 = x160 & x232;
  assign n2294 = n2292 & n2293;
  assign n2295 = x299 & ~n2294;
  assign n2296 = n2161 & ~n2295;
  assign n2297 = x109 & x145;
  assign n2298 = x180 & x181;
  assign n2299 = n2297 & n2298;
  assign n2300 = x182 & x232;
  assign n2301 = n2299 & n2300;
  assign n2302 = x109 & x299;
  assign n2303 = ~n2301 & ~n2302;
  assign n2304 = n2296 & ~n2303;
  assign n2305 = n2290 & ~n2304;
  assign n2306 = ~x228 & n2305;
  assign n2307 = n1530 & n1551;
  assign n2308 = ~x75 & x100;
  assign n2309 = n2225 & n2308;
  assign n2310 = n2307 & n2309;
  assign n2311 = n1560 & ~n2310;
  assign n2312 = x1093 & n2182;
  assign n2313 = x829 & x1092;
  assign n2314 = ~n1424 & n2313;
  assign n2315 = n2312 & ~n2314;
  assign n2316 = n2189 & n2315;
  assign n2317 = ~n1698 & ~n2235;
  assign n2318 = n2316 & ~n2317;
  assign n2319 = ~n2231 & ~n2236;
  assign n2320 = n2239 & ~n2319;
  assign n2321 = ~n2318 & ~n2320;
  assign n2322 = x39 & n1634;
  assign n2323 = ~n2321 & n2322;
  assign n2324 = n1521 & n2323;
  assign n2325 = ~x228 & ~n2324;
  assign n2326 = n2311 & n2325;
  assign n2327 = ~x30 & x228;
  assign n2328 = n1518 & ~n2327;
  assign n2329 = ~n2326 & n2328;
  assign n2330 = ~n2306 & ~n2329;
  assign n2331 = ~x299 & n2161;
  assign n2332 = ~n2330 & n2331;
  assign n2333 = x602 & n2332;
  assign n2334 = ~x228 & n2290;
  assign n2335 = ~x228 & n1560;
  assign n2336 = ~n1518 & ~n2327;
  assign n2337 = ~n2335 & n2336;
  assign n2338 = ~n2329 & ~n2337;
  assign n2339 = ~n2334 & n2338;
  assign n2340 = ~x299 & ~n2336;
  assign n2341 = x109 & ~x228;
  assign n2342 = n2294 & n2341;
  assign n2343 = n2161 & ~n2342;
  assign n2344 = ~n2340 & n2343;
  assign n2345 = x907 & n2344;
  assign n2346 = ~n2161 & n2175;
  assign n2347 = ~n2345 & ~n2346;
  assign n2348 = ~n2339 & ~n2347;
  assign n2349 = ~n2333 & ~n2348;
  assign n2350 = ~n2330 & ~n2331;
  assign n2351 = ~n2337 & ~n2350;
  assign n2352 = n2172 ^ x947;
  assign n2353 = ~n2161 & n2352;
  assign n2354 = n2353 ^ x947;
  assign n2355 = ~n2351 & n2354;
  assign n2356 = x587 & n2332;
  assign n2357 = ~n2355 & ~n2356;
  assign n2358 = x967 & n2332;
  assign n2359 = ~n2339 & n2344;
  assign n2360 = x970 & n2359;
  assign n2361 = ~n2358 & ~n2360;
  assign n2362 = x299 & x972;
  assign n2363 = ~x109 & n2362;
  assign n2364 = ~x299 & x961;
  assign n2365 = ~n2363 & ~n2364;
  assign n2366 = ~n2301 & ~n2365;
  assign n2367 = ~n2294 & n2362;
  assign n2368 = ~n2366 & ~n2367;
  assign n2369 = n2334 & ~n2368;
  assign n2370 = ~n2362 & ~n2364;
  assign n2371 = n2329 & ~n2370;
  assign n2372 = x972 & n2337;
  assign n2373 = ~n2371 & ~n2372;
  assign n2374 = ~n2369 & n2373;
  assign n2375 = n2161 & ~n2374;
  assign n2376 = x977 & n2332;
  assign n2377 = x960 & n2359;
  assign n2378 = ~n2376 & ~n2377;
  assign n2379 = x969 & n2332;
  assign n2380 = x963 & n2359;
  assign n2381 = ~n2379 & ~n2380;
  assign n2382 = x971 & n2332;
  assign n2383 = x975 & n2359;
  assign n2384 = ~n2382 & ~n2383;
  assign n2385 = x974 & n2332;
  assign n2386 = x978 & n2359;
  assign n2387 = ~n2385 & ~n2386;
  assign n2388 = ~x96 & n1265;
  assign n2389 = ~x90 & ~x93;
  assign n2390 = ~x35 & ~x70;
  assign n2391 = n2389 & n2390;
  assign n2392 = n2388 & n2391;
  assign n2393 = n1246 & n2392;
  assign n2394 = n1229 & n2393;
  assign n2395 = ~x92 & n1511;
  assign n2396 = n1518 & n2395;
  assign n2397 = n2394 & n2396;
  assign n2398 = x39 & ~x72;
  assign n2399 = n2397 & n2398;
  assign n2400 = ~x51 & ~x87;
  assign n2401 = n1232 & n2400;
  assign n2402 = n2399 & n2401;
  assign n2403 = ~n1656 & n1671;
  assign n2404 = n2234 & n2403;
  assign n2405 = n1518 & n1698;
  assign n2406 = ~n2179 & n2405;
  assign n2407 = ~n2404 & ~n2406;
  assign n2408 = n2316 & ~n2407;
  assign n2409 = ~n2240 & ~n2408;
  assign n2410 = n2402 & ~n2409;
  assign n2411 = n2311 & ~n2410;
  assign n2412 = ~n2305 & n2411;
  assign n2413 = n2412 ^ x24;
  assign n2414 = ~x954 & n2413;
  assign n2415 = n2414 ^ x24;
  assign n2416 = n1446 & n1598;
  assign n2417 = n1573 & ~n2416;
  assign n2418 = n1663 & ~n2417;
  assign n2419 = n2418 ^ x105;
  assign n2420 = ~x228 & ~n2419;
  assign n2421 = n2420 ^ x105;
  assign n2422 = ~x119 & ~x228;
  assign n2423 = x252 & ~x468;
  assign n2424 = n2422 & n2423;
  assign n2425 = x119 & ~x468;
  assign n2426 = ~x1056 & n2425;
  assign n2427 = ~n2424 & ~n2426;
  assign n2428 = ~x1077 & n2425;
  assign n2429 = ~n2424 & ~n2428;
  assign n2430 = ~x1073 & n2425;
  assign n2431 = ~n2424 & ~n2430;
  assign n2432 = ~x1041 & n2425;
  assign n2433 = ~n2424 & ~n2432;
  assign n2434 = n1249 & n1404;
  assign n2435 = x98 & n2434;
  assign n2436 = x51 & n2389;
  assign n2437 = ~x51 & ~x841;
  assign n2438 = x93 ^ x90;
  assign n2439 = n2437 & n2438;
  assign n2440 = ~n2436 & ~n2439;
  assign n2441 = n2390 & ~n2440;
  assign n2442 = n1247 & n2441;
  assign n2443 = ~n2435 & ~n2442;
  assign n2444 = ~x96 & n2443;
  assign n2445 = ~x98 & x1091;
  assign n2446 = n2221 & ~n2445;
  assign n2447 = ~x72 & ~n2446;
  assign n2448 = ~n2183 & n2447;
  assign n2449 = ~n2444 & n2448;
  assign n2450 = x91 & n1453;
  assign n2451 = ~x24 & ~x58;
  assign n2452 = n2450 & n2451;
  assign n2453 = ~n1416 & ~n2452;
  assign n2454 = ~x122 & n1431;
  assign n2455 = ~x72 & n1249;
  assign n2456 = n1252 & n2455;
  assign n2457 = n2454 & n2456;
  assign n2458 = ~n2453 & n2457;
  assign n2459 = ~n2449 & ~n2458;
  assign n2460 = n1249 & n1263;
  assign n2461 = ~x122 & x829;
  assign n2462 = ~x841 & n2461;
  assign n2463 = n1265 & n2462;
  assign n2464 = n2460 & n2463;
  assign n2465 = ~n2388 & ~n2464;
  assign n2466 = ~n2459 & ~n2465;
  assign n2467 = ~x39 & ~x72;
  assign n2468 = n2388 & n2467;
  assign n2469 = ~n2443 & n2468;
  assign n2470 = ~x87 & ~n2469;
  assign n2471 = ~n2183 & ~n2470;
  assign n2472 = ~x75 & ~n1565;
  assign n2473 = ~n2471 & n2472;
  assign n2474 = ~n2466 & n2473;
  assign n2475 = x299 & ~n1443;
  assign n2476 = x232 & n2161;
  assign n2477 = ~n2475 & n2476;
  assign n2478 = ~x299 & ~n1439;
  assign n2479 = n2477 & ~n2478;
  assign n2480 = ~n2213 & ~n2479;
  assign n2481 = x252 & n2480;
  assign n2482 = ~x24 & ~x100;
  assign n2483 = ~x87 & n2482;
  assign n2484 = n2454 & n2483;
  assign n2485 = n2481 & n2484;
  assign n2486 = n1521 & n2485;
  assign n2487 = x75 & ~n2486;
  assign n2488 = n1567 & n1633;
  assign n2489 = n1521 & n2488;
  assign n2490 = ~n2487 & n2489;
  assign n2491 = ~n1698 & ~n1701;
  assign n2492 = ~n2179 & ~n2491;
  assign n2493 = ~n1479 & n1480;
  assign n2494 = n2234 & n2493;
  assign n2495 = ~n2492 & ~n2494;
  assign n2496 = ~x224 & n1698;
  assign n2497 = ~x216 & n2235;
  assign n2498 = ~n2496 & ~n2497;
  assign n2499 = ~n2495 & ~n2498;
  assign n2500 = n2239 & n2499;
  assign n2501 = x39 & ~n2500;
  assign n2502 = n2454 & n2480;
  assign n2503 = x228 & n2502;
  assign n2504 = x100 & ~n2503;
  assign n2505 = n1512 & n1571;
  assign n2506 = ~n2504 & n2505;
  assign n2507 = ~n2501 & n2506;
  assign n2508 = n1521 & n2507;
  assign n2509 = ~n1514 & ~n2508;
  assign n2510 = ~n2490 & n2509;
  assign n2515 = x374 ^ x373;
  assign n2514 = x384 ^ x375;
  assign n2516 = n2515 ^ n2514;
  assign n2513 = x442 ^ x440;
  assign n2517 = n2516 ^ n2513;
  assign n2511 = x371 ^ x370;
  assign n2512 = n2511 ^ x369;
  assign n2518 = n2517 ^ n2512;
  assign n2519 = x1198 & n2518;
  assign n2524 = x386 ^ x380;
  assign n2523 = x372 ^ x363;
  assign n2525 = n2524 ^ n2523;
  assign n2522 = x388 ^ x387;
  assign n2526 = n2525 ^ n2522;
  assign n2520 = x339 ^ x338;
  assign n2521 = n2520 ^ x337;
  assign n2527 = n2526 ^ n2521;
  assign n2528 = x1196 & n2527;
  assign n2529 = ~n2519 & ~n2528;
  assign n2534 = x367 ^ x366;
  assign n2533 = x383 ^ x368;
  assign n2535 = n2534 ^ n2533;
  assign n2532 = x447 ^ x389;
  assign n2536 = n2535 ^ n2532;
  assign n2530 = x365 ^ x364;
  assign n2531 = n2530 ^ x336;
  assign n2537 = n2536 ^ n2531;
  assign n2538 = x1197 & n2537;
  assign n2539 = n2529 & ~n2538;
  assign n2544 = x379 ^ x378;
  assign n2543 = x439 ^ x385;
  assign n2545 = n2544 ^ n2543;
  assign n2542 = x382 ^ x381;
  assign n2546 = n2545 ^ n2542;
  assign n2540 = x377 ^ x376;
  assign n2541 = n2540 ^ x317;
  assign n2547 = n2546 ^ n2541;
  assign n2548 = x1199 & n2547;
  assign n2549 = ~x591 & ~n2548;
  assign n2550 = n2539 & n2549;
  assign n2551 = ~x590 & ~n2550;
  assign n2556 = x356 ^ x354;
  assign n2555 = x360 ^ x357;
  assign n2557 = n2556 ^ n2555;
  assign n2554 = x462 ^ x461;
  assign n2558 = n2557 ^ n2554;
  assign n2552 = x353 ^ x352;
  assign n2553 = n2552 ^ x351;
  assign n2559 = n2558 ^ n2553;
  assign n2560 = x1199 & n2559;
  assign n2565 = x441 ^ x361;
  assign n2564 = x460 ^ x458;
  assign n2566 = n2565 ^ n2564;
  assign n2563 = x455 ^ x452;
  assign n2567 = n2566 ^ n2563;
  assign n2561 = x355 ^ x342;
  assign n2562 = n2561 ^ x320;
  assign n2568 = n2567 ^ n2562;
  assign n2569 = x1196 & n2568;
  assign n2570 = ~n2560 & ~n2569;
  assign n2575 = x347 ^ x322;
  assign n2574 = x359 ^ x350;
  assign n2576 = n2575 ^ n2574;
  assign n2573 = x349 ^ x348;
  assign n2577 = n2576 ^ n2573;
  assign n2571 = x321 ^ x316;
  assign n2572 = n2571 ^ x315;
  assign n2578 = n2577 ^ n2572;
  assign n2579 = x1198 & n2578;
  assign n2584 = x345 ^ x344;
  assign n2583 = x358 ^ x346;
  assign n2585 = n2584 ^ n2583;
  assign n2582 = x450 ^ x362;
  assign n2586 = n2585 ^ n2582;
  assign n2580 = x343 ^ x327;
  assign n2581 = n2580 ^ x323;
  assign n2587 = n2586 ^ n2581;
  assign n2588 = x1197 & n2587;
  assign n2589 = ~n2579 & ~n2588;
  assign n2590 = n2570 & n2589;
  assign n2591 = ~x591 & ~x592;
  assign n2592 = ~n2590 & n2591;
  assign n2593 = ~n2551 & ~n2592;
  assign n2594 = ~x590 & ~x592;
  assign n2595 = ~x591 & n2594;
  assign n2596 = ~n2593 & ~n2595;
  assign n2597 = x588 & n2596;
  assign n2598 = ~x217 & ~n2597;
  assign n2603 = x424 ^ x423;
  assign n2602 = x432 ^ x425;
  assign n2604 = n2603 ^ n2602;
  assign n2601 = x459 ^ x454;
  assign n2605 = n2604 ^ n2601;
  assign n2599 = x421 ^ x420;
  assign n2600 = n2599 ^ x419;
  assign n2606 = n2605 ^ n2600;
  assign n2607 = x1198 & n2606;
  assign n2612 = x438 ^ x437;
  assign n2611 = x431 ^ x418;
  assign n2613 = n2612 ^ n2611;
  assign n2610 = x464 ^ x453;
  assign n2614 = n2613 ^ n2610;
  assign n2608 = x417 ^ x416;
  assign n2609 = n2608 ^ x415;
  assign n2615 = n2614 ^ n2609;
  assign n2616 = x1197 & n2615;
  assign n2617 = ~n2607 & ~n2616;
  assign n2622 = x448 ^ x445;
  assign n2621 = x433 ^ x430;
  assign n2623 = n2622 ^ n2621;
  assign n2620 = x451 ^ x449;
  assign n2624 = n2623 ^ n2620;
  assign n2618 = x428 ^ x427;
  assign n2619 = n2618 ^ x426;
  assign n2625 = n2624 ^ n2619;
  assign n2626 = x1199 & n2625;
  assign n2631 = x435 ^ x434;
  assign n2630 = x446 ^ x444;
  assign n2632 = n2631 ^ n2630;
  assign n2629 = x443 ^ x436;
  assign n2633 = n2632 ^ n2629;
  assign n2627 = x429 ^ x422;
  assign n2628 = n2627 ^ x414;
  assign n2634 = n2633 ^ n2628;
  assign n2635 = x1196 & n2634;
  assign n2636 = ~n2626 & ~n2635;
  assign n2637 = n2617 & n2636;
  assign n2638 = x588 & n2594;
  assign n2639 = ~n2637 & n2638;
  assign n2640 = ~n2596 & ~n2639;
  assign n2641 = n2598 & ~n2640;
  assign n2646 = x392 ^ x391;
  assign n2645 = x407 ^ x393;
  assign n2647 = n2646 ^ n2645;
  assign n2644 = x463 ^ x413;
  assign n2648 = n2647 ^ n2644;
  assign n2642 = x335 ^ x334;
  assign n2643 = n2642 ^ x333;
  assign n2649 = n2648 ^ n2643;
  assign n2650 = x1197 & n2649;
  assign n2655 = x396 ^ x395;
  assign n2654 = x408 ^ x400;
  assign n2656 = n2655 ^ n2654;
  assign n2653 = x399 ^ x398;
  assign n2657 = n2656 ^ n2653;
  assign n2651 = x394 ^ x329;
  assign n2652 = n2651 ^ x328;
  assign n2658 = n2657 ^ n2652;
  assign n2659 = x1198 & n2658;
  assign n2660 = ~n2650 & ~n2659;
  assign n2661 = ~x592 & ~n2660;
  assign n2662 = x591 & ~n2661;
  assign n2667 = x411 ^ x410;
  assign n2666 = x404 ^ x397;
  assign n2668 = n2667 ^ n2666;
  assign n2665 = x456 ^ x412;
  assign n2669 = n2668 ^ n2665;
  assign n2663 = x390 ^ x324;
  assign n2664 = n2663 ^ x319;
  assign n2670 = n2669 ^ n2664;
  assign n2671 = x1196 & n2670;
  assign n2676 = x402 ^ x401;
  assign n2675 = x409 ^ x406;
  assign n2677 = n2676 ^ n2675;
  assign n2674 = x405 ^ x403;
  assign n2678 = n2677 ^ n2674;
  assign n2672 = x326 ^ x325;
  assign n2673 = n2672 ^ x318;
  assign n2679 = n2678 ^ n2673;
  assign n2680 = x1199 & n2679;
  assign n2681 = ~n2671 & ~n2680;
  assign n2682 = n2594 & ~n2681;
  assign n2683 = x567 & n2682;
  assign n2684 = n2662 & ~n2683;
  assign n2685 = n2641 & ~n2684;
  assign n2686 = n1424 & n2685;
  assign n2687 = ~n2510 & ~n2686;
  assign n2688 = ~n2474 & n2687;
  assign n2689 = n2641 & ~n2662;
  assign n2690 = ~x286 & ~x289;
  assign n2691 = ~x285 & ~x288;
  assign n2692 = n2690 & n2691;
  assign n2693 = ~n2689 & ~n2692;
  assign n2694 = ~n2688 & ~n2693;
  assign n2695 = x1092 & x1093;
  assign n2696 = ~x98 & x567;
  assign n2697 = n2695 & ~n2696;
  assign n2698 = ~x1161 & ~x1162;
  assign n2699 = ~x1163 & n2698;
  assign n2700 = ~n2697 & n2699;
  assign n2701 = n1518 & n2700;
  assign n2702 = ~n2694 & n2701;
  assign n2703 = x567 & n2221;
  assign n2704 = ~x1199 & ~n2703;
  assign n2705 = ~x217 & ~x588;
  assign n2706 = x591 & ~x1091;
  assign n2707 = n2705 & n2706;
  assign n2708 = ~n2704 & n2707;
  assign n2709 = n2660 & n2708;
  assign n2710 = n2682 & n2709;
  assign n2711 = n1424 & n2181;
  assign n2712 = n2468 & n2711;
  assign n2713 = n2712 ^ n1565;
  assign n2714 = n2442 & n2713;
  assign n2715 = n2714 ^ n1565;
  assign n2716 = ~n2710 & n2715;
  assign n2717 = ~n2466 & ~n2716;
  assign n2718 = ~n2509 & ~n2717;
  assign n2719 = ~n1531 & ~n2183;
  assign n2720 = n2490 & n2719;
  assign n2721 = ~x122 & n2711;
  assign n2722 = ~x98 & n2721;
  assign n2723 = ~n2720 & ~n2722;
  assign n2724 = n2703 & n2710;
  assign n2725 = ~n2723 & ~n2724;
  assign n2726 = ~n2718 & ~n2725;
  assign n2727 = n2702 & ~n2726;
  assign n2728 = ~n2692 & n2721;
  assign n2729 = n2696 & n2698;
  assign n2730 = n2728 & n2729;
  assign n2731 = ~n1518 & n2730;
  assign n2732 = ~n2685 & n2731;
  assign n2733 = ~x31 & n2695;
  assign n2734 = x1161 & x1162;
  assign n2735 = n2733 & n2734;
  assign n2736 = ~n2732 & ~n2735;
  assign n2737 = ~x1163 & ~n2736;
  assign n2738 = ~n2727 & ~n2737;
  assign n2739 = x76 & n1333;
  assign n2740 = ~n1428 & ~n2692;
  assign n2741 = ~x137 & ~n1259;
  assign n2742 = ~x50 & n2741;
  assign n2743 = ~n2740 & n2742;
  assign n2744 = n2739 & n2743;
  assign n2745 = ~x24 & n1233;
  assign n2746 = x50 & n2745;
  assign n2747 = ~x841 & n1259;
  assign n2748 = x32 & ~x841;
  assign n2749 = ~x24 & n2748;
  assign n2750 = n2749 ^ x32;
  assign n2751 = ~n2747 & n2750;
  assign n2752 = ~n2746 & ~n2751;
  assign n2753 = ~n2744 & n2752;
  assign n2754 = n1662 & ~n2753;
  assign n2755 = n2221 ^ x129;
  assign n2756 = n2218 & n2755;
  assign n2757 = n2756 ^ x129;
  assign n2758 = n2308 & n2757;
  assign n2759 = ~n2223 & n2758;
  assign n2760 = x252 & ~n2480;
  assign n2761 = x75 & n2482;
  assign n2762 = ~n1428 & n2761;
  assign n2763 = ~n2760 & n2762;
  assign n2764 = ~n2759 & ~n2763;
  assign n2765 = n1446 & n2762;
  assign n2766 = n2480 & ~n2765;
  assign n2767 = ~x137 & ~n2766;
  assign n2768 = ~n2764 & n2767;
  assign n2769 = n2307 & n2768;
  assign n2770 = ~n2754 & ~n2769;
  assign n2771 = ~x70 & n1356;
  assign n2772 = ~n1410 & ~n2771;
  assign n2773 = n1403 & ~n2284;
  assign n2774 = ~n2772 & ~n2773;
  assign n2775 = x73 & n2273;
  assign n2776 = n1253 & n1264;
  assign n2777 = n2775 & n2776;
  assign n2778 = n2774 & ~n2777;
  assign n2779 = ~x195 & ~x196;
  assign n2780 = ~x138 & ~x139;
  assign n2781 = n2779 & n2780;
  assign n2782 = ~x79 & ~x118;
  assign n2783 = ~x33 & ~x34;
  assign n2784 = n2782 & n2783;
  assign n2785 = n2781 & n2784;
  assign n2786 = x954 ^ x33;
  assign n2787 = ~n2785 & ~n2786;
  assign n2788 = ~x63 & ~x107;
  assign n2789 = ~x40 & n2788;
  assign n2790 = ~n2787 & n2789;
  assign n2791 = x164 & x299;
  assign n2792 = x186 & ~x299;
  assign n2793 = ~n2791 & ~n2792;
  assign n2794 = n2476 & ~n2793;
  assign n2795 = ~n1510 & ~n2794;
  assign n2796 = n1540 & ~n2795;
  assign n2797 = n2790 & n2796;
  assign n2798 = n2778 & n2797;
  assign n2799 = ~n2169 & n2231;
  assign n2800 = ~x174 & n2799;
  assign n2801 = ~n2199 & n2236;
  assign n2802 = ~x152 & n2801;
  assign n2803 = ~n2800 & ~n2802;
  assign n2804 = n2316 & ~n2803;
  assign n2805 = x176 & n2799;
  assign n2806 = x154 & n2801;
  assign n2807 = ~n2805 & ~n2806;
  assign n2808 = n2239 & ~n2807;
  assign n2809 = ~n2804 & ~n2808;
  assign n2810 = n1521 & ~n2809;
  assign n2811 = x39 & ~n2810;
  assign n2812 = n2476 & ~n2811;
  assign n2813 = n1264 & n2275;
  assign n2814 = ~n2239 & ~n2316;
  assign n2815 = ~n2238 & ~n2814;
  assign n2816 = n2813 & n2815;
  assign n2817 = n1512 & n2816;
  assign n2818 = ~n2812 & n2817;
  assign n2819 = n1536 & n2813;
  assign n2820 = x92 & n2819;
  assign n2821 = x176 ^ x154;
  assign n2822 = ~x299 & n2821;
  assign n2823 = n2822 ^ x154;
  assign n2824 = n2476 & n2823;
  assign n2825 = n2789 & n2824;
  assign n2826 = n2820 & n2825;
  assign n2827 = ~n1513 & n2790;
  assign n2828 = ~n2819 & n2827;
  assign n2829 = ~n2826 & ~n2828;
  assign n2830 = ~n2818 & ~n2829;
  assign n2831 = n1512 & n2468;
  assign n2832 = n2460 & n2831;
  assign n2833 = x38 & ~n2832;
  assign n2834 = ~x54 & ~n2833;
  assign n2835 = ~n2830 & n2834;
  assign n2836 = ~x74 & ~n2795;
  assign n2837 = ~n2835 & n2836;
  assign n2838 = x191 ^ x169;
  assign n2839 = ~x299 & n2838;
  assign n2840 = n2839 ^ x169;
  assign n2841 = n2476 & n2840;
  assign n2842 = x74 & n2841;
  assign n2843 = n1508 & ~n2842;
  assign n2844 = ~n2837 & n2843;
  assign n2845 = ~n1508 & n2476;
  assign n2847 = x157 ^ x149;
  assign n2846 = x183 ^ x178;
  assign n2848 = n2847 ^ n2846;
  assign n2849 = ~x299 & n2848;
  assign n2850 = n2849 ^ n2847;
  assign n2851 = n2845 & n2850;
  assign n2852 = ~n2844 & ~n2851;
  assign n2853 = n1518 & ~n2852;
  assign n2854 = ~n2798 & n2853;
  assign n2855 = n1403 & n2282;
  assign n2856 = x193 ^ x172;
  assign n2857 = ~x299 & n2856;
  assign n2858 = n2857 ^ x172;
  assign n2859 = n2855 & n2858;
  assign n2860 = x180 ^ x158;
  assign n2861 = ~x299 & n2860;
  assign n2862 = n2861 ^ x158;
  assign n2863 = n1274 & n2862;
  assign n2864 = n1254 & n2863;
  assign n2865 = ~x198 & ~x299;
  assign n2866 = ~x841 & n1205;
  assign n2867 = n2865 & n2866;
  assign n2868 = n2275 & n2867;
  assign n2869 = ~x299 & ~n2771;
  assign n2870 = ~n2868 & ~n2869;
  assign n2871 = x183 & ~n2870;
  assign n2872 = ~x210 & n2748;
  assign n2873 = n2771 & ~n2872;
  assign n2874 = x149 & ~n2873;
  assign n2875 = ~x73 & ~n2874;
  assign n2876 = x73 & x152;
  assign n2877 = x299 & ~n2876;
  assign n2878 = x73 & ~x299;
  assign n2879 = ~x174 & n2878;
  assign n2880 = ~n2877 & ~n2879;
  assign n2881 = ~n2875 & ~n2880;
  assign n2882 = ~n2871 & ~n2881;
  assign n2883 = ~n2864 & n2882;
  assign n2884 = ~n2859 & n2883;
  assign n2885 = ~n1413 & ~n2884;
  assign n2886 = ~x39 & ~n2885;
  assign n2887 = n1634 & n2812;
  assign n2888 = ~n2886 & n2887;
  assign n2889 = n2854 & ~n2888;
  assign n2890 = n1510 & n1517;
  assign n2891 = n1509 & n2890;
  assign n2892 = n2789 & n2891;
  assign n2893 = n1515 & n1522;
  assign n2894 = x149 & n2476;
  assign n2895 = n2894 ^ n2787;
  assign n2896 = n2893 & ~n2895;
  assign n2897 = n2896 ^ n2787;
  assign n2898 = n2892 & ~n2897;
  assign n2899 = ~x74 & ~n2890;
  assign n2900 = x164 & n2899;
  assign n2901 = x74 & x169;
  assign n2902 = ~n2900 & ~n2901;
  assign n2903 = n2476 & ~n2902;
  assign n2904 = n1508 & ~n2903;
  assign n2905 = n2845 & n2847;
  assign n2906 = ~n2904 & ~n2905;
  assign n2907 = ~n1518 & ~n2906;
  assign n2908 = ~n2898 & n2907;
  assign n2909 = ~n2889 & ~n2908;
  assign n2910 = n1519 & n2778;
  assign n2911 = n1513 & n1515;
  assign n2912 = n2813 & n2911;
  assign n2913 = ~n1516 & ~n2912;
  assign n2914 = ~n2910 & ~n2913;
  assign n2915 = ~x33 & ~x954;
  assign n2916 = n2915 ^ x34;
  assign n2917 = n2785 & n2915;
  assign n2918 = n2916 & n2917;
  assign n2919 = n2918 ^ n2916;
  assign n2920 = ~n2914 & ~n2919;
  assign n2921 = ~n2820 & ~n2919;
  assign n2922 = x39 & n2817;
  assign n2923 = ~n2921 & ~n2922;
  assign n2924 = x177 ^ x155;
  assign n2925 = ~x299 & n2924;
  assign n2926 = n2925 ^ x155;
  assign n2927 = n2476 & n2926;
  assign n2928 = n2820 & n2927;
  assign n2929 = n2923 & ~n2928;
  assign n2930 = ~x144 & n2799;
  assign n2931 = ~x161 & n2801;
  assign n2932 = ~n2930 & ~n2931;
  assign n2933 = n2315 & ~n2932;
  assign n2934 = x177 & n2799;
  assign n2935 = x155 & n2801;
  assign n2936 = ~n2934 & ~n2935;
  assign n2937 = n1431 & ~n2936;
  assign n2938 = ~n2933 & ~n2937;
  assign n2939 = n2476 & ~n2938;
  assign n2940 = n2817 & ~n2939;
  assign n2941 = ~n1514 & n1516;
  assign n2942 = ~n2940 & n2941;
  assign n2943 = ~n2929 & n2942;
  assign n2944 = ~n2920 & ~n2943;
  assign n2945 = n2892 & ~n2944;
  assign n2946 = ~n1440 & ~n1444;
  assign n2947 = n2855 & ~n2946;
  assign n2948 = x140 & ~n2870;
  assign n2949 = x162 & x299;
  assign n2950 = ~n2873 & n2949;
  assign n2951 = x161 & x299;
  assign n2952 = x73 & ~n2951;
  assign n2953 = x144 & ~x299;
  assign n2954 = n2952 & ~n2953;
  assign n2955 = x181 ^ x159;
  assign n2956 = ~x299 & n2955;
  assign n2957 = n2956 ^ x159;
  assign n2958 = n2276 & n2957;
  assign n2959 = ~n2954 & ~n2958;
  assign n2960 = ~n2950 & n2959;
  assign n2961 = ~n2948 & n2960;
  assign n2962 = ~n2947 & n2961;
  assign n2963 = n1662 & ~n2962;
  assign n2964 = x188 ^ x167;
  assign n2965 = ~x299 & n2964;
  assign n2966 = n2965 ^ x167;
  assign n2967 = ~x74 & n2966;
  assign n2968 = ~n2834 & n2967;
  assign n2969 = x148 ^ x141;
  assign n2970 = x299 & n2969;
  assign n2971 = n2970 ^ x141;
  assign n2972 = x74 & n2971;
  assign n2973 = n1518 & ~n2972;
  assign n2974 = ~n2968 & n2973;
  assign n2975 = x167 & n2899;
  assign n2976 = x74 & x148;
  assign n2977 = ~n1518 & ~n2976;
  assign n2978 = ~n2975 & n2977;
  assign n2979 = n1508 & ~n2978;
  assign n2980 = ~n2974 & n2979;
  assign n2982 = ~x149 & ~x157;
  assign n2981 = x197 ^ x162;
  assign n2983 = n2982 ^ n2981;
  assign n2984 = ~n1656 & n2983;
  assign n2985 = ~n1508 & ~n2984;
  assign n2987 = ~x178 & ~x183;
  assign n2986 = x145 ^ x140;
  assign n2988 = n2987 ^ n2986;
  assign n2989 = n1656 & n2988;
  assign n2990 = n2985 & ~n2989;
  assign n2991 = ~n2980 & ~n2990;
  assign n2992 = ~n2963 & n2991;
  assign n2993 = n1576 & n2912;
  assign n2994 = x162 & n2993;
  assign n2995 = n2992 & ~n2994;
  assign n2996 = n2476 & ~n2995;
  assign n2997 = ~n2945 & ~n2996;
  assign n2998 = x24 & x59;
  assign n2999 = ~x55 & ~x74;
  assign n3000 = ~n2998 & n2999;
  assign n3001 = n1543 & n3000;
  assign n3002 = x841 ^ x93;
  assign n3003 = n1406 & n3002;
  assign n3004 = n2262 & ~n3003;
  assign n3005 = ~x122 & n2221;
  assign n3006 = ~n2740 & n3005;
  assign n3007 = x76 & ~n2741;
  assign n3008 = n3006 & n3007;
  assign n3009 = ~n1453 & ~n3008;
  assign n3010 = ~n3004 & ~n3009;
  assign n3011 = x40 & x1082;
  assign n3012 = ~n3010 & ~n3011;
  assign n3013 = ~n1413 & ~n3012;
  assign n3014 = n1544 & ~n2270;
  assign n3015 = x24 & ~x59;
  assign n3016 = ~n3014 & ~n3015;
  assign n3017 = ~n3013 & ~n3016;
  assign n3039 = ~n2832 & n2899;
  assign n3040 = n1539 & ~n3039;
  assign n3018 = x137 & ~n1428;
  assign n3019 = ~n2760 & ~n3018;
  assign n3020 = ~n1446 & ~n2213;
  assign n3021 = ~x38 & x75;
  assign n3022 = ~n3020 & n3021;
  assign n3023 = ~n3019 & n3022;
  assign n3024 = x38 & ~x75;
  assign n3025 = ~n3023 & ~n3024;
  assign n3026 = n2482 & ~n3025;
  assign n3027 = n2182 & n2480;
  assign n3028 = x683 & n3027;
  assign n3029 = x137 & n2760;
  assign n3030 = n3029 ^ x252;
  assign n3031 = ~n3028 & n3030;
  assign n3032 = ~x137 & ~n1446;
  assign n3033 = n1510 & ~n3032;
  assign n3034 = ~n3020 & n3033;
  assign n3035 = n2758 & n3034;
  assign n3036 = ~n3031 & n3035;
  assign n3037 = ~n3026 & ~n3036;
  assign n3038 = n2832 & ~n3037;
  assign n3041 = n3040 ^ n3038;
  assign n3042 = n3017 & n3041;
  assign n3043 = n3042 ^ n3040;
  assign n3044 = n3001 & n3043;
  assign n3045 = x36 & n1246;
  assign n3046 = n1333 & n3045;
  assign n3047 = ~n2452 & ~n3046;
  assign n3048 = n1252 & n2248;
  assign n3049 = ~n3047 & n3048;
  assign n3050 = ~n2221 & n3049;
  assign n3051 = n1246 & n3048;
  assign n3052 = n1333 & n3051;
  assign n3053 = ~x841 & n3052;
  assign n3054 = ~x70 & ~x89;
  assign n3055 = x332 & ~n3054;
  assign n3056 = n3053 & n3055;
  assign n3057 = n1354 & n3051;
  assign n3058 = x64 & n3057;
  assign n3059 = ~x841 & n3058;
  assign n3060 = ~n3056 & ~n3059;
  assign n3061 = x24 & n1535;
  assign n3062 = n3060 & ~n3061;
  assign n3063 = ~x986 & n2221;
  assign n3064 = x252 & ~n3063;
  assign n3065 = x108 & x314;
  assign n3066 = ~n3064 & n3065;
  assign n3067 = ~x35 & ~x48;
  assign n3068 = ~x47 & n3067;
  assign n3069 = ~n3066 & n3068;
  assign n3070 = x841 & ~n3067;
  assign n3071 = ~n3069 & ~n3070;
  assign n3072 = n2269 & n3071;
  assign n3073 = n1256 & n2747;
  assign n3074 = n1519 & n3073;
  assign n3075 = ~x287 & n2402;
  assign n3076 = ~x1093 & ~n2192;
  assign n3077 = x835 & ~n2201;
  assign n3078 = n2184 & n3077;
  assign n3079 = ~n3076 & n3078;
  assign n3080 = x835 & x984;
  assign n3081 = ~x979 & ~n3080;
  assign n3082 = ~n2187 & n3081;
  assign n3083 = x786 & ~x1082;
  assign n3084 = n3082 & n3083;
  assign n3085 = ~n3078 & n3084;
  assign n3086 = n3082 & ~n3085;
  assign n3087 = ~n3079 & n3086;
  assign n3088 = n3075 & n3087;
  assign n3089 = ~n3074 & ~n3088;
  assign n3090 = ~n3072 & n3089;
  assign n3091 = x102 ^ x40;
  assign n3092 = ~x102 & x1082;
  assign n3093 = n3091 & n3092;
  assign n3094 = n3093 ^ n3091;
  assign n3095 = n1662 & n3094;
  assign n3096 = ~n1248 & ~n1428;
  assign n3097 = ~n2444 & ~n3096;
  assign n3098 = n2308 & ~n2502;
  assign n3099 = ~n1531 & ~n3098;
  assign n3100 = x228 & ~n3099;
  assign n3101 = ~n2458 & n3100;
  assign n3102 = ~n3097 & n3101;
  assign n3103 = ~x250 & x252;
  assign n3104 = x901 & ~x959;
  assign n3105 = n3103 & n3104;
  assign n3106 = x94 & ~x110;
  assign n3107 = n3105 & n3106;
  assign n3108 = ~x94 & x110;
  assign n3109 = ~x480 & x949;
  assign n3110 = n3108 & n3109;
  assign n3111 = ~n3107 & ~n3110;
  assign n3112 = ~n2434 & ~n3111;
  assign n3113 = ~x87 & ~x100;
  assign n3114 = ~n1521 & ~n3113;
  assign n3115 = ~x228 & n3111;
  assign n3116 = x87 & x100;
  assign n3117 = n1633 & ~n3116;
  assign n3118 = n1518 & n3117;
  assign n3119 = ~n3115 & n3118;
  assign n3120 = ~n3114 & n3119;
  assign n3121 = ~n2487 & n3120;
  assign n3122 = ~n2465 & n3121;
  assign n3123 = ~n3112 & n3122;
  assign n3124 = ~n3102 & n3123;
  assign n3125 = ~x44 & n3124;
  assign n3126 = ~x101 & n3125;
  assign n3127 = n3126 ^ x41;
  assign n3128 = n2467 & ~n3127;
  assign n3129 = x287 & n2401;
  assign n3130 = n2397 & n3129;
  assign n3131 = n2476 & ~n3130;
  assign n3132 = x161 & ~n1656;
  assign n3133 = n1442 & n3132;
  assign n3134 = x144 & n1656;
  assign n3135 = n1438 & n3134;
  assign n3136 = ~n3133 & ~n3135;
  assign n3137 = n3131 & ~n3136;
  assign n3138 = n2398 & ~n3137;
  assign n3139 = ~n3128 & ~n3138;
  assign n3140 = n2206 & n3125;
  assign n3141 = n2210 & n3140;
  assign n3142 = ~x114 & n3141;
  assign n3143 = n3142 ^ x42;
  assign n3144 = n2467 & n3143;
  assign n3145 = ~x189 & n1656;
  assign n3146 = ~x166 & ~n1656;
  assign n3147 = ~n3145 & ~n3146;
  assign n3148 = n3131 & ~n3147;
  assign n3149 = n2398 & ~n3148;
  assign n3150 = ~x199 & ~x200;
  assign n3151 = ~x299 & ~n3150;
  assign n3152 = n1518 & n3151;
  assign n3153 = x207 & x208;
  assign n3154 = ~x199 & ~n3153;
  assign n3155 = n3152 & ~n3154;
  assign n3156 = x212 & x214;
  assign n3157 = x211 & n3156;
  assign n3158 = ~n1656 & n3157;
  assign n3159 = ~n3155 & ~n3158;
  assign n3160 = x219 & ~n1656;
  assign n3161 = n3159 & ~n3160;
  assign n3162 = n3149 & ~n3161;
  assign n3163 = ~n3144 & ~n3162;
  assign n3164 = ~x42 & n3142;
  assign n3165 = n3164 ^ x43;
  assign n3166 = n2467 & n3165;
  assign n3171 = n3150 ^ x200;
  assign n3172 = n3153 & n3171;
  assign n3173 = n3172 ^ x200;
  assign n3167 = ~x211 & ~x219;
  assign n3168 = n3167 ^ x211;
  assign n3169 = n3156 & n3168;
  assign n3170 = n3169 ^ x211;
  assign n3174 = n3173 ^ n3170;
  assign n3175 = ~n1656 & n3174;
  assign n3176 = n3175 ^ n3173;
  assign n3177 = n3149 & n3176;
  assign n3178 = ~n3166 & ~n3177;
  assign n3179 = n3124 ^ x44;
  assign n3180 = n2467 & n3179;
  assign n3181 = n2398 & n3131;
  assign n3182 = n1439 & n1656;
  assign n3183 = n1443 & ~n1656;
  assign n3184 = ~n3182 & ~n3183;
  assign n3185 = n3181 & ~n3184;
  assign n3186 = ~n3180 & ~n3185;
  assign n3187 = x979 & n3075;
  assign n3188 = x46 & ~x109;
  assign n3189 = n2248 & n3188;
  assign n3190 = n1380 & n3189;
  assign n3191 = n1403 & n3190;
  assign n3192 = x24 & n3191;
  assign n3193 = x61 & n3053;
  assign n3194 = ~n3192 & ~n3193;
  assign n3195 = ~n1428 & ~n2219;
  assign n3196 = n3049 & n3195;
  assign n3197 = ~n3052 & ~n3057;
  assign n3198 = ~x36 & ~x88;
  assign n3199 = ~x104 & n3198;
  assign n3200 = ~n2182 & ~n3199;
  assign n3201 = ~n3197 & n3200;
  assign n3202 = n3047 & n3201;
  assign n3203 = ~n3196 & ~n3202;
  assign n3204 = x841 & n3052;
  assign n3205 = x48 & n3204;
  assign n3206 = x74 & n2482;
  assign n3207 = n1558 & n3206;
  assign n3208 = x49 & n3204;
  assign n3209 = ~n3207 & ~n3208;
  assign n3210 = n1404 & n3048;
  assign n3211 = x24 & x50;
  assign n3212 = n3210 & n3211;
  assign n3213 = ~n2309 & ~n2762;
  assign n3214 = n3020 & ~n3213;
  assign n3215 = n2307 & n3214;
  assign n3216 = ~x58 & n3048;
  assign n3217 = ~x86 & n1236;
  assign n3218 = n1358 & n3217;
  assign n3219 = n3216 & n3218;
  assign n3220 = n1233 & n3219;
  assign n3221 = n3106 & n3220;
  assign n3222 = n2480 ^ n1428;
  assign n3223 = ~x252 & n3222;
  assign n3224 = n3223 ^ n1428;
  assign n3225 = n3221 & n3224;
  assign n3226 = ~n3215 & ~n3225;
  assign n3227 = ~n3212 & n3226;
  assign n3228 = n1286 & n1287;
  assign n3229 = n1331 & n3051;
  assign n3230 = n3228 & n3229;
  assign n3231 = x82 & ~x111;
  assign n3232 = n3230 & n3231;
  assign n3233 = n2212 & n3124;
  assign n3234 = n3233 ^ x52;
  assign n3235 = n2467 & n3234;
  assign n3236 = ~x211 & x219;
  assign n3237 = ~n1656 & ~n3236;
  assign n3238 = ~x219 & n3170;
  assign n3239 = x211 & ~x219;
  assign n3240 = ~n3238 & ~n3239;
  assign n3241 = n3237 & n3240;
  assign n3242 = ~x199 & x200;
  assign n3243 = ~x299 & ~n3242;
  assign n3244 = n1518 & n3243;
  assign n3245 = ~x200 & ~n3154;
  assign n3246 = n3244 & ~n3245;
  assign n3247 = ~n3241 & ~n3246;
  assign n3248 = n3161 & ~n3247;
  assign n3249 = n3149 & n3248;
  assign n3250 = ~n3235 & ~n3249;
  assign n3251 = ~x979 & n3080;
  assign n3252 = n3075 & n3251;
  assign n3253 = n1240 & n3216;
  assign n3254 = n2142 & n3253;
  assign n3255 = x53 & ~x60;
  assign n3256 = n3254 & n3255;
  assign n3257 = x24 & n3256;
  assign n3258 = ~n3252 & ~n3257;
  assign n3259 = x24 & n1559;
  assign n3260 = n1540 & n3259;
  assign n3261 = x106 & n3053;
  assign n3262 = ~n3260 & ~n3261;
  assign n3263 = x24 & n2993;
  assign n3264 = x45 & n3052;
  assign n3265 = ~n3263 & ~n3264;
  assign n3266 = ~x62 & x841;
  assign n3267 = n1562 & n3266;
  assign n3268 = x55 & ~x56;
  assign n3269 = ~x24 & ~x62;
  assign n3270 = n3268 & n3269;
  assign n3271 = ~n3267 & ~n3270;
  assign n3272 = n1523 & ~n3271;
  assign n3273 = ~x841 & n1563;
  assign n3274 = x62 & x924;
  assign n3275 = n3273 & ~n3274;
  assign n3276 = x24 & n1527;
  assign n3277 = ~n3275 & ~n3276;
  assign n3278 = n1247 & n2249;
  assign n3279 = ~x841 & n3278;
  assign n3280 = n3273 & n3274;
  assign n3281 = ~x57 & n1516;
  assign n3282 = n2998 & n3281;
  assign n3283 = n1522 & n3282;
  assign n3284 = ~n3280 & ~n3283;
  assign n3285 = n2187 & n3081;
  assign n3286 = n3075 & n3285;
  assign n3287 = ~x53 & x60;
  assign n3288 = n3254 & n3287;
  assign n3289 = x24 & n3288;
  assign n3290 = ~n3286 & ~n3289;
  assign n3291 = x61 & n3204;
  assign n3292 = ~x24 & n3288;
  assign n3293 = ~n3291 & ~n3292;
  assign n3294 = x62 & x841;
  assign n3295 = n3294 ^ n3269;
  assign n3296 = ~x57 & n3295;
  assign n3297 = n3296 ^ n3269;
  assign n3298 = ~n1575 & n3297;
  assign n3299 = ~x24 & n3191;
  assign n3300 = x63 & n3057;
  assign n3301 = x999 & n3300;
  assign n3302 = ~n3299 & ~n3301;
  assign n3303 = x841 & n3058;
  assign n3304 = x107 & n3057;
  assign n3305 = ~n3303 & ~n3304;
  assign n3306 = n3075 & n3085;
  assign n3307 = n1334 & n3051;
  assign n3308 = x81 & n1224;
  assign n3309 = x314 & n1226;
  assign n3310 = n3308 & n3309;
  assign n3311 = n3307 & n3310;
  assign n3312 = x219 ^ x199;
  assign n3313 = x299 & n3312;
  assign n3314 = n3313 ^ x199;
  assign n3315 = n3311 & n3314;
  assign n3316 = ~x69 & n1322;
  assign n3317 = n3229 & n3316;
  assign n3318 = x314 & n3317;
  assign n3319 = x83 & ~x103;
  assign n3320 = n3318 & n3319;
  assign n3321 = n2316 & n2402;
  assign n3322 = n1702 & ~n2179;
  assign n3323 = x299 & n1675;
  assign n3324 = n2234 & n3323;
  assign n3325 = ~n3322 & ~n3324;
  assign n3326 = n3321 & ~n3325;
  assign n3327 = x69 & ~x314;
  assign n3328 = ~x71 & ~n3327;
  assign n3329 = n3052 & ~n3328;
  assign n3330 = x24 & x70;
  assign n3331 = n2269 & n3330;
  assign n3332 = n2239 & n2402;
  assign n3333 = ~n3321 & ~n3332;
  assign n3334 = n1481 & n2234;
  assign n3335 = x210 & n3334;
  assign n3336 = n1485 & ~n2179;
  assign n3337 = x198 & n3336;
  assign n3338 = ~n3335 & ~n3337;
  assign n3339 = x589 & ~n3338;
  assign n3340 = ~n3333 & n3339;
  assign n3341 = ~x593 & n3340;
  assign n3342 = n2399 & n3129;
  assign n3343 = ~n3341 & ~n3342;
  assign n3344 = ~n3331 & n3343;
  assign n3345 = n3242 ^ n3239;
  assign n3346 = ~x299 & n3345;
  assign n3347 = n3346 ^ n3239;
  assign n3348 = n3311 & n3347;
  assign n3349 = ~n1296 & n3229;
  assign n3350 = x85 & n1284;
  assign n3351 = n1307 & n3350;
  assign n3352 = ~n1303 & n3351;
  assign n3353 = x314 & n3352;
  assign n3354 = n3349 & n3353;
  assign n3355 = ~n3348 & ~n3354;
  assign n3356 = x88 & n2312;
  assign n3357 = ~n1410 & n3356;
  assign n3358 = ~x38 & ~n3357;
  assign n3359 = x72 & n1272;
  assign n3360 = x24 & n3359;
  assign n3361 = n3358 & ~n3360;
  assign n3362 = n1519 & ~n3361;
  assign n3363 = n2499 & n3321;
  assign n3364 = ~n3362 & ~n3363;
  assign n3365 = x73 & n1662;
  assign n3366 = ~n2238 & n3321;
  assign n3367 = ~n3365 & ~n3366;
  assign n3368 = ~x314 & x1050;
  assign n3369 = ~x39 & ~n3368;
  assign n3370 = ~n3367 & ~n3369;
  assign n3371 = x479 & n1259;
  assign n3372 = n2221 & ~n3371;
  assign n3373 = ~x96 & ~n3372;
  assign n3374 = ~x479 & ~x841;
  assign n3375 = x96 & ~n3374;
  assign n3376 = ~n1428 & ~n3375;
  assign n3377 = n1519 & n3376;
  assign n3378 = ~n3373 & n3377;
  assign n3379 = ~n1420 & n3378;
  assign n3380 = x74 & n3259;
  assign n3381 = ~n3379 & ~n3380;
  assign n3382 = n1437 & n1519;
  assign n3383 = x75 & n3259;
  assign n3384 = ~n3382 & ~n3383;
  assign n3385 = n2692 & n2741;
  assign n3386 = ~n3006 & ~n3385;
  assign n3387 = n2739 & n3386;
  assign n3388 = x94 & ~n2480;
  assign n3389 = ~n3387 & ~n3388;
  assign n3390 = ~x94 & ~n2741;
  assign n3391 = n1428 & ~n3390;
  assign n3392 = x94 & ~x252;
  assign n3393 = n3391 & ~n3392;
  assign n3394 = ~n3389 & ~n3393;
  assign n3395 = n1662 & n3394;
  assign n3396 = x77 & x314;
  assign n3397 = ~n1237 & ~n3396;
  assign n3398 = n2269 & n3397;
  assign n3399 = x232 & n2425;
  assign n3427 = ~x34 & n2915;
  assign n3428 = n3427 ^ x79;
  assign n3429 = ~n2785 & n3428;
  assign n3400 = ~x166 & n2788;
  assign n3401 = n2775 & n3400;
  assign n3402 = ~x163 & x299;
  assign n3403 = ~n3401 & n3402;
  assign n3404 = ~n2855 & ~n3403;
  assign n3405 = x153 & n1390;
  assign n3406 = n2281 & n3405;
  assign n3407 = ~x40 & x95;
  assign n3408 = ~n3406 & ~n3407;
  assign n3409 = x299 & ~n3408;
  assign n3410 = n1453 & n3409;
  assign n3411 = x175 & ~x299;
  assign n3412 = ~n3410 & ~n3411;
  assign n3413 = ~n3404 & n3412;
  assign n3414 = x189 ^ x166;
  assign n3415 = ~x299 & n3414;
  assign n3416 = n3415 ^ x166;
  assign n3417 = n2777 & n3416;
  assign n3418 = n2476 & ~n3417;
  assign n3419 = x182 ^ x160;
  assign n3420 = ~x299 & n3419;
  assign n3421 = n3420 ^ x160;
  assign n3422 = n2277 & ~n3421;
  assign n3423 = n3418 & ~n3422;
  assign n3424 = ~x184 & ~n2870;
  assign n3425 = n3423 & ~n3424;
  assign n3426 = ~n3413 & n3425;
  assign n3430 = n3429 ^ n3426;
  assign n3431 = ~n2778 & ~n3430;
  assign n3432 = n3431 ^ n3429;
  assign n3433 = ~x39 & n3432;
  assign n3434 = ~n2816 & ~n3429;
  assign n3435 = ~x189 & n2799;
  assign n3436 = ~x166 & n2801;
  assign n3437 = ~n3435 & ~n3436;
  assign n3438 = n2316 & ~n3437;
  assign n3439 = x179 & n2799;
  assign n3440 = x156 & n2801;
  assign n3441 = ~n3439 & ~n3440;
  assign n3442 = n2239 & ~n3441;
  assign n3443 = ~n3438 & ~n3442;
  assign n3444 = n2476 & ~n3443;
  assign n3445 = n2813 & n3444;
  assign n3446 = x39 & ~n3445;
  assign n3447 = ~n3434 & n3446;
  assign n3448 = n1512 & n2788;
  assign n3449 = ~x38 & n3448;
  assign n3450 = ~n3447 & n3449;
  assign n3451 = ~n3433 & n3450;
  assign n3452 = ~n2820 & n3429;
  assign n3453 = n2788 & ~n3452;
  assign n3454 = x179 ^ x156;
  assign n3455 = ~x299 & n3454;
  assign n3456 = n3455 ^ x156;
  assign n3457 = n2476 & n3456;
  assign n3458 = n2820 & ~n3457;
  assign n3459 = n3453 & ~n3458;
  assign n3460 = n1511 & ~n3459;
  assign n3461 = ~n1532 & ~n3460;
  assign n3462 = ~x40 & ~n2833;
  assign n3463 = ~n3461 & n3462;
  assign n3464 = ~n3451 & n3463;
  assign n3469 = n2982 ^ x197;
  assign n3470 = n2981 & n3469;
  assign n3471 = n3470 ^ x162;
  assign n3472 = n3471 ^ x163;
  assign n3465 = n2987 ^ x145;
  assign n3466 = n2986 & n3465;
  assign n3467 = n3466 ^ x140;
  assign n3468 = n3467 ^ x184;
  assign n3473 = n3472 ^ n3468;
  assign n3474 = ~x299 & n3473;
  assign n3475 = n3474 ^ n3472;
  assign n3476 = n2845 & n3475;
  assign n3477 = n1509 & ~n1510;
  assign n3478 = x187 ^ x147;
  assign n3479 = ~x299 & n3478;
  assign n3480 = n3479 ^ x147;
  assign n3481 = n2476 & n3480;
  assign n3482 = n3477 & ~n3481;
  assign n3483 = ~n3476 & ~n3482;
  assign n3484 = ~n3464 & n3483;
  assign n3485 = n1518 & ~n3484;
  assign n3486 = x163 & n2476;
  assign n3487 = n3486 ^ n3429;
  assign n3488 = n2912 & ~n3487;
  assign n3489 = n3488 ^ n3429;
  assign n3490 = n2788 & ~n3489;
  assign n3491 = ~x40 & ~n1516;
  assign n3492 = n2891 & n3491;
  assign n3493 = ~n3490 & n3492;
  assign n3494 = n2845 & n3472;
  assign n3495 = x147 & n2476;
  assign n3496 = n1509 & ~n3495;
  assign n3497 = ~n3494 & ~n3496;
  assign n3498 = ~n1518 & ~n2891;
  assign n3499 = ~n3497 & n3498;
  assign n3500 = ~n3493 & ~n3499;
  assign n3501 = ~n3485 & n3500;
  assign n3502 = ~x63 & ~n2250;
  assign n3503 = n1575 & ~n3502;
  assign n3504 = ~x592 & ~n2681;
  assign n3505 = n2662 & ~n3504;
  assign n3506 = ~x588 & ~x590;
  assign n3507 = n2660 & ~n3506;
  assign n3508 = ~n2692 & ~n2721;
  assign n3509 = x590 & n2692;
  assign n3510 = x98 & ~x592;
  assign n3511 = x1199 & n3510;
  assign n3512 = ~n3509 & ~n3511;
  assign n3513 = ~n3508 & ~n3512;
  assign n3514 = ~n3507 & ~n3513;
  assign n3515 = n3505 & n3514;
  assign n3516 = n2396 & n2712;
  assign n3517 = ~n3515 & n3516;
  assign n3518 = ~n2470 & n3517;
  assign n3519 = ~n3503 & n3518;
  assign n3520 = n3505 & ~n3511;
  assign n3521 = n2728 & ~n3520;
  assign n3522 = ~n3519 & ~n3521;
  assign n3523 = n2641 & ~n3522;
  assign n3524 = ~n2697 & ~n3523;
  assign n3525 = ~x80 & n2699;
  assign n3526 = ~n3524 & n3525;
  assign n3527 = x81 & ~x314;
  assign n3528 = ~x68 & ~n3527;
  assign n3529 = ~n3197 & ~n3528;
  assign n3530 = x314 ^ x66;
  assign n3531 = x69 & n3530;
  assign n3532 = n3531 ^ x66;
  assign n3533 = n3052 & n3532;
  assign n3534 = ~x68 & x84;
  assign n3535 = n1229 & n3534;
  assign n3536 = n3349 & n3535;
  assign n3537 = ~x314 & n3319;
  assign n3538 = n3317 & n3537;
  assign n3539 = ~n3536 & ~n3538;
  assign n3540 = n3167 ^ n3150;
  assign n3541 = x299 & n3540;
  assign n3542 = n3541 ^ n3150;
  assign n3543 = n3311 & n3542;
  assign n3544 = ~x314 & n3352;
  assign n3545 = ~x67 & ~n3544;
  assign n3546 = n3349 & ~n3545;
  assign n3547 = ~n3325 & n3332;
  assign n3548 = n2260 & n3318;
  assign n3549 = x104 & n2182;
  assign n3550 = n3052 & n3549;
  assign n3551 = n2692 & n3550;
  assign n3552 = x88 & n2219;
  assign n3553 = n3057 & n3552;
  assign n3554 = ~n3551 & ~n3553;
  assign n3555 = x89 & x841;
  assign n3556 = ~x24 & x70;
  assign n3557 = ~n3555 & ~n3556;
  assign n3558 = n2269 & ~n3557;
  assign n3559 = ~x1050 & n3365;
  assign n3560 = x841 & n3278;
  assign n3561 = ~n3559 & ~n3560;
  assign n3562 = ~x24 & ~n1431;
  assign n3563 = n2450 & ~n3562;
  assign n3564 = n1431 & n3046;
  assign n3565 = ~n3563 & ~n3564;
  assign n3566 = n3216 & ~n3565;
  assign n3567 = n2402 & n2500;
  assign n3568 = ~n3566 & ~n3567;
  assign n3569 = ~x39 & x92;
  assign n3570 = n3368 & n3569;
  assign n3571 = ~n2241 & ~n3570;
  assign n3572 = n1573 & ~n3571;
  assign n3573 = n2145 & n2269;
  assign n3574 = n1551 & n1596;
  assign n3575 = ~x1050 & n3574;
  assign n3576 = ~n3573 & ~n3575;
  assign n3577 = x49 & n3053;
  assign n3578 = ~n1428 & n2481;
  assign n3579 = n3221 & n3578;
  assign n3580 = ~n3577 & ~n3579;
  assign n3581 = ~n3334 & ~n3336;
  assign n3582 = ~n3333 & ~n3581;
  assign n3583 = ~n3339 & n3582;
  assign n3584 = x89 & ~x332;
  assign n3585 = n3053 & n3584;
  assign n3586 = ~n3583 & ~n3585;
  assign n3587 = ~x32 & ~x40;
  assign n3588 = n1519 & n3587;
  assign n3589 = x95 & n3588;
  assign n3590 = n1254 & n3589;
  assign n3591 = x24 & n3590;
  assign n3592 = n3586 & ~n3591;
  assign n3593 = ~n1254 & n1410;
  assign n3594 = ~x95 & n3375;
  assign n3595 = ~n1429 & n3594;
  assign n3596 = ~x24 & x95;
  assign n3597 = ~x96 & n3596;
  assign n3598 = ~n3595 & ~n3597;
  assign n3599 = n3588 & ~n3598;
  assign n3600 = ~n3593 & n3599;
  assign n3601 = ~n1431 & ~n3372;
  assign n3602 = n3048 & n3601;
  assign n3603 = n1416 & n3602;
  assign n3604 = x593 & n3340;
  assign n3605 = ~n3603 & ~n3604;
  assign n3606 = ~n3365 & ~n3574;
  assign n3607 = x314 & x1050;
  assign n3608 = ~n3606 & n3607;
  assign n3609 = n2204 & n3125;
  assign n3610 = n3609 ^ x99;
  assign n3611 = n2467 & n3610;
  assign n3612 = x152 & n3146;
  assign n3613 = x161 & n3612;
  assign n3614 = x174 & n3145;
  assign n3615 = x144 & n3614;
  assign n3616 = ~n3613 & ~n3615;
  assign n3617 = n3181 & ~n3616;
  assign n3618 = ~n3611 & ~n3617;
  assign n3619 = n1446 & ~n2182;
  assign n3620 = x683 & ~n3619;
  assign n3621 = ~n2223 & ~n3620;
  assign n3622 = n2480 & n3621;
  assign n3623 = n2757 & ~n3622;
  assign n3624 = n2308 & ~n3623;
  assign n3625 = n1428 & n2761;
  assign n3626 = ~n2760 & n3625;
  assign n3627 = ~n3624 & ~n3626;
  assign n3628 = n2307 & ~n3627;
  assign n3629 = n3125 ^ x101;
  assign n3630 = n2467 & n3629;
  assign n3631 = ~x161 & n3612;
  assign n3632 = ~x144 & n3614;
  assign n3633 = ~n3631 & ~n3632;
  assign n3634 = n3181 & ~n3633;
  assign n3635 = ~n3630 & ~n3634;
  assign n3636 = x65 & n3057;
  assign n3637 = n1662 & ~n2265;
  assign n3638 = ~n2692 & n3550;
  assign n3639 = n3108 & n3220;
  assign n3640 = ~n3027 & n3639;
  assign n3641 = ~n3638 & ~n3640;
  assign n3642 = x106 & n3204;
  assign n3643 = ~x24 & n3256;
  assign n3644 = ~n3642 & ~n3643;
  assign n3645 = ~x999 & n3300;
  assign n3646 = ~n2400 & ~n3503;
  assign n3647 = x108 & ~n3066;
  assign n3648 = ~x98 & ~n3647;
  assign n3649 = n3210 & ~n3648;
  assign n3650 = ~n3646 & ~n3649;
  assign n3651 = n3210 & n3396;
  assign n3652 = n2260 & n3230;
  assign n3653 = x314 & n3652;
  assign n3654 = n3027 & n3639;
  assign n3655 = ~n3653 & ~n3654;
  assign n3656 = ~x24 & n1519;
  assign n3657 = n3359 & n3656;
  assign n3658 = ~x314 & n3652;
  assign n3659 = ~n3657 & ~n3658;
  assign n3660 = x124 & ~x468;
  assign n3661 = n2205 & n3125;
  assign n3662 = n3661 ^ x113;
  assign n3663 = n2467 & n3662;
  assign n3664 = n3141 ^ x114;
  assign n3665 = n2467 & n3664;
  assign n3666 = ~x116 & n3140;
  assign n3667 = n3666 ^ x115;
  assign n3668 = n2467 & n3667;
  assign n3669 = n3140 ^ x116;
  assign n3670 = n2467 & n3669;
  assign n3671 = x190 & n2316;
  assign n3672 = x178 & n2239;
  assign n3673 = ~n3671 & ~n3672;
  assign n3674 = n2799 & ~n3673;
  assign n3675 = x168 & n2316;
  assign n3676 = x157 & n2239;
  assign n3677 = ~n3675 & ~n3676;
  assign n3678 = n2801 & ~n3677;
  assign n3679 = ~n3674 & ~n3678;
  assign n3680 = x39 & ~x92;
  assign n3681 = ~n3679 & n3680;
  assign n3682 = x178 ^ x157;
  assign n3683 = ~x299 & n3682;
  assign n3684 = n3683 ^ x157;
  assign n3685 = n3569 & n3684;
  assign n3686 = ~n3681 & ~n3685;
  assign n3687 = ~x87 & n2476;
  assign n3688 = n2813 & n3687;
  assign n3689 = ~n3686 & n3688;
  assign n3690 = n2789 & ~n3689;
  assign n3691 = n1514 & ~n2778;
  assign n3711 = ~x38 & x39;
  assign n3712 = n2815 & n3711;
  assign n3713 = ~x92 & ~n1533;
  assign n3714 = ~n3712 & n3713;
  assign n3715 = ~x54 & n1509;
  assign n3716 = ~n1512 & ~n1537;
  assign n3717 = n3715 & ~n3716;
  assign n3718 = ~n3714 & n3717;
  assign n3719 = n1521 & n3718;
  assign n3720 = ~x954 & n2784;
  assign n3721 = ~n2781 & n3720;
  assign n3722 = ~x79 & n3427;
  assign n3723 = x118 & ~n3722;
  assign n3724 = ~n3721 & ~n3723;
  assign n3725 = n1511 & ~n3724;
  assign n3726 = ~n3719 & ~n3725;
  assign n3692 = x173 ^ x151;
  assign n3693 = ~x299 & n3692;
  assign n3694 = n3693 ^ x151;
  assign n3695 = n2855 & ~n3694;
  assign n3696 = n2476 & ~n3695;
  assign n3697 = ~n2277 & ~n3696;
  assign n3698 = ~x150 & ~n2873;
  assign n3699 = x73 & ~x168;
  assign n3700 = ~n3698 & ~n3699;
  assign n3701 = x299 & ~n3700;
  assign n3702 = ~x73 & x232;
  assign n3703 = n1205 & n3702;
  assign n3704 = n2873 & ~n3703;
  assign n3705 = ~x185 & ~x299;
  assign n3706 = ~n3704 & n3705;
  assign n3707 = ~x190 & n2878;
  assign n3708 = ~n3706 & ~n3707;
  assign n3709 = ~n3701 & n3708;
  assign n3710 = ~n3697 & n3709;
  assign n3727 = n3726 ^ n3710;
  assign n3728 = n3691 & n3727;
  assign n3729 = n3728 ^ n3726;
  assign n3730 = n3690 & ~n3729;
  assign n3731 = ~x163 & ~n3471;
  assign n3732 = n3731 ^ x150;
  assign n3733 = n2845 & ~n3732;
  assign n3734 = n1509 & ~n2890;
  assign n3735 = x165 & n2476;
  assign n3736 = n3734 & ~n3735;
  assign n3737 = ~n3733 & ~n3736;
  assign n3738 = ~n1656 & ~n3737;
  assign n3739 = ~n2476 & n3734;
  assign n3740 = n1516 & ~n3739;
  assign n3741 = ~n3738 & n3740;
  assign n3742 = ~x184 & ~n3467;
  assign n3743 = n3742 ^ x185;
  assign n3744 = n2845 & ~n3743;
  assign n3745 = ~x143 & n3477;
  assign n3746 = ~n3744 & ~n3745;
  assign n3747 = ~x299 & ~n3746;
  assign n3748 = n3741 & ~n3747;
  assign n3749 = ~n3730 & n3748;
  assign n3750 = x150 & n2476;
  assign n3751 = n3750 ^ n3724;
  assign n3752 = n2893 & n3751;
  assign n3753 = n3752 ^ n3724;
  assign n3754 = n2892 & ~n3753;
  assign n3755 = ~n1518 & n3737;
  assign n3756 = ~n3754 & n3755;
  assign n3757 = ~n3749 & ~n3756;
  assign n3758 = ~x109 & n1237;
  assign n3759 = n1385 & ~n3758;
  assign n3760 = ~n2304 & n3759;
  assign n3761 = n1390 & ~n1435;
  assign n3762 = ~n3760 & n3761;
  assign n3763 = n1662 & ~n3762;
  assign n3764 = n1618 & n2307;
  assign n3765 = ~n2495 & n3332;
  assign n3766 = ~n3574 & ~n3765;
  assign n3767 = ~n3764 & n3766;
  assign n3768 = ~n3763 & n3767;
  assign n3769 = n3768 ^ x128;
  assign n3770 = ~x228 & ~n3769;
  assign n3771 = n3770 ^ x128;
  assign n3772 = n1518 & ~n2510;
  assign n3773 = ~n2474 & n3772;
  assign n3774 = ~n2728 & ~n3773;
  assign n3775 = ~x31 & ~x80;
  assign n3776 = x818 & n3775;
  assign n3777 = x1093 & n3776;
  assign n3778 = x951 & x982;
  assign n3779 = n2695 & n3778;
  assign n3780 = n2699 & n3779;
  assign n3781 = ~n3777 & ~n3780;
  assign n3782 = ~x120 & n3781;
  assign n3783 = n3774 & ~n3782;
  assign n3784 = ~x24 & n3396;
  assign n3785 = n2862 & n3784;
  assign n3786 = n2269 & n3785;
  assign n3787 = x181 & n2231;
  assign n3788 = x159 & n2236;
  assign n3789 = ~n3787 & ~n3788;
  assign n3790 = n3075 & ~n3789;
  assign n3791 = ~n3132 & ~n3134;
  assign n3792 = n2400 & ~n3791;
  assign n3793 = ~n2401 & ~n3792;
  assign n3794 = x163 & ~n1656;
  assign n3795 = x87 & ~n3794;
  assign n3796 = x184 & n1656;
  assign n3797 = n3795 & ~n3796;
  assign n3798 = ~x146 & ~n1656;
  assign n3799 = n1440 & n1518;
  assign n3800 = x51 & ~x87;
  assign n3801 = ~n3799 & n3800;
  assign n3802 = ~n3798 & n3801;
  assign n3803 = ~n3797 & ~n3802;
  assign n3804 = n3793 & n3803;
  assign n3805 = ~n3790 & ~n3804;
  assign n3806 = ~n3786 & n3805;
  assign n3807 = n2476 & ~n3806;
  assign n3808 = x24 & x77;
  assign n3809 = ~x86 & ~n3808;
  assign n3810 = ~n3396 & n3809;
  assign n3811 = ~x39 & ~n3810;
  assign n3812 = n2396 & n3811;
  assign n3813 = n1418 & n3812;
  assign n3814 = n1379 & n3813;
  assign n3815 = n3457 & ~n3784;
  assign n3816 = n3814 & ~n3815;
  assign n3817 = n2401 & ~n3816;
  assign n3818 = x72 ^ x39;
  assign n3819 = n2397 & n3818;
  assign n3820 = x39 & n2317;
  assign n3821 = n3819 & ~n3820;
  assign n3822 = ~x125 & ~x133;
  assign n3823 = n3822 ^ x121;
  assign n3824 = ~x134 & ~x135;
  assign n3825 = ~x136 & n3824;
  assign n3826 = ~x130 & n3825;
  assign n3827 = ~x126 & ~x132;
  assign n3828 = n3826 & n3827;
  assign n3829 = n3822 & n3828;
  assign n3830 = n3823 & n3829;
  assign n3831 = n3830 ^ n3823;
  assign n3832 = ~n3821 & ~n3831;
  assign n3833 = ~n3814 & ~n3832;
  assign n3834 = n3817 & ~n3833;
  assign n3835 = ~n3807 & ~n3834;
  assign n3836 = ~x90 & ~x111;
  assign n3837 = ~x72 & n3836;
  assign n3838 = n2258 & n3837;
  assign n3839 = n2269 & ~n3838;
  assign n3840 = x39 & ~x110;
  assign n3841 = n2408 & n3840;
  assign n3842 = n2476 & ~n3184;
  assign n3843 = ~x39 & x110;
  assign n3844 = n2182 & n3843;
  assign n3845 = ~n2213 & n3844;
  assign n3846 = ~n3842 & n3845;
  assign n3847 = ~n3841 & ~n3846;
  assign n3848 = ~n3839 & n3847;
  assign n3849 = ~n1410 & ~n3810;
  assign n3850 = ~x39 & ~n3359;
  assign n3851 = ~n3849 & n3850;
  assign n3852 = n2395 & ~n3851;
  assign n3853 = ~x287 & n2476;
  assign n3854 = x158 & n1671;
  assign n3855 = n3853 & n3854;
  assign n3856 = n2498 & ~n3855;
  assign n3857 = n1521 & ~n3856;
  assign n3858 = ~x51 & ~n1232;
  assign n3859 = ~x152 & n3858;
  assign n3860 = x51 & x172;
  assign n3861 = ~n3859 & ~n3860;
  assign n3862 = x299 & n3861;
  assign n3863 = n2476 & ~n3862;
  assign n3864 = ~n3857 & ~n3863;
  assign n3865 = ~x72 & n2394;
  assign n3866 = x180 & ~x287;
  assign n3867 = n2161 & n3866;
  assign n3868 = x224 & ~n3867;
  assign n3869 = ~x51 & x222;
  assign n3870 = ~x223 & n3869;
  assign n3871 = n1232 & n3870;
  assign n3872 = ~n3868 & n3871;
  assign n3873 = n3865 & n3872;
  assign n3874 = ~x174 & n3858;
  assign n3875 = x51 & x193;
  assign n3876 = ~x299 & ~n3875;
  assign n3877 = ~n3874 & n3876;
  assign n3878 = ~n3873 & n3877;
  assign n3879 = ~n3864 & ~n3878;
  assign n3880 = x39 & ~n3879;
  assign n3881 = n3852 & ~n3880;
  assign n3882 = n3863 & ~n3877;
  assign n3883 = ~x121 & ~x125;
  assign n3884 = n3828 & n3883;
  assign n3885 = x133 ^ x125;
  assign n3886 = ~n3884 & ~n3885;
  assign n3887 = n2401 & ~n3886;
  assign n3888 = ~n3882 & ~n3887;
  assign n3889 = ~n3881 & n3888;
  assign n3890 = n1511 & n3680;
  assign n3891 = ~n2319 & n3890;
  assign n3892 = n3865 & n3891;
  assign n3893 = ~n3879 & n3892;
  assign n3894 = ~x87 & ~n3893;
  assign n3895 = ~n3889 & n3894;
  assign n3896 = x87 & n2476;
  assign n3897 = x162 ^ x140;
  assign n3898 = x299 & n3897;
  assign n3899 = n3898 ^ x140;
  assign n3900 = n3896 & n3899;
  assign n3901 = n1518 & ~n3900;
  assign n3902 = ~n3895 & n3901;
  assign n3903 = n1514 & n3814;
  assign n3904 = x197 ^ x145;
  assign n3905 = x299 & n3904;
  assign n3906 = n3905 ^ x145;
  assign n3907 = n3906 ^ n2926;
  assign n3908 = n3809 & n3907;
  assign n3909 = n3908 ^ n2926;
  assign n3910 = n2476 & n3909;
  assign n3911 = n3903 & ~n3910;
  assign n3912 = n3687 & ~n3861;
  assign n3913 = x162 & n3896;
  assign n3914 = ~n1518 & ~n3913;
  assign n3915 = ~n3912 & n3914;
  assign n3916 = ~n3887 & n3915;
  assign n3917 = ~n3911 & ~n3916;
  assign n3918 = ~n3902 & n3917;
  assign n3919 = ~x121 & n3822;
  assign n3920 = n3919 ^ x126;
  assign n3921 = n2401 & n3920;
  assign n3922 = ~n3828 & n3921;
  assign n3923 = ~n3903 & ~n3922;
  assign n3924 = ~n3821 & ~n3923;
  assign n3925 = x160 & n3853;
  assign n3926 = n2236 & ~n3925;
  assign n3927 = x182 & n3853;
  assign n3928 = n2231 & ~n3927;
  assign n3929 = ~n3926 & ~n3928;
  assign n3930 = n2399 & ~n3929;
  assign n3931 = x166 ^ x153;
  assign n3932 = ~x51 & ~n3931;
  assign n3933 = n3932 ^ x153;
  assign n3934 = n3687 & n3933;
  assign n3935 = ~n1518 & n3934;
  assign n3936 = ~n2401 & ~n3935;
  assign n3937 = ~n3930 & ~n3936;
  assign n3938 = ~n3924 & n3937;
  assign n3939 = n3684 ^ n2957;
  assign n3940 = ~n3809 & n3939;
  assign n3941 = n3940 ^ n2957;
  assign n3942 = n3903 & n3941;
  assign n3943 = ~n3416 & n3858;
  assign n3944 = x51 & n3411;
  assign n3945 = x51 & x153;
  assign n3946 = x299 & n3945;
  assign n3947 = ~n3944 & ~n3946;
  assign n3948 = ~n3943 & n3947;
  assign n3949 = ~x87 & n1518;
  assign n3950 = ~n3948 & n3949;
  assign n3951 = ~x150 & ~n1656;
  assign n3952 = n1518 & n3705;
  assign n3953 = x87 & ~n3952;
  assign n3954 = ~n3951 & n3953;
  assign n3955 = ~n3950 & ~n3954;
  assign n3956 = ~n3942 & n3955;
  assign n3957 = n2476 & ~n3956;
  assign n3958 = ~n3938 & ~n3957;
  assign n3959 = x250 & n2481;
  assign n3960 = x127 & ~n3959;
  assign n3961 = x94 & ~n3960;
  assign n3962 = n2221 & n3959;
  assign n3963 = n3961 & ~n3962;
  assign n3964 = x129 & ~n3963;
  assign n3965 = ~n3503 & n3964;
  assign n3966 = ~x100 & ~n2481;
  assign n3967 = ~x250 & ~n3966;
  assign n3968 = x129 & ~n3967;
  assign n3969 = ~n1508 & ~n3968;
  assign n3970 = n2221 & n3967;
  assign n3971 = n3969 & ~n3970;
  assign n3972 = ~n1575 & ~n3971;
  assign n3973 = ~n1662 & ~n3972;
  assign n3974 = x140 & n1698;
  assign n3975 = n1671 & n2949;
  assign n3976 = ~n3974 & ~n3975;
  assign n3977 = n3853 & ~n3976;
  assign n3978 = n2498 & ~n3977;
  assign n3979 = n1521 & ~n3978;
  assign n3980 = x39 & ~n3979;
  assign n3981 = n3852 & ~n3980;
  assign n3982 = n3827 & n3919;
  assign n3983 = ~x130 & n3982;
  assign n3984 = ~n3825 & n3983;
  assign n3985 = x130 & ~n3982;
  assign n3986 = n1232 & ~n3985;
  assign n3987 = ~n3984 & n3986;
  assign n3988 = ~n3892 & n3987;
  assign n3989 = ~n1232 & n2841;
  assign n3990 = ~n3988 & ~n3989;
  assign n3991 = n3949 & n3990;
  assign n3992 = ~n3981 & n3991;
  assign n3993 = ~n1232 & n2476;
  assign n3994 = x169 & n3993;
  assign n3995 = ~n1518 & ~n3896;
  assign n3996 = ~n3994 & n3995;
  assign n3997 = ~n3987 & n3996;
  assign n3998 = ~n3992 & ~n3997;
  assign n3999 = ~x51 & ~n3998;
  assign n4000 = ~x167 & ~n1656;
  assign n4001 = ~x188 & ~x299;
  assign n4002 = n1518 & n4001;
  assign n4003 = n2476 & ~n4002;
  assign n4004 = ~n4000 & n4003;
  assign n4005 = x87 & ~n4004;
  assign n4006 = ~n3999 & ~n4005;
  assign n4007 = ~n2319 & n2399;
  assign n4008 = n2401 & ~n4007;
  assign n4009 = ~n3814 & n4008;
  assign n4010 = n2476 & n3421;
  assign n4011 = ~x24 & x77;
  assign n4012 = ~n4010 & n4011;
  assign n4013 = x149 & n2235;
  assign n4014 = x183 & n1698;
  assign n4015 = ~n4013 & ~n4014;
  assign n4016 = ~n4012 & ~n4015;
  assign n4017 = n3853 & n4016;
  assign n4018 = n2401 & n4017;
  assign n4019 = ~n4009 & ~n4018;
  assign n4020 = ~n3826 & n3982;
  assign n4021 = ~x126 & n3919;
  assign n4022 = x132 & ~n4021;
  assign n4023 = ~n4020 & ~n4022;
  assign n4024 = ~n3821 & ~n4023;
  assign n4025 = ~n4019 & ~n4024;
  assign n4026 = n3903 & ~n4012;
  assign n4027 = ~x190 & n1656;
  assign n4028 = ~n1232 & ~n4027;
  assign n4029 = ~x168 & ~n1656;
  assign n4030 = n4028 & ~n4029;
  assign n4031 = n2400 & ~n4030;
  assign n4032 = x173 & n1656;
  assign n4033 = n3800 & ~n4032;
  assign n4034 = x151 & ~n1656;
  assign n4035 = n4033 & ~n4034;
  assign n4036 = x164 & ~n1656;
  assign n4037 = n1518 & n2792;
  assign n4038 = x87 & ~n4037;
  assign n4039 = ~n4036 & n4038;
  assign n4040 = n2476 & ~n4039;
  assign n4041 = ~n4035 & n4040;
  assign n4042 = ~n4031 & n4041;
  assign n4043 = ~n4026 & ~n4042;
  assign n4044 = ~n4025 & n4043;
  assign n4045 = x145 & n1698;
  assign n4046 = x197 & x299;
  assign n4047 = n1671 & n4046;
  assign n4048 = ~n4045 & ~n4047;
  assign n4049 = n3853 & ~n4048;
  assign n4050 = ~x72 & n2498;
  assign n4051 = ~n4049 & n4050;
  assign n4052 = n3818 & ~n4051;
  assign n4053 = ~n3503 & n4052;
  assign n4061 = ~x86 & n2745;
  assign n4062 = ~n2824 & ~n4061;
  assign n4054 = ~x133 & ~n3884;
  assign n4055 = n4008 & ~n4054;
  assign n4056 = ~x149 & ~n1656;
  assign n4057 = n3896 & ~n4056;
  assign n4058 = ~x183 & n1656;
  assign n4059 = n4057 & ~n4058;
  assign n4060 = ~n4055 & ~n4059;
  assign n4063 = n4062 ^ n4060;
  assign n4064 = ~n3903 & n4063;
  assign n4065 = n4064 ^ n4062;
  assign n4066 = ~n4053 & n4065;
  assign n4067 = n2400 & ~n3814;
  assign n4068 = ~x136 & n3983;
  assign n4069 = ~x135 & n4068;
  assign n4070 = x134 & ~n4069;
  assign n4071 = ~n3821 & ~n4070;
  assign n4072 = x186 & n1698;
  assign n4073 = n1671 & n2791;
  assign n4074 = ~n4072 & ~n4073;
  assign n4075 = n3853 & ~n4074;
  assign n4076 = n4050 & ~n4075;
  assign n4077 = n3819 & ~n4076;
  assign n4078 = ~n4071 & ~n4077;
  assign n4079 = n1232 & ~n4078;
  assign n4080 = x192 ^ x171;
  assign n4081 = n1656 & n4080;
  assign n4082 = n4081 ^ x171;
  assign n4083 = n3993 & n4082;
  assign n4084 = ~n4079 & ~n4083;
  assign n4085 = n4067 & n4084;
  assign n4086 = x150 & n2235;
  assign n4087 = x185 & n1698;
  assign n4088 = ~n4086 & ~n4087;
  assign n4089 = n3853 & ~n4088;
  assign n4090 = n4007 & ~n4089;
  assign n4091 = n1232 & ~n4090;
  assign n4092 = n4068 ^ x135;
  assign n4093 = n4068 & n4092;
  assign n4094 = ~x134 & n4093;
  assign n4095 = n4094 ^ n4092;
  assign n4096 = ~n3821 & n4095;
  assign n4097 = n4091 & ~n4096;
  assign n4098 = x194 ^ x170;
  assign n4099 = n1656 & n4098;
  assign n4100 = n4099 ^ x170;
  assign n4101 = n3993 & n4100;
  assign n4102 = ~n4097 & ~n4101;
  assign n4103 = n4067 & n4102;
  assign n4104 = x163 & n2235;
  assign n4105 = x184 & n1698;
  assign n4106 = ~n4104 & ~n4105;
  assign n4107 = n3853 & ~n4106;
  assign n4108 = n2498 & ~n4107;
  assign n4109 = n3865 & ~n4108;
  assign n4110 = x39 & n1232;
  assign n4111 = ~n4109 & n4110;
  assign n4112 = n2476 & n2971;
  assign n4113 = ~n1232 & ~n4112;
  assign n4114 = n2396 & ~n4113;
  assign n4115 = ~n4111 & n4114;
  assign n4116 = ~n3851 & n4115;
  assign n4117 = ~x148 & ~n1656;
  assign n4118 = n3993 & ~n4117;
  assign n4119 = ~x141 & n1656;
  assign n4120 = n4118 & ~n4119;
  assign n4121 = ~n3824 & n4068;
  assign n4122 = x136 & ~n3983;
  assign n4123 = n1232 & ~n4122;
  assign n4124 = ~n4121 & n4123;
  assign n4125 = ~n4120 & ~n4124;
  assign n4126 = ~n4007 & ~n4125;
  assign n4127 = n2400 & ~n4126;
  assign n4128 = ~n4116 & n4127;
  assign n4129 = ~x198 & n3182;
  assign n4130 = ~x210 & n3183;
  assign n4131 = ~n4129 & ~n4130;
  assign n4132 = x39 & n2476;
  assign n4133 = ~n4131 & n4132;
  assign n4134 = ~n3149 & n4133;
  assign n4135 = ~x39 & x137;
  assign n4136 = ~n4134 & ~n4135;
  assign n4137 = ~x39 & ~n2774;
  assign n4138 = n2241 & n2813;
  assign n4139 = ~n4137 & ~n4138;
  assign n4140 = n1512 & n1516;
  assign n4141 = ~n4139 & n4140;
  assign n4142 = n1560 & n2892;
  assign n4143 = ~n4141 & n4142;
  assign n4144 = n3367 & n4143;
  assign n4145 = n2780 & n3720;
  assign n4146 = ~n2779 & n4145;
  assign n4147 = ~x139 & n3720;
  assign n4148 = x138 & ~n4147;
  assign n4149 = ~n4146 & ~n4148;
  assign n4150 = n4144 & ~n4149;
  assign n4151 = ~n3367 & ~n4112;
  assign n4152 = ~n4150 & ~n4151;
  assign n4153 = n3720 ^ x139;
  assign n4154 = ~n2781 & n4153;
  assign n4155 = n4144 & n4154;
  assign n4156 = ~n2841 & ~n3367;
  assign n4157 = ~n4155 & ~n4156;
  assign n4158 = ~n2183 & n3073;
  assign n4159 = x35 & ~x93;
  assign n4160 = ~x841 & n4159;
  assign n4161 = n1405 & n4160;
  assign n4162 = ~x45 & ~x47;
  assign n4163 = ~x102 & n4162;
  assign n4164 = ~n3065 & n4163;
  assign n4165 = ~n4161 & n4164;
  assign n4166 = ~x47 & ~n1229;
  assign n4167 = ~x252 & ~n4166;
  assign n4168 = ~n4165 & ~n4167;
  assign n4169 = ~x40 & ~n4168;
  assign n4170 = ~n4158 & n4169;
  assign n4171 = n3358 & n4170;
  assign n4172 = ~n3503 & ~n4171;
  assign n4173 = ~n2495 & ~n3333;
  assign n4174 = ~x287 & ~n3082;
  assign n4175 = ~x120 & ~n4174;
  assign n4176 = ~n2202 & ~n4175;
  assign n4177 = n2402 & n4176;
  assign n4178 = ~n4173 & ~n4177;
  assign n4179 = ~n4172 & n4178;
  assign n4180 = n2695 & ~n4179;
  assign n4181 = x832 & n2695;
  assign n4182 = ~n4180 & ~n4181;
  assign n4183 = x1154 ^ x618;
  assign n4184 = x781 & n4183;
  assign n4185 = x1155 ^ x609;
  assign n4186 = x785 & n4185;
  assign n4187 = ~n4184 & ~n4186;
  assign n4188 = x1157 ^ x630;
  assign n4189 = x787 & n4188;
  assign n4190 = x1158 ^ x626;
  assign n4191 = x788 & n4190;
  assign n4192 = ~n4189 & ~n4191;
  assign n4193 = n4187 & n4192;
  assign n4194 = x1160 ^ x644;
  assign n4195 = x790 & n4194;
  assign n4196 = x603 & ~n4195;
  assign n4197 = n4193 & n4196;
  assign n4198 = x1159 ^ x619;
  assign n4199 = x789 & n4198;
  assign n4200 = x1153 ^ x608;
  assign n4201 = x778 & n4200;
  assign n4202 = ~n4199 & ~n4201;
  assign n4203 = x1156 ^ x629;
  assign n4204 = x792 & n4203;
  assign n4205 = n4202 & ~n4204;
  assign n4206 = n4197 & n4205;
  assign n4207 = x621 & x1091;
  assign n4208 = n4206 & ~n4207;
  assign n4209 = x1160 ^ x715;
  assign n4210 = x790 & n4209;
  assign n4211 = x1158 ^ x641;
  assign n4212 = x788 & n4211;
  assign n4213 = ~n4210 & ~n4212;
  assign n4214 = x1153 ^ x625;
  assign n4215 = x778 & n4214;
  assign n4216 = n4213 & ~n4215;
  assign n4217 = x1155 ^ x660;
  assign n4218 = x785 & n4217;
  assign n4219 = x680 & ~n4218;
  assign n4220 = x1154 ^ x627;
  assign n4221 = x781 & n4220;
  assign n4222 = x1157 ^ x647;
  assign n4223 = x787 & n4222;
  assign n4224 = ~n4221 & ~n4223;
  assign n4225 = n4219 & n4224;
  assign n4226 = n4216 & n4225;
  assign n4227 = x1156 ^ x628;
  assign n4228 = x792 & n4227;
  assign n4229 = x1159 ^ x648;
  assign n4230 = x789 & n4229;
  assign n4231 = ~n4228 & ~n4230;
  assign n4232 = n4226 & n4231;
  assign n4233 = x665 & x1091;
  assign n4234 = n4232 & ~n4233;
  assign n4235 = ~n4208 & n4234;
  assign n4236 = ~x738 & n4235;
  assign n4237 = ~x761 & n4208;
  assign n4238 = ~n4236 & ~n4237;
  assign n4239 = n4238 ^ x140;
  assign n4240 = ~n4182 & n4239;
  assign n4241 = n4240 ^ x140;
  assign n4242 = x706 & n4235;
  assign n4243 = x749 & n4208;
  assign n4244 = ~n4242 & ~n4243;
  assign n4245 = n4244 ^ x141;
  assign n4246 = ~n4182 & n4245;
  assign n4247 = n4246 ^ x141;
  assign n4248 = x735 & n4235;
  assign n4249 = x743 & n4208;
  assign n4250 = ~n4248 & ~n4249;
  assign n4251 = n4250 ^ x142;
  assign n4252 = ~n4182 & ~n4251;
  assign n4253 = n4252 ^ x142;
  assign n4254 = x687 & n4235;
  assign n4255 = ~x774 & n4208;
  assign n4256 = ~n4254 & ~n4255;
  assign n4257 = n4256 ^ x143;
  assign n4258 = ~n4182 & n4257;
  assign n4259 = n4258 ^ x143;
  assign n4260 = x736 & n4235;
  assign n4261 = x758 & n4208;
  assign n4262 = ~n4260 & ~n4261;
  assign n4263 = n4262 ^ x144;
  assign n4264 = ~n4182 & ~n4263;
  assign n4265 = n4264 ^ x144;
  assign n4266 = ~x698 & n4235;
  assign n4267 = ~x767 & n4208;
  assign n4268 = ~n4266 & ~n4267;
  assign n4269 = n4268 ^ x145;
  assign n4270 = ~n4182 & n4269;
  assign n4271 = n4270 ^ x145;
  assign n4272 = x907 & ~x947;
  assign n4273 = x735 & n4272;
  assign n4274 = x743 & x947;
  assign n4275 = ~n4273 & ~n4274;
  assign n4276 = n4275 ^ x146;
  assign n4277 = ~n4182 & ~n4276;
  assign n4278 = n4277 ^ x146;
  assign n4279 = x726 & n4272;
  assign n4280 = ~x770 & x947;
  assign n4281 = ~n4279 & ~n4280;
  assign n4282 = n4281 ^ x147;
  assign n4283 = ~n4182 & n4282;
  assign n4284 = n4283 ^ x147;
  assign n4285 = x706 & n4272;
  assign n4286 = x749 & x947;
  assign n4287 = ~n4285 & ~n4286;
  assign n4288 = n4287 ^ x148;
  assign n4289 = ~n4182 & n4288;
  assign n4290 = n4289 ^ x148;
  assign n4291 = ~n2192 & ~n4175;
  assign n4292 = n2190 & n2493;
  assign n4293 = n2492 & ~n2814;
  assign n4294 = ~n4292 & ~n4293;
  assign n4295 = ~n4291 & n4294;
  assign n4296 = n2402 & ~n4295;
  assign n4297 = ~n4172 & ~n4296;
  assign n4298 = n2695 & ~n4297;
  assign n4299 = ~n4181 & ~n4298;
  assign n4300 = ~x725 & n4272;
  assign n4301 = ~x755 & x947;
  assign n4302 = ~n4300 & ~n4301;
  assign n4303 = ~n4299 & ~n4302;
  assign n4304 = ~x149 & n4182;
  assign n4305 = ~n4303 & ~n4304;
  assign n4306 = ~x701 & n4272;
  assign n4307 = ~x751 & x947;
  assign n4308 = ~n4306 & ~n4307;
  assign n4309 = ~n4299 & ~n4308;
  assign n4310 = ~x150 & n4182;
  assign n4311 = ~n4309 & ~n4310;
  assign n4312 = ~x723 & n4272;
  assign n4313 = ~x745 & x947;
  assign n4314 = ~n4312 & ~n4313;
  assign n4315 = n4314 ^ x151;
  assign n4316 = ~n4182 & n4315;
  assign n4317 = n4316 ^ x151;
  assign n4318 = x696 & n4272;
  assign n4319 = x759 & x947;
  assign n4320 = ~n4318 & ~n4319;
  assign n4321 = n4320 ^ x152;
  assign n4322 = ~n4182 & ~n4321;
  assign n4323 = n4322 ^ x152;
  assign n4324 = x700 & n4272;
  assign n4325 = x766 & x947;
  assign n4326 = ~n4324 & ~n4325;
  assign n4327 = n4326 ^ x153;
  assign n4328 = ~n4182 & n4327;
  assign n4329 = n4328 ^ x153;
  assign n4330 = ~x704 & n4272;
  assign n4331 = ~x742 & x947;
  assign n4332 = ~n4330 & ~n4331;
  assign n4333 = ~n4299 & ~n4332;
  assign n4334 = ~x154 & n4182;
  assign n4335 = ~n4333 & ~n4334;
  assign n4336 = ~x686 & n4272;
  assign n4337 = ~x757 & x947;
  assign n4338 = ~n4336 & ~n4337;
  assign n4339 = ~n4299 & ~n4338;
  assign n4340 = ~x155 & n4182;
  assign n4341 = ~n4339 & ~n4340;
  assign n4342 = ~x724 & n4272;
  assign n4343 = ~x741 & x947;
  assign n4344 = ~n4342 & ~n4343;
  assign n4345 = ~n4299 & ~n4344;
  assign n4346 = ~x156 & n4182;
  assign n4347 = ~n4345 & ~n4346;
  assign n4348 = ~x688 & n4272;
  assign n4349 = ~x760 & x947;
  assign n4350 = ~n4348 & ~n4349;
  assign n4351 = n4350 ^ x157;
  assign n4352 = ~n4182 & n4351;
  assign n4353 = n4352 ^ x157;
  assign n4354 = ~x702 & n4272;
  assign n4355 = ~x753 & x947;
  assign n4356 = ~n4354 & ~n4355;
  assign n4357 = ~n4299 & ~n4356;
  assign n4358 = ~x158 & n4182;
  assign n4359 = ~n4357 & ~n4358;
  assign n4360 = ~x709 & n4272;
  assign n4361 = ~x754 & x947;
  assign n4362 = ~n4360 & ~n4361;
  assign n4363 = n4362 ^ x159;
  assign n4364 = ~n4182 & n4363;
  assign n4365 = n4364 ^ x159;
  assign n4366 = ~x734 & n4272;
  assign n4367 = ~x756 & x947;
  assign n4368 = ~n4366 & ~n4367;
  assign n4369 = n4368 ^ x160;
  assign n4370 = ~n4182 & n4369;
  assign n4371 = n4370 ^ x160;
  assign n4372 = x736 & n4272;
  assign n4373 = x758 & x947;
  assign n4374 = ~n4372 & ~n4373;
  assign n4375 = n4374 ^ x161;
  assign n4376 = ~n4182 & ~n4375;
  assign n4377 = n4376 ^ x161;
  assign n4378 = ~x738 & n4272;
  assign n4379 = ~x761 & x947;
  assign n4380 = ~n4378 & ~n4379;
  assign n4381 = n4380 ^ x162;
  assign n4382 = ~n4182 & n4381;
  assign n4383 = n4382 ^ x162;
  assign n4384 = ~x737 & n4272;
  assign n4385 = ~x777 & x947;
  assign n4386 = ~n4384 & ~n4385;
  assign n4387 = n4386 ^ x163;
  assign n4388 = ~n4182 & n4387;
  assign n4389 = n4388 ^ x163;
  assign n4390 = x703 & n4272;
  assign n4391 = ~x752 & x947;
  assign n4392 = ~n4390 & ~n4391;
  assign n4393 = n4392 ^ x164;
  assign n4394 = ~n4182 & n4393;
  assign n4395 = n4394 ^ x164;
  assign n4396 = x687 & n4272;
  assign n4397 = ~x774 & x947;
  assign n4398 = ~n4396 & ~n4397;
  assign n4399 = ~n4299 & ~n4398;
  assign n4400 = ~x165 & n4182;
  assign n4401 = ~n4399 & ~n4400;
  assign n4402 = x727 & n4272;
  assign n4403 = x772 & x947;
  assign n4404 = ~n4402 & ~n4403;
  assign n4405 = n4404 ^ x166;
  assign n4406 = ~n4182 & ~n4405;
  assign n4407 = n4406 ^ x166;
  assign n4408 = x705 & n4272;
  assign n4409 = ~x768 & x947;
  assign n4410 = ~n4408 & ~n4409;
  assign n4411 = n4410 ^ x167;
  assign n4412 = ~n4182 & n4411;
  assign n4413 = n4412 ^ x167;
  assign n4414 = x699 & n4272;
  assign n4415 = x763 & x947;
  assign n4416 = ~n4414 & ~n4415;
  assign n4417 = n4416 ^ x168;
  assign n4418 = ~n4182 & n4417;
  assign n4419 = n4418 ^ x168;
  assign n4420 = x729 & n4272;
  assign n4421 = x746 & x947;
  assign n4422 = ~n4420 & ~n4421;
  assign n4423 = n4422 ^ x169;
  assign n4424 = ~n4182 & n4423;
  assign n4425 = n4424 ^ x169;
  assign n4426 = x730 & n4272;
  assign n4427 = x748 & x947;
  assign n4428 = ~n4426 & ~n4427;
  assign n4429 = n4428 ^ x170;
  assign n4430 = ~n4182 & n4429;
  assign n4431 = n4430 ^ x170;
  assign n4432 = x691 & n4272;
  assign n4433 = x764 & x947;
  assign n4434 = ~n4432 & ~n4433;
  assign n4435 = n4434 ^ x171;
  assign n4436 = ~n4182 & n4435;
  assign n4437 = n4436 ^ x171;
  assign n4438 = x690 & n4272;
  assign n4439 = x739 & x947;
  assign n4440 = ~n4438 & ~n4439;
  assign n4441 = n4440 ^ x172;
  assign n4442 = ~n4182 & n4441;
  assign n4443 = n4442 ^ x172;
  assign n4444 = ~x723 & n4235;
  assign n4445 = ~x745 & n4208;
  assign n4446 = ~n4444 & ~n4445;
  assign n4447 = n4446 ^ x173;
  assign n4448 = ~n4182 & n4447;
  assign n4449 = n4448 ^ x173;
  assign n4450 = x696 & n4235;
  assign n4451 = x759 & n4208;
  assign n4452 = ~n4450 & ~n4451;
  assign n4453 = n4452 ^ x174;
  assign n4454 = ~n4182 & ~n4453;
  assign n4455 = n4454 ^ x174;
  assign n4456 = x700 & n4235;
  assign n4457 = x766 & n4208;
  assign n4458 = ~n4456 & ~n4457;
  assign n4459 = n4458 ^ x175;
  assign n4460 = ~n4182 & n4459;
  assign n4461 = n4460 ^ x175;
  assign n4462 = ~x704 & n4235;
  assign n4463 = ~x742 & n4208;
  assign n4464 = ~n4462 & ~n4463;
  assign n4465 = n4464 ^ x176;
  assign n4466 = ~n4182 & n4465;
  assign n4467 = n4466 ^ x176;
  assign n4468 = ~x686 & n4235;
  assign n4469 = ~x757 & n4208;
  assign n4470 = ~n4468 & ~n4469;
  assign n4471 = n4470 ^ x177;
  assign n4472 = ~n4182 & n4471;
  assign n4473 = n4472 ^ x177;
  assign n4474 = ~x688 & n4235;
  assign n4475 = ~x760 & n4208;
  assign n4476 = ~n4474 & ~n4475;
  assign n4477 = n4476 ^ x178;
  assign n4478 = ~n4182 & n4477;
  assign n4479 = n4478 ^ x178;
  assign n4480 = ~x724 & n4235;
  assign n4481 = ~x741 & n4208;
  assign n4482 = ~n4480 & ~n4481;
  assign n4483 = n4482 ^ x179;
  assign n4484 = ~n4182 & n4483;
  assign n4485 = n4484 ^ x179;
  assign n4486 = ~x702 & n4235;
  assign n4487 = ~x753 & n4208;
  assign n4488 = ~n4486 & ~n4487;
  assign n4489 = n4488 ^ x180;
  assign n4490 = ~n4182 & n4489;
  assign n4491 = n4490 ^ x180;
  assign n4492 = ~x709 & n4235;
  assign n4493 = ~x754 & n4208;
  assign n4494 = ~n4492 & ~n4493;
  assign n4495 = n4494 ^ x181;
  assign n4496 = ~n4182 & n4495;
  assign n4497 = n4496 ^ x181;
  assign n4498 = ~x734 & n4235;
  assign n4499 = ~x756 & n4208;
  assign n4500 = ~n4498 & ~n4499;
  assign n4501 = n4500 ^ x182;
  assign n4502 = ~n4182 & n4501;
  assign n4503 = n4502 ^ x182;
  assign n4504 = ~x725 & n4235;
  assign n4505 = ~x755 & n4208;
  assign n4506 = ~n4504 & ~n4505;
  assign n4507 = n4506 ^ x183;
  assign n4508 = ~n4182 & n4507;
  assign n4509 = n4508 ^ x183;
  assign n4510 = ~x737 & n4235;
  assign n4511 = ~x777 & n4208;
  assign n4512 = ~n4510 & ~n4511;
  assign n4513 = n4512 ^ x184;
  assign n4514 = ~n4182 & n4513;
  assign n4515 = n4514 ^ x184;
  assign n4516 = ~x701 & n4235;
  assign n4517 = ~x751 & n4208;
  assign n4518 = ~n4516 & ~n4517;
  assign n4519 = n4518 ^ x185;
  assign n4520 = ~n4182 & n4519;
  assign n4521 = n4520 ^ x185;
  assign n4522 = x703 & n4235;
  assign n4523 = ~x752 & n4208;
  assign n4524 = ~n4522 & ~n4523;
  assign n4525 = n4524 ^ x186;
  assign n4526 = ~n4182 & n4525;
  assign n4527 = n4526 ^ x186;
  assign n4528 = x726 & n4235;
  assign n4529 = ~x770 & n4208;
  assign n4530 = ~n4528 & ~n4529;
  assign n4531 = n4530 ^ x187;
  assign n4532 = ~n4182 & n4531;
  assign n4533 = n4532 ^ x187;
  assign n4534 = x705 & n4235;
  assign n4535 = ~x768 & n4208;
  assign n4536 = ~n4534 & ~n4535;
  assign n4537 = n4536 ^ x188;
  assign n4538 = ~n4182 & n4537;
  assign n4539 = n4538 ^ x188;
  assign n4540 = x727 & n4235;
  assign n4541 = x772 & n4208;
  assign n4542 = ~n4540 & ~n4541;
  assign n4543 = n4542 ^ x189;
  assign n4544 = ~n4182 & ~n4543;
  assign n4545 = n4544 ^ x189;
  assign n4546 = x699 & n4235;
  assign n4547 = x763 & n4208;
  assign n4548 = ~n4546 & ~n4547;
  assign n4549 = n4548 ^ x190;
  assign n4550 = ~n4182 & n4549;
  assign n4551 = n4550 ^ x190;
  assign n4552 = x729 & n4235;
  assign n4553 = x746 & n4208;
  assign n4554 = ~n4552 & ~n4553;
  assign n4555 = n4554 ^ x191;
  assign n4556 = ~n4182 & n4555;
  assign n4557 = n4556 ^ x191;
  assign n4558 = x691 & n4235;
  assign n4559 = x764 & n4208;
  assign n4560 = ~n4558 & ~n4559;
  assign n4561 = n4560 ^ x192;
  assign n4562 = ~n4182 & n4561;
  assign n4563 = n4562 ^ x192;
  assign n4564 = x690 & n4235;
  assign n4565 = x739 & n4208;
  assign n4566 = ~n4564 & ~n4565;
  assign n4567 = n4566 ^ x193;
  assign n4568 = ~n4182 & n4567;
  assign n4569 = n4568 ^ x193;
  assign n4570 = x730 & n4235;
  assign n4571 = x748 & n4208;
  assign n4572 = ~n4570 & ~n4571;
  assign n4573 = n4572 ^ x194;
  assign n4574 = ~n4182 & n4573;
  assign n4575 = n4574 ^ x194;
  assign n4576 = ~x196 & n4145;
  assign n4577 = x195 & ~n4576;
  assign n4578 = n4144 & n4577;
  assign n4579 = ~x299 & n4080;
  assign n4580 = n4579 ^ x171;
  assign n4581 = n2476 & n4580;
  assign n4582 = ~n3367 & ~n4581;
  assign n4583 = ~n4578 & ~n4582;
  assign n4584 = n4145 ^ x196;
  assign n4585 = n4145 & n4584;
  assign n4586 = ~x195 & n4585;
  assign n4587 = n4586 ^ n4584;
  assign n4588 = n4144 & n4587;
  assign n4589 = ~x299 & n4098;
  assign n4590 = n4589 ^ x170;
  assign n4591 = n2476 & n4590;
  assign n4592 = ~n3367 & ~n4591;
  assign n4593 = ~n4588 & ~n4592;
  assign n4594 = ~x698 & n4272;
  assign n4595 = ~x767 & x947;
  assign n4596 = ~n4594 & ~n4595;
  assign n4597 = n4596 ^ x197;
  assign n4598 = ~n4182 & n4597;
  assign n4599 = n4598 ^ x197;
  assign n4600 = x634 & n4235;
  assign n4601 = x633 & n4208;
  assign n4602 = ~n4600 & ~n4601;
  assign n4603 = n4602 ^ x198;
  assign n4604 = n4180 & ~n4603;
  assign n4605 = n4604 ^ x198;
  assign n4606 = x637 & n4235;
  assign n4607 = x617 & n4208;
  assign n4608 = ~n4606 & ~n4607;
  assign n4609 = n4608 ^ x199;
  assign n4610 = n4180 & ~n4609;
  assign n4611 = n4610 ^ x199;
  assign n4612 = x643 & n4235;
  assign n4613 = x606 & n4208;
  assign n4614 = ~n4612 & ~n4613;
  assign n4615 = n4614 ^ x200;
  assign n4616 = n4180 & ~n4615;
  assign n4617 = n4616 ^ x200;
  assign n4618 = ~n1241 & n3210;
  assign n4619 = ~x332 & ~n1548;
  assign n4620 = ~n4618 & n4619;
  assign n4621 = n1257 & ~n1656;
  assign n4622 = n4621 ^ x198;
  assign n4623 = x96 & n4622;
  assign n4624 = ~x32 & x70;
  assign n4625 = ~n4623 & n4624;
  assign n4626 = ~x70 & n2748;
  assign n4627 = ~n4622 & n4626;
  assign n4628 = ~n4625 & ~n4627;
  assign n4629 = x233 & ~n4628;
  assign n4630 = x237 & n4629;
  assign n4631 = n4620 & ~n4630;
  assign n4632 = n1656 & n2161;
  assign n4633 = ~n2354 & ~n4632;
  assign n4634 = ~n2161 & n2172;
  assign n4635 = ~x587 & ~n4634;
  assign n4636 = n1656 & n4635;
  assign n4637 = ~n4633 & ~n4636;
  assign n4638 = ~x332 & ~n4637;
  assign n4639 = ~n4631 & ~n4638;
  assign n4640 = ~x201 & ~n4639;
  assign n4641 = x237 & n4623;
  assign n4642 = x233 & n4637;
  assign n4643 = n4641 & n4642;
  assign n4644 = ~n4640 & ~n4643;
  assign n4645 = ~x233 & ~n4628;
  assign n4646 = x237 & n4645;
  assign n4647 = n4620 & ~n4646;
  assign n4648 = ~n4638 & ~n4647;
  assign n4649 = ~x202 & ~n4648;
  assign n4650 = ~x233 & n4637;
  assign n4651 = n4641 & n4650;
  assign n4652 = ~n4649 & ~n4651;
  assign n4653 = ~x237 & n4645;
  assign n4654 = n4620 & ~n4653;
  assign n4655 = ~n4638 & ~n4654;
  assign n4656 = ~x203 & ~n4655;
  assign n4657 = ~x237 & n4623;
  assign n4658 = n4650 & n4657;
  assign n4659 = ~n4656 & ~n4658;
  assign n4660 = ~x907 & ~n1656;
  assign n4661 = ~x602 & n4632;
  assign n4662 = n4661 ^ n2161;
  assign n4663 = ~n4660 & n4662;
  assign n4664 = ~n2346 & ~n4663;
  assign n4665 = ~x332 & n4664;
  assign n4666 = ~n4631 & ~n4665;
  assign n4667 = ~x204 & ~n4666;
  assign n4668 = n4641 & ~n4664;
  assign n4669 = x233 & n4668;
  assign n4670 = ~n4667 & ~n4669;
  assign n4671 = ~n4647 & ~n4665;
  assign n4672 = ~x205 & ~n4671;
  assign n4673 = ~x233 & n4668;
  assign n4674 = ~n4672 & ~n4673;
  assign n4675 = ~x237 & n4629;
  assign n4676 = n4620 & ~n4675;
  assign n4677 = ~n4665 & ~n4676;
  assign n4678 = ~x206 & ~n4677;
  assign n4679 = n4657 & ~n4664;
  assign n4680 = x233 & n4679;
  assign n4681 = ~n4678 & ~n4680;
  assign n4682 = x710 & n4235;
  assign n4683 = x623 & n4208;
  assign n4684 = ~n4682 & ~n4683;
  assign n4685 = n4684 ^ x207;
  assign n4686 = n4180 & n4685;
  assign n4687 = n4686 ^ x207;
  assign n4688 = x638 & n4235;
  assign n4689 = x607 & n4208;
  assign n4690 = ~n4688 & ~n4689;
  assign n4691 = n4690 ^ x208;
  assign n4692 = n4180 & n4691;
  assign n4693 = n4692 ^ x208;
  assign n4694 = x639 & n4235;
  assign n4695 = x622 & n4208;
  assign n4696 = ~n4694 & ~n4695;
  assign n4697 = n4696 ^ x209;
  assign n4698 = n4180 & n4697;
  assign n4699 = n4698 ^ x209;
  assign n4700 = x634 & n4272;
  assign n4701 = x633 & x947;
  assign n4702 = ~n4700 & ~n4701;
  assign n4703 = n4702 ^ x210;
  assign n4704 = n4180 & ~n4703;
  assign n4705 = n4704 ^ x210;
  assign n4706 = x643 & n4272;
  assign n4707 = x606 & x947;
  assign n4708 = ~n4706 & ~n4707;
  assign n4709 = n4708 ^ x211;
  assign n4710 = n4180 & ~n4709;
  assign n4711 = n4710 ^ x211;
  assign n4712 = ~x212 & ~n4180;
  assign n4713 = x638 & n4272;
  assign n4714 = x607 & x947;
  assign n4715 = ~n4713 & ~n4714;
  assign n4716 = n4298 & ~n4715;
  assign n4717 = ~n4712 & ~n4716;
  assign n4718 = ~x213 & ~n4180;
  assign n4719 = x639 & n4272;
  assign n4720 = x622 & x947;
  assign n4721 = ~n4719 & ~n4720;
  assign n4722 = n4298 & ~n4721;
  assign n4723 = ~n4718 & ~n4722;
  assign n4724 = x710 & n4272;
  assign n4725 = x623 & x947;
  assign n4726 = ~n4724 & ~n4725;
  assign n4727 = n4726 ^ x214;
  assign n4728 = n4180 & n4727;
  assign n4729 = n4728 ^ x214;
  assign n4730 = x681 & n4272;
  assign n4731 = x642 & x947;
  assign n4732 = ~n4730 & ~n4731;
  assign n4733 = n4732 ^ x215;
  assign n4734 = n4180 & ~n4733;
  assign n4735 = n4734 ^ x215;
  assign n4736 = x662 & n4272;
  assign n4737 = x614 & x947;
  assign n4738 = ~n4736 & ~n4737;
  assign n4739 = n4738 ^ x216;
  assign n4740 = n4180 & ~n4739;
  assign n4741 = n4740 ^ x216;
  assign n4742 = ~x695 & n4235;
  assign n4743 = x612 & n4208;
  assign n4744 = ~n4742 & ~n4743;
  assign n4745 = n4744 ^ x217;
  assign n4746 = n4180 & n4745;
  assign n4747 = n4746 ^ x217;
  assign n4748 = ~n4654 & ~n4665;
  assign n4749 = ~x218 & ~n4748;
  assign n4750 = ~x233 & n4679;
  assign n4751 = ~n4749 & ~n4750;
  assign n4752 = x219 & ~n4180;
  assign n4753 = x637 & n4272;
  assign n4754 = x617 & x947;
  assign n4755 = ~n4753 & ~n4754;
  assign n4756 = n4298 & ~n4755;
  assign n4757 = ~n4752 & ~n4756;
  assign n4758 = ~n4638 & ~n4676;
  assign n4759 = ~x220 & ~n4758;
  assign n4760 = n4642 & n4657;
  assign n4761 = ~n4759 & ~n4760;
  assign n4762 = x661 & n4272;
  assign n4763 = x616 & x947;
  assign n4764 = ~n4762 & ~n4763;
  assign n4765 = n4764 ^ x221;
  assign n4766 = n4180 & ~n4765;
  assign n4767 = n4766 ^ x221;
  assign n4768 = x661 & n4235;
  assign n4769 = x616 & n4208;
  assign n4770 = ~n4768 & ~n4769;
  assign n4771 = n4770 ^ x222;
  assign n4772 = n4180 & ~n4771;
  assign n4773 = n4772 ^ x222;
  assign n4774 = x681 & n4235;
  assign n4775 = x642 & n4208;
  assign n4776 = ~n4774 & ~n4775;
  assign n4777 = n4776 ^ x223;
  assign n4778 = n4180 & ~n4777;
  assign n4779 = n4778 ^ x223;
  assign n4780 = x662 & n4235;
  assign n4781 = x614 & n4208;
  assign n4782 = ~n4780 & ~n4781;
  assign n4783 = n4782 ^ x224;
  assign n4784 = n4180 & ~n4783;
  assign n4785 = n4784 ^ x224;
  assign n4786 = n1471 & n1519;
  assign n4787 = x70 & x332;
  assign n4788 = ~n1262 & ~n4787;
  assign n4789 = n1662 & ~n4788;
  assign n4790 = n1447 & n3764;
  assign n4791 = ~x55 & ~x137;
  assign n4792 = ~n4790 & n4791;
  assign n4793 = ~n1575 & ~n4792;
  assign n4794 = ~n4789 & ~n4793;
  assign n4795 = ~n4786 & n4794;
  assign n4796 = n1662 & n2156;
  assign n4797 = n1559 & ~n1570;
  assign n4798 = x479 & n3590;
  assign n4799 = n1574 & ~n4798;
  assign n4800 = ~n4797 & n4799;
  assign n4801 = ~n4796 & n4800;
  assign n4802 = n4801 ^ x231;
  assign n4803 = ~x228 & ~n4802;
  assign n4804 = n4803 ^ x231;
  assign n4805 = x1093 & n3046;
  assign n4806 = ~x58 & n1454;
  assign n4807 = n1393 & n4806;
  assign n4808 = ~x72 & ~n4807;
  assign n4809 = ~n3200 & n4808;
  assign n4810 = ~n4805 & n4809;
  assign n4811 = n1662 & ~n4810;
  assign n4812 = ~n3363 & ~n4811;
  assign n4813 = x36 & n1428;
  assign n4814 = ~n4812 & ~n4813;
  assign n4815 = ~n1421 & ~n2220;
  assign n4816 = n1518 & n1634;
  assign n4817 = ~n4815 & n4816;
  assign n4818 = ~n1420 & n4817;
  assign n4819 = ~x228 & ~n4818;
  assign n4820 = ~x39 & ~n4819;
  assign n4821 = x1091 & n3582;
  assign n4822 = ~n4820 & ~n4821;
  assign n4823 = ~x47 & ~n2221;
  assign n4824 = n1233 & n4823;
  assign n4825 = ~n2813 & n4824;
  assign n4826 = ~n4179 & ~n4825;
  assign n4827 = ~x64 & n2788;
  assign n4828 = x102 ^ x65;
  assign n4829 = n4827 & n4828;
  assign n4830 = n1336 & n4829;
  assign n4831 = ~n3011 & ~n4830;
  assign n4832 = ~n2250 & n4831;
  assign n4833 = ~n1575 & ~n3306;
  assign n4834 = ~n4832 & ~n4833;
  assign n4835 = x1155 & n3242;
  assign n4836 = x1156 & n3150;
  assign n4837 = ~n4835 & ~n4836;
  assign n4838 = x199 & ~x200;
  assign n4839 = x1154 & n4838;
  assign n4840 = n4837 & ~n4839;
  assign n4841 = ~x207 & x208;
  assign n4842 = ~n4840 & n4841;
  assign n4843 = x1155 & n4838;
  assign n4844 = x1156 & n3242;
  assign n4845 = ~n4843 & ~n4844;
  assign n4846 = x1157 & n3150;
  assign n4847 = n4845 & ~n4846;
  assign n4848 = x207 & ~x208;
  assign n4849 = ~n4847 & n4848;
  assign n4850 = ~n4842 & ~n4849;
  assign n4851 = ~x209 & n1656;
  assign n4852 = n4850 & n4851;
  assign n4853 = x1154 & n3242;
  assign n4854 = x1153 & n4838;
  assign n4855 = ~n4853 & ~n4854;
  assign n4856 = x1155 & n3150;
  assign n4857 = n4855 & ~n4856;
  assign n4858 = n3153 & ~n4857;
  assign n4859 = n4852 & ~n4858;
  assign n4860 = x208 ^ x207;
  assign n4861 = x1144 ^ x1143;
  assign n4862 = ~x200 & n4861;
  assign n4863 = n4862 ^ x1143;
  assign n4864 = n4860 & n4863;
  assign n4865 = ~x200 & n3153;
  assign n4866 = x1143 & n4865;
  assign n4867 = ~n4864 & ~n4866;
  assign n4868 = x1142 & ~n3150;
  assign n4869 = ~n3154 & n4868;
  assign n4870 = n4867 & ~n4869;
  assign n4871 = ~x207 & ~x208;
  assign n4872 = ~x200 & ~n4871;
  assign n4873 = x1142 & n4872;
  assign n4874 = x199 & ~n4873;
  assign n4875 = ~n4870 & ~n4874;
  assign n4876 = x209 & n1656;
  assign n4877 = ~n4875 & n4876;
  assign n4878 = x230 & ~n4877;
  assign n4879 = ~n4859 & n4878;
  assign n4880 = x1156 ^ x1154;
  assign n4881 = ~x219 & n4880;
  assign n4882 = n4881 ^ x1154;
  assign n4883 = ~x214 & ~n4882;
  assign n4884 = ~x211 & ~n4883;
  assign n4885 = x1155 ^ x1153;
  assign n4886 = ~x219 & n4885;
  assign n4887 = n4886 ^ x1153;
  assign n4888 = x214 & ~n4887;
  assign n4889 = n4884 & ~n4888;
  assign n4890 = ~x214 & ~x1155;
  assign n4891 = n3239 & ~n4890;
  assign n4892 = x214 & ~x1154;
  assign n4893 = n4891 & ~n4892;
  assign n4894 = ~n4889 & ~n4893;
  assign n4895 = x212 & ~n4894;
  assign n4896 = ~x213 & ~n1656;
  assign n4897 = x1157 ^ x1155;
  assign n4898 = ~x219 & n4897;
  assign n4899 = n4898 ^ x1155;
  assign n4900 = ~x211 & ~n4899;
  assign n4901 = ~x219 & x1156;
  assign n4902 = x211 & ~n4901;
  assign n4903 = ~x212 & x214;
  assign n4904 = ~n4902 & n4903;
  assign n4905 = ~n4900 & n4904;
  assign n4906 = n4896 & ~n4905;
  assign n4907 = ~n4895 & n4906;
  assign n4908 = ~x212 & ~x214;
  assign n4909 = n3238 & ~n4908;
  assign n4910 = x1143 & n4909;
  assign n4911 = n3156 & n3239;
  assign n4912 = n3236 & ~n4908;
  assign n4913 = ~n4911 & ~n4912;
  assign n4914 = x1142 & ~n4913;
  assign n4915 = x214 ^ x212;
  assign n4916 = n3167 & n4915;
  assign n4917 = x1144 & n4916;
  assign n4918 = ~n4914 & ~n4917;
  assign n4919 = ~n4910 & n4918;
  assign n4920 = x213 & ~n1656;
  assign n4921 = n4919 & n4920;
  assign n4922 = ~n4907 & ~n4921;
  assign n4923 = n4879 & n4922;
  assign n4924 = ~x230 & ~x233;
  assign n4925 = ~n4923 & ~n4924;
  assign n4926 = n4908 ^ n4871;
  assign n4927 = ~n1656 & n4926;
  assign n4928 = n4927 ^ n4871;
  assign n4929 = n3247 & ~n4928;
  assign n4930 = ~n3161 & n4929;
  assign n4931 = x1152 & n4930;
  assign n4932 = ~x1153 & n3247;
  assign n4933 = n3161 & ~n4928;
  assign n4934 = ~n4932 & n4933;
  assign n4935 = ~x1154 & ~n3247;
  assign n4936 = n4934 & ~n4935;
  assign n4937 = ~n4931 & ~n4936;
  assign n4938 = ~n4876 & ~n4920;
  assign n4939 = n4937 & n4938;
  assign n4940 = x1154 & n4930;
  assign n4941 = x1155 & n4909;
  assign n4942 = x1156 & n4916;
  assign n4943 = n4920 & ~n4942;
  assign n4944 = ~n4941 & n4943;
  assign n4945 = ~n4837 & n4860;
  assign n4946 = n3153 & n4856;
  assign n4947 = ~n4945 & ~n4946;
  assign n4948 = n4876 & n4947;
  assign n4949 = ~n4944 & ~n4948;
  assign n4950 = ~n4940 & ~n4949;
  assign n4951 = x230 & ~n4950;
  assign n4952 = ~n4939 & n4951;
  assign n4953 = ~x230 & x234;
  assign n4954 = ~n4952 & ~n4953;
  assign n4955 = n4857 ^ n4847;
  assign n4956 = ~x209 & n4955;
  assign n4957 = n4956 ^ n4847;
  assign n4958 = n4860 & ~n4957;
  assign n4959 = x1153 & n3242;
  assign n4960 = x1154 & n3150;
  assign n4961 = ~n4959 & ~n4960;
  assign n4962 = n4851 & n4961;
  assign n4963 = x209 & n4837;
  assign n4964 = n3153 & ~n4963;
  assign n4965 = n1656 & ~n4964;
  assign n4966 = ~n4962 & ~n4965;
  assign n4967 = ~n4958 & ~n4966;
  assign n4968 = x213 & n4880;
  assign n4969 = n4968 ^ x1154;
  assign n4970 = n4909 & n4969;
  assign n4971 = ~x213 & ~n4887;
  assign n4972 = ~x211 & n4915;
  assign n4973 = ~n4971 & n4972;
  assign n4974 = x213 & ~n4899;
  assign n4975 = n4973 & ~n4974;
  assign n4976 = x213 & n4885;
  assign n4977 = n4976 ^ x1153;
  assign n4978 = n4911 & n4977;
  assign n4979 = ~n1656 & ~n4978;
  assign n4980 = ~n4975 & n4979;
  assign n4981 = ~n4970 & n4980;
  assign n4982 = x230 & ~n4981;
  assign n4983 = ~n4967 & n4982;
  assign n4984 = ~x230 & x235;
  assign n4985 = ~n4983 & ~n4984;
  assign n4986 = n4899 ^ n4882;
  assign n4987 = ~x214 & n4986;
  assign n4988 = n4987 ^ n4882;
  assign n4989 = ~x211 & n4988;
  assign n4990 = x214 & ~x1155;
  assign n4991 = n3239 & ~n4990;
  assign n4992 = ~x214 & ~x1156;
  assign n4993 = n4991 & ~n4992;
  assign n4994 = ~n4989 & ~n4993;
  assign n4995 = x212 & ~n4994;
  assign n4996 = x1156 & n3236;
  assign n4997 = x1157 & n3239;
  assign n4998 = ~n4996 & ~n4997;
  assign n4999 = x1158 & n3167;
  assign n5000 = n4998 & ~n4999;
  assign n5001 = n4903 & ~n5000;
  assign n5002 = ~n4995 & ~n5001;
  assign n5003 = n4896 & ~n5002;
  assign n5004 = n4841 & ~n4847;
  assign n5005 = x1157 & n3242;
  assign n5006 = x1156 & n4838;
  assign n5007 = ~n5005 & ~n5006;
  assign n5008 = x1158 & n3150;
  assign n5009 = n5007 & ~n5008;
  assign n5010 = n4848 & ~n5009;
  assign n5011 = ~n5004 & ~n5010;
  assign n5012 = n3153 & ~n4840;
  assign n5013 = n5011 & ~n5012;
  assign n5014 = n4851 & ~n5013;
  assign n5015 = x1143 & ~n4913;
  assign n5016 = ~x219 & n4915;
  assign n5017 = x1145 ^ x1144;
  assign n5018 = ~x211 & n5017;
  assign n5019 = n5018 ^ x1144;
  assign n5020 = n5016 & n5019;
  assign n5021 = n3156 & n3167;
  assign n5022 = x1144 & n5021;
  assign n5023 = ~n5020 & ~n5022;
  assign n5024 = ~n5015 & n5023;
  assign n5025 = n4920 & ~n5024;
  assign n5026 = x230 & ~n5025;
  assign n5027 = ~n5014 & n5026;
  assign n5028 = ~n5003 & n5027;
  assign n5029 = n4860 ^ n3153;
  assign n5030 = x200 & n5029;
  assign n5031 = n5030 ^ n3153;
  assign n5032 = x1144 & n5031;
  assign n5033 = x200 & x1143;
  assign n5034 = n3153 & n5033;
  assign n5035 = ~n5032 & ~n5034;
  assign n5036 = ~x199 & ~n5035;
  assign n5037 = x1145 & n3154;
  assign n5038 = x199 & x1143;
  assign n5039 = ~n5037 & ~n5038;
  assign n5040 = n4872 & ~n5039;
  assign n5041 = ~n5036 & ~n5040;
  assign n5042 = n4876 & ~n5041;
  assign n5043 = n5028 & ~n5042;
  assign n5044 = ~x230 & x237;
  assign n5045 = ~n5043 & ~n5044;
  assign n5046 = x1151 & n4930;
  assign n5047 = ~x1152 & n3247;
  assign n5048 = n4933 & ~n5047;
  assign n5049 = ~x1153 & ~n3247;
  assign n5050 = n5048 & ~n5049;
  assign n5051 = ~n5046 & ~n5050;
  assign n5052 = n4938 & n5051;
  assign n5053 = n3153 & ~n4854;
  assign n5054 = ~n4871 & ~n5053;
  assign n5055 = ~n4857 & n5054;
  assign n5056 = n4876 & ~n5055;
  assign n5057 = n3153 & ~n4961;
  assign n5058 = n5056 & ~n5057;
  assign n5059 = x1153 & ~n4913;
  assign n5060 = x1154 & n5021;
  assign n5061 = x1155 ^ x1154;
  assign n5062 = ~x211 & n5061;
  assign n5063 = n5062 ^ x1154;
  assign n5064 = n5016 & n5063;
  assign n5065 = ~n5060 & ~n5064;
  assign n5066 = ~n5059 & n5065;
  assign n5067 = n4920 & n5066;
  assign n5068 = x230 & ~n5067;
  assign n5069 = ~n5058 & n5068;
  assign n5070 = ~n5052 & n5069;
  assign n5071 = ~x230 & x238;
  assign n5072 = ~n5070 & ~n5071;
  assign n5073 = ~x213 & n4994;
  assign n5074 = x213 & n5000;
  assign n5075 = ~n1656 & n4903;
  assign n5076 = ~n5074 & n5075;
  assign n5077 = ~n5073 & n5076;
  assign n5078 = n1656 & n4848;
  assign n5079 = n5009 ^ n4840;
  assign n5080 = x209 & n5079;
  assign n5081 = n5080 ^ n4840;
  assign n5082 = n5078 & ~n5081;
  assign n5083 = x230 & ~n5082;
  assign n5084 = ~n5077 & n5083;
  assign n5085 = ~x230 & ~x239;
  assign n5086 = ~n5084 & ~n5085;
  assign n5093 = x1145 & n4930;
  assign n5094 = ~x1147 & ~n3247;
  assign n5095 = n4933 & ~n5094;
  assign n5096 = ~x1146 & n3247;
  assign n5097 = n5095 & ~n5096;
  assign n5098 = ~n5093 & ~n5097;
  assign n5087 = x1147 & n4930;
  assign n5088 = ~x1149 & ~n3247;
  assign n5089 = n4933 & ~n5088;
  assign n5090 = ~x1148 & n3247;
  assign n5091 = n5089 & ~n5090;
  assign n5092 = ~n5087 & ~n5091;
  assign n5099 = n5098 ^ n5092;
  assign n5100 = ~n4938 & n5099;
  assign n5101 = n5100 ^ n5098;
  assign n5102 = n5101 ^ x240;
  assign n5103 = x230 & ~n5102;
  assign n5104 = n5103 ^ x240;
  assign n5105 = x1149 & n4930;
  assign n5106 = ~x1151 & ~n3247;
  assign n5107 = n4933 & ~n5106;
  assign n5108 = ~x1150 & n3247;
  assign n5109 = n5107 & ~n5108;
  assign n5110 = ~n5105 & ~n5109;
  assign n5111 = n5110 ^ n5051;
  assign n5112 = n4938 & n5111;
  assign n5113 = n5112 ^ n5051;
  assign n5114 = n5113 ^ x241;
  assign n5115 = x230 & ~n5114;
  assign n5116 = n5115 ^ x241;
  assign n5117 = x1144 & n4930;
  assign n5118 = ~x1145 & n3247;
  assign n5119 = n4933 & ~n5118;
  assign n5120 = ~x1146 & ~n3247;
  assign n5121 = n5119 & ~n5120;
  assign n5122 = ~n5117 & ~n5121;
  assign n5123 = ~n4938 & n5122;
  assign n5124 = n4896 & n4919;
  assign n5125 = n4851 & ~n4875;
  assign n5126 = x230 & ~n5125;
  assign n5127 = ~n5124 & n5126;
  assign n5128 = ~n5123 & n5127;
  assign n5129 = ~x230 & x242;
  assign n5130 = ~n5128 & ~n5129;
  assign n5131 = ~x230 & ~x1091;
  assign n5144 = x199 & ~x299;
  assign n5145 = n1518 & n5144;
  assign n5146 = x81 & ~n5145;
  assign n5147 = ~n3160 & n5146;
  assign n5148 = ~x83 & ~x85;
  assign n5149 = ~n5147 & n5148;
  assign n5150 = x314 & ~n5149;
  assign n5151 = x802 & n5150;
  assign n5152 = x276 & n5151;
  assign n5153 = x271 & n5152;
  assign n5154 = x273 & n5153;
  assign n5155 = x283 & n5154;
  assign n5156 = x272 & n5155;
  assign n5157 = x275 & n5156;
  assign n5158 = x268 & n5157;
  assign n5159 = x253 & n5158;
  assign n5160 = x254 & n5159;
  assign n5161 = x267 & n5160;
  assign n5162 = ~x263 & n5161;
  assign n5163 = n5162 ^ x243;
  assign n5132 = n4838 ^ n3236;
  assign n5133 = n1656 & n5132;
  assign n5134 = n5133 ^ n3236;
  assign n5135 = x1157 & n5134;
  assign n5136 = ~n1656 & ~n3167;
  assign n5137 = ~n3152 & ~n5136;
  assign n5138 = x1155 & n5137;
  assign n5139 = ~n5135 & ~n5138;
  assign n5140 = ~n1656 & ~n3239;
  assign n5141 = ~n3244 & ~n5140;
  assign n5142 = x1156 & n5141;
  assign n5143 = n5139 & ~n5142;
  assign n5164 = n5163 ^ n5143;
  assign n5165 = ~n5131 & n5164;
  assign n5166 = n5165 ^ n5163;
  assign n5167 = ~n4938 & n5098;
  assign n5168 = n4851 & n5041;
  assign n5169 = n4896 & n5024;
  assign n5170 = x230 & ~n5169;
  assign n5171 = ~n5168 & n5170;
  assign n5172 = ~n5167 & n5171;
  assign n5173 = ~x230 & x244;
  assign n5174 = ~n5172 & ~n5173;
  assign n5175 = x1146 & n4930;
  assign n5176 = ~x1148 & ~n3247;
  assign n5177 = n4933 & ~n5176;
  assign n5178 = ~x1147 & n3247;
  assign n5179 = n5177 & ~n5178;
  assign n5180 = ~n5175 & ~n5179;
  assign n5181 = n5180 ^ n5122;
  assign n5182 = ~n4938 & n5181;
  assign n5183 = n5182 ^ n5122;
  assign n5184 = n5183 ^ x245;
  assign n5185 = x230 & ~n5184;
  assign n5186 = n5185 ^ x245;
  assign n5187 = x1148 & n4930;
  assign n5188 = ~x1150 & ~n3247;
  assign n5189 = n4933 & ~n5188;
  assign n5190 = ~x1149 & n3247;
  assign n5191 = n5189 & ~n5190;
  assign n5192 = ~n5187 & ~n5191;
  assign n5193 = n5192 ^ n5180;
  assign n5194 = ~n4938 & n5193;
  assign n5195 = n5194 ^ n5180;
  assign n5196 = n5195 ^ x246;
  assign n5197 = x230 & ~n5196;
  assign n5198 = n5197 ^ x246;
  assign n5199 = n5110 ^ n5092;
  assign n5200 = ~n4938 & n5199;
  assign n5201 = n5200 ^ n5092;
  assign n5202 = n5201 ^ x247;
  assign n5203 = x230 & ~n5202;
  assign n5204 = n5203 ^ x247;
  assign n5205 = x1150 & n4930;
  assign n5206 = ~x1152 & ~n3247;
  assign n5207 = n4933 & ~n5206;
  assign n5208 = ~x1151 & n3247;
  assign n5209 = n5207 & ~n5208;
  assign n5210 = ~n5205 & ~n5209;
  assign n5211 = n5210 ^ n5192;
  assign n5212 = ~n4938 & n5211;
  assign n5213 = n5212 ^ n5192;
  assign n5214 = n5213 ^ x248;
  assign n5215 = x230 & ~n5214;
  assign n5216 = n5215 ^ x248;
  assign n5217 = n5210 ^ n4937;
  assign n5218 = n4938 & n5217;
  assign n5219 = n5218 ^ n4937;
  assign n5220 = n5219 ^ x249;
  assign n5221 = x230 & ~n5220;
  assign n5222 = n5221 ^ x249;
  assign n5223 = ~n3221 & ~n3764;
  assign n5224 = ~x250 & ~n5223;
  assign n5225 = x897 & n3150;
  assign n5226 = ~x476 & n3242;
  assign n5227 = ~n5225 & ~n5226;
  assign n5228 = x1053 ^ x1039;
  assign n5229 = ~x200 & n5228;
  assign n5230 = n5229 ^ x1039;
  assign n5231 = n5230 ^ x251;
  assign n5232 = ~n5227 & n5231;
  assign n5233 = n5232 ^ x251;
  assign n5234 = n2190 & ~n2201;
  assign n5235 = n2402 & n5234;
  assign n5236 = x1093 & ~n2699;
  assign n5237 = x252 & x1092;
  assign n5238 = ~n5236 & n5237;
  assign n5239 = ~n5235 & ~n5238;
  assign n5245 = n5158 ^ x253;
  assign n5240 = x1153 & n5134;
  assign n5241 = x1151 & n5137;
  assign n5242 = ~n5240 & ~n5241;
  assign n5243 = x1152 & n5141;
  assign n5244 = n5242 & ~n5243;
  assign n5246 = n5245 ^ n5244;
  assign n5247 = ~n5131 & ~n5246;
  assign n5248 = n5247 ^ n5245;
  assign n5254 = n5159 ^ x254;
  assign n5249 = x1153 & n5141;
  assign n5250 = x1152 & n5137;
  assign n5251 = ~n5249 & ~n5250;
  assign n5252 = x1154 & n5134;
  assign n5253 = n5251 & ~n5252;
  assign n5255 = n5254 ^ n5253;
  assign n5256 = ~n5131 & ~n5255;
  assign n5257 = n5256 ^ n5254;
  assign n5258 = x1049 ^ x1036;
  assign n5259 = ~x200 & n5258;
  assign n5260 = n5259 ^ x1036;
  assign n5261 = n5260 ^ x255;
  assign n5262 = ~n5227 & n5261;
  assign n5263 = n5262 ^ x255;
  assign n5264 = x1070 ^ x1048;
  assign n5265 = x200 & n5264;
  assign n5266 = n5265 ^ x1048;
  assign n5267 = n5266 ^ x256;
  assign n5268 = ~n5227 & n5267;
  assign n5269 = n5268 ^ x256;
  assign n5270 = x1084 ^ x1065;
  assign n5271 = ~x200 & n5270;
  assign n5272 = n5271 ^ x1065;
  assign n5273 = n5272 ^ x257;
  assign n5274 = ~n5227 & n5273;
  assign n5275 = n5274 ^ x257;
  assign n5276 = x1072 ^ x1062;
  assign n5277 = ~x200 & n5276;
  assign n5278 = n5277 ^ x1062;
  assign n5279 = n5278 ^ x258;
  assign n5280 = ~n5227 & n5279;
  assign n5281 = n5280 ^ x258;
  assign n5282 = x1069 ^ x1059;
  assign n5283 = x200 & n5282;
  assign n5284 = n5283 ^ x1059;
  assign n5285 = n5284 ^ x259;
  assign n5286 = ~n5227 & n5285;
  assign n5287 = n5286 ^ x259;
  assign n5288 = x1067 ^ x1044;
  assign n5289 = x200 & n5288;
  assign n5290 = n5289 ^ x1044;
  assign n5291 = n5290 ^ x260;
  assign n5292 = ~n5227 & n5291;
  assign n5293 = n5292 ^ x260;
  assign n5294 = x1040 ^ x1037;
  assign n5295 = x200 & n5294;
  assign n5296 = n5295 ^ x1037;
  assign n5297 = n5296 ^ x261;
  assign n5298 = ~n5227 & n5297;
  assign n5299 = n5298 ^ x261;
  assign n5300 = x1093 ^ x123;
  assign n5301 = ~x228 & ~n5300;
  assign n5302 = n5301 ^ x123;
  assign n5303 = n4933 & ~n5302;
  assign n5304 = x1142 & n5303;
  assign n5305 = ~x262 & n5302;
  assign n5306 = ~n5304 & ~n5305;
  assign n5312 = n5161 ^ x263;
  assign n5307 = x1156 & n5134;
  assign n5308 = x1154 & n5137;
  assign n5309 = ~n5307 & ~n5308;
  assign n5310 = x1155 & n5141;
  assign n5311 = n5309 & ~n5310;
  assign n5313 = n5312 ^ n5311;
  assign n5314 = ~n5131 & n5313;
  assign n5315 = n5314 ^ n5312;
  assign n5319 = x1141 & n5137;
  assign n5320 = x1143 & n5134;
  assign n5321 = ~n5319 & ~n5320;
  assign n5322 = x1142 & n5141;
  assign n5323 = n5321 & ~n5322;
  assign n5316 = x796 ^ x264;
  assign n5317 = n5150 & ~n5316;
  assign n5318 = n5317 ^ x264;
  assign n5324 = n5323 ^ n5318;
  assign n5325 = ~n5131 & n5324;
  assign n5326 = n5325 ^ n5318;
  assign n5330 = x1142 & n5137;
  assign n5331 = x1144 & n5134;
  assign n5332 = ~n5330 & ~n5331;
  assign n5333 = x1143 & n5141;
  assign n5334 = n5332 & ~n5333;
  assign n5327 = x819 ^ x265;
  assign n5328 = n5150 & ~n5327;
  assign n5329 = n5328 ^ x265;
  assign n5335 = n5334 ^ n5329;
  assign n5336 = ~n5131 & n5335;
  assign n5337 = n5336 ^ n5329;
  assign n5341 = x1134 & n5137;
  assign n5342 = x1136 & n5134;
  assign n5343 = ~n5341 & ~n5342;
  assign n5344 = x1135 & n5141;
  assign n5345 = n5343 & ~n5344;
  assign n5338 = x948 ^ x266;
  assign n5339 = n5150 & n5338;
  assign n5340 = n5339 ^ x266;
  assign n5346 = n5345 ^ n5340;
  assign n5347 = ~n5131 & ~n5346;
  assign n5348 = n5347 ^ n5340;
  assign n5354 = n5160 ^ x267;
  assign n5349 = x1154 & n5141;
  assign n5350 = x1153 & n5137;
  assign n5351 = ~n5349 & ~n5350;
  assign n5352 = x1155 & n5134;
  assign n5353 = n5351 & ~n5352;
  assign n5355 = n5354 ^ n5353;
  assign n5356 = ~n5131 & ~n5355;
  assign n5357 = n5356 ^ n5354;
  assign n5363 = n5157 ^ x268;
  assign n5358 = x1152 & n5134;
  assign n5359 = x1150 & n5137;
  assign n5360 = ~n5358 & ~n5359;
  assign n5361 = x1151 & n5141;
  assign n5362 = n5360 & ~n5361;
  assign n5364 = n5363 ^ n5362;
  assign n5365 = ~n5131 & ~n5364;
  assign n5366 = n5365 ^ n5363;
  assign n5370 = x1136 & n5137;
  assign n5371 = x1138 & n5134;
  assign n5372 = ~n5370 & ~n5371;
  assign n5373 = x1137 & n5141;
  assign n5374 = n5372 & ~n5373;
  assign n5367 = x817 ^ x269;
  assign n5368 = n5150 & ~n5367;
  assign n5369 = n5368 ^ x269;
  assign n5375 = n5374 ^ n5369;
  assign n5376 = ~n5131 & n5375;
  assign n5377 = n5376 ^ n5369;
  assign n5381 = x1139 & n5137;
  assign n5382 = x1141 & n5134;
  assign n5383 = ~n5381 & ~n5382;
  assign n5384 = x1140 & n5141;
  assign n5385 = n5383 & ~n5384;
  assign n5378 = x805 ^ x270;
  assign n5379 = n5150 & ~n5378;
  assign n5380 = n5379 ^ x270;
  assign n5386 = n5385 ^ n5380;
  assign n5387 = ~n5131 & n5386;
  assign n5388 = n5387 ^ n5380;
  assign n5394 = n5152 ^ x271;
  assign n5389 = x1146 & n5141;
  assign n5390 = x1145 & n5137;
  assign n5391 = ~n5389 & ~n5390;
  assign n5392 = x1147 & n5134;
  assign n5393 = n5391 & ~n5392;
  assign n5395 = n5394 ^ n5393;
  assign n5396 = ~n5131 & ~n5395;
  assign n5397 = n5396 ^ n5394;
  assign n5403 = n5155 ^ x272;
  assign n5398 = x1150 & n5134;
  assign n5399 = x1148 & n5137;
  assign n5400 = ~n5398 & ~n5399;
  assign n5401 = x1149 & n5141;
  assign n5402 = n5400 & ~n5401;
  assign n5404 = n5403 ^ n5402;
  assign n5405 = ~n5131 & ~n5404;
  assign n5406 = n5405 ^ n5403;
  assign n5412 = n5153 ^ x273;
  assign n5407 = x1146 & n5137;
  assign n5408 = x1148 & n5134;
  assign n5409 = ~n5407 & ~n5408;
  assign n5410 = x1147 & n5141;
  assign n5411 = n5409 & ~n5410;
  assign n5413 = n5412 ^ n5411;
  assign n5414 = ~n5131 & ~n5413;
  assign n5415 = n5414 ^ n5412;
  assign n5419 = x1145 & n5134;
  assign n5420 = x1143 & n5137;
  assign n5421 = ~n5419 & ~n5420;
  assign n5422 = x1144 & n5141;
  assign n5423 = n5421 & ~n5422;
  assign n5416 = x659 ^ x274;
  assign n5417 = n5150 & ~n5416;
  assign n5418 = n5417 ^ x274;
  assign n5424 = n5423 ^ n5418;
  assign n5425 = ~n5131 & n5424;
  assign n5426 = n5425 ^ n5418;
  assign n5432 = n5156 ^ x275;
  assign n5427 = x1151 & n5134;
  assign n5428 = x1149 & n5137;
  assign n5429 = ~n5427 & ~n5428;
  assign n5430 = x1150 & n5141;
  assign n5431 = n5429 & ~n5430;
  assign n5433 = n5432 ^ n5431;
  assign n5434 = ~n5131 & ~n5433;
  assign n5435 = n5434 ^ n5432;
  assign n5441 = n5151 ^ x276;
  assign n5436 = x1146 & n5134;
  assign n5437 = x1144 & n5137;
  assign n5438 = ~n5436 & ~n5437;
  assign n5439 = x1145 & n5141;
  assign n5440 = n5438 & ~n5439;
  assign n5442 = n5441 ^ n5440;
  assign n5443 = ~n5131 & ~n5442;
  assign n5444 = n5443 ^ n5441;
  assign n5448 = x1140 & n5137;
  assign n5449 = x1142 & n5134;
  assign n5450 = ~n5448 & ~n5449;
  assign n5451 = x1141 & n5141;
  assign n5452 = n5450 & ~n5451;
  assign n5445 = x820 ^ x277;
  assign n5446 = n5150 & ~n5445;
  assign n5447 = n5446 ^ x277;
  assign n5453 = n5452 ^ n5447;
  assign n5454 = ~n5131 & n5453;
  assign n5455 = n5454 ^ n5447;
  assign n5459 = x1132 & n5137;
  assign n5460 = x1134 & n5134;
  assign n5461 = ~n5459 & ~n5460;
  assign n5462 = x1133 & n5141;
  assign n5463 = n5461 & ~n5462;
  assign n5456 = x976 ^ x278;
  assign n5457 = n5150 & n5456;
  assign n5458 = n5457 ^ x278;
  assign n5464 = n5463 ^ n5458;
  assign n5465 = ~n5131 & ~n5464;
  assign n5466 = n5465 ^ n5458;
  assign n5470 = x1133 & n5137;
  assign n5471 = x1135 & n5134;
  assign n5472 = ~n5470 & ~n5471;
  assign n5473 = x1134 & n5141;
  assign n5474 = n5472 & ~n5473;
  assign n5467 = x958 ^ x279;
  assign n5468 = n5150 & n5467;
  assign n5469 = n5468 ^ x279;
  assign n5475 = n5474 ^ n5469;
  assign n5476 = ~n5131 & ~n5475;
  assign n5477 = n5476 ^ n5469;
  assign n5481 = x1135 & n5137;
  assign n5482 = x1137 & n5134;
  assign n5483 = ~n5481 & ~n5482;
  assign n5484 = x1136 & n5141;
  assign n5485 = n5483 & ~n5484;
  assign n5478 = x914 ^ x280;
  assign n5479 = n5150 & ~n5478;
  assign n5480 = n5479 ^ x280;
  assign n5486 = n5485 ^ n5480;
  assign n5487 = ~n5131 & n5486;
  assign n5488 = n5487 ^ n5480;
  assign n5492 = x1137 & n5137;
  assign n5493 = x1139 & n5134;
  assign n5494 = ~n5492 & ~n5493;
  assign n5495 = x1138 & n5141;
  assign n5496 = n5494 & ~n5495;
  assign n5489 = x830 ^ x281;
  assign n5490 = n5150 & ~n5489;
  assign n5491 = n5490 ^ x281;
  assign n5497 = n5496 ^ n5491;
  assign n5498 = ~n5131 & n5497;
  assign n5499 = n5498 ^ n5491;
  assign n5503 = x1138 & n5137;
  assign n5504 = x1140 & n5134;
  assign n5505 = ~n5503 & ~n5504;
  assign n5506 = x1139 & n5141;
  assign n5507 = n5505 & ~n5506;
  assign n5500 = x836 ^ x282;
  assign n5501 = n5150 & ~n5500;
  assign n5502 = n5501 ^ x282;
  assign n5508 = n5507 ^ n5502;
  assign n5509 = ~n5131 & n5508;
  assign n5510 = n5509 ^ n5502;
  assign n5516 = n5154 ^ x283;
  assign n5511 = x1149 & n5134;
  assign n5512 = x1147 & n5137;
  assign n5513 = ~n5511 & ~n5512;
  assign n5514 = x1148 & n5141;
  assign n5515 = n5513 & ~n5514;
  assign n5517 = n5516 ^ n5515;
  assign n5518 = ~n5131 & ~n5517;
  assign n5519 = n5518 ^ n5516;
  assign n5520 = x1143 & ~n3247;
  assign n5521 = n5303 & n5520;
  assign n5522 = ~x284 & n5302;
  assign n5523 = ~n5521 & ~n5522;
  assign n5524 = ~n3111 & n3220;
  assign n5525 = ~n2721 & n5524;
  assign n5526 = x289 & n5525;
  assign n5527 = x286 & x288;
  assign n5528 = n5526 & n5527;
  assign n5529 = n5528 ^ x285;
  assign n5530 = ~x288 & n2721;
  assign n5531 = ~n5524 & n5530;
  assign n5532 = x285 & n2690;
  assign n5533 = n5531 & n5532;
  assign n5534 = ~x793 & ~n5533;
  assign n5535 = n5529 & n5534;
  assign n5536 = x288 & n5525;
  assign n5537 = ~n5531 & ~n5536;
  assign n5538 = x286 & ~n5537;
  assign n5539 = ~x793 & ~n5538;
  assign n5540 = ~n2692 & n5531;
  assign n5541 = ~n5536 & ~n5540;
  assign n5542 = ~x286 & n5541;
  assign n5543 = n5539 & ~n5542;
  assign n5544 = ~x287 & x457;
  assign n5545 = ~x332 & ~n5544;
  assign n5546 = n2728 ^ x288;
  assign n5547 = n5546 ^ n5524;
  assign n5548 = ~x793 & n5547;
  assign n5549 = ~x289 & ~n5536;
  assign n5550 = x286 & ~n5526;
  assign n5551 = ~n5549 & n5550;
  assign n5552 = x289 & ~n5527;
  assign n5553 = n5552 ^ n5532;
  assign n5554 = ~n5531 & n5553;
  assign n5555 = n5554 ^ n5532;
  assign n5556 = ~n5551 & ~n5555;
  assign n5557 = ~x793 & ~n5556;
  assign n5558 = x1048 ^ x290;
  assign n5559 = ~x476 & n5558;
  assign n5560 = n5559 ^ x290;
  assign n5561 = x1049 ^ x291;
  assign n5562 = ~x476 & n5561;
  assign n5563 = n5562 ^ x291;
  assign n5564 = x1084 ^ x292;
  assign n5565 = ~x476 & n5564;
  assign n5566 = n5565 ^ x292;
  assign n5567 = x1059 ^ x293;
  assign n5568 = ~x476 & n5567;
  assign n5569 = n5568 ^ x293;
  assign n5570 = x1072 ^ x294;
  assign n5571 = ~x476 & n5570;
  assign n5572 = n5571 ^ x294;
  assign n5573 = x1053 ^ x295;
  assign n5574 = ~x476 & n5573;
  assign n5575 = n5574 ^ x295;
  assign n5576 = x1037 ^ x296;
  assign n5577 = ~x476 & n5576;
  assign n5578 = n5577 ^ x296;
  assign n5579 = x1044 ^ x297;
  assign n5580 = ~x476 & n5579;
  assign n5581 = n5580 ^ x297;
  assign n5582 = x1044 ^ x298;
  assign n5583 = ~x478 & n5582;
  assign n5584 = n5583 ^ x298;
  assign n5585 = x106 & n3052;
  assign n5586 = x39 & ~x287;
  assign n5587 = n3251 & n5586;
  assign n5588 = ~n3256 & ~n5587;
  assign n5589 = ~n5585 & n5588;
  assign n5590 = n1518 & n1548;
  assign n5591 = n5589 & ~n5590;
  assign n5592 = ~x24 & n1526;
  assign n5593 = ~x312 & n5592;
  assign n5594 = n5593 ^ x300;
  assign n5595 = ~x55 & ~n5594;
  assign n5596 = ~x300 & ~x312;
  assign n5597 = n5592 & n5596;
  assign n5598 = n5597 ^ x301;
  assign n5599 = ~x55 & ~n5598;
  assign n5600 = n1699 ^ n1672;
  assign n5601 = n1656 & n5600;
  assign n5602 = n5601 ^ n1672;
  assign n5603 = x937 & n5602;
  assign n5604 = n1488 & ~n1656;
  assign n5605 = ~n2062 & ~n5604;
  assign n5606 = ~x237 & ~n5605;
  assign n5607 = ~n5603 & ~n5606;
  assign n5608 = n1702 ^ n1675;
  assign n5609 = n1656 & n5608;
  assign n5610 = n5609 ^ n1675;
  assign n5611 = x273 & n5610;
  assign n5612 = x1148 & ~n2139;
  assign n5613 = ~n5611 & ~n5612;
  assign n5614 = n5607 & n5613;
  assign n5615 = x1049 ^ x303;
  assign n5616 = ~x478 & n5615;
  assign n5617 = n5616 ^ x303;
  assign n5618 = x1048 ^ x304;
  assign n5619 = ~x478 & n5618;
  assign n5620 = n5619 ^ x304;
  assign n5621 = x1084 ^ x305;
  assign n5622 = ~x478 & n5621;
  assign n5623 = n5622 ^ x305;
  assign n5624 = x1059 ^ x306;
  assign n5625 = ~x478 & n5624;
  assign n5626 = n5625 ^ x306;
  assign n5627 = x1053 ^ x307;
  assign n5628 = ~x478 & n5627;
  assign n5629 = n5628 ^ x307;
  assign n5630 = x1037 ^ x308;
  assign n5631 = ~x478 & n5630;
  assign n5632 = n5631 ^ x308;
  assign n5633 = x1072 ^ x309;
  assign n5634 = ~x478 & n5633;
  assign n5635 = n5634 ^ x309;
  assign n5636 = x271 & n5610;
  assign n5637 = ~x233 & ~n5605;
  assign n5638 = ~n5636 & ~n5637;
  assign n5639 = x1147 & ~n2139;
  assign n5640 = x934 & n5602;
  assign n5641 = ~n5639 & ~n5640;
  assign n5642 = n5638 & n5641;
  assign n5643 = x301 & n5596;
  assign n5644 = n5592 & n5643;
  assign n5645 = n5644 ^ x311;
  assign n5646 = ~x55 & ~n5645;
  assign n5647 = n5592 ^ x312;
  assign n5648 = ~x55 & n5647;
  assign n5649 = ~n3639 & ~n3652;
  assign n5650 = n2221 & ~n5649;
  assign n5651 = ~n3658 & ~n5650;
  assign n5652 = n5651 ^ x313;
  assign n5653 = ~x954 & n5652;
  assign n5654 = n5653 ^ x313;
  assign n5655 = n3825 & n3983;
  assign n5656 = n4009 & n5655;
  assign n5657 = ~x340 & n5524;
  assign n5658 = x1080 ^ x315;
  assign n5659 = n5657 & n5658;
  assign n5660 = n5659 ^ x315;
  assign n5661 = x1047 ^ x316;
  assign n5662 = n5657 & n5661;
  assign n5663 = n5662 ^ x316;
  assign n5664 = ~x330 & n5524;
  assign n5665 = x1078 ^ x317;
  assign n5666 = n5664 & n5665;
  assign n5667 = n5666 ^ x317;
  assign n5668 = ~x341 & n5524;
  assign n5669 = x1074 ^ x318;
  assign n5670 = n5668 & n5669;
  assign n5671 = n5670 ^ x318;
  assign n5672 = x1072 ^ x319;
  assign n5673 = n5668 & n5672;
  assign n5674 = n5673 ^ x319;
  assign n5675 = x1048 ^ x320;
  assign n5676 = n5657 & n5675;
  assign n5677 = n5676 ^ x320;
  assign n5678 = x1058 ^ x321;
  assign n5679 = n5657 & n5678;
  assign n5680 = n5679 ^ x321;
  assign n5681 = x1051 ^ x322;
  assign n5682 = n5657 & n5681;
  assign n5683 = n5682 ^ x322;
  assign n5684 = x1065 ^ x323;
  assign n5685 = n5657 & n5684;
  assign n5686 = n5685 ^ x323;
  assign n5687 = x1086 ^ x324;
  assign n5688 = n5668 & n5687;
  assign n5689 = n5688 ^ x324;
  assign n5690 = x1063 ^ x325;
  assign n5691 = n5668 & n5690;
  assign n5692 = n5691 ^ x325;
  assign n5693 = x1057 ^ x326;
  assign n5694 = n5668 & n5693;
  assign n5695 = n5694 ^ x326;
  assign n5696 = x1040 ^ x327;
  assign n5697 = n5657 & n5696;
  assign n5698 = n5697 ^ x327;
  assign n5699 = x1058 ^ x328;
  assign n5700 = n5668 & n5699;
  assign n5701 = n5700 ^ x328;
  assign n5702 = x1043 ^ x329;
  assign n5703 = n5668 & n5702;
  assign n5704 = n5703 ^ x329;
  assign n5705 = x1092 & ~n1421;
  assign n5706 = x340 ^ x330;
  assign n5707 = n5524 & n5706;
  assign n5708 = n5707 ^ x330;
  assign n5709 = n5705 & ~n5708;
  assign n5710 = x341 ^ x331;
  assign n5711 = n5524 & n5710;
  assign n5712 = n5711 ^ x331;
  assign n5713 = n5705 & ~n5712;
  assign n5714 = n1662 & n3055;
  assign n5715 = ~n3191 & ~n3342;
  assign n5716 = ~n1535 & n5715;
  assign n5717 = ~n5714 & n5716;
  assign n5718 = x1040 ^ x333;
  assign n5719 = n5668 & n5718;
  assign n5720 = n5719 ^ x333;
  assign n5721 = x1065 ^ x334;
  assign n5722 = n5668 & n5721;
  assign n5723 = n5722 ^ x334;
  assign n5724 = x1069 ^ x335;
  assign n5725 = n5668 & n5724;
  assign n5726 = n5725 ^ x335;
  assign n5727 = x1070 ^ x336;
  assign n5728 = n5664 & n5727;
  assign n5729 = n5728 ^ x336;
  assign n5730 = x1044 ^ x337;
  assign n5731 = n5664 & n5730;
  assign n5732 = n5731 ^ x337;
  assign n5733 = x1072 ^ x338;
  assign n5734 = n5664 & n5733;
  assign n5735 = n5734 ^ x338;
  assign n5736 = x1086 ^ x339;
  assign n5737 = n5664 & n5736;
  assign n5738 = n5737 ^ x339;
  assign n5739 = ~x340 & ~n5524;
  assign n5740 = n5705 & ~n5739;
  assign n5741 = ~x331 & n5524;
  assign n5742 = n5740 & ~n5741;
  assign n5743 = x341 ^ x330;
  assign n5744 = ~n5524 & n5743;
  assign n5745 = n5744 ^ x330;
  assign n5746 = n5705 & ~n5745;
  assign n5747 = x1049 ^ x342;
  assign n5748 = n5657 & n5747;
  assign n5749 = n5748 ^ x342;
  assign n5750 = x1062 ^ x343;
  assign n5751 = n5657 & n5750;
  assign n5752 = n5751 ^ x343;
  assign n5753 = x1069 ^ x344;
  assign n5754 = n5657 & n5753;
  assign n5755 = n5754 ^ x344;
  assign n5756 = x1039 ^ x345;
  assign n5757 = n5657 & n5756;
  assign n5758 = n5757 ^ x345;
  assign n5759 = x1067 ^ x346;
  assign n5760 = n5657 & n5759;
  assign n5761 = n5760 ^ x346;
  assign n5762 = x1055 ^ x347;
  assign n5763 = n5657 & n5762;
  assign n5764 = n5763 ^ x347;
  assign n5765 = x1087 ^ x348;
  assign n5766 = n5657 & n5765;
  assign n5767 = n5766 ^ x348;
  assign n5768 = x1043 ^ x349;
  assign n5769 = n5657 & n5768;
  assign n5770 = n5769 ^ x349;
  assign n5771 = x1035 ^ x350;
  assign n5772 = n5657 & n5771;
  assign n5773 = n5772 ^ x350;
  assign n5774 = x1079 ^ x351;
  assign n5775 = n5657 & n5774;
  assign n5776 = n5775 ^ x351;
  assign n5777 = x1078 ^ x352;
  assign n5778 = n5657 & n5777;
  assign n5779 = n5778 ^ x352;
  assign n5780 = x1063 ^ x353;
  assign n5781 = n5657 & n5780;
  assign n5782 = n5781 ^ x353;
  assign n5783 = x1045 ^ x354;
  assign n5784 = n5657 & n5783;
  assign n5785 = n5784 ^ x354;
  assign n5786 = x1084 ^ x355;
  assign n5787 = n5657 & n5786;
  assign n5788 = n5787 ^ x355;
  assign n5789 = x1081 ^ x356;
  assign n5790 = n5657 & n5789;
  assign n5791 = n5790 ^ x356;
  assign n5792 = x1076 ^ x357;
  assign n5793 = n5657 & n5792;
  assign n5794 = n5793 ^ x357;
  assign n5795 = x1071 ^ x358;
  assign n5796 = n5657 & n5795;
  assign n5797 = n5796 ^ x358;
  assign n5798 = x1068 ^ x359;
  assign n5799 = n5657 & n5798;
  assign n5800 = n5799 ^ x359;
  assign n5801 = x1042 ^ x360;
  assign n5802 = n5657 & n5801;
  assign n5803 = n5802 ^ x360;
  assign n5804 = x1059 ^ x361;
  assign n5805 = n5657 & n5804;
  assign n5806 = n5805 ^ x361;
  assign n5807 = x1070 ^ x362;
  assign n5808 = n5657 & n5807;
  assign n5809 = n5808 ^ x362;
  assign n5810 = x1049 ^ x363;
  assign n5811 = n5664 & n5810;
  assign n5812 = n5811 ^ x363;
  assign n5813 = x1062 ^ x364;
  assign n5814 = n5664 & n5813;
  assign n5815 = n5814 ^ x364;
  assign n5816 = x1065 ^ x365;
  assign n5817 = n5664 & n5816;
  assign n5818 = n5817 ^ x365;
  assign n5819 = x1069 ^ x366;
  assign n5820 = n5664 & n5819;
  assign n5821 = n5820 ^ x366;
  assign n5822 = x1039 ^ x367;
  assign n5823 = n5664 & n5822;
  assign n5824 = n5823 ^ x367;
  assign n5825 = x1067 ^ x368;
  assign n5826 = n5664 & n5825;
  assign n5827 = n5826 ^ x368;
  assign n5828 = x1080 ^ x369;
  assign n5829 = n5664 & n5828;
  assign n5830 = n5829 ^ x369;
  assign n5831 = x1055 ^ x370;
  assign n5832 = n5664 & n5831;
  assign n5833 = n5832 ^ x370;
  assign n5834 = x1051 ^ x371;
  assign n5835 = n5664 & n5834;
  assign n5836 = n5835 ^ x371;
  assign n5837 = x1048 ^ x372;
  assign n5838 = n5664 & n5837;
  assign n5839 = n5838 ^ x372;
  assign n5840 = x1087 ^ x373;
  assign n5841 = n5664 & n5840;
  assign n5842 = n5841 ^ x373;
  assign n5843 = x1035 ^ x374;
  assign n5844 = n5664 & n5843;
  assign n5845 = n5844 ^ x374;
  assign n5846 = x1047 ^ x375;
  assign n5847 = n5664 & n5846;
  assign n5848 = n5847 ^ x375;
  assign n5849 = x1079 ^ x376;
  assign n5850 = n5664 & n5849;
  assign n5851 = n5850 ^ x376;
  assign n5852 = x1074 ^ x377;
  assign n5853 = n5664 & n5852;
  assign n5854 = n5853 ^ x377;
  assign n5855 = x1063 ^ x378;
  assign n5856 = n5664 & n5855;
  assign n5857 = n5856 ^ x378;
  assign n5858 = x1045 ^ x379;
  assign n5859 = n5664 & n5858;
  assign n5860 = n5859 ^ x379;
  assign n5861 = x1084 ^ x380;
  assign n5862 = n5664 & n5861;
  assign n5863 = n5862 ^ x380;
  assign n5864 = x1081 ^ x381;
  assign n5865 = n5664 & n5864;
  assign n5866 = n5865 ^ x381;
  assign n5867 = x1076 ^ x382;
  assign n5868 = n5664 & n5867;
  assign n5869 = n5868 ^ x382;
  assign n5870 = x1071 ^ x383;
  assign n5871 = n5664 & n5870;
  assign n5872 = n5871 ^ x383;
  assign n5873 = x1068 ^ x384;
  assign n5874 = n5664 & n5873;
  assign n5875 = n5874 ^ x384;
  assign n5876 = x1042 ^ x385;
  assign n5877 = n5664 & n5876;
  assign n5878 = n5877 ^ x385;
  assign n5879 = x1059 ^ x386;
  assign n5880 = n5664 & n5879;
  assign n5881 = n5880 ^ x386;
  assign n5882 = x1053 ^ x387;
  assign n5883 = n5664 & n5882;
  assign n5884 = n5883 ^ x387;
  assign n5885 = x1037 ^ x388;
  assign n5886 = n5664 & n5885;
  assign n5887 = n5886 ^ x388;
  assign n5888 = x1036 ^ x389;
  assign n5889 = n5664 & n5888;
  assign n5890 = n5889 ^ x389;
  assign n5891 = x1049 ^ x390;
  assign n5892 = n5668 & n5891;
  assign n5893 = n5892 ^ x390;
  assign n5894 = x1062 ^ x391;
  assign n5895 = n5668 & n5894;
  assign n5896 = n5895 ^ x391;
  assign n5897 = x1039 ^ x392;
  assign n5898 = n5668 & n5897;
  assign n5899 = n5898 ^ x392;
  assign n5900 = x1067 ^ x393;
  assign n5901 = n5668 & n5900;
  assign n5902 = n5901 ^ x393;
  assign n5903 = x1080 ^ x394;
  assign n5904 = n5668 & n5903;
  assign n5905 = n5904 ^ x394;
  assign n5906 = x1055 ^ x395;
  assign n5907 = n5668 & n5906;
  assign n5908 = n5907 ^ x395;
  assign n5909 = x1051 ^ x396;
  assign n5910 = n5668 & n5909;
  assign n5911 = n5910 ^ x396;
  assign n5912 = x1048 ^ x397;
  assign n5913 = n5668 & n5912;
  assign n5914 = n5913 ^ x397;
  assign n5915 = x1087 ^ x398;
  assign n5916 = n5668 & n5915;
  assign n5917 = n5916 ^ x398;
  assign n5918 = x1047 ^ x399;
  assign n5919 = n5668 & n5918;
  assign n5920 = n5919 ^ x399;
  assign n5921 = x1035 ^ x400;
  assign n5922 = n5668 & n5921;
  assign n5923 = n5922 ^ x400;
  assign n5924 = x1079 ^ x401;
  assign n5925 = n5668 & n5924;
  assign n5926 = n5925 ^ x401;
  assign n5927 = x1078 ^ x402;
  assign n5928 = n5668 & n5927;
  assign n5929 = n5928 ^ x402;
  assign n5930 = x1045 ^ x403;
  assign n5931 = n5668 & n5930;
  assign n5932 = n5931 ^ x403;
  assign n5933 = x1084 ^ x404;
  assign n5934 = n5668 & n5933;
  assign n5935 = n5934 ^ x404;
  assign n5936 = x1081 ^ x405;
  assign n5937 = n5668 & n5936;
  assign n5938 = n5937 ^ x405;
  assign n5939 = x1076 ^ x406;
  assign n5940 = n5668 & n5939;
  assign n5941 = n5940 ^ x406;
  assign n5942 = x1071 ^ x407;
  assign n5943 = n5668 & n5942;
  assign n5944 = n5943 ^ x407;
  assign n5945 = x1068 ^ x408;
  assign n5946 = n5668 & n5945;
  assign n5947 = n5946 ^ x408;
  assign n5948 = x1042 ^ x409;
  assign n5949 = n5668 & n5948;
  assign n5950 = n5949 ^ x409;
  assign n5951 = x1059 ^ x410;
  assign n5952 = n5668 & n5951;
  assign n5953 = n5952 ^ x410;
  assign n5954 = x1053 ^ x411;
  assign n5955 = n5668 & n5954;
  assign n5956 = n5955 ^ x411;
  assign n5957 = x1037 ^ x412;
  assign n5958 = n5668 & n5957;
  assign n5959 = n5958 ^ x412;
  assign n5960 = x1036 ^ x413;
  assign n5961 = n5668 & n5960;
  assign n5962 = n5961 ^ x413;
  assign n5963 = x1049 ^ x414;
  assign n5964 = n5741 & n5963;
  assign n5965 = n5964 ^ x414;
  assign n5966 = x1062 ^ x415;
  assign n5967 = n5741 & n5966;
  assign n5968 = n5967 ^ x415;
  assign n5969 = x1069 ^ x416;
  assign n5970 = n5741 & n5969;
  assign n5971 = n5970 ^ x416;
  assign n5972 = x1039 ^ x417;
  assign n5973 = n5741 & n5972;
  assign n5974 = n5973 ^ x417;
  assign n5975 = x1067 ^ x418;
  assign n5976 = n5741 & n5975;
  assign n5977 = n5976 ^ x418;
  assign n5978 = x1080 ^ x419;
  assign n5979 = n5741 & n5978;
  assign n5980 = n5979 ^ x419;
  assign n5981 = x1055 ^ x420;
  assign n5982 = n5741 & n5981;
  assign n5983 = n5982 ^ x420;
  assign n5984 = x1051 ^ x421;
  assign n5985 = n5741 & n5984;
  assign n5986 = n5985 ^ x421;
  assign n5987 = x1048 ^ x422;
  assign n5988 = n5741 & n5987;
  assign n5989 = n5988 ^ x422;
  assign n5990 = x1087 ^ x423;
  assign n5991 = n5741 & n5990;
  assign n5992 = n5991 ^ x423;
  assign n5993 = x1047 ^ x424;
  assign n5994 = n5741 & n5993;
  assign n5995 = n5994 ^ x424;
  assign n5996 = x1035 ^ x425;
  assign n5997 = n5741 & n5996;
  assign n5998 = n5997 ^ x425;
  assign n5999 = x1079 ^ x426;
  assign n6000 = n5741 & n5999;
  assign n6001 = n6000 ^ x426;
  assign n6002 = x1078 ^ x427;
  assign n6003 = n5741 & n6002;
  assign n6004 = n6003 ^ x427;
  assign n6005 = x1045 ^ x428;
  assign n6006 = n5741 & n6005;
  assign n6007 = n6006 ^ x428;
  assign n6008 = x1084 ^ x429;
  assign n6009 = n5741 & n6008;
  assign n6010 = n6009 ^ x429;
  assign n6011 = x1076 ^ x430;
  assign n6012 = n5741 & n6011;
  assign n6013 = n6012 ^ x430;
  assign n6014 = x1071 ^ x431;
  assign n6015 = n5741 & n6014;
  assign n6016 = n6015 ^ x431;
  assign n6017 = x1068 ^ x432;
  assign n6018 = n5741 & n6017;
  assign n6019 = n6018 ^ x432;
  assign n6020 = x1042 ^ x433;
  assign n6021 = n5741 & n6020;
  assign n6022 = n6021 ^ x433;
  assign n6023 = x1059 ^ x434;
  assign n6024 = n5741 & n6023;
  assign n6025 = n6024 ^ x434;
  assign n6026 = x1053 ^ x435;
  assign n6027 = n5741 & n6026;
  assign n6028 = n6027 ^ x435;
  assign n6029 = x1037 ^ x436;
  assign n6030 = n5741 & n6029;
  assign n6031 = n6030 ^ x436;
  assign n6032 = x1070 ^ x437;
  assign n6033 = n5741 & n6032;
  assign n6034 = n6033 ^ x437;
  assign n6035 = x1036 ^ x438;
  assign n6036 = n5741 & n6035;
  assign n6037 = n6036 ^ x438;
  assign n6038 = x1057 ^ x439;
  assign n6039 = n5664 & n6038;
  assign n6040 = n6039 ^ x439;
  assign n6041 = x1043 ^ x440;
  assign n6042 = n5664 & n6041;
  assign n6043 = n6042 ^ x440;
  assign n6044 = x1044 ^ x441;
  assign n6045 = n5657 & n6044;
  assign n6046 = n6045 ^ x441;
  assign n6047 = x1058 ^ x442;
  assign n6048 = n5664 & n6047;
  assign n6049 = n6048 ^ x442;
  assign n6050 = x1044 ^ x443;
  assign n6051 = n5741 & n6050;
  assign n6052 = n6051 ^ x443;
  assign n6053 = x1072 ^ x444;
  assign n6054 = n5741 & n6053;
  assign n6055 = n6054 ^ x444;
  assign n6056 = x1081 ^ x445;
  assign n6057 = n5741 & n6056;
  assign n6058 = n6057 ^ x445;
  assign n6059 = x1086 ^ x446;
  assign n6060 = n5741 & n6059;
  assign n6061 = n6060 ^ x446;
  assign n6062 = x1040 ^ x447;
  assign n6063 = n5664 & n6062;
  assign n6064 = n6063 ^ x447;
  assign n6065 = x1074 ^ x448;
  assign n6066 = n5741 & n6065;
  assign n6067 = n6066 ^ x448;
  assign n6068 = x1057 ^ x449;
  assign n6069 = n5741 & n6068;
  assign n6070 = n6069 ^ x449;
  assign n6071 = x1036 ^ x450;
  assign n6072 = n5657 & n6071;
  assign n6073 = n6072 ^ x450;
  assign n6074 = x1063 ^ x451;
  assign n6075 = n5741 & n6074;
  assign n6076 = n6075 ^ x451;
  assign n6077 = x1053 ^ x452;
  assign n6078 = n5657 & n6077;
  assign n6079 = n6078 ^ x452;
  assign n6080 = x1040 ^ x453;
  assign n6081 = n5741 & n6080;
  assign n6082 = n6081 ^ x453;
  assign n6083 = x1043 ^ x454;
  assign n6084 = n5741 & n6083;
  assign n6085 = n6084 ^ x454;
  assign n6086 = x1037 ^ x455;
  assign n6087 = n5657 & n6086;
  assign n6088 = n6087 ^ x455;
  assign n6089 = x1044 ^ x456;
  assign n6090 = n5668 & n6089;
  assign n6091 = n6090 ^ x456;
  assign n6092 = x599 & x815;
  assign n6093 = x810 & ~n6092;
  assign n6094 = x596 & ~n6093;
  assign n6095 = x804 & ~n6094;
  assign n6096 = x594 & x600;
  assign n6097 = x597 & x601;
  assign n6098 = n6096 & n6097;
  assign n6099 = ~x804 & ~x810;
  assign n6100 = ~x595 & ~n6099;
  assign n6101 = n6098 & ~n6100;
  assign n6102 = ~n6095 & n6101;
  assign n6103 = ~x601 & ~n6099;
  assign n6104 = ~x815 & ~n6103;
  assign n6105 = x600 & ~x810;
  assign n6106 = x804 & ~n6105;
  assign n6107 = n6104 & ~n6106;
  assign n6108 = ~n6102 & ~n6107;
  assign n6109 = x605 & ~n6108;
  assign n6110 = ~x815 & x990;
  assign n6111 = n6096 & n6110;
  assign n6112 = n6106 & n6111;
  assign n6113 = ~n6109 & ~n6112;
  assign n6114 = x821 & ~n6113;
  assign n6115 = x1072 ^ x458;
  assign n6116 = n5657 & n6115;
  assign n6117 = n6116 ^ x458;
  assign n6118 = x1058 ^ x459;
  assign n6119 = n5741 & n6118;
  assign n6120 = n6119 ^ x459;
  assign n6121 = x1086 ^ x460;
  assign n6122 = n5657 & n6121;
  assign n6123 = n6122 ^ x460;
  assign n6124 = x1057 ^ x461;
  assign n6125 = n5657 & n6124;
  assign n6126 = n6125 ^ x461;
  assign n6127 = x1074 ^ x462;
  assign n6128 = n5657 & n6127;
  assign n6129 = n6128 ^ x462;
  assign n6130 = x1070 ^ x463;
  assign n6131 = n5668 & n6130;
  assign n6132 = n6131 ^ x463;
  assign n6133 = x1065 ^ x464;
  assign n6134 = n5741 & n6133;
  assign n6135 = n6134 ^ x464;
  assign n6136 = ~x243 & n5610;
  assign n6137 = x926 & n5602;
  assign n6138 = ~n6136 & ~n6137;
  assign n6139 = x1157 & ~n2139;
  assign n6140 = n6138 & ~n6139;
  assign n6141 = x275 & n5610;
  assign n6142 = x943 & n5602;
  assign n6143 = ~n6141 & ~n6142;
  assign n6144 = x1151 & ~n2139;
  assign n6145 = n6143 & ~n6144;
  assign n6146 = n3307 & n4830;
  assign n6147 = x40 & x1001;
  assign n6148 = n2186 & n6147;
  assign n6149 = n2183 & n6148;
  assign n6150 = ~n6146 & ~n6149;
  assign n6151 = ~x24 & n1535;
  assign n6152 = x468 & ~n6151;
  assign n6153 = ~n3286 & ~n6152;
  assign n6154 = x942 & n5602;
  assign n6155 = ~x263 & n5610;
  assign n6156 = ~n6154 & ~n6155;
  assign n6157 = x1156 & ~n2139;
  assign n6158 = n6156 & ~n6157;
  assign n6159 = x925 & n5602;
  assign n6160 = x267 & n5610;
  assign n6161 = ~n6159 & ~n6160;
  assign n6162 = x1155 & ~n2139;
  assign n6163 = n6161 & ~n6162;
  assign n6164 = x941 & n5602;
  assign n6165 = x253 & n5610;
  assign n6166 = ~n6164 & ~n6165;
  assign n6167 = x1153 & ~n2139;
  assign n6168 = n6166 & ~n6167;
  assign n6169 = x254 & n5610;
  assign n6170 = x923 & n5602;
  assign n6171 = ~n6169 & ~n6170;
  assign n6172 = x1154 & ~n2139;
  assign n6173 = n6171 & ~n6172;
  assign n6174 = x922 & n5602;
  assign n6175 = x268 & n5610;
  assign n6176 = ~n6174 & ~n6175;
  assign n6177 = x1152 & ~n2139;
  assign n6178 = n6176 & ~n6177;
  assign n6179 = x931 & n5602;
  assign n6180 = x272 & n5610;
  assign n6181 = ~n6179 & ~n6180;
  assign n6182 = x1150 & ~n2139;
  assign n6183 = n6181 & ~n6182;
  assign n6184 = x936 & n5602;
  assign n6185 = x283 & n5610;
  assign n6186 = ~n6184 & ~n6185;
  assign n6187 = x1149 & ~n2139;
  assign n6188 = n6186 & ~n6187;
  assign n6189 = x71 & n5141;
  assign n6190 = ~n3536 & ~n6189;
  assign n6191 = x71 & n5137;
  assign n6192 = x481 ^ x248;
  assign n6193 = ~n4643 & n6192;
  assign n6194 = n6193 ^ x248;
  assign n6195 = x482 ^ x249;
  assign n6196 = ~n4658 & n6195;
  assign n6197 = n6196 ^ x249;
  assign n6198 = x483 ^ x242;
  assign n6199 = ~n4680 & n6198;
  assign n6200 = n6199 ^ x242;
  assign n6201 = x484 ^ x249;
  assign n6202 = ~n4680 & n6201;
  assign n6203 = n6202 ^ x249;
  assign n6204 = x485 ^ x234;
  assign n6205 = ~n4750 & n6204;
  assign n6206 = n6205 ^ x234;
  assign n6207 = x486 ^ x244;
  assign n6208 = ~n4750 & n6207;
  assign n6209 = n6208 ^ x244;
  assign n6210 = x487 ^ x246;
  assign n6211 = ~n4643 & n6210;
  assign n6212 = n6211 ^ x246;
  assign n6213 = x488 ^ x239;
  assign n6214 = ~n4643 & ~n6213;
  assign n6215 = n6214 ^ x239;
  assign n6216 = x489 ^ x242;
  assign n6217 = ~n4750 & n6216;
  assign n6218 = n6217 ^ x242;
  assign n6219 = x490 ^ x241;
  assign n6220 = ~n4680 & n6219;
  assign n6221 = n6220 ^ x241;
  assign n6222 = x491 ^ x238;
  assign n6223 = ~n4680 & n6222;
  assign n6224 = n6223 ^ x238;
  assign n6225 = x492 ^ x240;
  assign n6226 = ~n4680 & n6225;
  assign n6227 = n6226 ^ x240;
  assign n6228 = x493 ^ x244;
  assign n6229 = ~n4680 & n6228;
  assign n6230 = n6229 ^ x244;
  assign n6231 = x494 ^ x239;
  assign n6232 = ~n4680 & ~n6231;
  assign n6233 = n6232 ^ x239;
  assign n6234 = x495 ^ x235;
  assign n6235 = ~n4680 & n6234;
  assign n6236 = n6235 ^ x235;
  assign n6237 = x496 ^ x249;
  assign n6238 = ~n4673 & n6237;
  assign n6239 = n6238 ^ x249;
  assign n6240 = x497 ^ x239;
  assign n6241 = ~n4673 & ~n6240;
  assign n6242 = n6241 ^ x239;
  assign n6243 = x498 ^ x238;
  assign n6244 = ~n4658 & n6243;
  assign n6245 = n6244 ^ x238;
  assign n6246 = x499 ^ x246;
  assign n6247 = ~n4673 & n6246;
  assign n6248 = n6247 ^ x246;
  assign n6249 = x500 ^ x241;
  assign n6250 = ~n4673 & n6249;
  assign n6251 = n6250 ^ x241;
  assign n6252 = x501 ^ x248;
  assign n6253 = ~n4673 & n6252;
  assign n6254 = n6253 ^ x248;
  assign n6255 = x502 ^ x247;
  assign n6256 = ~n4673 & n6255;
  assign n6257 = n6256 ^ x247;
  assign n6258 = x503 ^ x245;
  assign n6259 = ~n4673 & n6258;
  assign n6260 = n6259 ^ x245;
  assign n6261 = x504 ^ x242;
  assign n6262 = ~n4669 & n6261;
  assign n6263 = n6262 ^ x242;
  assign n6264 = x505 ^ x234;
  assign n6265 = ~n4673 & n6264;
  assign n6266 = n6265 ^ x234;
  assign n6267 = x506 ^ x241;
  assign n6268 = ~n4669 & n6267;
  assign n6269 = n6268 ^ x241;
  assign n6270 = x507 ^ x238;
  assign n6271 = ~n4669 & n6270;
  assign n6272 = n6271 ^ x238;
  assign n6273 = x508 ^ x247;
  assign n6274 = ~n4669 & n6273;
  assign n6275 = n6274 ^ x247;
  assign n6276 = x509 ^ x245;
  assign n6277 = ~n4669 & n6276;
  assign n6278 = n6277 ^ x245;
  assign n6279 = x510 ^ x242;
  assign n6280 = ~n4643 & n6279;
  assign n6281 = n6280 ^ x242;
  assign n6282 = x511 ^ x234;
  assign n6283 = ~n4643 & n6282;
  assign n6284 = n6283 ^ x234;
  assign n6285 = x512 ^ x235;
  assign n6286 = ~n4643 & n6285;
  assign n6287 = n6286 ^ x235;
  assign n6288 = x513 ^ x244;
  assign n6289 = ~n4643 & n6288;
  assign n6290 = n6289 ^ x244;
  assign n6291 = x514 ^ x245;
  assign n6292 = ~n4643 & n6291;
  assign n6293 = n6292 ^ x245;
  assign n6294 = x515 ^ x240;
  assign n6295 = ~n4643 & n6294;
  assign n6296 = n6295 ^ x240;
  assign n6297 = x516 ^ x247;
  assign n6298 = ~n4643 & n6297;
  assign n6299 = n6298 ^ x247;
  assign n6300 = x517 ^ x238;
  assign n6301 = ~n4643 & n6300;
  assign n6302 = n6301 ^ x238;
  assign n6303 = x518 ^ x234;
  assign n6304 = ~n4651 & n6303;
  assign n6305 = n6304 ^ x234;
  assign n6306 = x519 ^ x239;
  assign n6307 = ~n4651 & ~n6306;
  assign n6308 = n6307 ^ x239;
  assign n6309 = x520 ^ x246;
  assign n6310 = ~n4651 & n6309;
  assign n6311 = n6310 ^ x246;
  assign n6312 = x521 ^ x248;
  assign n6313 = ~n4651 & n6312;
  assign n6314 = n6313 ^ x248;
  assign n6315 = x522 ^ x238;
  assign n6316 = ~n4651 & n6315;
  assign n6317 = n6316 ^ x238;
  assign n6318 = x523 ^ x234;
  assign n6319 = ~n4760 & n6318;
  assign n6320 = n6319 ^ x234;
  assign n6321 = x524 ^ x239;
  assign n6322 = ~n4760 & ~n6321;
  assign n6323 = n6322 ^ x239;
  assign n6324 = x525 ^ x245;
  assign n6325 = ~n4760 & n6324;
  assign n6326 = n6325 ^ x245;
  assign n6327 = x526 ^ x246;
  assign n6328 = ~n4760 & n6327;
  assign n6329 = n6328 ^ x246;
  assign n6330 = x527 ^ x247;
  assign n6331 = ~n4760 & n6330;
  assign n6332 = n6331 ^ x247;
  assign n6333 = x528 ^ x249;
  assign n6334 = ~n4760 & n6333;
  assign n6335 = n6334 ^ x249;
  assign n6336 = x529 ^ x238;
  assign n6337 = ~n4760 & n6336;
  assign n6338 = n6337 ^ x238;
  assign n6339 = x530 ^ x240;
  assign n6340 = ~n4760 & n6339;
  assign n6341 = n6340 ^ x240;
  assign n6342 = x531 ^ x235;
  assign n6343 = ~n4658 & n6342;
  assign n6344 = n6343 ^ x235;
  assign n6345 = x532 ^ x247;
  assign n6346 = ~n4658 & n6345;
  assign n6347 = n6346 ^ x247;
  assign n6348 = x533 ^ x235;
  assign n6349 = ~n4669 & n6348;
  assign n6350 = n6349 ^ x235;
  assign n6351 = x534 ^ x239;
  assign n6352 = ~n4669 & ~n6351;
  assign n6353 = n6352 ^ x239;
  assign n6354 = x535 ^ x240;
  assign n6355 = ~n4669 & n6354;
  assign n6356 = n6355 ^ x240;
  assign n6357 = x536 ^ x246;
  assign n6358 = ~n4669 & n6357;
  assign n6359 = n6358 ^ x246;
  assign n6360 = x537 ^ x248;
  assign n6361 = ~n4669 & n6360;
  assign n6362 = n6361 ^ x248;
  assign n6363 = x538 ^ x249;
  assign n6364 = ~n4669 & n6363;
  assign n6365 = n6364 ^ x249;
  assign n6366 = x539 ^ x242;
  assign n6367 = ~n4673 & n6366;
  assign n6368 = n6367 ^ x242;
  assign n6369 = x540 ^ x235;
  assign n6370 = ~n4673 & n6369;
  assign n6371 = n6370 ^ x235;
  assign n6372 = x541 ^ x244;
  assign n6373 = ~n4673 & n6372;
  assign n6374 = n6373 ^ x244;
  assign n6375 = x542 ^ x240;
  assign n6376 = ~n4673 & n6375;
  assign n6377 = n6376 ^ x240;
  assign n6378 = x543 ^ x238;
  assign n6379 = ~n4673 & n6378;
  assign n6380 = n6379 ^ x238;
  assign n6381 = x544 ^ x234;
  assign n6382 = ~n4680 & n6381;
  assign n6383 = n6382 ^ x234;
  assign n6384 = x545 ^ x245;
  assign n6385 = ~n4680 & n6384;
  assign n6386 = n6385 ^ x245;
  assign n6387 = x546 ^ x246;
  assign n6388 = ~n4680 & n6387;
  assign n6389 = n6388 ^ x246;
  assign n6390 = x547 ^ x247;
  assign n6391 = ~n4680 & n6390;
  assign n6392 = n6391 ^ x247;
  assign n6393 = x548 ^ x248;
  assign n6394 = ~n4680 & n6393;
  assign n6395 = n6394 ^ x248;
  assign n6396 = x549 ^ x235;
  assign n6397 = ~n4750 & n6396;
  assign n6398 = n6397 ^ x235;
  assign n6399 = x550 ^ x239;
  assign n6400 = ~n4750 & ~n6399;
  assign n6401 = n6400 ^ x239;
  assign n6402 = x551 ^ x240;
  assign n6403 = ~n4750 & n6402;
  assign n6404 = n6403 ^ x240;
  assign n6405 = x552 ^ x247;
  assign n6406 = ~n4750 & n6405;
  assign n6407 = n6406 ^ x247;
  assign n6408 = x553 ^ x241;
  assign n6409 = ~n4750 & n6408;
  assign n6410 = n6409 ^ x241;
  assign n6411 = x554 ^ x248;
  assign n6412 = ~n4750 & n6411;
  assign n6413 = n6412 ^ x248;
  assign n6414 = x555 ^ x249;
  assign n6415 = ~n4750 & n6414;
  assign n6416 = n6415 ^ x249;
  assign n6417 = x556 ^ x242;
  assign n6418 = ~n4658 & n6417;
  assign n6419 = n6418 ^ x242;
  assign n6420 = x557 ^ x234;
  assign n6421 = ~n4669 & n6420;
  assign n6422 = n6421 ^ x234;
  assign n6423 = x558 ^ x244;
  assign n6424 = ~n4669 & n6423;
  assign n6425 = n6424 ^ x244;
  assign n6426 = x559 ^ x241;
  assign n6427 = ~n4643 & n6426;
  assign n6428 = n6427 ^ x241;
  assign n6429 = x560 ^ x240;
  assign n6430 = ~n4658 & n6429;
  assign n6431 = n6430 ^ x240;
  assign n6432 = x561 ^ x247;
  assign n6433 = ~n4651 & n6432;
  assign n6434 = n6433 ^ x247;
  assign n6435 = x562 ^ x241;
  assign n6436 = ~n4658 & n6435;
  assign n6437 = n6436 ^ x241;
  assign n6438 = x563 ^ x246;
  assign n6439 = ~n4750 & n6438;
  assign n6440 = n6439 ^ x246;
  assign n6441 = x564 ^ x246;
  assign n6442 = ~n4658 & n6441;
  assign n6443 = n6442 ^ x246;
  assign n6444 = x565 ^ x248;
  assign n6445 = ~n4658 & n6444;
  assign n6446 = n6445 ^ x248;
  assign n6447 = x566 ^ x244;
  assign n6448 = ~n4658 & n6447;
  assign n6449 = n6448 ^ x244;
  assign n6450 = x665 & n4232;
  assign n6451 = x621 & n4206;
  assign n6452 = ~n6450 & ~n6451;
  assign n6453 = x230 & x1093;
  assign n6454 = x1091 & n6453;
  assign n6455 = ~n6452 & n6454;
  assign n6456 = ~x567 & ~n6453;
  assign n6457 = ~n6455 & ~n6456;
  assign n6458 = x1092 & ~n6457;
  assign n6459 = x568 ^ x245;
  assign n6460 = ~n4658 & n6459;
  assign n6461 = n6460 ^ x245;
  assign n6462 = x569 ^ x239;
  assign n6463 = ~n4658 & ~n6462;
  assign n6464 = n6463 ^ x239;
  assign n6465 = x570 ^ x234;
  assign n6466 = ~n4658 & n6465;
  assign n6467 = n6466 ^ x234;
  assign n6468 = x571 ^ x241;
  assign n6469 = ~n4760 & n6468;
  assign n6470 = n6469 ^ x241;
  assign n6471 = x572 ^ x244;
  assign n6472 = ~n4760 & n6471;
  assign n6473 = n6472 ^ x244;
  assign n6474 = x573 ^ x242;
  assign n6475 = ~n4760 & n6474;
  assign n6476 = n6475 ^ x242;
  assign n6477 = x574 ^ x241;
  assign n6478 = ~n4651 & n6477;
  assign n6479 = n6478 ^ x241;
  assign n6480 = x575 ^ x235;
  assign n6481 = ~n4760 & n6480;
  assign n6482 = n6481 ^ x235;
  assign n6483 = x576 ^ x248;
  assign n6484 = ~n4760 & n6483;
  assign n6485 = n6484 ^ x248;
  assign n6486 = x577 ^ x238;
  assign n6487 = ~n4750 & n6486;
  assign n6488 = n6487 ^ x238;
  assign n6489 = x578 ^ x249;
  assign n6490 = ~n4651 & n6489;
  assign n6491 = n6490 ^ x249;
  assign n6492 = x579 ^ x249;
  assign n6493 = ~n4643 & n6492;
  assign n6494 = n6493 ^ x249;
  assign n6495 = x580 ^ x245;
  assign n6496 = ~n4750 & n6495;
  assign n6497 = n6496 ^ x245;
  assign n6498 = x581 ^ x235;
  assign n6499 = ~n4651 & n6498;
  assign n6500 = n6499 ^ x235;
  assign n6501 = x582 ^ x240;
  assign n6502 = ~n4651 & n6501;
  assign n6503 = n6502 ^ x240;
  assign n6504 = x584 ^ x245;
  assign n6505 = ~n4651 & n6504;
  assign n6506 = n6505 ^ x245;
  assign n6507 = x585 ^ x244;
  assign n6508 = ~n4651 & n6507;
  assign n6509 = n6508 ^ x244;
  assign n6510 = x586 ^ x242;
  assign n6511 = ~n4651 & n6510;
  assign n6512 = n6511 ^ x242;
  assign n6513 = n4208 ^ x587;
  assign n6514 = x230 & n6513;
  assign n6515 = n6514 ^ x587;
  assign n6516 = ~x123 & x824;
  assign n6517 = x950 & n6516;
  assign n6518 = ~x588 & ~n6517;
  assign n6519 = n5705 & ~n6518;
  assign n6520 = ~x591 & n6517;
  assign n6521 = n6519 & ~n6520;
  assign n6522 = x204 & x237;
  assign n6523 = x233 & ~n6522;
  assign n6524 = x206 & ~x237;
  assign n6525 = n6523 & ~n6524;
  assign n6526 = x218 ^ x205;
  assign n6527 = ~x237 & n6526;
  assign n6528 = n6527 ^ x205;
  assign n6529 = ~x233 & ~n6528;
  assign n6530 = ~n6525 & ~n6529;
  assign n6531 = ~n4664 & ~n6530;
  assign n6532 = x201 & x237;
  assign n6533 = x233 & ~n6532;
  assign n6534 = x220 & ~x237;
  assign n6535 = n6533 & ~n6534;
  assign n6536 = x203 ^ x202;
  assign n6537 = ~x237 & n6536;
  assign n6538 = n6537 ^ x202;
  assign n6539 = ~x233 & ~n6538;
  assign n6540 = ~n6535 & ~n6539;
  assign n6541 = n4637 & ~n6540;
  assign n6542 = ~n6531 & ~n6541;
  assign n6543 = x588 & n6517;
  assign n6544 = n5705 & ~n6543;
  assign n6545 = x590 & ~n6517;
  assign n6546 = n6544 & ~n6545;
  assign n6547 = ~x591 & ~n6517;
  assign n6548 = n5705 & ~n6547;
  assign n6549 = ~x592 & n6517;
  assign n6550 = n6548 & ~n6549;
  assign n6551 = ~x592 & ~n6517;
  assign n6552 = n5705 & ~n6551;
  assign n6553 = ~x590 & n6517;
  assign n6554 = n6552 & ~n6553;
  assign n6594 = ~x238 & x507;
  assign n6595 = x233 & ~n6594;
  assign n6596 = ~n6363 & n6595;
  assign n6597 = ~n6261 & ~n6348;
  assign n6598 = n6596 & n6597;
  assign n6599 = x238 & ~x507;
  assign n6600 = ~n6273 & ~n6599;
  assign n6601 = n6598 & n6600;
  assign n6602 = ~n6354 & ~n6420;
  assign n6603 = ~n6267 & ~n6423;
  assign n6604 = n6602 & n6603;
  assign n6605 = ~n6276 & ~n6360;
  assign n6606 = n6351 & ~n6357;
  assign n6607 = n6605 & n6606;
  assign n6608 = n6604 & n6607;
  assign n6609 = n6601 & n6608;
  assign n6610 = ~x245 & x503;
  assign n6611 = ~x246 & x499;
  assign n6612 = ~n6610 & ~n6611;
  assign n6613 = x241 & ~x500;
  assign n6614 = ~n6366 & ~n6613;
  assign n6615 = n6612 & n6614;
  assign n6616 = ~x233 & ~n6237;
  assign n6617 = n6615 & n6616;
  assign n6618 = x246 & ~x499;
  assign n6619 = ~x241 & x500;
  assign n6620 = ~n6618 & ~n6619;
  assign n6621 = x245 & ~x503;
  assign n6622 = n6620 & ~n6621;
  assign n6623 = n6617 & n6622;
  assign n6624 = ~n6252 & ~n6378;
  assign n6625 = ~n6255 & ~n6369;
  assign n6626 = n6624 & n6625;
  assign n6627 = ~n6264 & ~n6372;
  assign n6628 = n6240 & ~n6375;
  assign n6629 = n6627 & n6628;
  assign n6630 = n6626 & n6629;
  assign n6631 = n6623 & n6630;
  assign n6632 = ~n6609 & ~n6631;
  assign n6555 = x248 & ~x554;
  assign n6556 = ~x247 & x552;
  assign n6557 = ~n6555 & ~n6556;
  assign n6558 = ~x240 & x551;
  assign n6559 = ~n6216 & ~n6558;
  assign n6560 = n6557 & n6559;
  assign n6561 = ~x233 & ~n6207;
  assign n6562 = n6560 & n6561;
  assign n6563 = x240 & ~x551;
  assign n6564 = ~x248 & x554;
  assign n6565 = ~n6563 & ~n6564;
  assign n6566 = x247 & ~x552;
  assign n6567 = n6565 & ~n6566;
  assign n6568 = n6562 & n6567;
  assign n6569 = ~n6438 & ~n6486;
  assign n6570 = ~n6204 & ~n6495;
  assign n6571 = n6569 & n6570;
  assign n6572 = ~n6396 & ~n6414;
  assign n6573 = n6399 & ~n6408;
  assign n6574 = n6572 & n6573;
  assign n6575 = n6571 & n6574;
  assign n6576 = n6568 & n6575;
  assign n6577 = ~x241 & x490;
  assign n6578 = x233 & ~n6577;
  assign n6579 = ~n6390 & n6578;
  assign n6580 = ~n6198 & ~n6384;
  assign n6581 = n6579 & n6580;
  assign n6582 = x241 & ~x490;
  assign n6583 = ~n6222 & ~n6582;
  assign n6584 = n6581 & n6583;
  assign n6585 = ~n6201 & ~n6387;
  assign n6586 = ~n6228 & ~n6393;
  assign n6587 = n6585 & n6586;
  assign n6588 = ~n6225 & ~n6381;
  assign n6589 = n6231 & ~n6234;
  assign n6590 = n6588 & n6589;
  assign n6591 = n6587 & n6590;
  assign n6592 = n6584 & n6591;
  assign n6593 = ~n6576 & ~n6592;
  assign n6633 = n6632 ^ n6593;
  assign n6634 = ~x237 & n6633;
  assign n6635 = n6634 ^ n6632;
  assign n6636 = ~n4664 & ~n6635;
  assign n6637 = ~x245 & x514;
  assign n6638 = ~n6492 & ~n6637;
  assign n6639 = x233 & n6638;
  assign n6640 = ~n6297 & ~n6426;
  assign n6641 = n6639 & n6640;
  assign n6642 = x245 & ~x514;
  assign n6643 = ~n6192 & ~n6642;
  assign n6644 = n6641 & n6643;
  assign n6645 = ~n6282 & ~n6288;
  assign n6646 = ~n6279 & ~n6294;
  assign n6647 = n6645 & n6646;
  assign n6648 = n6213 & ~n6285;
  assign n6649 = ~n6210 & ~n6300;
  assign n6650 = n6648 & n6649;
  assign n6651 = n6647 & n6650;
  assign n6652 = n6644 & n6651;
  assign n6653 = x237 & ~n6652;
  assign n6654 = ~x248 & x521;
  assign n6655 = ~x233 & ~n6654;
  assign n6656 = ~n6477 & n6655;
  assign n6657 = ~n6315 & ~n6489;
  assign n6658 = n6656 & n6657;
  assign n6659 = x248 & ~x521;
  assign n6660 = ~n6507 & ~n6659;
  assign n6661 = n6658 & n6660;
  assign n6662 = n6306 & ~n6504;
  assign n6663 = ~n6303 & ~n6309;
  assign n6664 = n6662 & n6663;
  assign n6665 = ~n6432 & ~n6510;
  assign n6666 = ~n6498 & ~n6501;
  assign n6667 = n6665 & n6666;
  assign n6668 = n6664 & n6667;
  assign n6669 = n6661 & n6668;
  assign n6670 = n6653 & ~n6669;
  assign n6671 = n4637 & ~n6670;
  assign n6672 = n6321 & ~n6324;
  assign n6673 = ~n6333 & ~n6336;
  assign n6674 = n6672 & n6673;
  assign n6675 = ~n6327 & ~n6480;
  assign n6676 = ~n6318 & ~n6474;
  assign n6677 = n6675 & n6676;
  assign n6678 = n6674 & n6677;
  assign n6679 = ~x244 & x572;
  assign n6680 = ~x247 & x527;
  assign n6681 = ~n6679 & ~n6680;
  assign n6682 = ~n6483 & n6681;
  assign n6683 = x247 & ~x527;
  assign n6684 = x233 & ~n6683;
  assign n6685 = ~n6468 & n6684;
  assign n6686 = n6682 & n6685;
  assign n6687 = n6678 & n6686;
  assign n6688 = x244 & ~x572;
  assign n6689 = ~n6339 & ~n6688;
  assign n6690 = n6687 & n6689;
  assign n6691 = ~n6444 & ~n6465;
  assign n6692 = ~n6429 & ~n6441;
  assign n6693 = n6691 & n6692;
  assign n6694 = ~n6345 & ~n6459;
  assign n6695 = ~n6243 & n6462;
  assign n6696 = n6694 & n6695;
  assign n6697 = n6693 & n6696;
  assign n6698 = ~x249 & x482;
  assign n6699 = ~x233 & ~n6698;
  assign n6700 = ~n6435 & n6699;
  assign n6701 = ~n6342 & ~n6447;
  assign n6702 = n6700 & n6701;
  assign n6703 = n6697 & n6702;
  assign n6704 = x249 & ~x482;
  assign n6705 = ~n6417 & ~n6704;
  assign n6706 = n6703 & n6705;
  assign n6707 = ~n6690 & ~n6706;
  assign n6708 = ~x237 & n6707;
  assign n6709 = n6671 & ~n6708;
  assign n6710 = ~n6636 & ~n6709;
  assign n6711 = ~x806 & x990;
  assign n6712 = x600 & n6711;
  assign n6713 = n6712 ^ x594;
  assign n6714 = ~x332 & n6713;
  assign n6715 = x605 & ~x806;
  assign n6716 = n6098 & n6715;
  assign n6717 = n6716 ^ x595;
  assign n6718 = ~x332 & n6717;
  assign n6719 = n6096 & n6711;
  assign n6720 = x595 & x597;
  assign n6721 = n6719 & n6720;
  assign n6722 = n6721 ^ x596;
  assign n6723 = ~x332 & n6722;
  assign n6724 = n6719 ^ x597;
  assign n6725 = ~x332 & n6724;
  assign n6726 = ~x882 & n1518;
  assign n6727 = x947 & n6726;
  assign n6728 = x598 & ~n6727;
  assign n6729 = x740 & x780;
  assign n6730 = n2172 & n6729;
  assign n6731 = ~n6728 & ~n6730;
  assign n6732 = x596 & n6721;
  assign n6733 = n6732 ^ x599;
  assign n6734 = ~x332 & n6733;
  assign n6735 = n6711 ^ x600;
  assign n6736 = ~x332 & n6735;
  assign n6737 = ~x601 & x806;
  assign n6738 = ~x332 & ~n6737;
  assign n6739 = ~x806 & ~x989;
  assign n6740 = n6738 & ~n6739;
  assign n6741 = n4234 ^ x602;
  assign n6742 = x230 & n6741;
  assign n6743 = n6742 ^ x602;
  assign n6744 = x832 & ~x980;
  assign n6745 = x1060 & n6744;
  assign n6746 = x1038 & ~x1061;
  assign n6747 = n6745 & n6746;
  assign n6748 = x952 & n6747;
  assign n6749 = x603 & ~n6748;
  assign n6750 = ~x966 & ~n6749;
  assign n6751 = x1100 & n6748;
  assign n6752 = n6750 & ~n6751;
  assign n6753 = ~x871 & x966;
  assign n6754 = ~x872 & n6753;
  assign n6755 = ~n6752 & ~n6754;
  assign n6756 = x823 & n2174;
  assign n6757 = ~x299 & x983;
  assign n6758 = x907 & n6757;
  assign n6759 = x604 & ~n6758;
  assign n6760 = n6759 ^ x779;
  assign n6761 = ~n6756 & ~n6760;
  assign n6762 = n6761 ^ x779;
  assign n6763 = x806 ^ x605;
  assign n6764 = ~x332 & ~n6763;
  assign n6765 = ~x606 & ~n6748;
  assign n6766 = ~x966 & ~n6765;
  assign n6767 = ~x1104 & n6748;
  assign n6768 = n6766 & ~n6767;
  assign n6769 = x837 & x966;
  assign n6770 = ~n6768 & ~n6769;
  assign n6771 = ~x1107 & n6748;
  assign n6772 = ~x966 & ~n6771;
  assign n6773 = ~x607 & ~n6748;
  assign n6774 = n6772 & ~n6773;
  assign n6775 = ~x1116 & n6748;
  assign n6776 = ~x966 & ~n6775;
  assign n6777 = ~x608 & ~n6748;
  assign n6778 = n6776 & ~n6777;
  assign n6779 = ~x1118 & n6748;
  assign n6780 = ~x966 & ~n6779;
  assign n6781 = ~x609 & ~n6748;
  assign n6782 = n6780 & ~n6781;
  assign n6783 = ~x1113 & n6748;
  assign n6784 = ~x966 & ~n6783;
  assign n6785 = ~x610 & ~n6748;
  assign n6786 = n6784 & ~n6785;
  assign n6787 = ~x1114 & n6748;
  assign n6788 = ~x966 & ~n6787;
  assign n6789 = ~x611 & ~n6748;
  assign n6790 = n6788 & ~n6789;
  assign n6791 = ~x1111 & n6748;
  assign n6792 = ~x966 & ~n6791;
  assign n6793 = ~x612 & ~n6748;
  assign n6794 = n6792 & ~n6793;
  assign n6795 = ~x1115 & n6748;
  assign n6796 = ~x966 & ~n6795;
  assign n6797 = ~x613 & ~n6748;
  assign n6798 = n6796 & ~n6797;
  assign n6799 = x1102 ^ x614;
  assign n6800 = n6748 & n6799;
  assign n6801 = n6800 ^ x614;
  assign n6802 = n6801 ^ x871;
  assign n6803 = ~x966 & n6802;
  assign n6804 = n6803 ^ x871;
  assign n6805 = x907 & n6726;
  assign n6806 = ~x615 & ~n6805;
  assign n6807 = x779 & x797;
  assign n6808 = n2175 & n6807;
  assign n6809 = ~n6806 & ~n6808;
  assign n6810 = ~x616 & ~n6748;
  assign n6811 = ~x966 & ~n6810;
  assign n6812 = ~x1101 & n6748;
  assign n6813 = n6811 & ~n6812;
  assign n6814 = x872 & x966;
  assign n6815 = ~n6813 & ~n6814;
  assign n6816 = ~x617 & ~n6748;
  assign n6817 = ~x966 & ~n6816;
  assign n6818 = ~x1105 & n6748;
  assign n6819 = n6817 & ~n6818;
  assign n6820 = x850 & x966;
  assign n6821 = ~n6819 & ~n6820;
  assign n6822 = ~x1117 & n6748;
  assign n6823 = ~x966 & ~n6822;
  assign n6824 = ~x618 & ~n6748;
  assign n6825 = n6823 & ~n6824;
  assign n6826 = ~x1122 & n6748;
  assign n6827 = ~x966 & ~n6826;
  assign n6828 = ~x619 & ~n6748;
  assign n6829 = n6827 & ~n6828;
  assign n6830 = ~x1112 & n6748;
  assign n6831 = ~x966 & ~n6830;
  assign n6832 = ~x620 & ~n6748;
  assign n6833 = n6831 & ~n6832;
  assign n6834 = ~x1108 & n6748;
  assign n6835 = ~x966 & ~n6834;
  assign n6836 = ~x621 & ~n6748;
  assign n6837 = n6835 & ~n6836;
  assign n6838 = ~x1109 & n6748;
  assign n6839 = ~x966 & ~n6838;
  assign n6840 = ~x622 & ~n6748;
  assign n6841 = n6839 & ~n6840;
  assign n6842 = ~x1106 & n6748;
  assign n6843 = ~x966 & ~n6842;
  assign n6844 = ~x623 & ~n6748;
  assign n6845 = n6843 & ~n6844;
  assign n6846 = x831 & n2171;
  assign n6847 = x947 & n6757;
  assign n6848 = x624 & ~n6847;
  assign n6849 = n6848 ^ x780;
  assign n6850 = ~n6846 & ~n6849;
  assign n6851 = n6850 ^ x780;
  assign n6852 = x1066 & x1088;
  assign n6853 = ~x973 & ~x1054;
  assign n6854 = n6852 & n6853;
  assign n6855 = x832 & n6854;
  assign n6856 = ~x953 & n6855;
  assign n6857 = ~x1116 & n6856;
  assign n6858 = ~x962 & ~n6857;
  assign n6859 = ~x625 & ~n6856;
  assign n6860 = n6858 & ~n6859;
  assign n6861 = ~x1121 & n6748;
  assign n6862 = ~x966 & ~n6861;
  assign n6863 = ~x626 & ~n6748;
  assign n6864 = n6862 & ~n6863;
  assign n6865 = ~x1117 & n6856;
  assign n6866 = ~x962 & ~n6865;
  assign n6867 = ~x627 & ~n6856;
  assign n6868 = n6866 & ~n6867;
  assign n6869 = ~x1119 & n6856;
  assign n6870 = ~x962 & ~n6869;
  assign n6871 = ~x628 & ~n6856;
  assign n6872 = n6870 & ~n6871;
  assign n6873 = ~x1119 & n6748;
  assign n6874 = ~x966 & ~n6873;
  assign n6875 = ~x629 & ~n6748;
  assign n6876 = n6874 & ~n6875;
  assign n6877 = ~x1120 & n6748;
  assign n6878 = ~x966 & ~n6877;
  assign n6879 = ~x630 & ~n6748;
  assign n6880 = n6878 & ~n6879;
  assign n6881 = ~x1113 & n6856;
  assign n6882 = ~x962 & ~n6881;
  assign n6883 = x631 & ~n6856;
  assign n6884 = n6882 & ~n6883;
  assign n6885 = ~x1115 & n6856;
  assign n6886 = ~x962 & ~n6885;
  assign n6887 = x632 & ~n6856;
  assign n6888 = n6886 & ~n6887;
  assign n6889 = ~x1110 & n6748;
  assign n6890 = ~x966 & ~n6889;
  assign n6891 = ~x633 & ~n6748;
  assign n6892 = n6890 & ~n6891;
  assign n6893 = ~x1110 & n6856;
  assign n6894 = ~x962 & ~n6893;
  assign n6895 = ~x634 & ~n6856;
  assign n6896 = n6894 & ~n6895;
  assign n6897 = ~x1112 & n6856;
  assign n6898 = ~x962 & ~n6897;
  assign n6899 = x635 & ~n6856;
  assign n6900 = n6898 & ~n6899;
  assign n6901 = ~x1127 & n6748;
  assign n6902 = ~x966 & ~n6901;
  assign n6903 = ~x636 & ~n6748;
  assign n6904 = n6902 & ~n6903;
  assign n6905 = ~x1105 & n6856;
  assign n6906 = ~x962 & ~n6905;
  assign n6907 = ~x637 & ~n6856;
  assign n6908 = n6906 & ~n6907;
  assign n6909 = ~x1107 & n6856;
  assign n6910 = ~x962 & ~n6909;
  assign n6911 = ~x638 & ~n6856;
  assign n6912 = n6910 & ~n6911;
  assign n6913 = ~x1109 & n6856;
  assign n6914 = ~x962 & ~n6913;
  assign n6915 = ~x639 & ~n6856;
  assign n6916 = n6914 & ~n6915;
  assign n6917 = ~x1128 & n6748;
  assign n6918 = ~x966 & ~n6917;
  assign n6919 = ~x640 & ~n6748;
  assign n6920 = n6918 & ~n6919;
  assign n6921 = ~x1121 & n6856;
  assign n6922 = ~x962 & ~n6921;
  assign n6923 = ~x641 & ~n6856;
  assign n6924 = n6922 & ~n6923;
  assign n6925 = ~x1103 & n6748;
  assign n6926 = ~x966 & ~n6925;
  assign n6927 = ~x642 & ~n6748;
  assign n6928 = n6926 & ~n6927;
  assign n6929 = ~x1104 & n6856;
  assign n6930 = ~x962 & ~n6929;
  assign n6931 = ~x643 & ~n6856;
  assign n6932 = n6930 & ~n6931;
  assign n6933 = ~x1123 & n6748;
  assign n6934 = ~x966 & ~n6933;
  assign n6935 = ~x644 & ~n6748;
  assign n6936 = n6934 & ~n6935;
  assign n6937 = ~x1125 & n6748;
  assign n6938 = ~x966 & ~n6937;
  assign n6939 = ~x645 & ~n6748;
  assign n6940 = n6938 & ~n6939;
  assign n6941 = ~x1114 & n6856;
  assign n6942 = ~x962 & ~n6941;
  assign n6943 = x646 & ~n6856;
  assign n6944 = n6942 & ~n6943;
  assign n6945 = ~x1120 & n6856;
  assign n6946 = ~x962 & ~n6945;
  assign n6947 = ~x647 & ~n6856;
  assign n6948 = n6946 & ~n6947;
  assign n6949 = ~x1122 & n6856;
  assign n6950 = ~x962 & ~n6949;
  assign n6951 = ~x648 & ~n6856;
  assign n6952 = n6950 & ~n6951;
  assign n6953 = ~x1126 & n6856;
  assign n6954 = ~x962 & ~n6953;
  assign n6955 = x649 & ~n6856;
  assign n6956 = n6954 & ~n6955;
  assign n6957 = ~x1127 & n6856;
  assign n6958 = ~x962 & ~n6957;
  assign n6959 = x650 & ~n6856;
  assign n6960 = n6958 & ~n6959;
  assign n6961 = ~x1130 & n6748;
  assign n6962 = ~x966 & ~n6961;
  assign n6963 = ~x651 & ~n6748;
  assign n6964 = n6962 & ~n6963;
  assign n6965 = ~x1131 & n6748;
  assign n6966 = ~x966 & ~n6965;
  assign n6967 = ~x652 & ~n6748;
  assign n6968 = n6966 & ~n6967;
  assign n6969 = ~x1129 & n6748;
  assign n6970 = ~x966 & ~n6969;
  assign n6971 = ~x653 & ~n6748;
  assign n6972 = n6970 & ~n6971;
  assign n6973 = ~x1130 & n6856;
  assign n6974 = ~x962 & ~n6973;
  assign n6975 = x654 & ~n6856;
  assign n6976 = n6974 & ~n6975;
  assign n6977 = ~x1124 & n6856;
  assign n6978 = ~x962 & ~n6977;
  assign n6979 = x655 & ~n6856;
  assign n6980 = n6978 & ~n6979;
  assign n6981 = ~x1126 & n6748;
  assign n6982 = ~x966 & ~n6981;
  assign n6983 = ~x656 & ~n6748;
  assign n6984 = n6982 & ~n6983;
  assign n6985 = ~x1131 & n6856;
  assign n6986 = ~x962 & ~n6985;
  assign n6987 = x657 & ~n6856;
  assign n6988 = n6986 & ~n6987;
  assign n6989 = ~x1124 & n6748;
  assign n6990 = ~x966 & ~n6989;
  assign n6991 = ~x658 & ~n6748;
  assign n6992 = n6990 & ~n6991;
  assign n6993 = x266 & x992;
  assign n6994 = ~x280 & n6993;
  assign n6995 = ~x269 & n6994;
  assign n6996 = ~x281 & ~x282;
  assign n6997 = n6995 & n6996;
  assign n6998 = ~x270 & ~x277;
  assign n6999 = ~x264 & n6998;
  assign n7000 = n6997 & n6999;
  assign n7001 = ~x265 & n7000;
  assign n7002 = n7001 ^ x274;
  assign n7003 = ~x1118 & n6856;
  assign n7004 = ~x962 & ~n7003;
  assign n7005 = ~x660 & ~n6856;
  assign n7006 = n7004 & ~n7005;
  assign n7007 = ~x1101 & n6856;
  assign n7008 = ~x962 & ~n7007;
  assign n7009 = ~x661 & ~n6856;
  assign n7010 = n7008 & ~n7009;
  assign n7011 = ~x1102 & n6856;
  assign n7012 = ~x962 & ~n7011;
  assign n7013 = ~x662 & ~n6856;
  assign n7014 = n7012 & ~n7013;
  assign n7015 = x591 & ~x592;
  assign n7016 = x334 & n7015;
  assign n7017 = ~x591 & x592;
  assign n7018 = x365 & n7017;
  assign n7019 = ~n7016 & ~n7018;
  assign n7020 = n3506 & ~n7019;
  assign n7021 = x588 & n2595;
  assign n7022 = x464 & n7021;
  assign n7023 = ~n7020 & ~n7022;
  assign n7024 = n1483 & n7023;
  assign n7025 = ~x588 & ~n2595;
  assign n7026 = n2591 & n7025;
  assign n7027 = x323 & n7026;
  assign n7028 = n7024 & ~n7027;
  assign n7029 = x1065 ^ x257;
  assign n7030 = x199 & n7029;
  assign n7031 = n7030 ^ x257;
  assign n7032 = ~n1483 & ~n7031;
  assign n7033 = n2699 & ~n7032;
  assign n7034 = ~n7028 & n7033;
  assign n7038 = x815 ^ x633;
  assign n7039 = ~x1136 & n7038;
  assign n7040 = n7039 ^ x633;
  assign n7035 = x855 ^ x766;
  assign n7036 = ~x1136 & n7035;
  assign n7037 = n7036 ^ x766;
  assign n7041 = n7040 ^ n7037;
  assign n7042 = x1134 & n7041;
  assign n7043 = n7042 ^ n7040;
  assign n7044 = ~x1135 & ~n7043;
  assign n7045 = x784 ^ x634;
  assign n7046 = ~x1136 & n7045;
  assign n7047 = n7046 ^ x634;
  assign n7048 = ~x1134 & n7047;
  assign n7049 = x1134 & x1136;
  assign n7050 = x700 & n7049;
  assign n7051 = x1135 & ~n7050;
  assign n7052 = ~n7048 & n7051;
  assign n7053 = ~x1137 & ~x1138;
  assign n7054 = ~n2699 & n7053;
  assign n7055 = ~n7052 & n7054;
  assign n7056 = ~n7044 & n7055;
  assign n7057 = ~n7034 & ~n7056;
  assign n7058 = x404 & n7015;
  assign n7059 = x380 & n7017;
  assign n7060 = ~n7058 & ~n7059;
  assign n7061 = n3506 & ~n7060;
  assign n7062 = x429 & n7021;
  assign n7063 = ~n7061 & ~n7062;
  assign n7064 = n1483 & n7063;
  assign n7065 = x355 & n7026;
  assign n7066 = n7064 & ~n7065;
  assign n7067 = x199 & n5564;
  assign n7068 = n7067 ^ x292;
  assign n7069 = ~n1483 & ~n7068;
  assign n7070 = n2699 & ~n7069;
  assign n7071 = ~n7066 & n7070;
  assign n7075 = x811 ^ x614;
  assign n7076 = ~x1136 & n7075;
  assign n7077 = n7076 ^ x614;
  assign n7072 = x872 ^ x772;
  assign n7073 = ~x1136 & n7072;
  assign n7074 = n7073 ^ x772;
  assign n7078 = n7077 ^ n7074;
  assign n7079 = x1134 & n7078;
  assign n7080 = n7079 ^ n7077;
  assign n7081 = ~x1135 & ~n7080;
  assign n7082 = x785 ^ x662;
  assign n7083 = ~x1136 & n7082;
  assign n7084 = n7083 ^ x662;
  assign n7085 = ~x1134 & n7084;
  assign n7086 = x727 & n7049;
  assign n7087 = x1135 & ~n7086;
  assign n7088 = ~n7085 & n7087;
  assign n7089 = n7054 & ~n7088;
  assign n7090 = ~n7081 & n7089;
  assign n7091 = ~n7071 & ~n7090;
  assign n7092 = ~x1108 & n6856;
  assign n7093 = ~x962 & ~n7092;
  assign n7094 = ~x665 & ~n6856;
  assign n7095 = n7093 & ~n7094;
  assign n7096 = x456 & n7015;
  assign n7097 = x337 & n7017;
  assign n7098 = ~n7096 & ~n7097;
  assign n7099 = n3506 & ~n7098;
  assign n7100 = x443 & n7021;
  assign n7101 = ~n7099 & ~n7100;
  assign n7102 = n1483 & n7101;
  assign n7103 = x441 & n7026;
  assign n7104 = n7102 & ~n7103;
  assign n7105 = x199 & n5579;
  assign n7106 = n7105 ^ x297;
  assign n7107 = ~n1483 & ~n7106;
  assign n7108 = n2699 & ~n7107;
  assign n7109 = ~n7104 & n7108;
  assign n7110 = x799 ^ x607;
  assign n7111 = ~x1136 & ~n7110;
  assign n7112 = n7111 ^ x607;
  assign n7113 = ~x1134 & n7112;
  assign n7114 = ~x873 & ~x1136;
  assign n7115 = ~x764 & n7049;
  assign n7116 = n7115 ^ x1134;
  assign n7117 = ~n7114 & n7116;
  assign n7118 = ~n7113 & ~n7117;
  assign n7119 = ~x1135 & n7118;
  assign n7120 = x790 ^ x638;
  assign n7121 = ~x1136 & n7120;
  assign n7122 = n7121 ^ x638;
  assign n7123 = ~x1134 & n7122;
  assign n7124 = x691 & n7049;
  assign n7125 = x1135 & ~n7124;
  assign n7126 = ~n7123 & n7125;
  assign n7127 = n7054 & ~n7126;
  assign n7128 = ~n7119 & n7127;
  assign n7129 = ~n7109 & ~n7128;
  assign n7130 = x458 & n7026;
  assign n7131 = x319 & n7015;
  assign n7132 = x338 & n7017;
  assign n7133 = ~n7131 & ~n7132;
  assign n7134 = n3506 & ~n7133;
  assign n7135 = x444 & n7021;
  assign n7136 = ~n7134 & ~n7135;
  assign n7137 = ~n7130 & n7136;
  assign n7138 = n1483 & n7137;
  assign n7139 = x199 & n5570;
  assign n7140 = n7139 ^ x294;
  assign n7141 = ~n1483 & ~n7140;
  assign n7142 = n2699 & ~n7141;
  assign n7143 = ~n7138 & n7142;
  assign n7144 = x809 ^ x642;
  assign n7145 = ~x1136 & ~n7144;
  assign n7146 = n7145 ^ x642;
  assign n7147 = ~x1134 & n7146;
  assign n7148 = ~x871 & ~x1136;
  assign n7149 = ~x763 & n7049;
  assign n7150 = n7149 ^ x1134;
  assign n7151 = ~n7148 & n7150;
  assign n7152 = ~n7147 & ~n7151;
  assign n7153 = ~x1135 & n7152;
  assign n7154 = x792 ^ x681;
  assign n7155 = ~x1136 & n7154;
  assign n7156 = n7155 ^ x681;
  assign n7157 = ~x1134 & n7156;
  assign n7158 = x699 & n7049;
  assign n7159 = x1135 & ~n7158;
  assign n7160 = ~n7157 & n7159;
  assign n7161 = n7054 & ~n7160;
  assign n7162 = ~n7153 & n7161;
  assign n7163 = ~n7143 & ~n7162;
  assign n7164 = x342 & n7026;
  assign n7165 = x390 & n7015;
  assign n7166 = x363 & n7017;
  assign n7167 = ~n7165 & ~n7166;
  assign n7168 = n3506 & ~n7167;
  assign n7169 = x414 & n7021;
  assign n7170 = ~n7168 & ~n7169;
  assign n7171 = ~n7164 & n7170;
  assign n7172 = n1483 & n7171;
  assign n7173 = x199 & n5561;
  assign n7174 = n7173 ^ x291;
  assign n7175 = ~n1483 & ~n7174;
  assign n7176 = n2699 & ~n7175;
  assign n7177 = ~n7172 & n7176;
  assign n7181 = x981 ^ x603;
  assign n7182 = ~x1136 & n7181;
  assign n7183 = n7182 ^ x603;
  assign n7178 = x837 ^ x759;
  assign n7179 = ~x1136 & n7178;
  assign n7180 = n7179 ^ x759;
  assign n7184 = n7183 ^ n7180;
  assign n7185 = x1134 & n7184;
  assign n7186 = n7185 ^ n7183;
  assign n7187 = ~x1135 & ~n7186;
  assign n7188 = x778 ^ x680;
  assign n7189 = ~x1136 & n7188;
  assign n7190 = n7189 ^ x680;
  assign n7191 = ~x1134 & n7190;
  assign n7192 = x696 & n7049;
  assign n7193 = x1135 & ~n7192;
  assign n7194 = ~n7191 & n7193;
  assign n7195 = n7054 & ~n7194;
  assign n7196 = ~n7187 & n7195;
  assign n7197 = ~n7177 & ~n7196;
  assign n7198 = ~x1125 & n6856;
  assign n7199 = ~x962 & ~n7198;
  assign n7200 = x669 & ~n6856;
  assign n7201 = n7199 & ~n7200;
  assign n7202 = x723 & x1135;
  assign n7203 = x1134 & ~n7202;
  assign n7204 = x745 & ~x1135;
  assign n7205 = n7203 & ~n7204;
  assign n7206 = ~x612 & ~x1135;
  assign n7207 = ~x1134 & ~n7206;
  assign n7208 = x695 & x1135;
  assign n7209 = n7207 & ~n7208;
  assign n7210 = ~n7205 & ~n7209;
  assign n7211 = x1136 & ~n7210;
  assign n7212 = ~x1135 & ~x1136;
  assign n7213 = x1134 & n7212;
  assign n7214 = x852 & n7213;
  assign n7215 = ~n7211 & ~n7214;
  assign n7216 = n7054 & ~n7215;
  assign n7217 = x415 & n7021;
  assign n7218 = n1483 & ~n7217;
  assign n7219 = x391 & n2594;
  assign n7220 = x364 & ~x590;
  assign n7221 = ~x591 & n7220;
  assign n7222 = ~n7219 & ~n7221;
  assign n7223 = x343 & n2591;
  assign n7224 = n7222 & ~n7223;
  assign n7225 = n7025 & ~n7224;
  assign n7226 = n7218 & ~n7225;
  assign n7227 = x1062 ^ x258;
  assign n7228 = x199 & n7227;
  assign n7229 = n7228 ^ x258;
  assign n7230 = ~n1483 & ~n7229;
  assign n7231 = n2699 & ~n7230;
  assign n7232 = ~n7226 & n7231;
  assign n7233 = ~n7216 & ~n7232;
  assign n7234 = x333 & n7015;
  assign n7235 = x447 & n7017;
  assign n7236 = ~n7234 & ~n7235;
  assign n7237 = n3506 & ~n7236;
  assign n7238 = x453 & n7021;
  assign n7239 = ~n7237 & ~n7238;
  assign n7240 = n1483 & n7239;
  assign n7241 = x327 & n7026;
  assign n7242 = n7240 & ~n7241;
  assign n7243 = x1040 ^ x261;
  assign n7244 = x199 & n7243;
  assign n7245 = n7244 ^ x261;
  assign n7246 = ~n1483 & ~n7245;
  assign n7247 = n2699 & ~n7246;
  assign n7248 = ~n7242 & n7247;
  assign n7249 = x724 & x1135;
  assign n7250 = x1134 & ~n7249;
  assign n7251 = x741 & ~x1135;
  assign n7252 = n7250 & ~n7251;
  assign n7253 = ~x611 & ~x1135;
  assign n7254 = ~x1134 & ~n7253;
  assign n7255 = x646 & x1135;
  assign n7256 = n7254 & ~n7255;
  assign n7257 = ~n7252 & ~n7256;
  assign n7258 = x1136 & ~n7257;
  assign n7259 = x865 & n7213;
  assign n7260 = ~n7258 & ~n7259;
  assign n7261 = n7054 & ~n7260;
  assign n7262 = ~n7248 & ~n7261;
  assign n7263 = x320 & n7026;
  assign n7264 = x397 & n7015;
  assign n7265 = x372 & n7017;
  assign n7266 = ~n7264 & ~n7265;
  assign n7267 = n3506 & ~n7266;
  assign n7268 = x422 & n7021;
  assign n7269 = ~n7267 & ~n7268;
  assign n7270 = ~n7263 & n7269;
  assign n7271 = n1483 & n7270;
  assign n7272 = x199 & n5558;
  assign n7273 = n7272 ^ x290;
  assign n7274 = ~n1483 & ~n7273;
  assign n7275 = n2699 & ~n7274;
  assign n7276 = ~n7271 & n7275;
  assign n7280 = x808 ^ x616;
  assign n7281 = ~x1136 & n7280;
  assign n7282 = n7281 ^ x616;
  assign n7277 = x850 ^ x758;
  assign n7278 = ~x1136 & n7277;
  assign n7279 = n7278 ^ x758;
  assign n7283 = n7282 ^ n7279;
  assign n7284 = x1134 & n7283;
  assign n7285 = n7284 ^ n7282;
  assign n7286 = ~x1135 & ~n7285;
  assign n7287 = x781 ^ x661;
  assign n7288 = ~x1136 & n7287;
  assign n7289 = n7288 ^ x661;
  assign n7290 = ~x1134 & n7289;
  assign n7291 = x736 & n7049;
  assign n7292 = x1135 & ~n7291;
  assign n7293 = ~n7290 & n7292;
  assign n7294 = n7054 & ~n7293;
  assign n7295 = ~n7286 & n7294;
  assign n7296 = ~n7276 & ~n7295;
  assign n7297 = x411 & n7015;
  assign n7298 = x387 & n7017;
  assign n7299 = ~n7297 & ~n7298;
  assign n7300 = n3506 & ~n7299;
  assign n7301 = x435 & n7021;
  assign n7302 = ~n7300 & ~n7301;
  assign n7303 = n1483 & n7302;
  assign n7304 = x452 & n7026;
  assign n7305 = n7303 & ~n7304;
  assign n7306 = x199 & n5573;
  assign n7307 = n7306 ^ x295;
  assign n7308 = ~n1483 & ~n7307;
  assign n7309 = n2699 & ~n7308;
  assign n7310 = ~n7305 & n7309;
  assign n7314 = x866 ^ x749;
  assign n7315 = ~x1136 & n7314;
  assign n7316 = n7315 ^ x749;
  assign n7311 = x814 ^ x617;
  assign n7312 = ~x1136 & ~n7311;
  assign n7313 = n7312 ^ x617;
  assign n7317 = n7316 ^ n7313;
  assign n7318 = ~x1134 & n7317;
  assign n7319 = n7318 ^ n7316;
  assign n7320 = ~x1135 & ~n7319;
  assign n7321 = x788 ^ x637;
  assign n7322 = ~x1136 & n7321;
  assign n7323 = n7322 ^ x637;
  assign n7324 = ~x1134 & n7323;
  assign n7325 = x706 & n7049;
  assign n7326 = x1135 & ~n7325;
  assign n7327 = ~n7324 & n7326;
  assign n7328 = n7054 & ~n7327;
  assign n7329 = ~n7320 & n7328;
  assign n7330 = ~n7310 & ~n7329;
  assign n7331 = x362 & n7026;
  assign n7332 = x463 & n7015;
  assign n7333 = x336 & n7017;
  assign n7334 = ~n7332 & ~n7333;
  assign n7335 = n3506 & ~n7334;
  assign n7336 = x437 & n7021;
  assign n7337 = ~n7335 & ~n7336;
  assign n7338 = ~n7331 & n7337;
  assign n7339 = n1483 & n7338;
  assign n7340 = x1070 ^ x256;
  assign n7341 = x199 & n7340;
  assign n7342 = n7341 ^ x256;
  assign n7343 = ~n1483 & ~n7342;
  assign n7344 = n2699 & ~n7343;
  assign n7345 = ~n7339 & n7344;
  assign n7349 = x804 ^ x622;
  assign n7350 = ~x1136 & n7349;
  assign n7351 = n7350 ^ x622;
  assign n7346 = x859 ^ x743;
  assign n7347 = ~x1136 & n7346;
  assign n7348 = n7347 ^ x743;
  assign n7352 = n7351 ^ n7348;
  assign n7353 = x1134 & n7352;
  assign n7354 = n7353 ^ n7351;
  assign n7355 = ~x1135 & ~n7354;
  assign n7356 = x783 ^ x639;
  assign n7357 = ~x1136 & n7356;
  assign n7358 = n7357 ^ x639;
  assign n7359 = ~x1134 & n7358;
  assign n7360 = x735 & n7049;
  assign n7361 = x1135 & ~n7360;
  assign n7362 = ~n7359 & n7361;
  assign n7363 = n7054 & ~n7362;
  assign n7364 = ~n7355 & n7363;
  assign n7365 = ~n7345 & ~n7364;
  assign n7366 = x412 & n7015;
  assign n7367 = x388 & n7017;
  assign n7368 = ~n7366 & ~n7367;
  assign n7369 = n3506 & ~n7368;
  assign n7370 = x436 & n7021;
  assign n7371 = ~n7369 & ~n7370;
  assign n7372 = n1483 & n7371;
  assign n7373 = x455 & n7026;
  assign n7374 = n7372 & ~n7373;
  assign n7375 = x199 & n5576;
  assign n7376 = n7375 ^ x296;
  assign n7377 = ~n1483 & ~n7376;
  assign n7378 = n2699 & ~n7377;
  assign n7379 = ~n7374 & n7378;
  assign n7380 = x803 ^ x623;
  assign n7381 = ~x1136 & ~n7380;
  assign n7382 = n7381 ^ x623;
  assign n7383 = ~x1134 & n7382;
  assign n7384 = ~x876 & ~x1136;
  assign n7385 = ~x748 & n7049;
  assign n7386 = n7385 ^ x1134;
  assign n7387 = ~n7384 & n7386;
  assign n7388 = ~n7383 & ~n7387;
  assign n7389 = ~x1135 & n7388;
  assign n7390 = x789 ^ x710;
  assign n7391 = ~x1136 & n7390;
  assign n7392 = n7391 ^ x710;
  assign n7393 = ~x1134 & n7392;
  assign n7394 = x730 & n7049;
  assign n7395 = x1135 & ~n7394;
  assign n7396 = ~n7393 & n7395;
  assign n7397 = n7054 & ~n7396;
  assign n7398 = ~n7389 & n7397;
  assign n7399 = ~n7379 & ~n7398;
  assign n7400 = x361 & n7026;
  assign n7401 = x410 & n7015;
  assign n7402 = x386 & n7017;
  assign n7403 = ~n7401 & ~n7402;
  assign n7404 = n3506 & ~n7403;
  assign n7405 = x434 & n7021;
  assign n7406 = ~n7404 & ~n7405;
  assign n7407 = ~n7400 & n7406;
  assign n7408 = n1483 & n7407;
  assign n7409 = x199 & n5567;
  assign n7410 = n7409 ^ x293;
  assign n7411 = ~n1483 & ~n7410;
  assign n7412 = n2699 & ~n7411;
  assign n7413 = ~n7408 & n7412;
  assign n7417 = x881 ^ x746;
  assign n7418 = ~x1136 & n7417;
  assign n7419 = n7418 ^ x746;
  assign n7414 = x812 ^ x606;
  assign n7415 = ~x1136 & ~n7414;
  assign n7416 = n7415 ^ x606;
  assign n7420 = n7419 ^ n7416;
  assign n7421 = ~x1134 & n7420;
  assign n7422 = n7421 ^ n7419;
  assign n7423 = ~x1135 & ~n7422;
  assign n7424 = x787 ^ x643;
  assign n7425 = ~x1136 & n7424;
  assign n7426 = n7425 ^ x643;
  assign n7427 = ~x1134 & n7426;
  assign n7428 = x729 & n7049;
  assign n7429 = x1135 & ~n7428;
  assign n7430 = ~n7427 & n7429;
  assign n7431 = n7054 & ~n7430;
  assign n7432 = ~n7423 & n7431;
  assign n7433 = ~n7413 & ~n7432;
  assign n7434 = x344 & n7026;
  assign n7435 = x335 & n7015;
  assign n7436 = x366 & n7017;
  assign n7437 = ~n7435 & ~n7436;
  assign n7438 = n3506 & ~n7437;
  assign n7439 = x416 & n7021;
  assign n7440 = ~n7438 & ~n7439;
  assign n7441 = ~n7434 & n7440;
  assign n7442 = n1483 & n7441;
  assign n7443 = x1069 ^ x259;
  assign n7444 = x199 & n7443;
  assign n7445 = n7444 ^ x259;
  assign n7446 = ~n1483 & ~n7445;
  assign n7447 = n2699 & ~n7446;
  assign n7448 = ~n7442 & n7447;
  assign n7449 = x742 ^ x704;
  assign n7450 = ~x1135 & n7449;
  assign n7451 = n7450 ^ x704;
  assign n7452 = x1134 & n7451;
  assign n7453 = x1136 & ~n7452;
  assign n7454 = x635 ^ x620;
  assign n7455 = x1135 & ~n7454;
  assign n7456 = n7455 ^ x620;
  assign n7457 = ~x1134 & ~n7456;
  assign n7458 = n7453 & ~n7457;
  assign n7459 = x870 & n7213;
  assign n7460 = ~n7458 & ~n7459;
  assign n7461 = n7054 & ~n7460;
  assign n7462 = ~n7448 & ~n7461;
  assign n7463 = x688 & x1135;
  assign n7464 = x1134 & ~n7463;
  assign n7465 = x760 & ~x1135;
  assign n7466 = n7464 & ~n7465;
  assign n7467 = ~x613 & ~x1135;
  assign n7468 = ~x1134 & ~n7467;
  assign n7469 = x632 & x1135;
  assign n7470 = n7468 & ~n7469;
  assign n7471 = ~n7466 & ~n7470;
  assign n7472 = x1136 & ~n7471;
  assign n7473 = x856 & n7213;
  assign n7474 = ~n7472 & ~n7473;
  assign n7475 = n7054 & ~n7474;
  assign n7476 = x393 & n2594;
  assign n7477 = x346 & n2591;
  assign n7478 = ~n7476 & ~n7477;
  assign n7479 = x368 & ~x590;
  assign n7480 = ~x591 & n7479;
  assign n7481 = n7478 & ~n7480;
  assign n7482 = n7025 & ~n7481;
  assign n7483 = x418 & n7021;
  assign n7484 = n1483 & ~n7483;
  assign n7485 = ~n7482 & n7484;
  assign n7486 = x1067 ^ x260;
  assign n7487 = x199 & n7486;
  assign n7488 = n7487 ^ x260;
  assign n7489 = ~n1483 & ~n7488;
  assign n7490 = n2699 & ~n7489;
  assign n7491 = ~n7485 & n7490;
  assign n7492 = ~n7475 & ~n7491;
  assign n7493 = x413 & n7015;
  assign n7494 = x389 & n7017;
  assign n7495 = ~n7493 & ~n7494;
  assign n7496 = n3506 & ~n7495;
  assign n7497 = x438 & n7021;
  assign n7498 = ~n7496 & ~n7497;
  assign n7499 = n1483 & n7498;
  assign n7500 = x450 & n7026;
  assign n7501 = n7499 & ~n7500;
  assign n7502 = x1036 ^ x255;
  assign n7503 = x199 & n7502;
  assign n7504 = n7503 ^ x255;
  assign n7505 = ~n1483 & ~n7504;
  assign n7506 = n2699 & ~n7505;
  assign n7507 = ~n7501 & n7506;
  assign n7511 = x810 ^ x621;
  assign n7512 = ~x1136 & n7511;
  assign n7513 = n7512 ^ x621;
  assign n7508 = x874 ^ x739;
  assign n7509 = ~x1136 & n7508;
  assign n7510 = n7509 ^ x739;
  assign n7514 = n7513 ^ n7510;
  assign n7515 = x1134 & n7514;
  assign n7516 = n7515 ^ n7513;
  assign n7517 = ~x1135 & ~n7516;
  assign n7518 = x791 ^ x665;
  assign n7519 = ~x1136 & n7518;
  assign n7520 = n7519 ^ x665;
  assign n7521 = ~x1134 & n7520;
  assign n7522 = x690 & n7049;
  assign n7523 = x1135 & ~n7522;
  assign n7524 = ~n7521 & n7523;
  assign n7525 = n7054 & ~n7524;
  assign n7526 = ~n7517 & n7525;
  assign n7527 = ~n7507 & ~n7526;
  assign n7528 = ~x1100 & n6856;
  assign n7529 = ~x962 & ~n7528;
  assign n7530 = ~x680 & ~n6856;
  assign n7531 = n7529 & ~n7530;
  assign n7532 = ~x1103 & n6856;
  assign n7533 = ~x962 & ~n7532;
  assign n7534 = ~x681 & ~n6856;
  assign n7535 = n7533 & ~n7534;
  assign n7536 = x392 & n7015;
  assign n7537 = x367 & n7017;
  assign n7538 = ~n7536 & ~n7537;
  assign n7539 = n3506 & ~n7538;
  assign n7540 = x417 & n7021;
  assign n7541 = ~n7539 & ~n7540;
  assign n7542 = n1483 & n7541;
  assign n7543 = x345 & n7026;
  assign n7544 = n7542 & ~n7543;
  assign n7545 = x1039 ^ x251;
  assign n7546 = x199 & n7545;
  assign n7547 = n7546 ^ x251;
  assign n7548 = ~n1483 & ~n7547;
  assign n7549 = n2699 & ~n7548;
  assign n7550 = ~n7544 & n7549;
  assign n7551 = x686 & x1135;
  assign n7552 = x1134 & ~n7551;
  assign n7553 = x757 & ~x1135;
  assign n7554 = n7552 & ~n7553;
  assign n7555 = ~x610 & ~x1135;
  assign n7556 = ~x1134 & ~n7555;
  assign n7557 = x631 & x1135;
  assign n7558 = n7556 & ~n7557;
  assign n7559 = ~n7554 & ~n7558;
  assign n7560 = x1136 & ~n7559;
  assign n7561 = x848 & n7213;
  assign n7562 = ~n7560 & ~n7561;
  assign n7563 = n7054 & ~n7562;
  assign n7564 = ~n7550 & ~n7563;
  assign n7565 = x953 & n6855;
  assign n7566 = ~x1130 & n7565;
  assign n7567 = ~x962 & ~n7566;
  assign n7568 = x684 & ~n7565;
  assign n7569 = n7567 & ~n7568;
  assign n7570 = x406 & n7015;
  assign n7571 = x382 & n7017;
  assign n7572 = ~n7570 & ~n7571;
  assign n7573 = n3506 & ~n7572;
  assign n7574 = x430 & n7021;
  assign n7575 = ~n7573 & ~n7574;
  assign n7576 = n1483 & n7575;
  assign n7577 = x357 & n7026;
  assign n7578 = n7576 & ~n7577;
  assign n7579 = ~x199 & n5290;
  assign n7580 = x199 & x1076;
  assign n7581 = ~n1483 & ~n7580;
  assign n7582 = ~n7579 & n7581;
  assign n7583 = n2699 & ~n7582;
  assign n7584 = ~n7578 & n7583;
  assign n7585 = x728 & x1135;
  assign n7586 = x1134 & ~n7585;
  assign n7587 = x744 & ~x1135;
  assign n7588 = n7586 & ~n7587;
  assign n7589 = ~x652 & ~x1135;
  assign n7590 = ~x1134 & ~n7589;
  assign n7591 = x657 & x1135;
  assign n7592 = n7590 & ~n7591;
  assign n7593 = ~n7588 & ~n7592;
  assign n7594 = x1136 & ~n7593;
  assign n7595 = ~x813 & ~x1134;
  assign n7596 = n7212 & ~n7595;
  assign n7597 = ~x860 & x1134;
  assign n7598 = n7596 & ~n7597;
  assign n7599 = ~n7594 & ~n7598;
  assign n7600 = n7054 & ~n7599;
  assign n7601 = ~n7584 & ~n7600;
  assign n7602 = ~x1113 & n7565;
  assign n7603 = ~x962 & ~n7602;
  assign n7604 = x686 & ~n7565;
  assign n7605 = n7603 & ~n7604;
  assign n7606 = ~x1127 & n7565;
  assign n7607 = ~x962 & ~n7606;
  assign n7608 = ~x687 & ~n7565;
  assign n7609 = n7607 & ~n7608;
  assign n7610 = ~x1115 & n7565;
  assign n7611 = ~x962 & ~n7610;
  assign n7612 = x688 & ~n7565;
  assign n7613 = n7611 & ~n7612;
  assign n7614 = x351 & n7026;
  assign n7615 = x401 & n7015;
  assign n7616 = x376 & n7017;
  assign n7617 = ~n7615 & ~n7616;
  assign n7618 = n3506 & ~n7617;
  assign n7619 = x426 & n7021;
  assign n7620 = ~n7618 & ~n7619;
  assign n7621 = ~n7614 & n7620;
  assign n7622 = n1483 & n7621;
  assign n7623 = ~x199 & n5260;
  assign n7624 = x199 & x1079;
  assign n7625 = ~n1483 & ~n7624;
  assign n7626 = ~n7623 & n7625;
  assign n7627 = n2699 & ~n7626;
  assign n7628 = ~n7622 & n7627;
  assign n7632 = x752 ^ x703;
  assign n7633 = ~x1135 & ~n7632;
  assign n7634 = n7633 ^ x703;
  assign n7629 = x658 ^ x655;
  assign n7630 = ~x1135 & ~n7629;
  assign n7631 = n7630 ^ x655;
  assign n7635 = n7634 ^ n7631;
  assign n7636 = ~x1134 & ~n7635;
  assign n7637 = n7636 ^ n7634;
  assign n7638 = x1136 & n7637;
  assign n7639 = ~x798 & ~x1134;
  assign n7640 = n7212 & ~n7639;
  assign n7641 = ~x843 & x1134;
  assign n7642 = n7640 & ~n7641;
  assign n7643 = ~n7638 & ~n7642;
  assign n7644 = n7054 & ~n7643;
  assign n7645 = ~n7628 & ~n7644;
  assign n7646 = ~x1108 & n7565;
  assign n7647 = ~x962 & ~n7646;
  assign n7648 = ~x690 & ~n7565;
  assign n7649 = n7647 & ~n7648;
  assign n7650 = ~x1107 & n7565;
  assign n7651 = ~x962 & ~n7650;
  assign n7652 = ~x691 & ~n7565;
  assign n7653 = n7651 & ~n7652;
  assign n7654 = x402 & n7015;
  assign n7655 = x317 & n7017;
  assign n7656 = ~n7654 & ~n7655;
  assign n7657 = n3506 & ~n7656;
  assign n7658 = x427 & n7021;
  assign n7659 = ~n7657 & ~n7658;
  assign n7660 = n1483 & n7659;
  assign n7661 = x352 & n7026;
  assign n7662 = n7660 & ~n7661;
  assign n7663 = ~x199 & n5272;
  assign n7664 = x199 & x1078;
  assign n7665 = ~n1483 & ~n7664;
  assign n7666 = ~n7663 & n7665;
  assign n7667 = n2699 & ~n7666;
  assign n7668 = ~n7662 & n7667;
  assign n7672 = x770 ^ x726;
  assign n7673 = ~x1135 & ~n7672;
  assign n7674 = n7673 ^ x726;
  assign n7669 = x656 ^ x649;
  assign n7670 = ~x1135 & ~n7669;
  assign n7671 = n7670 ^ x649;
  assign n7675 = n7674 ^ n7671;
  assign n7676 = ~x1134 & ~n7675;
  assign n7677 = n7676 ^ n7674;
  assign n7678 = x1136 & n7677;
  assign n7679 = ~x801 & ~x1134;
  assign n7680 = n7212 & ~n7679;
  assign n7681 = ~x844 & x1134;
  assign n7682 = n7680 & ~n7681;
  assign n7683 = ~n7678 & ~n7682;
  assign n7684 = n7054 & ~n7683;
  assign n7685 = ~n7668 & ~n7684;
  assign n7686 = ~x1129 & n6856;
  assign n7687 = ~x962 & ~n7686;
  assign n7688 = x693 & ~n6856;
  assign n7689 = n7687 & ~n7688;
  assign n7690 = ~x1128 & n7565;
  assign n7691 = ~x962 & ~n7690;
  assign n7692 = x694 & ~n7565;
  assign n7693 = n7691 & ~n7692;
  assign n7694 = ~x1111 & n6856;
  assign n7695 = ~x962 & ~n7694;
  assign n7696 = x695 & ~n6856;
  assign n7697 = n7695 & ~n7696;
  assign n7698 = ~x1100 & n7565;
  assign n7699 = ~x962 & ~n7698;
  assign n7700 = ~x696 & ~n7565;
  assign n7701 = n7699 & ~n7700;
  assign n7702 = ~x1129 & n7565;
  assign n7703 = ~x962 & ~n7702;
  assign n7704 = x697 & ~n7565;
  assign n7705 = n7703 & ~n7704;
  assign n7706 = ~x1116 & n7565;
  assign n7707 = ~x962 & ~n7706;
  assign n7708 = x698 & ~n7565;
  assign n7709 = n7707 & ~n7708;
  assign n7710 = ~x1103 & n7565;
  assign n7711 = ~x962 & ~n7710;
  assign n7712 = ~x699 & ~n7565;
  assign n7713 = n7711 & ~n7712;
  assign n7714 = ~x1110 & n7565;
  assign n7715 = ~x962 & ~n7714;
  assign n7716 = ~x700 & ~n7565;
  assign n7717 = n7715 & ~n7716;
  assign n7718 = ~x1123 & n7565;
  assign n7719 = ~x962 & ~n7718;
  assign n7720 = x701 & ~n7565;
  assign n7721 = n7719 & ~n7720;
  assign n7722 = ~x1117 & n7565;
  assign n7723 = ~x962 & ~n7722;
  assign n7724 = x702 & ~n7565;
  assign n7725 = n7723 & ~n7724;
  assign n7726 = ~x1124 & n7565;
  assign n7727 = ~x962 & ~n7726;
  assign n7728 = ~x703 & ~n7565;
  assign n7729 = n7727 & ~n7728;
  assign n7730 = ~x1112 & n7565;
  assign n7731 = ~x962 & ~n7730;
  assign n7732 = x704 & ~n7565;
  assign n7733 = n7731 & ~n7732;
  assign n7734 = ~x1125 & n7565;
  assign n7735 = ~x962 & ~n7734;
  assign n7736 = ~x705 & ~n7565;
  assign n7737 = n7735 & ~n7736;
  assign n7738 = ~x1105 & n7565;
  assign n7739 = ~x962 & ~n7738;
  assign n7740 = ~x706 & ~n7565;
  assign n7741 = n7739 & ~n7740;
  assign n7742 = x395 & n7015;
  assign n7743 = x370 & n7017;
  assign n7744 = ~n7742 & ~n7743;
  assign n7745 = n3506 & ~n7744;
  assign n7746 = x420 & n7021;
  assign n7747 = ~n7745 & ~n7746;
  assign n7748 = n1483 & n7747;
  assign n7749 = x347 & n7026;
  assign n7750 = n7748 & ~n7749;
  assign n7751 = ~x304 & n3150;
  assign n7752 = x199 & ~x1055;
  assign n7753 = ~n7751 & ~n7752;
  assign n7754 = ~x1048 & n3242;
  assign n7755 = n7753 & ~n7754;
  assign n7756 = ~n1483 & ~n7755;
  assign n7757 = n2699 & ~n7756;
  assign n7758 = ~n7750 & n7757;
  assign n7759 = x753 ^ x702;
  assign n7760 = ~x1135 & n7759;
  assign n7761 = n7760 ^ x702;
  assign n7762 = x1134 & n7761;
  assign n7763 = x1136 & ~n7762;
  assign n7764 = x627 ^ x618;
  assign n7765 = x1135 & n7764;
  assign n7766 = n7765 ^ x618;
  assign n7767 = ~x1134 & ~n7766;
  assign n7768 = n7763 & ~n7767;
  assign n7769 = x847 & n7213;
  assign n7770 = ~n7768 & ~n7769;
  assign n7771 = n7054 & ~n7770;
  assign n7772 = ~n7758 & ~n7771;
  assign n7773 = x321 & n7026;
  assign n7774 = x328 & n7015;
  assign n7775 = x442 & n7017;
  assign n7776 = ~n7774 & ~n7775;
  assign n7777 = n3506 & ~n7776;
  assign n7778 = x459 & n7021;
  assign n7779 = ~n7777 & ~n7778;
  assign n7780 = ~n7773 & n7779;
  assign n7781 = n1483 & n7780;
  assign n7782 = ~x305 & n3150;
  assign n7783 = x199 & ~x1058;
  assign n7784 = ~n7782 & ~n7783;
  assign n7785 = ~x1084 & n3242;
  assign n7786 = n7784 & ~n7785;
  assign n7787 = ~n1483 & ~n7786;
  assign n7788 = n2699 & ~n7787;
  assign n7789 = ~n7781 & n7788;
  assign n7790 = x754 ^ x709;
  assign n7791 = ~x1135 & n7790;
  assign n7792 = n7791 ^ x709;
  assign n7793 = x1134 & n7792;
  assign n7794 = x1136 & ~n7793;
  assign n7795 = x660 ^ x609;
  assign n7796 = x1135 & n7795;
  assign n7797 = n7796 ^ x609;
  assign n7798 = ~x1134 & ~n7797;
  assign n7799 = n7794 & ~n7798;
  assign n7800 = x857 & n7213;
  assign n7801 = ~n7799 & ~n7800;
  assign n7802 = n7054 & ~n7801;
  assign n7803 = ~n7789 & ~n7802;
  assign n7804 = ~x1118 & n7565;
  assign n7805 = ~x962 & ~n7804;
  assign n7806 = x709 & ~n7565;
  assign n7807 = n7805 & ~n7806;
  assign n7808 = ~x1106 & n6856;
  assign n7809 = ~x962 & ~n7808;
  assign n7810 = ~x710 & ~n6856;
  assign n7811 = n7809 & ~n7810;
  assign n7812 = x398 & n7015;
  assign n7813 = x373 & n7017;
  assign n7814 = ~n7812 & ~n7813;
  assign n7815 = n3506 & ~n7814;
  assign n7816 = x423 & n7021;
  assign n7817 = ~n7815 & ~n7816;
  assign n7818 = n1483 & n7817;
  assign n7819 = x348 & n7026;
  assign n7820 = n7818 & ~n7819;
  assign n7821 = ~x306 & n3150;
  assign n7822 = x199 & ~x1087;
  assign n7823 = ~n7821 & ~n7822;
  assign n7824 = ~x1059 & n3242;
  assign n7825 = n7823 & ~n7824;
  assign n7826 = ~n1483 & ~n7825;
  assign n7827 = n2699 & ~n7826;
  assign n7828 = ~n7820 & n7827;
  assign n7829 = x755 ^ x725;
  assign n7830 = ~x1135 & n7829;
  assign n7831 = n7830 ^ x725;
  assign n7832 = x1134 & n7831;
  assign n7833 = x1136 & ~n7832;
  assign n7834 = x647 ^ x630;
  assign n7835 = x1135 & n7834;
  assign n7836 = n7835 ^ x630;
  assign n7837 = ~x1134 & ~n7836;
  assign n7838 = n7833 & ~n7837;
  assign n7839 = x858 & n7213;
  assign n7840 = ~n7838 & ~n7839;
  assign n7841 = n7054 & ~n7840;
  assign n7842 = ~n7828 & ~n7841;
  assign n7843 = x400 & n7015;
  assign n7844 = x374 & n7017;
  assign n7845 = ~n7843 & ~n7844;
  assign n7846 = n3506 & ~n7845;
  assign n7847 = x425 & n7021;
  assign n7848 = ~n7846 & ~n7847;
  assign n7849 = n1483 & n7848;
  assign n7850 = x350 & n7026;
  assign n7851 = n7849 & ~n7850;
  assign n7852 = ~x298 & n3150;
  assign n7853 = x199 & ~x1035;
  assign n7854 = ~n7852 & ~n7853;
  assign n7855 = ~x1044 & n3242;
  assign n7856 = n7854 & ~n7855;
  assign n7857 = ~n1483 & ~n7856;
  assign n7858 = n2699 & ~n7857;
  assign n7859 = ~n7851 & n7858;
  assign n7860 = x751 ^ x701;
  assign n7861 = ~x1135 & n7860;
  assign n7862 = n7861 ^ x701;
  assign n7863 = x1134 & n7862;
  assign n7864 = x1136 & ~n7863;
  assign n7865 = x715 ^ x644;
  assign n7866 = x1135 & n7865;
  assign n7867 = n7866 ^ x644;
  assign n7868 = ~x1134 & ~n7867;
  assign n7869 = n7864 & ~n7868;
  assign n7870 = x842 & n7213;
  assign n7871 = ~n7869 & ~n7870;
  assign n7872 = n7054 & ~n7871;
  assign n7873 = ~n7859 & ~n7872;
  assign n7874 = x396 & n7015;
  assign n7875 = x371 & n7017;
  assign n7876 = ~n7874 & ~n7875;
  assign n7877 = n3506 & ~n7876;
  assign n7878 = x421 & n7021;
  assign n7879 = ~n7877 & ~n7878;
  assign n7880 = n1483 & n7879;
  assign n7881 = x322 & n7026;
  assign n7882 = n7880 & ~n7881;
  assign n7883 = ~x309 & n3150;
  assign n7884 = x199 & ~x1051;
  assign n7885 = ~n7883 & ~n7884;
  assign n7886 = ~x1072 & n3242;
  assign n7887 = n7885 & ~n7886;
  assign n7888 = ~n1483 & ~n7887;
  assign n7889 = n2699 & ~n7888;
  assign n7890 = ~n7882 & n7889;
  assign n7891 = x756 ^ x734;
  assign n7892 = ~x1135 & n7891;
  assign n7893 = n7892 ^ x734;
  assign n7894 = x1134 & n7893;
  assign n7895 = x1136 & ~n7894;
  assign n7896 = x629 ^ x628;
  assign n7897 = ~x1135 & n7896;
  assign n7898 = n7897 ^ x628;
  assign n7899 = ~x1134 & ~n7898;
  assign n7900 = n7895 & ~n7899;
  assign n7901 = x854 & n7213;
  assign n7902 = ~n7900 & ~n7901;
  assign n7903 = n7054 & ~n7902;
  assign n7904 = ~n7890 & ~n7903;
  assign n7905 = x461 & n7026;
  assign n7906 = x326 & n7015;
  assign n7907 = x439 & n7017;
  assign n7908 = ~n7906 & ~n7907;
  assign n7909 = n3506 & ~n7908;
  assign n7910 = x449 & n7021;
  assign n7911 = ~n7909 & ~n7910;
  assign n7912 = ~n7905 & n7911;
  assign n7913 = n1483 & n7912;
  assign n7914 = ~x199 & n5230;
  assign n7915 = x199 & x1057;
  assign n7916 = ~n1483 & ~n7915;
  assign n7917 = ~n7914 & n7916;
  assign n7918 = n2699 & ~n7917;
  assign n7919 = ~n7913 & n7918;
  assign n7920 = x697 & x1135;
  assign n7921 = x1134 & ~n7920;
  assign n7922 = x762 & ~x1135;
  assign n7923 = n7921 & ~n7922;
  assign n7924 = ~x653 & ~x1135;
  assign n7925 = ~x1134 & ~n7924;
  assign n7926 = x693 & x1135;
  assign n7927 = n7925 & ~n7926;
  assign n7928 = ~n7923 & ~n7927;
  assign n7929 = x1136 & ~n7928;
  assign n7930 = ~x816 & ~x1134;
  assign n7931 = n7212 & ~n7930;
  assign n7932 = ~x867 & x1134;
  assign n7933 = n7931 & ~n7932;
  assign n7934 = ~n7929 & ~n7933;
  assign n7935 = n7054 & ~n7934;
  assign n7936 = ~n7919 & ~n7935;
  assign n7937 = ~x1123 & n6856;
  assign n7938 = ~x962 & ~n7937;
  assign n7939 = ~x715 & ~n6856;
  assign n7940 = n7938 & ~n7939;
  assign n7941 = x349 & n7026;
  assign n7942 = x329 & n7015;
  assign n7943 = x440 & n7017;
  assign n7944 = ~n7942 & ~n7943;
  assign n7945 = n3506 & ~n7944;
  assign n7946 = ~n7941 & ~n7945;
  assign n7947 = x454 & n7021;
  assign n7948 = n1483 & ~n7947;
  assign n7949 = n7946 & n7948;
  assign n7950 = ~x1053 & n3242;
  assign n7951 = ~x307 & n3150;
  assign n7952 = ~n7950 & ~n7951;
  assign n7953 = x199 & ~x1043;
  assign n7954 = n7952 & ~n7953;
  assign n7955 = ~n1483 & ~n7954;
  assign n7956 = n2699 & ~n7955;
  assign n7957 = ~n7949 & n7956;
  assign n7958 = x761 ^ x738;
  assign n7959 = ~x1135 & n7958;
  assign n7960 = n7959 ^ x738;
  assign n7961 = x1134 & n7960;
  assign n7962 = x1136 & ~n7961;
  assign n7963 = x641 ^ x626;
  assign n7964 = x1135 & n7963;
  assign n7965 = n7964 ^ x626;
  assign n7966 = ~x1134 & ~n7965;
  assign n7967 = n7962 & ~n7966;
  assign n7968 = x845 & n7213;
  assign n7969 = ~n7967 & ~n7968;
  assign n7970 = n7054 & ~n7969;
  assign n7971 = ~n7957 & ~n7970;
  assign n7972 = x462 & n7026;
  assign n7973 = x318 & n7015;
  assign n7974 = x377 & n7017;
  assign n7975 = ~n7973 & ~n7974;
  assign n7976 = n3506 & ~n7975;
  assign n7977 = x448 & n7021;
  assign n7978 = ~n7976 & ~n7977;
  assign n7979 = ~n7972 & n7978;
  assign n7980 = n1483 & n7979;
  assign n7981 = ~x199 & n5266;
  assign n7982 = x199 & x1074;
  assign n7983 = ~n1483 & ~n7982;
  assign n7984 = ~n7981 & n7983;
  assign n7985 = n2699 & ~n7984;
  assign n7986 = ~n7980 & n7985;
  assign n7987 = x768 ^ x705;
  assign n7988 = ~x1135 & ~n7987;
  assign n7989 = n7988 ^ x705;
  assign n7990 = x1134 & ~n7989;
  assign n7991 = x1136 & ~n7990;
  assign n7992 = x669 ^ x645;
  assign n7993 = x1135 & ~n7992;
  assign n7994 = n7993 ^ x645;
  assign n7995 = ~x1134 & ~n7994;
  assign n7996 = n7991 & ~n7995;
  assign n7997 = ~x800 & ~x1134;
  assign n7998 = n7212 & ~n7997;
  assign n7999 = ~x839 & x1134;
  assign n8000 = n7998 & ~n7999;
  assign n8001 = ~n7996 & ~n8000;
  assign n8002 = n7054 & ~n8001;
  assign n8003 = ~n7986 & ~n8002;
  assign n8004 = x315 & n7026;
  assign n8005 = x419 & n7021;
  assign n8006 = ~n8004 & ~n8005;
  assign n8007 = x394 & n7015;
  assign n8008 = x369 & n7017;
  assign n8009 = ~n8007 & ~n8008;
  assign n8010 = n3506 & ~n8009;
  assign n8011 = n1483 & ~n8010;
  assign n8012 = n8006 & n8011;
  assign n8013 = ~x303 & n3150;
  assign n8014 = x199 & ~x1080;
  assign n8015 = ~n8013 & ~n8014;
  assign n8016 = ~x1049 & n3242;
  assign n8017 = n8015 & ~n8016;
  assign n8018 = ~n1483 & ~n8017;
  assign n8019 = n2699 & ~n8018;
  assign n8020 = ~n8012 & n8019;
  assign n8021 = x767 ^ x698;
  assign n8022 = ~x1135 & n8021;
  assign n8023 = n8022 ^ x698;
  assign n8024 = x1134 & n8023;
  assign n8025 = x1136 & ~n8024;
  assign n8026 = x625 ^ x608;
  assign n8027 = x1135 & n8026;
  assign n8028 = n8027 ^ x608;
  assign n8029 = ~x1134 & ~n8028;
  assign n8030 = n8025 & ~n8029;
  assign n8031 = x853 & n7213;
  assign n8032 = ~n8030 & ~n8031;
  assign n8033 = n7054 & ~n8032;
  assign n8034 = ~n8020 & ~n8033;
  assign n8035 = x353 & n7026;
  assign n8036 = x325 & n7015;
  assign n8037 = x378 & n7017;
  assign n8038 = ~n8036 & ~n8037;
  assign n8039 = n3506 & ~n8038;
  assign n8040 = x451 & n7021;
  assign n8041 = ~n8039 & ~n8040;
  assign n8042 = ~n8035 & n8041;
  assign n8043 = n1483 & n8042;
  assign n8044 = ~x199 & n5278;
  assign n8045 = x199 & x1063;
  assign n8046 = ~n1483 & ~n8045;
  assign n8047 = ~n8044 & n8046;
  assign n8048 = n2699 & ~n8047;
  assign n8049 = ~n8043 & n8048;
  assign n8050 = x774 & ~x1135;
  assign n8051 = x1134 & ~n8050;
  assign n8052 = ~x687 & x1135;
  assign n8053 = n8051 & ~n8052;
  assign n8054 = ~x636 & ~x1135;
  assign n8055 = ~x1134 & ~n8054;
  assign n8056 = x650 & x1135;
  assign n8057 = n8055 & ~n8056;
  assign n8058 = ~n8053 & ~n8057;
  assign n8059 = x1136 & ~n8058;
  assign n8060 = ~x807 & ~x1134;
  assign n8061 = n7212 & ~n8060;
  assign n8062 = ~x868 & x1134;
  assign n8063 = n8061 & ~n8062;
  assign n8064 = ~n8059 & ~n8063;
  assign n8065 = n7054 & ~n8064;
  assign n8066 = ~n8049 & ~n8065;
  assign n8067 = x356 & n7026;
  assign n8068 = x405 & n7015;
  assign n8069 = x381 & n7017;
  assign n8070 = ~n8068 & ~n8069;
  assign n8071 = n3506 & ~n8070;
  assign n8072 = x445 & n7021;
  assign n8073 = ~n8071 & ~n8072;
  assign n8074 = ~n8067 & n8073;
  assign n8075 = n1483 & n8074;
  assign n8076 = ~x199 & n5296;
  assign n8077 = x199 & x1081;
  assign n8078 = ~n1483 & ~n8077;
  assign n8079 = ~n8076 & n8078;
  assign n8080 = n2699 & ~n8079;
  assign n8081 = ~n8075 & n8080;
  assign n8082 = x684 & x1135;
  assign n8083 = x1134 & ~n8082;
  assign n8084 = x750 & ~x1135;
  assign n8085 = n8083 & ~n8084;
  assign n8086 = ~x651 & ~x1135;
  assign n8087 = ~x1134 & ~n8086;
  assign n8088 = x654 & x1135;
  assign n8089 = n8087 & ~n8088;
  assign n8090 = ~n8085 & ~n8089;
  assign n8091 = x1136 & ~n8090;
  assign n8092 = ~x794 & ~x1134;
  assign n8093 = n7212 & ~n8092;
  assign n8094 = ~x880 & x1134;
  assign n8095 = n8093 & ~n8094;
  assign n8096 = ~n8091 & ~n8095;
  assign n8097 = n7054 & ~n8096;
  assign n8098 = ~n8081 & ~n8097;
  assign n8099 = x747 & x773;
  assign n8100 = x731 & ~x945;
  assign n8101 = n8099 & n8100;
  assign n8102 = x775 & x988;
  assign n8103 = n8101 & n8102;
  assign n8104 = x769 & n8103;
  assign n8105 = n8104 ^ x721;
  assign n8106 = x798 ^ x765;
  assign n8107 = x800 ^ x771;
  assign n8108 = ~n8106 & ~n8107;
  assign n8109 = x807 ^ x747;
  assign n8110 = x816 ^ x775;
  assign n8111 = ~n8109 & ~n8110;
  assign n8112 = n8108 & n8111;
  assign n8113 = x794 ^ x769;
  assign n8114 = x801 ^ x773;
  assign n8115 = ~n8113 & ~n8114;
  assign n8116 = x813 ^ x721;
  assign n8117 = x795 ^ x731;
  assign n8118 = ~n8116 & ~n8117;
  assign n8119 = n8115 & n8118;
  assign n8120 = n8112 & n8119;
  assign n8121 = n8105 & ~n8120;
  assign n8122 = x403 & n7015;
  assign n8123 = x379 & n7017;
  assign n8124 = ~n8122 & ~n8123;
  assign n8125 = n3506 & ~n8124;
  assign n8126 = x428 & n7021;
  assign n8127 = ~n8125 & ~n8126;
  assign n8128 = n1483 & n8127;
  assign n8129 = x354 & n7026;
  assign n8130 = n8128 & ~n8129;
  assign n8131 = ~x199 & n5284;
  assign n8132 = x199 & x1045;
  assign n8133 = ~n1483 & ~n8132;
  assign n8134 = ~n8131 & n8133;
  assign n8135 = n2699 & ~n8134;
  assign n8136 = ~n8130 & n8135;
  assign n8137 = x694 & x1135;
  assign n8138 = x1134 & ~n8137;
  assign n8139 = x776 & ~x1135;
  assign n8140 = n8138 & ~n8139;
  assign n8141 = ~x640 & ~x1135;
  assign n8142 = ~x1134 & ~n8141;
  assign n8143 = x732 & x1135;
  assign n8144 = n8142 & ~n8143;
  assign n8145 = ~n8140 & ~n8144;
  assign n8146 = x1136 & ~n8145;
  assign n8147 = ~x795 & ~x1134;
  assign n8148 = n7212 & ~n8147;
  assign n8149 = ~x851 & x1134;
  assign n8150 = n8148 & ~n8149;
  assign n8151 = ~n8146 & ~n8150;
  assign n8152 = n7054 & ~n8151;
  assign n8153 = ~n8136 & ~n8152;
  assign n8154 = ~x1111 & n7565;
  assign n8155 = ~x962 & ~n8154;
  assign n8156 = x723 & ~n7565;
  assign n8157 = n8155 & ~n8156;
  assign n8158 = ~x1114 & n7565;
  assign n8159 = ~x962 & ~n8158;
  assign n8160 = x724 & ~n7565;
  assign n8161 = n8159 & ~n8160;
  assign n8162 = ~x1120 & n7565;
  assign n8163 = ~x962 & ~n8162;
  assign n8164 = x725 & ~n7565;
  assign n8165 = n8163 & ~n8164;
  assign n8166 = ~x1126 & n7565;
  assign n8167 = ~x962 & ~n8166;
  assign n8168 = ~x726 & ~n7565;
  assign n8169 = n8167 & ~n8168;
  assign n8170 = ~x1102 & n7565;
  assign n8171 = ~x962 & ~n8170;
  assign n8172 = ~x727 & ~n7565;
  assign n8173 = n8171 & ~n8172;
  assign n8174 = ~x1131 & n7565;
  assign n8175 = ~x962 & ~n8174;
  assign n8176 = x728 & ~n7565;
  assign n8177 = n8175 & ~n8176;
  assign n8178 = ~x1104 & n7565;
  assign n8179 = ~x962 & ~n8178;
  assign n8180 = ~x729 & ~n7565;
  assign n8181 = n8179 & ~n8180;
  assign n8182 = ~x1106 & n7565;
  assign n8183 = ~x962 & ~n8182;
  assign n8184 = ~x730 & ~n7565;
  assign n8185 = n8183 & ~n8184;
  assign n8186 = ~x945 & x988;
  assign n8187 = n8099 & n8186;
  assign n8188 = n8187 ^ x731;
  assign n8189 = ~n8120 & n8188;
  assign n8190 = ~x1128 & n6856;
  assign n8191 = ~x962 & ~n8190;
  assign n8192 = x732 & ~n6856;
  assign n8193 = n8191 & ~n8192;
  assign n8194 = x316 & n7026;
  assign n8195 = x399 & n7015;
  assign n8196 = x375 & n7017;
  assign n8197 = ~n8195 & ~n8196;
  assign n8198 = n3506 & ~n8197;
  assign n8199 = x424 & n7021;
  assign n8200 = ~n8198 & ~n8199;
  assign n8201 = ~n8194 & n8200;
  assign n8202 = n1483 & n8201;
  assign n8203 = ~x308 & n3150;
  assign n8204 = x199 & ~x1047;
  assign n8205 = ~n8203 & ~n8204;
  assign n8206 = ~x1037 & n3242;
  assign n8207 = n8205 & ~n8206;
  assign n8208 = ~n1483 & ~n8207;
  assign n8209 = n2699 & ~n8208;
  assign n8210 = ~n8202 & n8209;
  assign n8211 = x777 ^ x737;
  assign n8212 = ~x1135 & n8211;
  assign n8213 = n8212 ^ x737;
  assign n8214 = x1134 & n8213;
  assign n8215 = x1136 & ~n8214;
  assign n8216 = x648 ^ x619;
  assign n8217 = x1135 & n8216;
  assign n8218 = n8217 ^ x619;
  assign n8219 = ~x1134 & ~n8218;
  assign n8220 = n8215 & ~n8219;
  assign n8221 = x838 & n7213;
  assign n8222 = ~n8220 & ~n8221;
  assign n8223 = n7054 & ~n8222;
  assign n8224 = ~n8210 & ~n8223;
  assign n8225 = ~x1119 & n7565;
  assign n8226 = ~x962 & ~n8225;
  assign n8227 = x734 & ~n7565;
  assign n8228 = n8226 & ~n8227;
  assign n8229 = ~x1109 & n7565;
  assign n8230 = ~x962 & ~n8229;
  assign n8231 = ~x735 & ~n7565;
  assign n8232 = n8230 & ~n8231;
  assign n8233 = ~x1101 & n7565;
  assign n8234 = ~x962 & ~n8233;
  assign n8235 = ~x736 & ~n7565;
  assign n8236 = n8234 & ~n8235;
  assign n8237 = ~x1122 & n7565;
  assign n8238 = ~x962 & ~n8237;
  assign n8239 = x737 & ~n7565;
  assign n8240 = n8238 & ~n8239;
  assign n8241 = ~x1121 & n7565;
  assign n8242 = ~x962 & ~n8241;
  assign n8243 = x738 & ~n7565;
  assign n8244 = n8242 & ~n8243;
  assign n8245 = ~x952 & n6747;
  assign n8246 = x739 & ~n8245;
  assign n8247 = ~x966 & ~n8246;
  assign n8248 = x1108 & n8245;
  assign n8249 = n8247 & ~n8248;
  assign n8250 = ~x741 & ~n8245;
  assign n8251 = ~x966 & ~n8250;
  assign n8252 = x1114 & n8245;
  assign n8253 = n8251 & ~n8252;
  assign n8254 = ~x742 & ~n8245;
  assign n8255 = ~x966 & ~n8254;
  assign n8256 = x1112 & n8245;
  assign n8257 = n8255 & ~n8256;
  assign n8258 = x743 & ~n8245;
  assign n8259 = ~x966 & ~n8258;
  assign n8260 = x1109 & n8245;
  assign n8261 = n8259 & ~n8260;
  assign n8262 = ~x744 & ~n8245;
  assign n8263 = ~x966 & ~n8262;
  assign n8264 = x1131 & n8245;
  assign n8265 = n8263 & ~n8264;
  assign n8266 = ~x745 & ~n8245;
  assign n8267 = ~x966 & ~n8266;
  assign n8268 = x1111 & n8245;
  assign n8269 = n8267 & ~n8268;
  assign n8270 = x746 & ~n8245;
  assign n8271 = ~x966 & ~n8270;
  assign n8272 = x1104 & n8245;
  assign n8273 = n8271 & ~n8272;
  assign n8274 = x773 & n8186;
  assign n8275 = n8274 ^ x747;
  assign n8276 = ~n8120 & n8275;
  assign n8277 = x748 & ~n8245;
  assign n8278 = ~x966 & ~n8277;
  assign n8279 = x1106 & n8245;
  assign n8280 = n8278 & ~n8279;
  assign n8281 = x749 & ~n8245;
  assign n8282 = ~x966 & ~n8281;
  assign n8283 = x1105 & n8245;
  assign n8284 = n8282 & ~n8283;
  assign n8285 = ~x750 & ~n8245;
  assign n8286 = ~x966 & ~n8285;
  assign n8287 = x1130 & n8245;
  assign n8288 = n8286 & ~n8287;
  assign n8289 = ~x751 & ~n8245;
  assign n8290 = ~x966 & ~n8289;
  assign n8291 = x1123 & n8245;
  assign n8292 = n8290 & ~n8291;
  assign n8293 = ~x752 & ~n8245;
  assign n8294 = ~x966 & ~n8293;
  assign n8295 = x1124 & n8245;
  assign n8296 = n8294 & ~n8295;
  assign n8297 = ~x753 & ~n8245;
  assign n8298 = ~x966 & ~n8297;
  assign n8299 = x1117 & n8245;
  assign n8300 = n8298 & ~n8299;
  assign n8301 = ~x754 & ~n8245;
  assign n8302 = ~x966 & ~n8301;
  assign n8303 = x1118 & n8245;
  assign n8304 = n8302 & ~n8303;
  assign n8305 = ~x755 & ~n8245;
  assign n8306 = ~x966 & ~n8305;
  assign n8307 = x1120 & n8245;
  assign n8308 = n8306 & ~n8307;
  assign n8309 = ~x756 & ~n8245;
  assign n8310 = ~x966 & ~n8309;
  assign n8311 = x1119 & n8245;
  assign n8312 = n8310 & ~n8311;
  assign n8313 = ~x757 & ~n8245;
  assign n8314 = ~x966 & ~n8313;
  assign n8315 = x1113 & n8245;
  assign n8316 = n8314 & ~n8315;
  assign n8317 = x758 & ~n8245;
  assign n8318 = ~x966 & ~n8317;
  assign n8319 = x1101 & n8245;
  assign n8320 = n8318 & ~n8319;
  assign n8321 = x759 & ~n8245;
  assign n8322 = ~x966 & ~n8321;
  assign n8323 = x1100 & n8245;
  assign n8324 = n8322 & ~n8323;
  assign n8325 = ~x760 & ~n8245;
  assign n8326 = ~x966 & ~n8325;
  assign n8327 = x1115 & n8245;
  assign n8328 = n8326 & ~n8327;
  assign n8329 = ~x761 & ~n8245;
  assign n8330 = ~x966 & ~n8329;
  assign n8331 = x1121 & n8245;
  assign n8332 = n8330 & ~n8331;
  assign n8333 = ~x762 & ~n8245;
  assign n8334 = ~x966 & ~n8333;
  assign n8335 = x1129 & n8245;
  assign n8336 = n8334 & ~n8335;
  assign n8337 = x763 & ~n8245;
  assign n8338 = ~x966 & ~n8337;
  assign n8339 = x1103 & n8245;
  assign n8340 = n8338 & ~n8339;
  assign n8341 = x764 & ~n8245;
  assign n8342 = ~x966 & ~n8341;
  assign n8343 = x1107 & n8245;
  assign n8344 = n8342 & ~n8343;
  assign n8345 = ~x773 & ~x794;
  assign n8346 = ~x795 & ~x816;
  assign n8347 = n8345 & n8346;
  assign n8348 = ~x721 & ~x747;
  assign n8349 = ~x765 & ~x771;
  assign n8350 = n8348 & n8349;
  assign n8351 = n8347 & n8350;
  assign n8352 = n8120 & ~n8351;
  assign n8353 = x945 ^ x765;
  assign n8354 = ~n8352 & ~n8353;
  assign n8355 = x766 & ~n8245;
  assign n8356 = ~x966 & ~n8355;
  assign n8357 = x1110 & n8245;
  assign n8358 = n8356 & ~n8357;
  assign n8359 = ~x767 & ~n8245;
  assign n8360 = ~x966 & ~n8359;
  assign n8361 = x1116 & n8245;
  assign n8362 = n8360 & ~n8361;
  assign n8363 = ~x768 & ~n8245;
  assign n8364 = ~x966 & ~n8363;
  assign n8365 = x1125 & n8245;
  assign n8366 = n8364 & ~n8365;
  assign n8367 = n8103 ^ x769;
  assign n8368 = ~n8120 & n8367;
  assign n8369 = ~x770 & ~n8245;
  assign n8370 = ~x966 & ~n8369;
  assign n8371 = x1126 & n8245;
  assign n8372 = n8370 & ~n8371;
  assign n8373 = x987 ^ x771;
  assign n8374 = ~x945 & n8373;
  assign n8375 = n8374 ^ x771;
  assign n8376 = ~n8352 & n8375;
  assign n8377 = x772 & ~n8245;
  assign n8378 = ~x966 & ~n8377;
  assign n8379 = x1102 & n8245;
  assign n8380 = n8378 & ~n8379;
  assign n8381 = n8186 ^ x773;
  assign n8382 = ~n8352 & n8381;
  assign n8383 = ~x774 & ~n8245;
  assign n8384 = ~x966 & ~n8383;
  assign n8385 = x1127 & n8245;
  assign n8386 = n8384 & ~n8385;
  assign n8387 = x765 & x771;
  assign n8388 = n8101 & n8387;
  assign n8389 = n8388 ^ x775;
  assign n8390 = ~n8120 & n8389;
  assign n8391 = ~x776 & ~n8245;
  assign n8392 = ~x966 & ~n8391;
  assign n8393 = x1128 & n8245;
  assign n8394 = n8392 & ~n8393;
  assign n8395 = ~x777 & ~n8245;
  assign n8396 = ~x966 & ~n8395;
  assign n8397 = x1122 & n8245;
  assign n8398 = n8396 & ~n8397;
  assign n8399 = x832 & x956;
  assign n8400 = ~x1083 & x1085;
  assign n8401 = n8399 & n8400;
  assign n8402 = ~x1046 & n8401;
  assign n8403 = ~x968 & n8402;
  assign n8404 = x1100 ^ x778;
  assign n8405 = n8403 & n8404;
  assign n8406 = n8405 ^ x778;
  assign n8407 = x779 & ~n6805;
  assign n8408 = x780 & ~n6727;
  assign n8409 = x1101 ^ x781;
  assign n8410 = n8403 & n8409;
  assign n8411 = n8410 ^ x781;
  assign n8412 = ~n2185 & ~n6757;
  assign n8413 = ~n6726 & n8412;
  assign n8414 = x1109 ^ x783;
  assign n8415 = n8403 & n8414;
  assign n8416 = n8415 ^ x783;
  assign n8417 = x1110 ^ x784;
  assign n8418 = n8403 & n8417;
  assign n8419 = n8418 ^ x784;
  assign n8420 = x1102 ^ x785;
  assign n8421 = n8403 & n8420;
  assign n8422 = n8421 ^ x785;
  assign n8423 = x786 ^ x24;
  assign n8424 = x954 & n8423;
  assign n8425 = n8424 ^ x24;
  assign n8426 = x1104 ^ x787;
  assign n8427 = n8403 & n8426;
  assign n8428 = n8427 ^ x787;
  assign n8429 = x1105 ^ x788;
  assign n8430 = n8403 & n8429;
  assign n8431 = n8430 ^ x788;
  assign n8432 = x1106 ^ x789;
  assign n8433 = n8403 & n8432;
  assign n8434 = n8433 ^ x789;
  assign n8435 = x1107 ^ x790;
  assign n8436 = n8403 & n8435;
  assign n8437 = n8436 ^ x790;
  assign n8438 = x1108 ^ x791;
  assign n8439 = n8403 & n8438;
  assign n8440 = n8439 ^ x791;
  assign n8441 = x1103 ^ x792;
  assign n8442 = n8403 & n8441;
  assign n8443 = n8442 ^ x792;
  assign n8444 = x968 & n8402;
  assign n8445 = x1130 ^ x794;
  assign n8446 = n8444 & n8445;
  assign n8447 = n8446 ^ x794;
  assign n8448 = x1128 ^ x795;
  assign n8449 = n8444 & n8448;
  assign n8450 = n8449 ^ x795;
  assign n8451 = x266 & ~x269;
  assign n8452 = x279 & n8451;
  assign n8453 = x278 & ~x280;
  assign n8454 = n8452 & n8453;
  assign n8455 = n6996 & n6998;
  assign n8456 = n8454 & n8455;
  assign n8457 = n8456 ^ x264;
  assign n8458 = x1124 ^ x798;
  assign n8459 = n8444 & n8458;
  assign n8460 = n8459 ^ x798;
  assign n8461 = x1107 ^ x799;
  assign n8462 = n8444 & ~n8461;
  assign n8463 = n8462 ^ x799;
  assign n8464 = x1125 ^ x800;
  assign n8465 = n8444 & n8464;
  assign n8466 = n8465 ^ x800;
  assign n8467 = x1126 ^ x801;
  assign n8468 = n8444 & n8467;
  assign n8469 = n8468 ^ x801;
  assign n8470 = ~x274 & n7001;
  assign n8471 = x1106 ^ x803;
  assign n8472 = n8444 & ~n8471;
  assign n8473 = n8472 ^ x803;
  assign n8474 = x1109 ^ x804;
  assign n8475 = n8444 & n8474;
  assign n8476 = n8475 ^ x804;
  assign n8477 = n6997 ^ x270;
  assign n8478 = x1127 ^ x807;
  assign n8479 = n8444 & n8478;
  assign n8480 = n8479 ^ x807;
  assign n8481 = x1101 ^ x808;
  assign n8482 = n8444 & n8481;
  assign n8483 = n8482 ^ x808;
  assign n8484 = x1103 ^ x809;
  assign n8485 = n8444 & ~n8484;
  assign n8486 = n8485 ^ x809;
  assign n8487 = x1108 ^ x810;
  assign n8488 = n8444 & n8487;
  assign n8489 = n8488 ^ x810;
  assign n8490 = x1102 ^ x811;
  assign n8491 = n8444 & n8490;
  assign n8492 = n8491 ^ x811;
  assign n8493 = x1104 ^ x812;
  assign n8494 = n8444 & ~n8493;
  assign n8495 = n8494 ^ x812;
  assign n8496 = x1131 ^ x813;
  assign n8497 = n8444 & n8496;
  assign n8498 = n8497 ^ x813;
  assign n8499 = x1105 ^ x814;
  assign n8500 = n8444 & ~n8499;
  assign n8501 = n8500 ^ x814;
  assign n8502 = x1110 ^ x815;
  assign n8503 = n8444 & n8502;
  assign n8504 = n8503 ^ x815;
  assign n8505 = x1129 ^ x816;
  assign n8506 = n8444 & n8505;
  assign n8507 = n8506 ^ x816;
  assign n8508 = n6994 ^ x269;
  assign n8509 = ~n3776 & ~n3780;
  assign n8510 = n7000 ^ x265;
  assign n8511 = ~x270 & n6997;
  assign n8512 = n8511 ^ x277;
  assign n8513 = ~x811 & ~x893;
  assign n8514 = n1424 & n2699;
  assign n8515 = ~x982 & ~n1423;
  assign n8516 = ~n8514 & ~n8515;
  assign n8517 = n1426 & ~n8516;
  assign n8518 = x123 & n1484;
  assign n8523 = x1127 ^ x1126;
  assign n8522 = x1125 ^ x1124;
  assign n8524 = n8523 ^ n8522;
  assign n8520 = x1129 ^ x1128;
  assign n8519 = x1131 ^ x1130;
  assign n8521 = n8520 ^ n8519;
  assign n8525 = n8524 ^ n8521;
  assign n8526 = n8525 ^ x825;
  assign n8527 = ~n8518 & ~n8526;
  assign n8528 = n8527 ^ x825;
  assign n8533 = x1119 ^ x1118;
  assign n8532 = x1117 ^ x1116;
  assign n8534 = n8533 ^ n8532;
  assign n8530 = x1121 ^ x1120;
  assign n8529 = x1123 ^ x1122;
  assign n8531 = n8530 ^ n8529;
  assign n8535 = n8534 ^ n8531;
  assign n8536 = n8535 ^ x826;
  assign n8537 = ~n8518 & ~n8536;
  assign n8538 = n8537 ^ x826;
  assign n8543 = x1101 ^ x1100;
  assign n8542 = x1103 ^ x1102;
  assign n8544 = n8543 ^ n8542;
  assign n8540 = x1105 ^ x1104;
  assign n8539 = x1107 ^ x1106;
  assign n8541 = n8540 ^ n8539;
  assign n8545 = n8544 ^ n8541;
  assign n8546 = n8545 ^ x827;
  assign n8547 = ~n8518 & ~n8546;
  assign n8548 = n8547 ^ x827;
  assign n8553 = x1115 ^ x1114;
  assign n8552 = x1113 ^ x1112;
  assign n8554 = n8553 ^ n8552;
  assign n8550 = x1111 ^ x1110;
  assign n8549 = x1109 ^ x1108;
  assign n8551 = n8550 ^ n8549;
  assign n8555 = n8554 ^ n8551;
  assign n8556 = n8555 ^ x828;
  assign n8557 = ~n8518 & ~n8556;
  assign n8558 = n8557 ^ x828;
  assign n8559 = x1091 & n2695;
  assign n8560 = n2699 & n8559;
  assign n8561 = ~x951 & x1092;
  assign n8562 = ~n8560 & ~n8561;
  assign n8563 = n8454 ^ x281;
  assign n8564 = ~x832 & ~x1163;
  assign n8565 = n2734 & n8564;
  assign n8566 = n8559 & n8565;
  assign n8567 = x1091 ^ x833;
  assign n8568 = n2695 & n8567;
  assign n8569 = n8568 ^ x833;
  assign n8570 = x946 & n2695;
  assign n8571 = ~x281 & n6995;
  assign n8572 = n8571 ^ x282;
  assign n8573 = x1049 ^ x837;
  assign n8574 = ~x955 & n8573;
  assign n8575 = n8574 ^ x837;
  assign n8576 = x1047 ^ x838;
  assign n8577 = ~x955 & n8576;
  assign n8578 = n8577 ^ x838;
  assign n8579 = x1074 ^ x839;
  assign n8580 = ~x955 & n8579;
  assign n8581 = n8580 ^ x839;
  assign n8582 = x1196 ^ x840;
  assign n8583 = n2695 & n8582;
  assign n8584 = n8583 ^ x840;
  assign n8585 = x1035 ^ x842;
  assign n8586 = ~x955 & n8585;
  assign n8587 = n8586 ^ x842;
  assign n8588 = x1079 ^ x843;
  assign n8589 = ~x955 & n8588;
  assign n8590 = n8589 ^ x843;
  assign n8591 = x1078 ^ x844;
  assign n8592 = ~x955 & n8591;
  assign n8593 = n8592 ^ x844;
  assign n8594 = x1043 ^ x845;
  assign n8595 = ~x955 & n8594;
  assign n8596 = n8595 ^ x845;
  assign n8597 = x1134 ^ x846;
  assign n8598 = ~n5302 & n8597;
  assign n8599 = n8598 ^ x846;
  assign n8600 = x1055 ^ x847;
  assign n8601 = ~x955 & n8600;
  assign n8602 = n8601 ^ x847;
  assign n8603 = x1039 ^ x848;
  assign n8604 = ~x955 & n8603;
  assign n8605 = n8604 ^ x848;
  assign n8606 = x1198 ^ x849;
  assign n8607 = n2695 & n8606;
  assign n8608 = n8607 ^ x849;
  assign n8609 = x1048 ^ x850;
  assign n8610 = ~x955 & n8609;
  assign n8611 = n8610 ^ x850;
  assign n8612 = x1045 ^ x851;
  assign n8613 = ~x955 & n8612;
  assign n8614 = n8613 ^ x851;
  assign n8615 = x1062 ^ x852;
  assign n8616 = ~x955 & n8615;
  assign n8617 = n8616 ^ x852;
  assign n8618 = x1080 ^ x853;
  assign n8619 = ~x955 & n8618;
  assign n8620 = n8619 ^ x853;
  assign n8621 = x1051 ^ x854;
  assign n8622 = ~x955 & n8621;
  assign n8623 = n8622 ^ x854;
  assign n8624 = x1065 ^ x855;
  assign n8625 = ~x955 & n8624;
  assign n8626 = n8625 ^ x855;
  assign n8627 = x1067 ^ x856;
  assign n8628 = ~x955 & n8627;
  assign n8629 = n8628 ^ x856;
  assign n8630 = x1058 ^ x857;
  assign n8631 = ~x955 & n8630;
  assign n8632 = n8631 ^ x857;
  assign n8633 = x1087 ^ x858;
  assign n8634 = ~x955 & n8633;
  assign n8635 = n8634 ^ x858;
  assign n8636 = x1070 ^ x859;
  assign n8637 = ~x955 & n8636;
  assign n8638 = n8637 ^ x859;
  assign n8639 = x1076 ^ x860;
  assign n8640 = ~x955 & n8639;
  assign n8641 = n8640 ^ x860;
  assign n8642 = x1141 ^ x861;
  assign n8643 = ~n5302 & n8642;
  assign n8644 = n8643 ^ x861;
  assign n8645 = x1139 ^ x862;
  assign n8646 = ~n5302 & n8645;
  assign n8647 = n8646 ^ x862;
  assign n8648 = x1199 ^ x863;
  assign n8649 = n2695 & n8648;
  assign n8650 = n8649 ^ x863;
  assign n8651 = x1197 ^ x864;
  assign n8652 = n2695 & n8651;
  assign n8653 = n8652 ^ x864;
  assign n8654 = x1040 ^ x865;
  assign n8655 = ~x955 & n8654;
  assign n8656 = n8655 ^ x865;
  assign n8657 = x1053 ^ x866;
  assign n8658 = ~x955 & n8657;
  assign n8659 = n8658 ^ x866;
  assign n8660 = x1057 ^ x867;
  assign n8661 = ~x955 & n8660;
  assign n8662 = n8661 ^ x867;
  assign n8663 = x1063 ^ x868;
  assign n8664 = ~x955 & n8663;
  assign n8665 = n8664 ^ x868;
  assign n8666 = x1140 ^ x869;
  assign n8667 = ~n5302 & n8666;
  assign n8668 = n8667 ^ x869;
  assign n8669 = x1069 ^ x870;
  assign n8670 = ~x955 & n8669;
  assign n8671 = n8670 ^ x870;
  assign n8672 = x1072 ^ x871;
  assign n8673 = ~x955 & n8672;
  assign n8674 = n8673 ^ x871;
  assign n8675 = x1084 ^ x872;
  assign n8676 = ~x955 & n8675;
  assign n8677 = n8676 ^ x872;
  assign n8678 = x1044 ^ x873;
  assign n8679 = ~x955 & n8678;
  assign n8680 = n8679 ^ x873;
  assign n8681 = x1036 ^ x874;
  assign n8682 = ~x955 & n8681;
  assign n8683 = n8682 ^ x874;
  assign n8684 = x1136 ^ x875;
  assign n8685 = ~n5302 & n8684;
  assign n8686 = n8685 ^ x875;
  assign n8687 = x1037 ^ x876;
  assign n8688 = ~x955 & n8687;
  assign n8689 = n8688 ^ x876;
  assign n8690 = x1138 ^ x877;
  assign n8691 = ~n5302 & n8690;
  assign n8692 = n8691 ^ x877;
  assign n8693 = x1137 ^ x878;
  assign n8694 = ~n5302 & n8693;
  assign n8695 = n8694 ^ x878;
  assign n8696 = x1135 ^ x879;
  assign n8697 = ~n5302 & n8696;
  assign n8698 = n8697 ^ x879;
  assign n8699 = x1081 ^ x880;
  assign n8700 = ~x955 & n8699;
  assign n8701 = n8700 ^ x880;
  assign n8702 = x1059 ^ x881;
  assign n8703 = ~x955 & n8702;
  assign n8704 = n8703 ^ x881;
  assign n8705 = x1107 ^ x883;
  assign n8706 = ~n8518 & ~n8705;
  assign n8707 = n8706 ^ x883;
  assign n8708 = x1124 ^ x884;
  assign n8709 = ~n8518 & ~n8708;
  assign n8710 = n8709 ^ x884;
  assign n8711 = x1125 ^ x885;
  assign n8712 = ~n8518 & ~n8711;
  assign n8713 = n8712 ^ x885;
  assign n8714 = x1109 ^ x886;
  assign n8715 = ~n8518 & ~n8714;
  assign n8716 = n8715 ^ x886;
  assign n8717 = x1100 ^ x887;
  assign n8718 = ~n8518 & ~n8717;
  assign n8719 = n8718 ^ x887;
  assign n8720 = x1120 ^ x888;
  assign n8721 = ~n8518 & ~n8720;
  assign n8722 = n8721 ^ x888;
  assign n8723 = x1103 ^ x889;
  assign n8724 = ~n8518 & ~n8723;
  assign n8725 = n8724 ^ x889;
  assign n8726 = x1126 ^ x890;
  assign n8727 = ~n8518 & ~n8726;
  assign n8728 = n8727 ^ x890;
  assign n8729 = x1116 ^ x891;
  assign n8730 = ~n8518 & ~n8729;
  assign n8731 = n8730 ^ x891;
  assign n8732 = x1101 ^ x892;
  assign n8733 = ~n8518 & ~n8732;
  assign n8734 = n8733 ^ x892;
  assign n8735 = x1119 ^ x894;
  assign n8736 = ~n8518 & ~n8735;
  assign n8737 = n8736 ^ x894;
  assign n8738 = x1113 ^ x895;
  assign n8739 = ~n8518 & ~n8738;
  assign n8740 = n8739 ^ x895;
  assign n8741 = x1118 ^ x896;
  assign n8742 = ~n8518 & ~n8741;
  assign n8743 = n8742 ^ x896;
  assign n8744 = x1129 ^ x898;
  assign n8745 = ~n8518 & ~n8744;
  assign n8746 = n8745 ^ x898;
  assign n8747 = x1115 ^ x899;
  assign n8748 = ~n8518 & ~n8747;
  assign n8749 = n8748 ^ x899;
  assign n8750 = x1110 ^ x900;
  assign n8751 = ~n8518 & ~n8750;
  assign n8752 = n8751 ^ x900;
  assign n8753 = x1111 ^ x902;
  assign n8754 = ~n8518 & ~n8753;
  assign n8755 = n8754 ^ x902;
  assign n8756 = x1121 ^ x903;
  assign n8757 = ~n8518 & ~n8756;
  assign n8758 = n8757 ^ x903;
  assign n8759 = x1127 ^ x904;
  assign n8760 = ~n8518 & ~n8759;
  assign n8761 = n8760 ^ x904;
  assign n8762 = x1131 ^ x905;
  assign n8763 = ~n8518 & ~n8762;
  assign n8764 = n8763 ^ x905;
  assign n8765 = x1128 ^ x906;
  assign n8766 = ~n8518 & ~n8765;
  assign n8767 = n8766 ^ x906;
  assign n8768 = ~x624 & ~x979;
  assign n8769 = x604 & n8768;
  assign n8770 = ~x598 & x979;
  assign n8771 = ~x615 & n8770;
  assign n8772 = ~n8769 & ~n8771;
  assign n8773 = n8772 ^ x907;
  assign n8774 = x782 & ~n8773;
  assign n8775 = n8774 ^ x907;
  assign n8776 = x1122 ^ x908;
  assign n8777 = ~n8518 & ~n8776;
  assign n8778 = n8777 ^ x908;
  assign n8779 = x1105 ^ x909;
  assign n8780 = ~n8518 & ~n8779;
  assign n8781 = n8780 ^ x909;
  assign n8782 = x1117 ^ x910;
  assign n8783 = ~n8518 & ~n8782;
  assign n8784 = n8783 ^ x910;
  assign n8785 = x1130 ^ x911;
  assign n8786 = ~n8518 & ~n8785;
  assign n8787 = n8786 ^ x911;
  assign n8788 = x1114 ^ x912;
  assign n8789 = ~n8518 & ~n8788;
  assign n8790 = n8789 ^ x912;
  assign n8791 = x1106 ^ x913;
  assign n8792 = ~n8518 & ~n8791;
  assign n8793 = n8792 ^ x913;
  assign n8794 = n6993 ^ x280;
  assign n8795 = x1108 ^ x915;
  assign n8796 = ~n8518 & ~n8795;
  assign n8797 = n8796 ^ x915;
  assign n8798 = x1123 ^ x916;
  assign n8799 = ~n8518 & ~n8798;
  assign n8800 = n8799 ^ x916;
  assign n8801 = x1112 ^ x917;
  assign n8802 = ~n8518 & ~n8801;
  assign n8803 = n8802 ^ x917;
  assign n8804 = x1104 ^ x918;
  assign n8805 = ~n8518 & ~n8804;
  assign n8806 = n8805 ^ x918;
  assign n8807 = x1102 ^ x919;
  assign n8808 = ~n8518 & ~n8807;
  assign n8809 = n8808 ^ x919;
  assign n8810 = x1139 ^ x920;
  assign n8811 = x1093 & n8810;
  assign n8812 = n8811 ^ x920;
  assign n8813 = x1140 ^ x921;
  assign n8814 = x1093 & n8813;
  assign n8815 = n8814 ^ x921;
  assign n8816 = x1152 ^ x922;
  assign n8817 = x1093 & n8816;
  assign n8818 = n8817 ^ x922;
  assign n8819 = x1154 ^ x923;
  assign n8820 = x1093 & n8819;
  assign n8821 = n8820 ^ x923;
  assign n8822 = x311 & n5643;
  assign n8823 = x1155 ^ x925;
  assign n8824 = x1093 & n8823;
  assign n8825 = n8824 ^ x925;
  assign n8826 = x1157 ^ x926;
  assign n8827 = x1093 & n8826;
  assign n8828 = n8827 ^ x926;
  assign n8829 = x1145 ^ x927;
  assign n8830 = x1093 & n8829;
  assign n8831 = n8830 ^ x927;
  assign n8832 = x1136 ^ x928;
  assign n8833 = x1093 & n8832;
  assign n8834 = n8833 ^ x928;
  assign n8835 = x1144 ^ x929;
  assign n8836 = x1093 & n8835;
  assign n8837 = n8836 ^ x929;
  assign n8838 = x1134 ^ x930;
  assign n8839 = x1093 & n8838;
  assign n8840 = n8839 ^ x930;
  assign n8841 = x1150 ^ x931;
  assign n8842 = x1093 & n8841;
  assign n8843 = n8842 ^ x931;
  assign n8844 = x1142 ^ x932;
  assign n8845 = x1093 & n8844;
  assign n8846 = n8845 ^ x932;
  assign n8847 = x1137 ^ x933;
  assign n8848 = x1093 & n8847;
  assign n8849 = n8848 ^ x933;
  assign n8850 = x1147 ^ x934;
  assign n8851 = x1093 & n8850;
  assign n8852 = n8851 ^ x934;
  assign n8853 = x1141 ^ x935;
  assign n8854 = x1093 & n8853;
  assign n8855 = n8854 ^ x935;
  assign n8856 = x1149 ^ x936;
  assign n8857 = x1093 & n8856;
  assign n8858 = n8857 ^ x936;
  assign n8859 = x1148 ^ x937;
  assign n8860 = x1093 & n8859;
  assign n8861 = n8860 ^ x937;
  assign n8862 = x1135 ^ x938;
  assign n8863 = x1093 & n8862;
  assign n8864 = n8863 ^ x938;
  assign n8865 = x1146 ^ x939;
  assign n8866 = x1093 & n8865;
  assign n8867 = n8866 ^ x939;
  assign n8868 = x1138 ^ x940;
  assign n8869 = x1093 & n8868;
  assign n8870 = n8869 ^ x940;
  assign n8871 = x1153 ^ x941;
  assign n8872 = x1093 & n8871;
  assign n8873 = n8872 ^ x941;
  assign n8874 = x1156 ^ x942;
  assign n8875 = x1093 & n8874;
  assign n8876 = n8875 ^ x942;
  assign n8877 = x1151 ^ x943;
  assign n8878 = x1093 & n8877;
  assign n8879 = n8878 ^ x943;
  assign n8880 = x1143 ^ x944;
  assign n8881 = x1093 & n8880;
  assign n8882 = n8881 ^ x944;
  assign n8883 = x230 & n2695;
  assign n8884 = ~n8768 & ~n8770;
  assign n8885 = n8884 ^ x947;
  assign n8886 = x782 & n8885;
  assign n8887 = n8886 ^ x947;
  assign n8888 = x992 ^ x266;
  assign n8889 = x949 ^ x313;
  assign n8890 = x954 & ~n8889;
  assign n8891 = n8890 ^ x313;
  assign n8892 = x1092 & n1423;
  assign n8893 = x957 & x1092;
  assign n8894 = ~x31 & ~n8893;
  assign n8895 = ~x782 & x960;
  assign n8896 = ~x230 & x961;
  assign n8897 = ~x782 & x963;
  assign n8898 = ~x230 & x967;
  assign n8899 = ~x230 & x969;
  assign n8900 = ~x782 & x970;
  assign n8901 = ~x230 & x971;
  assign n8902 = ~x782 & x972;
  assign n8903 = ~x230 & x974;
  assign n8904 = ~x782 & x975;
  assign n8905 = ~x230 & x977;
  assign n8906 = ~x782 & x978;
  assign n8907 = ~x598 & x615;
  assign n8908 = x824 & x1092;
  assign n8909 = ~x604 & ~x624;
  assign y0 = x668;
  assign y1 = x672;
  assign y2 = x664;
  assign y3 = x667;
  assign y4 = x676;
  assign y5 = x673;
  assign y6 = x675;
  assign y7 = x666;
  assign y8 = x679;
  assign y9 = x674;
  assign y10 = x663;
  assign y11 = x670;
  assign y12 = x677;
  assign y13 = x682;
  assign y14 = x671;
  assign y15 = x678;
  assign y16 = x718;
  assign y17 = x707;
  assign y18 = x708;
  assign y19 = x713;
  assign y20 = x711;
  assign y21 = x716;
  assign y22 = x733;
  assign y23 = x712;
  assign y24 = x689;
  assign y25 = x717;
  assign y26 = x692;
  assign y27 = x719;
  assign y28 = x722;
  assign y29 = x714;
  assign y30 = x720;
  assign y31 = x685;
  assign y32 = x837;
  assign y33 = x850;
  assign y34 = x872;
  assign y35 = x871;
  assign y36 = x881;
  assign y37 = x866;
  assign y38 = x876;
  assign y39 = x873;
  assign y40 = x874;
  assign y41 = x859;
  assign y42 = x855;
  assign y43 = x852;
  assign y44 = x870;
  assign y45 = x848;
  assign y46 = x865;
  assign y47 = x856;
  assign y48 = x853;
  assign y49 = x847;
  assign y50 = x857;
  assign y51 = x854;
  assign y52 = x858;
  assign y53 = x845;
  assign y54 = x838;
  assign y55 = x842;
  assign y56 = x843;
  assign y57 = x839;
  assign y58 = x844;
  assign y59 = x868;
  assign y60 = x851;
  assign y61 = x867;
  assign y62 = x880;
  assign y63 = x860;
  assign y64 = x1030;
  assign y65 = x1034;
  assign y66 = x1015;
  assign y67 = x1020;
  assign y68 = x1025;
  assign y69 = x1005;
  assign y70 = x996;
  assign y71 = x1012;
  assign y72 = x993;
  assign y73 = x1016;
  assign y74 = x1021;
  assign y75 = x1010;
  assign y76 = x1027;
  assign y77 = x1018;
  assign y78 = x1017;
  assign y79 = x1024;
  assign y80 = x1009;
  assign y81 = x1032;
  assign y82 = x1003;
  assign y83 = x997;
  assign y84 = x1013;
  assign y85 = x1011;
  assign y86 = x1008;
  assign y87 = x1019;
  assign y88 = x1031;
  assign y89 = x1022;
  assign y90 = x1000;
  assign y91 = x1023;
  assign y92 = x1002;
  assign y93 = x1026;
  assign y94 = x1006;
  assign y95 = x998;
  assign y96 = x31;
  assign y97 = x80;
  assign y98 = x893;
  assign y99 = x467;
  assign y100 = x78;
  assign y101 = x112;
  assign y102 = x13;
  assign y103 = x25;
  assign y104 = x226;
  assign y105 = x127;
  assign y106 = x822;
  assign y107 = x808;
  assign y108 = x227;
  assign y109 = x477;
  assign y110 = x834;
  assign y111 = x229;
  assign y112 = x12;
  assign y113 = x11;
  assign y114 = x10;
  assign y115 = x9;
  assign y116 = x8;
  assign y117 = x7;
  assign y118 = x6;
  assign y119 = x5;
  assign y120 = x4;
  assign y121 = x3;
  assign y122 = x0;
  assign y123 = x2;
  assign y124 = x1;
  assign y125 = x310;
  assign y126 = x302;
  assign y127 = x475;
  assign y128 = x474;
  assign y129 = x466;
  assign y130 = x473;
  assign y131 = x471;
  assign y132 = x472;
  assign y133 = x470;
  assign y134 = x469;
  assign y135 = x465;
  assign y136 = x1028;
  assign y137 = x1033;
  assign y138 = x995;
  assign y139 = x994;
  assign y140 = x28;
  assign y141 = x27;
  assign y142 = x26;
  assign y143 = x29;
  assign y144 = x15;
  assign y145 = x14;
  assign y146 = x21;
  assign y147 = x20;
  assign y148 = x19;
  assign y149 = x18;
  assign y150 = x17;
  assign y151 = x16;
  assign y152 = x1096;
  assign y153 = ~n1661;
  assign y154 = ~n1708;
  assign y155 = ~n1728;
  assign y156 = ~n1772;
  assign y157 = ~n1823;
  assign y158 = n1864;
  assign y159 = ~n1902;
  assign y160 = ~n1942;
  assign y161 = n1984;
  assign y162 = n2032;
  assign y163 = n2073;
  assign y164 = n2108;
  assign y165 = n2141;
  assign y166 = ~1'b0;
  assign y167 = ~n2247;
  assign y168 = x228;
  assign y169 = x22;
  assign y170 = ~x1090;
  assign y171 = n2349;
  assign y172 = n2357;
  assign y173 = n2361;
  assign y174 = ~n2375;
  assign y175 = n2378;
  assign y176 = n2381;
  assign y177 = n2384;
  assign y178 = n2387;
  assign y179 = x1089;
  assign y180 = x23;
  assign y181 = ~n2247;
  assign y182 = ~n2415;
  assign y183 = n2421;
  assign y184 = n2427;
  assign y185 = n2429;
  assign y186 = n2431;
  assign y187 = n2433;
  assign y188 = x37;
  assign y189 = ~n2738;
  assign y190 = ~n2770;
  assign y191 = ~n2909;
  assign y192 = n2997;
  assign y193 = n3044;
  assign y194 = n3050;
  assign y195 = ~n2412;
  assign y196 = ~n3062;
  assign y197 = ~n3090;
  assign y198 = n3095;
  assign y199 = n3139;
  assign y200 = ~n3163;
  assign y201 = ~n3178;
  assign y202 = ~n3186;
  assign y203 = n3187;
  assign y204 = ~n3194;
  assign y205 = ~n3203;
  assign y206 = n3205;
  assign y207 = ~n3209;
  assign y208 = ~n3227;
  assign y209 = n3232;
  assign y210 = ~n3250;
  assign y211 = ~n3258;
  assign y212 = ~n3262;
  assign y213 = ~n3265;
  assign y214 = n3272;
  assign y215 = ~n3277;
  assign y216 = n3279;
  assign y217 = ~n3284;
  assign y218 = ~n3290;
  assign y219 = ~n3293;
  assign y220 = n3298;
  assign y221 = ~n3302;
  assign y222 = ~n3305;
  assign y223 = n3306;
  assign y224 = n3315;
  assign y225 = n3320;
  assign y226 = n3326;
  assign y227 = n3329;
  assign y228 = ~n3344;
  assign y229 = ~n3355;
  assign y230 = ~n3364;
  assign y231 = n3370;
  assign y232 = ~n3381;
  assign y233 = ~n3384;
  assign y234 = n3395;
  assign y235 = n3398;
  assign y236 = n3399;
  assign y237 = ~n3501;
  assign y238 = n3526;
  assign y239 = n3529;
  assign y240 = n3533;
  assign y241 = ~n3539;
  assign y242 = n3543;
  assign y243 = n3546;
  assign y244 = n3547;
  assign y245 = n3548;
  assign y246 = ~n3554;
  assign y247 = n3558;
  assign y248 = ~n3561;
  assign y249 = ~n3568;
  assign y250 = n3572;
  assign y251 = ~n3576;
  assign y252 = ~n3580;
  assign y253 = ~n3592;
  assign y254 = n3600;
  assign y255 = ~n3605;
  assign y256 = n3608;
  assign y257 = ~n3618;
  assign y258 = n3628;
  assign y259 = ~n3635;
  assign y260 = n3636;
  assign y261 = n3637;
  assign y262 = ~n3641;
  assign y263 = x117;
  assign y264 = ~n3644;
  assign y265 = n3645;
  assign y266 = ~n3650;
  assign y267 = n3651;
  assign y268 = ~n3655;
  assign y269 = ~n3659;
  assign y270 = ~n3660;
  assign y271 = n3663;
  assign y272 = n3665;
  assign y273 = n3668;
  assign y274 = n3670;
  assign y275 = ~n2418;
  assign y276 = n3757;
  assign y277 = n3771;
  assign y278 = n3783;
  assign y279 = n3835;
  assign y280 = ~n3774;
  assign y281 = n3848;
  assign y282 = ~n3918;
  assign y283 = n3958;
  assign y284 = n3965;
  assign y285 = x131;
  assign y286 = ~n3973;
  assign y287 = ~n4006;
  assign y288 = ~n3768;
  assign y289 = n4044;
  assign y290 = n4066;
  assign y291 = n4085;
  assign y292 = n4103;
  assign y293 = n4128;
  assign y294 = ~n4136;
  assign y295 = ~n4152;
  assign y296 = ~n4157;
  assign y297 = ~n4241;
  assign y298 = ~n4247;
  assign y299 = n4253;
  assign y300 = ~n4259;
  assign y301 = n4265;
  assign y302 = ~n4271;
  assign y303 = n4278;
  assign y304 = ~n4284;
  assign y305 = ~n4290;
  assign y306 = ~n4305;
  assign y307 = ~n4311;
  assign y308 = ~n4317;
  assign y309 = n4323;
  assign y310 = ~n4329;
  assign y311 = ~n4335;
  assign y312 = ~n4341;
  assign y313 = ~n4347;
  assign y314 = ~n4353;
  assign y315 = ~n4359;
  assign y316 = ~n4365;
  assign y317 = ~n4371;
  assign y318 = n4377;
  assign y319 = ~n4383;
  assign y320 = ~n4389;
  assign y321 = ~n4395;
  assign y322 = ~n4401;
  assign y323 = n4407;
  assign y324 = ~n4413;
  assign y325 = ~n4419;
  assign y326 = ~n4425;
  assign y327 = ~n4431;
  assign y328 = ~n4437;
  assign y329 = ~n4443;
  assign y330 = ~n4449;
  assign y331 = n4455;
  assign y332 = ~n4461;
  assign y333 = ~n4467;
  assign y334 = ~n4473;
  assign y335 = ~n4479;
  assign y336 = ~n4485;
  assign y337 = ~n4491;
  assign y338 = ~n4497;
  assign y339 = ~n4503;
  assign y340 = ~n4509;
  assign y341 = ~n4515;
  assign y342 = ~n4521;
  assign y343 = ~n4527;
  assign y344 = ~n4533;
  assign y345 = ~n4539;
  assign y346 = n4545;
  assign y347 = ~n4551;
  assign y348 = ~n4557;
  assign y349 = ~n4563;
  assign y350 = ~n4569;
  assign y351 = ~n4575;
  assign y352 = ~n4583;
  assign y353 = ~n4593;
  assign y354 = ~n4599;
  assign y355 = n4605;
  assign y356 = n4611;
  assign y357 = n4617;
  assign y358 = ~n4644;
  assign y359 = ~n4652;
  assign y360 = ~n4659;
  assign y361 = ~n4670;
  assign y362 = ~n4674;
  assign y363 = ~n4681;
  assign y364 = ~n4687;
  assign y365 = ~n4693;
  assign y366 = ~n4699;
  assign y367 = n4705;
  assign y368 = n4711;
  assign y369 = ~n4717;
  assign y370 = ~n4723;
  assign y371 = ~n4729;
  assign y372 = n4735;
  assign y373 = n4741;
  assign y374 = ~n4747;
  assign y375 = ~n4751;
  assign y376 = ~n4757;
  assign y377 = ~n4761;
  assign y378 = n4767;
  assign y379 = n4773;
  assign y380 = n4779;
  assign y381 = n4785;
  assign y382 = ~n4795;
  assign y383 = n4804;
  assign y384 = ~n4814;
  assign y385 = ~n4822;
  assign y386 = x232;
  assign y387 = n4826;
  assign y388 = x236;
  assign y389 = ~n4834;
  assign y390 = ~n4925;
  assign y391 = ~n4954;
  assign y392 = ~n4985;
  assign y393 = ~n4801;
  assign y394 = n5045;
  assign y395 = ~n5072;
  assign y396 = n5086;
  assign y397 = n5104;
  assign y398 = n5116;
  assign y399 = ~n5130;
  assign y400 = ~n5166;
  assign y401 = ~n5174;
  assign y402 = n5186;
  assign y403 = n5198;
  assign y404 = n5204;
  assign y405 = n5216;
  assign y406 = n5222;
  assign y407 = n5224;
  assign y408 = n5233;
  assign y409 = ~n5239;
  assign y410 = n5248;
  assign y411 = n5257;
  assign y412 = n5263;
  assign y413 = n5269;
  assign y414 = n5275;
  assign y415 = n5281;
  assign y416 = n5287;
  assign y417 = n5293;
  assign y418 = n5299;
  assign y419 = ~n5306;
  assign y420 = ~n5315;
  assign y421 = ~n5326;
  assign y422 = ~n5337;
  assign y423 = n5348;
  assign y424 = n5357;
  assign y425 = n5366;
  assign y426 = ~n5377;
  assign y427 = ~n5388;
  assign y428 = n5397;
  assign y429 = n5406;
  assign y430 = n5415;
  assign y431 = ~n5426;
  assign y432 = n5435;
  assign y433 = n5444;
  assign y434 = ~n5455;
  assign y435 = n5466;
  assign y436 = n5477;
  assign y437 = ~n5488;
  assign y438 = ~n5499;
  assign y439 = ~n5510;
  assign y440 = n5519;
  assign y441 = ~n5523;
  assign y442 = n5535;
  assign y443 = n5543;
  assign y444 = n5545;
  assign y445 = n5548;
  assign y446 = n5557;
  assign y447 = n5560;
  assign y448 = n5563;
  assign y449 = n5566;
  assign y450 = n5569;
  assign y451 = n5572;
  assign y452 = n5575;
  assign y453 = n5578;
  assign y454 = n5581;
  assign y455 = n5584;
  assign y456 = ~n5591;
  assign y457 = ~n5595;
  assign y458 = n5599;
  assign y459 = ~n5614;
  assign y460 = n5617;
  assign y461 = n5620;
  assign y462 = n5623;
  assign y463 = n5626;
  assign y464 = n5629;
  assign y465 = n5632;
  assign y466 = n5635;
  assign y467 = ~n5642;
  assign y468 = n5646;
  assign y469 = n5648;
  assign y470 = ~n5654;
  assign y471 = n5656;
  assign y472 = n5660;
  assign y473 = n5663;
  assign y474 = n5667;
  assign y475 = n5671;
  assign y476 = n5674;
  assign y477 = n5677;
  assign y478 = n5680;
  assign y479 = n5683;
  assign y480 = n5686;
  assign y481 = n5689;
  assign y482 = n5692;
  assign y483 = n5695;
  assign y484 = n5698;
  assign y485 = n5701;
  assign y486 = n5704;
  assign y487 = n5709;
  assign y488 = n5713;
  assign y489 = ~n5717;
  assign y490 = n5720;
  assign y491 = n5723;
  assign y492 = n5726;
  assign y493 = n5729;
  assign y494 = n5732;
  assign y495 = n5735;
  assign y496 = n5738;
  assign y497 = ~n5742;
  assign y498 = n5746;
  assign y499 = n5749;
  assign y500 = n5752;
  assign y501 = n5755;
  assign y502 = n5758;
  assign y503 = n5761;
  assign y504 = n5764;
  assign y505 = n5767;
  assign y506 = n5770;
  assign y507 = n5773;
  assign y508 = n5776;
  assign y509 = n5779;
  assign y510 = n5782;
  assign y511 = n5785;
  assign y512 = n5788;
  assign y513 = n5791;
  assign y514 = n5794;
  assign y515 = n5797;
  assign y516 = n5800;
  assign y517 = n5803;
  assign y518 = n5806;
  assign y519 = n5809;
  assign y520 = n5812;
  assign y521 = n5815;
  assign y522 = n5818;
  assign y523 = n5821;
  assign y524 = n5824;
  assign y525 = n5827;
  assign y526 = n5830;
  assign y527 = n5833;
  assign y528 = n5836;
  assign y529 = n5839;
  assign y530 = n5842;
  assign y531 = n5845;
  assign y532 = n5848;
  assign y533 = n5851;
  assign y534 = n5854;
  assign y535 = n5857;
  assign y536 = n5860;
  assign y537 = n5863;
  assign y538 = n5866;
  assign y539 = n5869;
  assign y540 = n5872;
  assign y541 = n5875;
  assign y542 = n5878;
  assign y543 = n5881;
  assign y544 = n5884;
  assign y545 = n5887;
  assign y546 = n5890;
  assign y547 = n5893;
  assign y548 = n5896;
  assign y549 = n5899;
  assign y550 = n5902;
  assign y551 = n5905;
  assign y552 = n5908;
  assign y553 = n5911;
  assign y554 = n5914;
  assign y555 = n5917;
  assign y556 = n5920;
  assign y557 = n5923;
  assign y558 = n5926;
  assign y559 = n5929;
  assign y560 = n5932;
  assign y561 = n5935;
  assign y562 = n5938;
  assign y563 = n5941;
  assign y564 = n5944;
  assign y565 = n5947;
  assign y566 = n5950;
  assign y567 = n5953;
  assign y568 = n5956;
  assign y569 = n5959;
  assign y570 = n5962;
  assign y571 = n5965;
  assign y572 = n5968;
  assign y573 = n5971;
  assign y574 = n5974;
  assign y575 = n5977;
  assign y576 = n5980;
  assign y577 = n5983;
  assign y578 = n5986;
  assign y579 = n5989;
  assign y580 = n5992;
  assign y581 = n5995;
  assign y582 = n5998;
  assign y583 = n6001;
  assign y584 = n6004;
  assign y585 = n6007;
  assign y586 = n6010;
  assign y587 = n6013;
  assign y588 = n6016;
  assign y589 = n6019;
  assign y590 = n6022;
  assign y591 = n6025;
  assign y592 = n6028;
  assign y593 = n6031;
  assign y594 = n6034;
  assign y595 = n6037;
  assign y596 = n6040;
  assign y597 = n6043;
  assign y598 = n6046;
  assign y599 = n6049;
  assign y600 = n6052;
  assign y601 = n6055;
  assign y602 = n6058;
  assign y603 = n6061;
  assign y604 = n6064;
  assign y605 = n6067;
  assign y606 = n6070;
  assign y607 = n6073;
  assign y608 = n6076;
  assign y609 = n6079;
  assign y610 = n6082;
  assign y611 = n6085;
  assign y612 = n6088;
  assign y613 = n6091;
  assign y614 = n6114;
  assign y615 = n6117;
  assign y616 = n6120;
  assign y617 = n6123;
  assign y618 = n6126;
  assign y619 = n6129;
  assign y620 = n6132;
  assign y621 = n6135;
  assign y622 = ~n6140;
  assign y623 = ~n6145;
  assign y624 = ~n6150;
  assign y625 = ~n6153;
  assign y626 = ~n6158;
  assign y627 = ~n6163;
  assign y628 = ~n6168;
  assign y629 = ~n6173;
  assign y630 = ~n6178;
  assign y631 = ~n6183;
  assign y632 = ~n6188;
  assign y633 = ~n6190;
  assign y634 = n5651;
  assign y635 = n6191;
  assign y636 = x583;
  assign y637 = n5524;
  assign y638 = n6194;
  assign y639 = n6197;
  assign y640 = n6200;
  assign y641 = n6203;
  assign y642 = n6206;
  assign y643 = n6209;
  assign y644 = n6212;
  assign y645 = n6215;
  assign y646 = n6218;
  assign y647 = n6221;
  assign y648 = n6224;
  assign y649 = n6227;
  assign y650 = n6230;
  assign y651 = n6233;
  assign y652 = n6236;
  assign y653 = n6239;
  assign y654 = n6242;
  assign y655 = n6245;
  assign y656 = n6248;
  assign y657 = n6251;
  assign y658 = n6254;
  assign y659 = n6257;
  assign y660 = n6260;
  assign y661 = n6263;
  assign y662 = n6266;
  assign y663 = n6269;
  assign y664 = n6272;
  assign y665 = n6275;
  assign y666 = n6278;
  assign y667 = n6281;
  assign y668 = n6284;
  assign y669 = n6287;
  assign y670 = n6290;
  assign y671 = n6293;
  assign y672 = n6296;
  assign y673 = n6299;
  assign y674 = n6302;
  assign y675 = n6305;
  assign y676 = n6308;
  assign y677 = n6311;
  assign y678 = n6314;
  assign y679 = n6317;
  assign y680 = n6320;
  assign y681 = n6323;
  assign y682 = n6326;
  assign y683 = n6329;
  assign y684 = n6332;
  assign y685 = n6335;
  assign y686 = n6338;
  assign y687 = n6341;
  assign y688 = n6344;
  assign y689 = n6347;
  assign y690 = n6350;
  assign y691 = n6353;
  assign y692 = n6356;
  assign y693 = n6359;
  assign y694 = n6362;
  assign y695 = n6365;
  assign y696 = n6368;
  assign y697 = n6371;
  assign y698 = n6374;
  assign y699 = n6377;
  assign y700 = n6380;
  assign y701 = n6383;
  assign y702 = n6386;
  assign y703 = n6389;
  assign y704 = n6392;
  assign y705 = n6395;
  assign y706 = n6398;
  assign y707 = n6401;
  assign y708 = n6404;
  assign y709 = n6407;
  assign y710 = n6410;
  assign y711 = n6413;
  assign y712 = n6416;
  assign y713 = n6419;
  assign y714 = n6422;
  assign y715 = n6425;
  assign y716 = n6428;
  assign y717 = n6431;
  assign y718 = n6434;
  assign y719 = n6437;
  assign y720 = n6440;
  assign y721 = n6443;
  assign y722 = n6446;
  assign y723 = n6449;
  assign y724 = n6458;
  assign y725 = n6461;
  assign y726 = n6464;
  assign y727 = n6467;
  assign y728 = n6470;
  assign y729 = n6473;
  assign y730 = n6476;
  assign y731 = n6479;
  assign y732 = n6482;
  assign y733 = n6485;
  assign y734 = n6488;
  assign y735 = n6491;
  assign y736 = n6494;
  assign y737 = n6497;
  assign y738 = n6500;
  assign y739 = n6503;
  assign y740 = ~n2221;
  assign y741 = n6506;
  assign y742 = n6509;
  assign y743 = n6512;
  assign y744 = n6515;
  assign y745 = n6521;
  assign y746 = ~n6542;
  assign y747 = ~n6546;
  assign y748 = n6550;
  assign y749 = n6554;
  assign y750 = ~n6710;
  assign y751 = n6714;
  assign y752 = n6718;
  assign y753 = n6723;
  assign y754 = n6725;
  assign y755 = ~n6731;
  assign y756 = n6734;
  assign y757 = n6736;
  assign y758 = n6740;
  assign y759 = n6743;
  assign y760 = n6755;
  assign y761 = ~n6762;
  assign y762 = n6764;
  assign y763 = ~n6770;
  assign y764 = n6774;
  assign y765 = n6778;
  assign y766 = n6782;
  assign y767 = n6786;
  assign y768 = n6790;
  assign y769 = n6794;
  assign y770 = n6798;
  assign y771 = n6804;
  assign y772 = ~n6809;
  assign y773 = ~n6815;
  assign y774 = ~n6821;
  assign y775 = n6825;
  assign y776 = n6829;
  assign y777 = n6833;
  assign y778 = n6837;
  assign y779 = n6841;
  assign y780 = n6845;
  assign y781 = ~n6851;
  assign y782 = n6860;
  assign y783 = n6864;
  assign y784 = n6868;
  assign y785 = n6872;
  assign y786 = n6876;
  assign y787 = n6880;
  assign y788 = n6884;
  assign y789 = n6888;
  assign y790 = n6892;
  assign y791 = n6896;
  assign y792 = n6900;
  assign y793 = n6904;
  assign y794 = n6908;
  assign y795 = n6912;
  assign y796 = n6916;
  assign y797 = n6920;
  assign y798 = n6924;
  assign y799 = n6928;
  assign y800 = n6932;
  assign y801 = n6936;
  assign y802 = n6940;
  assign y803 = n6944;
  assign y804 = n6948;
  assign y805 = n6952;
  assign y806 = n6956;
  assign y807 = n6960;
  assign y808 = n6964;
  assign y809 = n6968;
  assign y810 = n6972;
  assign y811 = n6976;
  assign y812 = n6980;
  assign y813 = n6984;
  assign y814 = n6988;
  assign y815 = n6992;
  assign y816 = ~n7002;
  assign y817 = n7006;
  assign y818 = n7010;
  assign y819 = n7014;
  assign y820 = ~n7057;
  assign y821 = ~n7091;
  assign y822 = n7095;
  assign y823 = ~n7129;
  assign y824 = ~n7163;
  assign y825 = ~n7197;
  assign y826 = n7201;
  assign y827 = ~n7233;
  assign y828 = ~n7262;
  assign y829 = ~n7296;
  assign y830 = ~n7330;
  assign y831 = ~n7365;
  assign y832 = ~n7399;
  assign y833 = ~n7433;
  assign y834 = ~n7462;
  assign y835 = ~n7492;
  assign y836 = ~n7527;
  assign y837 = n7531;
  assign y838 = n7535;
  assign y839 = ~n7564;
  assign y840 = n1428;
  assign y841 = n7569;
  assign y842 = ~n7601;
  assign y843 = n7605;
  assign y844 = n7609;
  assign y845 = n7613;
  assign y846 = ~n7645;
  assign y847 = n7649;
  assign y848 = n7653;
  assign y849 = ~n7685;
  assign y850 = n7689;
  assign y851 = n7693;
  assign y852 = n7697;
  assign y853 = n7701;
  assign y854 = n7705;
  assign y855 = n7709;
  assign y856 = n7713;
  assign y857 = n7717;
  assign y858 = n7721;
  assign y859 = n7725;
  assign y860 = n7729;
  assign y861 = n7733;
  assign y862 = n7737;
  assign y863 = n7741;
  assign y864 = ~n7772;
  assign y865 = ~n7803;
  assign y866 = n7807;
  assign y867 = n7811;
  assign y868 = ~n7842;
  assign y869 = ~n7873;
  assign y870 = ~n7904;
  assign y871 = ~n7936;
  assign y872 = n7940;
  assign y873 = ~n7971;
  assign y874 = ~n8003;
  assign y875 = ~n8034;
  assign y876 = ~n8066;
  assign y877 = ~n8098;
  assign y878 = n8121;
  assign y879 = ~n8153;
  assign y880 = n8157;
  assign y881 = n8161;
  assign y882 = n8165;
  assign y883 = n8169;
  assign y884 = n8173;
  assign y885 = n8177;
  assign y886 = n8181;
  assign y887 = n8185;
  assign y888 = n8189;
  assign y889 = n8193;
  assign y890 = ~n8224;
  assign y891 = n8228;
  assign y892 = n8232;
  assign y893 = n8236;
  assign y894 = n8240;
  assign y895 = n8244;
  assign y896 = ~n8249;
  assign y897 = n6748;
  assign y898 = ~n8253;
  assign y899 = ~n8257;
  assign y900 = ~n8261;
  assign y901 = ~n8265;
  assign y902 = ~n8269;
  assign y903 = ~n8273;
  assign y904 = n8276;
  assign y905 = ~n8280;
  assign y906 = ~n8284;
  assign y907 = ~n8288;
  assign y908 = ~n8292;
  assign y909 = ~n8296;
  assign y910 = ~n8300;
  assign y911 = ~n8304;
  assign y912 = ~n8308;
  assign y913 = ~n8312;
  assign y914 = ~n8316;
  assign y915 = ~n8320;
  assign y916 = ~n8324;
  assign y917 = ~n8328;
  assign y918 = ~n8332;
  assign y919 = ~n8336;
  assign y920 = ~n8340;
  assign y921 = ~n8344;
  assign y922 = n8354;
  assign y923 = ~n8358;
  assign y924 = ~n8362;
  assign y925 = ~n8366;
  assign y926 = n8368;
  assign y927 = ~n8372;
  assign y928 = n8376;
  assign y929 = ~n8380;
  assign y930 = n8382;
  assign y931 = ~n8386;
  assign y932 = n8390;
  assign y933 = ~n8394;
  assign y934 = ~n8398;
  assign y935 = n8406;
  assign y936 = ~n8407;
  assign y937 = ~n8408;
  assign y938 = n8411;
  assign y939 = ~n8413;
  assign y940 = n8416;
  assign y941 = n8419;
  assign y942 = n8422;
  assign y943 = ~n8425;
  assign y944 = n8428;
  assign y945 = n8431;
  assign y946 = n8434;
  assign y947 = n8437;
  assign y948 = n8440;
  assign y949 = n8443;
  assign y950 = n2183;
  assign y951 = n8447;
  assign y952 = n8450;
  assign y953 = ~n8457;
  assign y954 = n6856;
  assign y955 = n8460;
  assign y956 = ~n8463;
  assign y957 = n8466;
  assign y958 = n8469;
  assign y959 = n8470;
  assign y960 = ~n8473;
  assign y961 = n8476;
  assign y962 = ~n8477;
  assign y963 = n8352;
  assign y964 = n8480;
  assign y965 = n8483;
  assign y966 = ~n8486;
  assign y967 = n8489;
  assign y968 = n8492;
  assign y969 = ~n8495;
  assign y970 = n8498;
  assign y971 = ~n8501;
  assign y972 = n8504;
  assign y973 = n8507;
  assign y974 = ~n8508;
  assign y975 = ~n8509;
  assign y976 = ~n8510;
  assign y977 = ~n8512;
  assign y978 = n8120;
  assign y979 = n8513;
  assign y980 = n7565;
  assign y981 = n8517;
  assign y982 = ~n8528;
  assign y983 = ~n8538;
  assign y984 = ~n8548;
  assign y985 = ~n8558;
  assign y986 = ~n8562;
  assign y987 = ~n8563;
  assign y988 = n8245;
  assign y989 = n8566;
  assign y990 = n8569;
  assign y991 = n8570;
  assign y992 = ~n8572;
  assign y993 = n8575;
  assign y994 = n8578;
  assign y995 = n8581;
  assign y996 = n8584;
  assign y997 = n2785;
  assign y998 = n8587;
  assign y999 = n8590;
  assign y1000 = n8593;
  assign y1001 = n8596;
  assign y1002 = n8599;
  assign y1003 = n8602;
  assign y1004 = n8605;
  assign y1005 = n8608;
  assign y1006 = n8611;
  assign y1007 = n8614;
  assign y1008 = n8617;
  assign y1009 = n8620;
  assign y1010 = n8623;
  assign y1011 = n8626;
  assign y1012 = n8629;
  assign y1013 = n8632;
  assign y1014 = n8635;
  assign y1015 = n8638;
  assign y1016 = n8641;
  assign y1017 = n8644;
  assign y1018 = n8647;
  assign y1019 = n8650;
  assign y1020 = n8653;
  assign y1021 = n8656;
  assign y1022 = n8659;
  assign y1023 = n8662;
  assign y1024 = n8665;
  assign y1025 = n8668;
  assign y1026 = n8671;
  assign y1027 = n8674;
  assign y1028 = n8677;
  assign y1029 = n8680;
  assign y1030 = n8683;
  assign y1031 = n8686;
  assign y1032 = n8689;
  assign y1033 = n8692;
  assign y1034 = n8695;
  assign y1035 = n8698;
  assign y1036 = n8701;
  assign y1037 = n8704;
  assign y1038 = ~n1518;
  assign y1039 = ~n8707;
  assign y1040 = ~n8710;
  assign y1041 = ~n8713;
  assign y1042 = ~n8716;
  assign y1043 = ~n8719;
  assign y1044 = ~n8722;
  assign y1045 = ~n8725;
  assign y1046 = ~n8728;
  assign y1047 = ~n8731;
  assign y1048 = ~n8734;
  assign y1049 = ~n4827;
  assign y1050 = ~n8737;
  assign y1051 = ~n8740;
  assign y1052 = ~n8743;
  assign y1053 = x67;
  assign y1054 = ~n8746;
  assign y1055 = ~n8749;
  assign y1056 = ~n8752;
  assign y1057 = ~n2213;
  assign y1058 = ~n8755;
  assign y1059 = ~n8758;
  assign y1060 = ~n8761;
  assign y1061 = ~n8764;
  assign y1062 = ~n8767;
  assign y1063 = n8775;
  assign y1064 = ~n8778;
  assign y1065 = ~n8781;
  assign y1066 = ~n8784;
  assign y1067 = ~n8787;
  assign y1068 = ~n8790;
  assign y1069 = ~n8793;
  assign y1070 = ~n8794;
  assign y1071 = ~n8797;
  assign y1072 = ~n8800;
  assign y1073 = ~n8803;
  assign y1074 = ~n8806;
  assign y1075 = ~n8809;
  assign y1076 = n8812;
  assign y1077 = n8815;
  assign y1078 = n8818;
  assign y1079 = n8821;
  assign y1080 = n8822;
  assign y1081 = n8825;
  assign y1082 = n8828;
  assign y1083 = n8831;
  assign y1084 = n8834;
  assign y1085 = n8837;
  assign y1086 = n8840;
  assign y1087 = n8843;
  assign y1088 = n8846;
  assign y1089 = n8849;
  assign y1090 = n8852;
  assign y1091 = n8855;
  assign y1092 = n8858;
  assign y1093 = n8861;
  assign y1094 = n8864;
  assign y1095 = n8867;
  assign y1096 = n8870;
  assign y1097 = n8873;
  assign y1098 = n8876;
  assign y1099 = n8879;
  assign y1100 = n8882;
  assign y1101 = ~n2176;
  assign y1102 = n8883;
  assign y1103 = n8887;
  assign y1104 = n8888;
  assign y1105 = ~n8891;
  assign y1106 = n8892;
  assign y1107 = n2314;
  assign y1108 = x1134;
  assign y1109 = x964;
  assign y1110 = ~x954;
  assign y1111 = x965;
  assign y1112 = ~n8894;
  assign y1113 = x991;
  assign y1114 = x985;
  assign y1115 = n8895;
  assign y1116 = n8896;
  assign y1117 = x1014;
  assign y1118 = n8897;
  assign y1119 = x1029;
  assign y1120 = x1004;
  assign y1121 = x1007;
  assign y1122 = n8898;
  assign y1123 = x1135;
  assign y1124 = n8899;
  assign y1125 = n8900;
  assign y1126 = n8901;
  assign y1127 = n8902;
  assign y1128 = n8903;
  assign y1129 = n8904;
  assign y1130 = ~x278;
  assign y1131 = n8905;
  assign y1132 = n8906;
  assign y1133 = ~n8907;
  assign y1134 = x1064;
  assign y1135 = n8908;
  assign y1136 = x299;
  assign y1137 = ~n8909;
  assign y1138 = x1075;
  assign y1139 = x1052;
  assign y1140 = x771;
  assign y1141 = x765;
  assign y1142 = x605;
  assign y1143 = x601;
  assign y1144 = x278;
  assign y1145 = x279;
  assign y1146 = ~x915;
  assign y1147 = ~x825;
  assign y1148 = ~x826;
  assign y1149 = ~x913;
  assign y1150 = ~x894;
  assign y1151 = ~x905;
  assign y1152 = x1095;
  assign y1153 = ~x890;
  assign y1154 = x1094;
  assign y1155 = ~x906;
  assign y1156 = ~x896;
  assign y1157 = ~x909;
  assign y1158 = ~x911;
  assign y1159 = ~x908;
  assign y1160 = ~x891;
  assign y1161 = ~x902;
  assign y1162 = ~x903;
  assign y1163 = ~x883;
  assign y1164 = ~x888;
  assign y1165 = ~x919;
  assign y1166 = ~x886;
  assign y1167 = ~x912;
  assign y1168 = ~x895;
  assign y1169 = ~x916;
  assign y1170 = ~x889;
  assign y1171 = ~x900;
  assign y1172 = ~x885;
  assign y1173 = ~x904;
  assign y1174 = ~x899;
  assign y1175 = ~x918;
  assign y1176 = ~x898;
  assign y1177 = ~x917;
  assign y1178 = ~x827;
  assign y1179 = ~x887;
  assign y1180 = ~x884;
  assign y1181 = ~x910;
  assign y1182 = ~x828;
  assign y1183 = ~x892;
  assign y1184 = x1187;
  assign y1185 = x1172;
  assign y1186 = x1170;
  assign y1187 = x1138;
  assign y1188 = x1177;
  assign y1189 = x1178;
  assign y1190 = x863;
  assign y1191 = x1203;
  assign y1192 = x1185;
  assign y1193 = x1171;
  assign y1194 = x1192;
  assign y1195 = x1137;
  assign y1196 = x1186;
  assign y1197 = x1165;
  assign y1198 = x1164;
  assign y1199 = x1098;
  assign y1200 = x1183;
  assign y1201 = x230;
  assign y1202 = x1169;
  assign y1203 = x1136;
  assign y1204 = x1181;
  assign y1205 = x849;
  assign y1206 = x1193;
  assign y1207 = x1182;
  assign y1208 = x1168;
  assign y1209 = x1175;
  assign y1210 = x1191;
  assign y1211 = x1099;
  assign y1212 = x1174;
  assign y1213 = x1179;
  assign y1214 = x1202;
  assign y1215 = x1176;
  assign y1216 = x1173;
  assign y1217 = x1201;
  assign y1218 = x1167;
  assign y1219 = x840;
  assign y1220 = x1189;
  assign y1221 = x1195;
  assign y1222 = x864;
  assign y1223 = x1190;
  assign y1224 = x1188;
  assign y1225 = x1180;
  assign y1226 = x1194;
  assign y1227 = x1097;
  assign y1228 = x1166;
  assign y1229 = x1200;
  assign y1230 = x1184;
endmodule
