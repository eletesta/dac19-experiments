module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129;
  wire n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199;
  assign n513 = ~x376 & x504;
  assign n514 = ~x373 & x501;
  assign n515 = x367 & ~x495;
  assign n516 = x364 & ~x492;
  assign n517 = ~x362 & x490;
  assign n518 = x360 & ~x488;
  assign n519 = x355 & ~x483;
  assign n520 = ~x349 & x477;
  assign n521 = ~x346 & x474;
  assign n522 = x344 & ~x472;
  assign n523 = x339 & ~x467;
  assign n524 = ~x335 & x463;
  assign n525 = ~x332 & x460;
  assign n526 = ~x329 & x457;
  assign n527 = ~x322 & x450;
  assign n528 = x315 & ~x443;
  assign n529 = ~x309 & x437;
  assign n530 = ~x294 & x422;
  assign n531 = x292 & ~x420;
  assign n532 = x287 & ~x415;
  assign n533 = ~x283 & x411;
  assign n534 = x277 & ~x405;
  assign n535 = x274 & ~x402;
  assign n536 = ~x272 & x400;
  assign n537 = x270 & ~x398;
  assign n538 = ~x268 & x396;
  assign n539 = ~x261 & x389;
  assign n540 = x257 & ~x385;
  assign n541 = x256 & ~x384;
  assign n542 = ~n540 & ~n541;
  assign n543 = ~x258 & x386;
  assign n544 = ~x257 & x385;
  assign n545 = ~n543 & ~n544;
  assign n546 = ~n542 & n545;
  assign n547 = x259 & ~x387;
  assign n548 = x258 & ~x386;
  assign n549 = ~n547 & ~n548;
  assign n550 = ~n546 & n549;
  assign n551 = ~x260 & x388;
  assign n552 = ~x259 & x387;
  assign n553 = ~n551 & ~n552;
  assign n554 = ~n550 & n553;
  assign n555 = x260 & ~x388;
  assign n556 = ~n554 & ~n555;
  assign n557 = ~n539 & ~n556;
  assign n558 = x262 & ~x390;
  assign n559 = x261 & ~x389;
  assign n560 = ~n558 & ~n559;
  assign n561 = ~n557 & n560;
  assign n562 = ~x263 & x391;
  assign n563 = ~x262 & x390;
  assign n564 = ~n562 & ~n563;
  assign n565 = ~n561 & n564;
  assign n566 = x264 & ~x392;
  assign n567 = x263 & ~x391;
  assign n568 = ~n566 & ~n567;
  assign n569 = ~n565 & n568;
  assign n570 = ~x265 & x393;
  assign n571 = ~x264 & x392;
  assign n572 = ~n570 & ~n571;
  assign n573 = ~n569 & n572;
  assign n574 = x266 & ~x394;
  assign n575 = x265 & ~x393;
  assign n576 = ~n574 & ~n575;
  assign n577 = ~n573 & n576;
  assign n578 = ~x267 & x395;
  assign n579 = ~x266 & x394;
  assign n580 = ~n578 & ~n579;
  assign n581 = ~n577 & n580;
  assign n582 = x267 & ~x395;
  assign n583 = ~n581 & ~n582;
  assign n584 = ~n538 & ~n583;
  assign n585 = x269 & ~x397;
  assign n586 = x268 & ~x396;
  assign n587 = ~n585 & ~n586;
  assign n588 = ~n584 & n587;
  assign n589 = ~x269 & x397;
  assign n590 = ~n588 & ~n589;
  assign n591 = ~n537 & ~n590;
  assign n592 = ~x271 & x399;
  assign n593 = ~x270 & x398;
  assign n594 = ~n592 & ~n593;
  assign n595 = ~n591 & n594;
  assign n596 = x271 & ~x399;
  assign n597 = ~n595 & ~n596;
  assign n598 = ~n536 & ~n597;
  assign n599 = x273 & ~x401;
  assign n600 = x272 & ~x400;
  assign n601 = ~n599 & ~n600;
  assign n602 = ~n598 & n601;
  assign n603 = ~x273 & x401;
  assign n604 = ~n602 & ~n603;
  assign n605 = ~n535 & ~n604;
  assign n606 = ~x275 & x403;
  assign n607 = ~x274 & x402;
  assign n608 = ~n606 & ~n607;
  assign n609 = ~n605 & n608;
  assign n610 = x276 & ~x404;
  assign n611 = x275 & ~x403;
  assign n612 = ~n610 & ~n611;
  assign n613 = ~n609 & n612;
  assign n614 = ~x276 & x404;
  assign n615 = ~n613 & ~n614;
  assign n616 = ~n534 & ~n615;
  assign n617 = ~x278 & x406;
  assign n618 = ~x277 & x405;
  assign n619 = ~n617 & ~n618;
  assign n620 = ~n616 & n619;
  assign n621 = x279 & ~x407;
  assign n622 = x278 & ~x406;
  assign n623 = ~n621 & ~n622;
  assign n624 = ~n620 & n623;
  assign n625 = ~x280 & x408;
  assign n626 = ~x279 & x407;
  assign n627 = ~n625 & ~n626;
  assign n628 = ~n624 & n627;
  assign n629 = x281 & ~x409;
  assign n630 = x280 & ~x408;
  assign n631 = ~n629 & ~n630;
  assign n632 = ~n628 & n631;
  assign n633 = ~x282 & x410;
  assign n634 = ~x281 & x409;
  assign n635 = ~n633 & ~n634;
  assign n636 = ~n632 & n635;
  assign n637 = x282 & ~x410;
  assign n638 = ~n636 & ~n637;
  assign n639 = ~n533 & ~n638;
  assign n640 = x284 & ~x412;
  assign n641 = x283 & ~x411;
  assign n642 = ~n640 & ~n641;
  assign n643 = ~n639 & n642;
  assign n644 = ~x285 & x413;
  assign n645 = ~x284 & x412;
  assign n646 = ~n644 & ~n645;
  assign n647 = ~n643 & n646;
  assign n648 = x286 & ~x414;
  assign n649 = x285 & ~x413;
  assign n650 = ~n648 & ~n649;
  assign n651 = ~n647 & n650;
  assign n652 = ~x286 & x414;
  assign n653 = ~n651 & ~n652;
  assign n654 = ~n532 & ~n653;
  assign n655 = ~x288 & x416;
  assign n656 = ~x287 & x415;
  assign n657 = ~n655 & ~n656;
  assign n658 = ~n654 & n657;
  assign n659 = x289 & ~x417;
  assign n660 = x288 & ~x416;
  assign n661 = ~n659 & ~n660;
  assign n662 = ~n658 & n661;
  assign n663 = ~x290 & x418;
  assign n664 = ~x289 & x417;
  assign n665 = ~n663 & ~n664;
  assign n666 = ~n662 & n665;
  assign n667 = x291 & ~x419;
  assign n668 = x290 & ~x418;
  assign n669 = ~n667 & ~n668;
  assign n670 = ~n666 & n669;
  assign n671 = ~x291 & x419;
  assign n672 = ~n670 & ~n671;
  assign n673 = ~n531 & ~n672;
  assign n674 = ~x293 & x421;
  assign n675 = ~x292 & x420;
  assign n676 = ~n674 & ~n675;
  assign n677 = ~n673 & n676;
  assign n678 = x293 & ~x421;
  assign n679 = ~n677 & ~n678;
  assign n680 = ~n530 & ~n679;
  assign n681 = x295 & ~x423;
  assign n682 = x294 & ~x422;
  assign n683 = ~n681 & ~n682;
  assign n684 = ~n680 & n683;
  assign n685 = ~x297 & x425;
  assign n686 = ~x298 & x426;
  assign n687 = ~n685 & ~n686;
  assign n688 = ~x295 & x423;
  assign n689 = ~x296 & x424;
  assign n690 = ~n688 & ~n689;
  assign n691 = n687 & n690;
  assign n692 = ~n684 & n691;
  assign n693 = x297 & ~x425;
  assign n694 = x296 & ~x424;
  assign n695 = ~n693 & ~n694;
  assign n696 = n687 & ~n695;
  assign n697 = x299 & ~x427;
  assign n698 = x298 & ~x426;
  assign n699 = ~n697 & ~n698;
  assign n700 = ~n696 & n699;
  assign n701 = ~n692 & n700;
  assign n702 = ~x302 & x430;
  assign n703 = ~x301 & x429;
  assign n704 = ~n702 & ~n703;
  assign n705 = ~x299 & x427;
  assign n706 = ~x300 & x428;
  assign n707 = ~n705 & ~n706;
  assign n708 = n704 & n707;
  assign n709 = ~n701 & n708;
  assign n710 = x301 & ~x429;
  assign n711 = x300 & ~x428;
  assign n712 = ~n710 & ~n711;
  assign n713 = n704 & ~n712;
  assign n714 = x302 & ~x430;
  assign n715 = x303 & ~x431;
  assign n716 = ~n714 & ~n715;
  assign n717 = ~n713 & n716;
  assign n718 = ~n709 & n717;
  assign n719 = ~x304 & x432;
  assign n720 = ~x303 & x431;
  assign n721 = ~n719 & ~n720;
  assign n722 = ~n718 & n721;
  assign n723 = x305 & ~x433;
  assign n724 = x304 & ~x432;
  assign n725 = ~n723 & ~n724;
  assign n726 = ~n722 & n725;
  assign n727 = ~x306 & x434;
  assign n728 = ~x305 & x433;
  assign n729 = ~n727 & ~n728;
  assign n730 = ~n726 & n729;
  assign n731 = x307 & ~x435;
  assign n732 = x306 & ~x434;
  assign n733 = ~n731 & ~n732;
  assign n734 = ~n730 & n733;
  assign n735 = ~x308 & x436;
  assign n736 = ~x307 & x435;
  assign n737 = ~n735 & ~n736;
  assign n738 = ~n734 & n737;
  assign n739 = x308 & ~x436;
  assign n740 = ~n738 & ~n739;
  assign n741 = ~n529 & ~n740;
  assign n742 = x310 & ~x438;
  assign n743 = x309 & ~x437;
  assign n744 = ~n742 & ~n743;
  assign n745 = ~n741 & n744;
  assign n746 = ~x311 & x439;
  assign n747 = ~x310 & x438;
  assign n748 = ~n746 & ~n747;
  assign n749 = ~n745 & n748;
  assign n750 = x312 & ~x440;
  assign n751 = x311 & ~x439;
  assign n752 = ~n750 & ~n751;
  assign n753 = ~n749 & n752;
  assign n754 = ~x313 & x441;
  assign n755 = ~x312 & x440;
  assign n756 = ~n754 & ~n755;
  assign n757 = ~n753 & n756;
  assign n758 = x314 & ~x442;
  assign n759 = x313 & ~x441;
  assign n760 = ~n758 & ~n759;
  assign n761 = ~n757 & n760;
  assign n762 = ~x314 & x442;
  assign n763 = ~n761 & ~n762;
  assign n764 = ~n528 & ~n763;
  assign n765 = ~x315 & x443;
  assign n766 = ~x316 & x444;
  assign n767 = ~n765 & ~n766;
  assign n768 = ~x318 & x446;
  assign n769 = ~x317 & x445;
  assign n770 = ~n768 & ~n769;
  assign n771 = ~x319 & x447;
  assign n772 = n770 & ~n771;
  assign n773 = n767 & n772;
  assign n774 = ~n764 & n773;
  assign n775 = x317 & ~x445;
  assign n776 = x316 & ~x444;
  assign n777 = ~n775 & ~n776;
  assign n778 = n772 & ~n777;
  assign n779 = x320 & ~x448;
  assign n780 = x447 ^ x319;
  assign n781 = x318 & ~x446;
  assign n782 = n781 ^ x447;
  assign n783 = ~n780 & n782;
  assign n784 = n783 ^ x319;
  assign n785 = ~n779 & ~n784;
  assign n786 = ~n778 & n785;
  assign n787 = ~n774 & n786;
  assign n788 = ~x321 & x449;
  assign n789 = ~x320 & x448;
  assign n790 = ~n788 & ~n789;
  assign n791 = ~n787 & n790;
  assign n792 = x321 & ~x449;
  assign n793 = ~n791 & ~n792;
  assign n794 = ~n527 & ~n793;
  assign n795 = x323 & ~x451;
  assign n796 = x322 & ~x450;
  assign n797 = ~n795 & ~n796;
  assign n798 = ~n794 & n797;
  assign n799 = ~x325 & x453;
  assign n800 = ~x326 & x454;
  assign n801 = ~n799 & ~n800;
  assign n802 = ~x323 & x451;
  assign n803 = ~x324 & x452;
  assign n804 = ~n802 & ~n803;
  assign n805 = n801 & n804;
  assign n806 = ~n798 & n805;
  assign n807 = x325 & ~x453;
  assign n808 = x324 & ~x452;
  assign n809 = ~n807 & ~n808;
  assign n810 = n801 & ~n809;
  assign n811 = x327 & ~x455;
  assign n812 = x326 & ~x454;
  assign n813 = ~n811 & ~n812;
  assign n814 = ~n810 & n813;
  assign n815 = ~n806 & n814;
  assign n816 = ~x328 & x456;
  assign n817 = ~x327 & x455;
  assign n818 = ~n816 & ~n817;
  assign n819 = ~n815 & n818;
  assign n820 = x328 & ~x456;
  assign n821 = ~n819 & ~n820;
  assign n822 = ~n526 & ~n821;
  assign n823 = x330 & ~x458;
  assign n824 = x329 & ~x457;
  assign n825 = ~n823 & ~n824;
  assign n826 = ~n822 & n825;
  assign n827 = ~x331 & x459;
  assign n828 = ~x330 & x458;
  assign n829 = ~n827 & ~n828;
  assign n830 = ~n826 & n829;
  assign n831 = x331 & ~x459;
  assign n832 = ~n830 & ~n831;
  assign n833 = ~n525 & ~n832;
  assign n834 = x333 & ~x461;
  assign n835 = x332 & ~x460;
  assign n836 = ~n834 & ~n835;
  assign n837 = ~n833 & n836;
  assign n838 = ~x334 & x462;
  assign n839 = ~x333 & x461;
  assign n840 = ~n838 & ~n839;
  assign n841 = ~n837 & n840;
  assign n842 = x334 & ~x462;
  assign n843 = ~n841 & ~n842;
  assign n844 = ~n524 & ~n843;
  assign n845 = x336 & ~x464;
  assign n846 = x335 & ~x463;
  assign n847 = ~n845 & ~n846;
  assign n848 = ~n844 & n847;
  assign n849 = ~x337 & x465;
  assign n850 = ~x336 & x464;
  assign n851 = ~n849 & ~n850;
  assign n852 = ~n848 & n851;
  assign n853 = x338 & ~x466;
  assign n854 = x337 & ~x465;
  assign n855 = ~n853 & ~n854;
  assign n856 = ~n852 & n855;
  assign n857 = ~x338 & x466;
  assign n858 = ~n856 & ~n857;
  assign n859 = ~n523 & ~n858;
  assign n860 = ~x340 & x468;
  assign n861 = ~x339 & x467;
  assign n862 = ~n860 & ~n861;
  assign n863 = ~n859 & n862;
  assign n864 = x341 & ~x469;
  assign n865 = x340 & ~x468;
  assign n866 = ~n864 & ~n865;
  assign n867 = ~n863 & n866;
  assign n868 = ~x342 & x470;
  assign n869 = ~x341 & x469;
  assign n870 = ~n868 & ~n869;
  assign n871 = ~n867 & n870;
  assign n872 = x343 & ~x471;
  assign n873 = x342 & ~x470;
  assign n874 = ~n872 & ~n873;
  assign n875 = ~n871 & n874;
  assign n876 = ~x343 & x471;
  assign n877 = ~n875 & ~n876;
  assign n878 = ~n522 & ~n877;
  assign n879 = ~x345 & x473;
  assign n880 = ~x344 & x472;
  assign n881 = ~n879 & ~n880;
  assign n882 = ~n878 & n881;
  assign n883 = x345 & ~x473;
  assign n884 = ~n882 & ~n883;
  assign n885 = ~n521 & ~n884;
  assign n886 = x347 & ~x475;
  assign n887 = x346 & ~x474;
  assign n888 = ~n886 & ~n887;
  assign n889 = ~n885 & n888;
  assign n890 = ~x348 & x476;
  assign n891 = ~x347 & x475;
  assign n892 = ~n890 & ~n891;
  assign n893 = ~n889 & n892;
  assign n894 = x348 & ~x476;
  assign n895 = ~n893 & ~n894;
  assign n896 = ~n520 & ~n895;
  assign n897 = x350 & ~x478;
  assign n898 = x349 & ~x477;
  assign n899 = ~n897 & ~n898;
  assign n900 = ~n896 & n899;
  assign n901 = ~x351 & x479;
  assign n902 = ~x350 & x478;
  assign n903 = ~n901 & ~n902;
  assign n904 = ~n900 & n903;
  assign n905 = x352 & ~x480;
  assign n906 = x351 & ~x479;
  assign n907 = ~n905 & ~n906;
  assign n908 = ~n904 & n907;
  assign n909 = ~x353 & x481;
  assign n910 = ~x352 & x480;
  assign n911 = ~n909 & ~n910;
  assign n912 = ~n908 & n911;
  assign n913 = x354 & ~x482;
  assign n914 = x353 & ~x481;
  assign n915 = ~n913 & ~n914;
  assign n916 = ~n912 & n915;
  assign n917 = ~x354 & x482;
  assign n918 = ~n916 & ~n917;
  assign n919 = ~n519 & ~n918;
  assign n920 = ~x356 & x484;
  assign n921 = ~x355 & x483;
  assign n922 = ~n920 & ~n921;
  assign n923 = ~n919 & n922;
  assign n924 = x357 & ~x485;
  assign n925 = x356 & ~x484;
  assign n926 = ~n924 & ~n925;
  assign n927 = ~n923 & n926;
  assign n928 = ~x358 & x486;
  assign n929 = ~x357 & x485;
  assign n930 = ~n928 & ~n929;
  assign n931 = ~n927 & n930;
  assign n932 = x359 & ~x487;
  assign n933 = x358 & ~x486;
  assign n934 = ~n932 & ~n933;
  assign n935 = ~n931 & n934;
  assign n936 = ~x359 & x487;
  assign n937 = ~n935 & ~n936;
  assign n938 = ~n518 & ~n937;
  assign n939 = ~x361 & x489;
  assign n940 = ~x360 & x488;
  assign n941 = ~n939 & ~n940;
  assign n942 = ~n938 & n941;
  assign n943 = x361 & ~x489;
  assign n944 = ~n942 & ~n943;
  assign n945 = ~n517 & ~n944;
  assign n946 = x363 & ~x491;
  assign n947 = x362 & ~x490;
  assign n948 = ~n946 & ~n947;
  assign n949 = ~n945 & n948;
  assign n950 = ~x363 & x491;
  assign n951 = ~n949 & ~n950;
  assign n952 = ~n516 & ~n951;
  assign n953 = ~x365 & x493;
  assign n954 = ~x364 & x492;
  assign n955 = ~n953 & ~n954;
  assign n956 = ~n952 & n955;
  assign n957 = x366 & ~x494;
  assign n958 = x365 & ~x493;
  assign n959 = ~n957 & ~n958;
  assign n960 = ~n956 & n959;
  assign n961 = ~x366 & x494;
  assign n962 = ~n960 & ~n961;
  assign n963 = ~n515 & ~n962;
  assign n964 = ~x368 & x496;
  assign n965 = ~x367 & x495;
  assign n966 = ~n964 & ~n965;
  assign n967 = ~n963 & n966;
  assign n968 = x369 & ~x497;
  assign n969 = x368 & ~x496;
  assign n970 = ~n968 & ~n969;
  assign n971 = ~n967 & n970;
  assign n972 = ~x370 & x498;
  assign n973 = ~x369 & x497;
  assign n974 = ~n972 & ~n973;
  assign n975 = ~n971 & n974;
  assign n976 = x371 & ~x499;
  assign n977 = x370 & ~x498;
  assign n978 = ~n976 & ~n977;
  assign n979 = ~n975 & n978;
  assign n980 = ~x372 & x500;
  assign n981 = ~x371 & x499;
  assign n982 = ~n980 & ~n981;
  assign n983 = ~n979 & n982;
  assign n984 = x372 & ~x500;
  assign n985 = ~n983 & ~n984;
  assign n986 = ~n514 & ~n985;
  assign n987 = x374 & ~x502;
  assign n988 = x373 & ~x501;
  assign n989 = ~n987 & ~n988;
  assign n990 = ~n986 & n989;
  assign n991 = ~x375 & x503;
  assign n992 = ~x374 & x502;
  assign n993 = ~n991 & ~n992;
  assign n994 = ~n990 & n993;
  assign n995 = x375 & ~x503;
  assign n996 = ~n994 & ~n995;
  assign n997 = ~n513 & ~n996;
  assign n998 = x377 & ~x505;
  assign n999 = x376 & ~x504;
  assign n1000 = ~n998 & ~n999;
  assign n1001 = ~n997 & n1000;
  assign n1002 = ~x378 & x506;
  assign n1003 = ~x377 & x505;
  assign n1004 = ~n1002 & ~n1003;
  assign n1005 = ~n1001 & n1004;
  assign n1006 = x379 & ~x507;
  assign n1007 = x378 & ~x506;
  assign n1008 = ~n1006 & ~n1007;
  assign n1009 = ~n1005 & n1008;
  assign n1010 = ~x381 & x509;
  assign n1011 = ~x382 & x510;
  assign n1012 = ~n1010 & ~n1011;
  assign n1013 = ~x379 & x507;
  assign n1014 = ~x380 & x508;
  assign n1015 = ~n1013 & ~n1014;
  assign n1016 = n1012 & n1015;
  assign n1017 = ~n1009 & n1016;
  assign n1018 = x381 & ~x509;
  assign n1019 = x380 & ~x508;
  assign n1020 = ~n1018 & ~n1019;
  assign n1021 = n1012 & ~n1020;
  assign n1022 = ~x383 & x511;
  assign n1023 = x382 & ~x510;
  assign n1024 = ~n1022 & ~n1023;
  assign n1025 = ~n1021 & n1024;
  assign n1026 = ~n1017 & n1025;
  assign n1027 = x383 & ~x511;
  assign n1028 = ~n1026 & ~n1027;
  assign n1029 = x506 ^ x378;
  assign n1030 = ~n1028 & n1029;
  assign n1031 = n1030 ^ x378;
  assign n1032 = ~x122 & x250;
  assign n1033 = x120 & ~x248;
  assign n1034 = x117 & ~x245;
  assign n1035 = x114 & ~x242;
  assign n1036 = ~x110 & x238;
  assign n1037 = x106 & ~x234;
  assign n1038 = ~x102 & x230;
  assign n1039 = x98 & ~x226;
  assign n1040 = x95 & ~x223;
  assign n1041 = ~x93 & x221;
  assign n1042 = x91 & ~x219;
  assign n1043 = x82 & ~x210;
  assign n1044 = ~x65 & x193;
  assign n1045 = x57 & ~x185;
  assign n1046 = x50 & ~x178;
  assign n1047 = x39 & ~x167;
  assign n1048 = ~x33 & x161;
  assign n1049 = ~x30 & x158;
  assign n1050 = ~x27 & x155;
  assign n1051 = x19 & ~x147;
  assign n1052 = x16 & ~x144;
  assign n1053 = ~x14 & x142;
  assign n1054 = x12 & ~x140;
  assign n1055 = x9 & ~x137;
  assign n1056 = x6 & ~x134;
  assign n1057 = x1 & ~x129;
  assign n1058 = x0 & ~x128;
  assign n1059 = ~n1057 & ~n1058;
  assign n1060 = ~x2 & x130;
  assign n1061 = ~x1 & x129;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = ~n1059 & n1062;
  assign n1064 = x3 & ~x131;
  assign n1065 = x2 & ~x130;
  assign n1066 = ~n1064 & ~n1065;
  assign n1067 = ~n1063 & n1066;
  assign n1068 = ~x4 & x132;
  assign n1069 = ~x3 & x131;
  assign n1070 = ~n1068 & ~n1069;
  assign n1071 = ~n1067 & n1070;
  assign n1072 = x5 & ~x133;
  assign n1073 = x4 & ~x132;
  assign n1074 = ~n1072 & ~n1073;
  assign n1075 = ~n1071 & n1074;
  assign n1076 = ~x5 & x133;
  assign n1077 = ~n1075 & ~n1076;
  assign n1078 = ~n1056 & ~n1077;
  assign n1079 = ~x7 & x135;
  assign n1080 = ~x6 & x134;
  assign n1081 = ~n1079 & ~n1080;
  assign n1082 = ~n1078 & n1081;
  assign n1083 = x8 & ~x136;
  assign n1084 = x7 & ~x135;
  assign n1085 = ~n1083 & ~n1084;
  assign n1086 = ~n1082 & n1085;
  assign n1087 = ~x8 & x136;
  assign n1088 = ~n1086 & ~n1087;
  assign n1089 = ~n1055 & ~n1088;
  assign n1090 = ~x10 & x138;
  assign n1091 = ~x9 & x137;
  assign n1092 = ~n1090 & ~n1091;
  assign n1093 = ~n1089 & n1092;
  assign n1094 = x11 & ~x139;
  assign n1095 = x10 & ~x138;
  assign n1096 = ~n1094 & ~n1095;
  assign n1097 = ~n1093 & n1096;
  assign n1098 = ~x11 & x139;
  assign n1099 = ~n1097 & ~n1098;
  assign n1100 = ~n1054 & ~n1099;
  assign n1101 = ~x13 & x141;
  assign n1102 = ~x12 & x140;
  assign n1103 = ~n1101 & ~n1102;
  assign n1104 = ~n1100 & n1103;
  assign n1105 = x13 & ~x141;
  assign n1106 = ~n1104 & ~n1105;
  assign n1107 = ~n1053 & ~n1106;
  assign n1108 = x15 & ~x143;
  assign n1109 = x14 & ~x142;
  assign n1110 = ~n1108 & ~n1109;
  assign n1111 = ~n1107 & n1110;
  assign n1112 = ~x15 & x143;
  assign n1113 = ~n1111 & ~n1112;
  assign n1114 = ~n1052 & ~n1113;
  assign n1115 = ~x17 & x145;
  assign n1116 = ~x16 & x144;
  assign n1117 = ~n1115 & ~n1116;
  assign n1118 = ~n1114 & n1117;
  assign n1119 = x18 & ~x146;
  assign n1120 = x17 & ~x145;
  assign n1121 = ~n1119 & ~n1120;
  assign n1122 = ~n1118 & n1121;
  assign n1123 = ~x18 & x146;
  assign n1124 = ~n1122 & ~n1123;
  assign n1125 = ~n1051 & ~n1124;
  assign n1126 = ~x20 & x148;
  assign n1127 = ~x19 & x147;
  assign n1128 = ~n1126 & ~n1127;
  assign n1129 = ~n1125 & n1128;
  assign n1130 = x21 & ~x149;
  assign n1131 = x20 & ~x148;
  assign n1132 = ~n1130 & ~n1131;
  assign n1133 = ~n1129 & n1132;
  assign n1134 = ~x22 & x150;
  assign n1135 = ~x21 & x149;
  assign n1136 = ~n1134 & ~n1135;
  assign n1137 = ~n1133 & n1136;
  assign n1138 = x23 & ~x151;
  assign n1139 = x22 & ~x150;
  assign n1140 = ~n1138 & ~n1139;
  assign n1141 = ~n1137 & n1140;
  assign n1142 = ~x24 & x152;
  assign n1143 = ~x23 & x151;
  assign n1144 = ~n1142 & ~n1143;
  assign n1145 = ~n1141 & n1144;
  assign n1146 = x25 & ~x153;
  assign n1147 = x24 & ~x152;
  assign n1148 = ~n1146 & ~n1147;
  assign n1149 = ~n1145 & n1148;
  assign n1150 = ~x26 & x154;
  assign n1151 = ~x25 & x153;
  assign n1152 = ~n1150 & ~n1151;
  assign n1153 = ~n1149 & n1152;
  assign n1154 = x26 & ~x154;
  assign n1155 = ~n1153 & ~n1154;
  assign n1156 = ~n1050 & ~n1155;
  assign n1157 = x28 & ~x156;
  assign n1158 = x27 & ~x155;
  assign n1159 = ~n1157 & ~n1158;
  assign n1160 = ~n1156 & n1159;
  assign n1161 = ~x29 & x157;
  assign n1162 = ~x28 & x156;
  assign n1163 = ~n1161 & ~n1162;
  assign n1164 = ~n1160 & n1163;
  assign n1165 = x29 & ~x157;
  assign n1166 = ~n1164 & ~n1165;
  assign n1167 = ~n1049 & ~n1166;
  assign n1168 = x31 & ~x159;
  assign n1169 = x30 & ~x158;
  assign n1170 = ~n1168 & ~n1169;
  assign n1171 = ~n1167 & n1170;
  assign n1172 = ~x32 & x160;
  assign n1173 = ~x31 & x159;
  assign n1174 = ~n1172 & ~n1173;
  assign n1175 = ~n1171 & n1174;
  assign n1176 = x32 & ~x160;
  assign n1177 = ~n1175 & ~n1176;
  assign n1178 = ~n1048 & ~n1177;
  assign n1179 = x34 & ~x162;
  assign n1180 = x33 & ~x161;
  assign n1181 = ~n1179 & ~n1180;
  assign n1182 = ~n1178 & n1181;
  assign n1183 = ~x35 & x163;
  assign n1184 = ~x34 & x162;
  assign n1185 = ~n1183 & ~n1184;
  assign n1186 = ~n1182 & n1185;
  assign n1187 = x36 & ~x164;
  assign n1188 = x35 & ~x163;
  assign n1189 = ~n1187 & ~n1188;
  assign n1190 = ~n1186 & n1189;
  assign n1191 = ~x37 & x165;
  assign n1192 = ~x36 & x164;
  assign n1193 = ~n1191 & ~n1192;
  assign n1194 = ~n1190 & n1193;
  assign n1195 = x38 & ~x166;
  assign n1196 = x37 & ~x165;
  assign n1197 = ~n1195 & ~n1196;
  assign n1198 = ~n1194 & n1197;
  assign n1199 = ~x38 & x166;
  assign n1200 = ~n1198 & ~n1199;
  assign n1201 = ~n1047 & ~n1200;
  assign n1202 = ~x41 & x169;
  assign n1203 = ~x42 & x170;
  assign n1204 = ~n1202 & ~n1203;
  assign n1205 = ~x39 & x167;
  assign n1206 = ~x40 & x168;
  assign n1207 = ~n1205 & ~n1206;
  assign n1208 = n1204 & n1207;
  assign n1209 = ~n1201 & n1208;
  assign n1210 = x41 & ~x169;
  assign n1211 = x40 & ~x168;
  assign n1212 = ~n1210 & ~n1211;
  assign n1213 = n1204 & ~n1212;
  assign n1214 = x43 & ~x171;
  assign n1215 = x42 & ~x170;
  assign n1216 = ~n1214 & ~n1215;
  assign n1217 = ~n1213 & n1216;
  assign n1218 = ~n1209 & n1217;
  assign n1219 = ~x46 & x174;
  assign n1220 = ~x45 & x173;
  assign n1221 = ~n1219 & ~n1220;
  assign n1222 = ~x43 & x171;
  assign n1223 = ~x44 & x172;
  assign n1224 = ~n1222 & ~n1223;
  assign n1225 = n1221 & n1224;
  assign n1226 = ~n1218 & n1225;
  assign n1227 = x45 & ~x173;
  assign n1228 = x44 & ~x172;
  assign n1229 = ~n1227 & ~n1228;
  assign n1230 = n1221 & ~n1229;
  assign n1231 = x46 & ~x174;
  assign n1232 = x47 & ~x175;
  assign n1233 = ~n1231 & ~n1232;
  assign n1234 = ~n1230 & n1233;
  assign n1235 = ~n1226 & n1234;
  assign n1236 = ~x48 & x176;
  assign n1237 = ~x47 & x175;
  assign n1238 = ~n1236 & ~n1237;
  assign n1239 = ~n1235 & n1238;
  assign n1240 = x49 & ~x177;
  assign n1241 = x48 & ~x176;
  assign n1242 = ~n1240 & ~n1241;
  assign n1243 = ~n1239 & n1242;
  assign n1244 = ~x49 & x177;
  assign n1245 = ~n1243 & ~n1244;
  assign n1246 = ~n1046 & ~n1245;
  assign n1247 = ~x51 & x179;
  assign n1248 = ~x50 & x178;
  assign n1249 = ~n1247 & ~n1248;
  assign n1250 = ~n1246 & n1249;
  assign n1251 = x52 & ~x180;
  assign n1252 = x51 & ~x179;
  assign n1253 = ~n1251 & ~n1252;
  assign n1254 = ~n1250 & n1253;
  assign n1255 = ~x53 & x181;
  assign n1256 = ~x52 & x180;
  assign n1257 = ~n1255 & ~n1256;
  assign n1258 = ~n1254 & n1257;
  assign n1259 = x54 & ~x182;
  assign n1260 = x53 & ~x181;
  assign n1261 = ~n1259 & ~n1260;
  assign n1262 = ~n1258 & n1261;
  assign n1263 = ~x55 & x183;
  assign n1264 = ~x54 & x182;
  assign n1265 = ~n1263 & ~n1264;
  assign n1266 = ~n1262 & n1265;
  assign n1267 = x56 & ~x184;
  assign n1268 = x55 & ~x183;
  assign n1269 = ~n1267 & ~n1268;
  assign n1270 = ~n1266 & n1269;
  assign n1271 = ~x56 & x184;
  assign n1272 = ~n1270 & ~n1271;
  assign n1273 = ~n1045 & ~n1272;
  assign n1274 = ~x58 & x186;
  assign n1275 = ~x57 & x185;
  assign n1276 = ~n1274 & ~n1275;
  assign n1277 = ~n1273 & n1276;
  assign n1278 = x59 & ~x187;
  assign n1279 = x58 & ~x186;
  assign n1280 = ~n1278 & ~n1279;
  assign n1281 = ~n1277 & n1280;
  assign n1282 = ~x62 & x190;
  assign n1283 = ~x61 & x189;
  assign n1284 = ~n1282 & ~n1283;
  assign n1285 = ~x59 & x187;
  assign n1286 = ~x60 & x188;
  assign n1287 = ~n1285 & ~n1286;
  assign n1288 = n1284 & n1287;
  assign n1289 = ~n1281 & n1288;
  assign n1290 = x61 & ~x189;
  assign n1291 = x60 & ~x188;
  assign n1292 = ~n1290 & ~n1291;
  assign n1293 = n1284 & ~n1292;
  assign n1294 = x63 & ~x191;
  assign n1295 = x62 & ~x190;
  assign n1296 = ~n1294 & ~n1295;
  assign n1297 = ~n1293 & n1296;
  assign n1298 = ~n1289 & n1297;
  assign n1299 = ~x64 & x192;
  assign n1300 = ~x63 & x191;
  assign n1301 = ~n1299 & ~n1300;
  assign n1302 = ~n1298 & n1301;
  assign n1303 = x64 & ~x192;
  assign n1304 = ~n1302 & ~n1303;
  assign n1305 = ~n1044 & ~n1304;
  assign n1306 = x66 & ~x194;
  assign n1307 = x65 & ~x193;
  assign n1308 = ~n1306 & ~n1307;
  assign n1309 = ~n1305 & n1308;
  assign n1310 = ~x67 & x195;
  assign n1311 = ~x66 & x194;
  assign n1312 = ~n1310 & ~n1311;
  assign n1313 = ~n1309 & n1312;
  assign n1314 = x67 & ~x195;
  assign n1315 = ~n1313 & ~n1314;
  assign n1316 = ~x70 & x198;
  assign n1317 = ~x69 & x197;
  assign n1318 = ~n1316 & ~n1317;
  assign n1319 = ~x68 & x196;
  assign n1320 = n1318 & ~n1319;
  assign n1321 = ~n1315 & n1320;
  assign n1322 = x69 & ~x197;
  assign n1323 = x68 & ~x196;
  assign n1324 = ~n1322 & ~n1323;
  assign n1325 = n1318 & ~n1324;
  assign n1326 = x70 & ~x198;
  assign n1327 = x71 & ~x199;
  assign n1328 = ~n1326 & ~n1327;
  assign n1329 = ~n1325 & n1328;
  assign n1330 = ~n1321 & n1329;
  assign n1331 = ~x72 & x200;
  assign n1332 = ~x71 & x199;
  assign n1333 = ~n1331 & ~n1332;
  assign n1334 = ~n1330 & n1333;
  assign n1335 = x73 & ~x201;
  assign n1336 = x72 & ~x200;
  assign n1337 = ~n1335 & ~n1336;
  assign n1338 = ~n1334 & n1337;
  assign n1339 = ~x74 & x202;
  assign n1340 = ~x73 & x201;
  assign n1341 = ~n1339 & ~n1340;
  assign n1342 = ~n1338 & n1341;
  assign n1343 = x75 & ~x203;
  assign n1344 = x74 & ~x202;
  assign n1345 = ~n1343 & ~n1344;
  assign n1346 = ~n1342 & n1345;
  assign n1347 = ~x76 & x204;
  assign n1348 = ~x75 & x203;
  assign n1349 = ~n1347 & ~n1348;
  assign n1350 = ~n1346 & n1349;
  assign n1351 = x77 & ~x205;
  assign n1352 = x76 & ~x204;
  assign n1353 = ~n1351 & ~n1352;
  assign n1354 = ~n1350 & n1353;
  assign n1355 = ~x78 & x206;
  assign n1356 = ~x77 & x205;
  assign n1357 = ~n1355 & ~n1356;
  assign n1358 = ~n1354 & n1357;
  assign n1359 = x79 & ~x207;
  assign n1360 = x78 & ~x206;
  assign n1361 = ~n1359 & ~n1360;
  assign n1362 = ~n1358 & n1361;
  assign n1363 = ~x80 & x208;
  assign n1364 = ~x79 & x207;
  assign n1365 = ~n1363 & ~n1364;
  assign n1366 = ~n1362 & n1365;
  assign n1367 = x81 & ~x209;
  assign n1368 = x80 & ~x208;
  assign n1369 = ~n1367 & ~n1368;
  assign n1370 = ~n1366 & n1369;
  assign n1371 = ~x81 & x209;
  assign n1372 = ~n1370 & ~n1371;
  assign n1373 = ~n1043 & ~n1372;
  assign n1374 = ~x83 & x211;
  assign n1375 = ~x82 & x210;
  assign n1376 = ~n1374 & ~n1375;
  assign n1377 = ~n1373 & n1376;
  assign n1378 = x84 & ~x212;
  assign n1379 = x83 & ~x211;
  assign n1380 = ~n1378 & ~n1379;
  assign n1381 = ~n1377 & n1380;
  assign n1382 = ~x85 & x213;
  assign n1383 = ~x84 & x212;
  assign n1384 = ~n1382 & ~n1383;
  assign n1385 = ~n1381 & n1384;
  assign n1386 = x86 & ~x214;
  assign n1387 = x85 & ~x213;
  assign n1388 = ~n1386 & ~n1387;
  assign n1389 = ~n1385 & n1388;
  assign n1390 = ~x87 & x215;
  assign n1391 = ~x86 & x214;
  assign n1392 = ~n1390 & ~n1391;
  assign n1393 = ~n1389 & n1392;
  assign n1394 = x88 & ~x216;
  assign n1395 = x87 & ~x215;
  assign n1396 = ~n1394 & ~n1395;
  assign n1397 = ~n1393 & n1396;
  assign n1398 = ~x89 & x217;
  assign n1399 = ~x88 & x216;
  assign n1400 = ~n1398 & ~n1399;
  assign n1401 = ~n1397 & n1400;
  assign n1402 = x90 & ~x218;
  assign n1403 = x89 & ~x217;
  assign n1404 = ~n1402 & ~n1403;
  assign n1405 = ~n1401 & n1404;
  assign n1406 = ~x90 & x218;
  assign n1407 = ~n1405 & ~n1406;
  assign n1408 = ~n1042 & ~n1407;
  assign n1409 = ~x92 & x220;
  assign n1410 = ~x91 & x219;
  assign n1411 = ~n1409 & ~n1410;
  assign n1412 = ~n1408 & n1411;
  assign n1413 = x92 & ~x220;
  assign n1414 = ~n1412 & ~n1413;
  assign n1415 = ~n1041 & ~n1414;
  assign n1416 = x94 & ~x222;
  assign n1417 = x93 & ~x221;
  assign n1418 = ~n1416 & ~n1417;
  assign n1419 = ~n1415 & n1418;
  assign n1420 = ~x94 & x222;
  assign n1421 = ~n1419 & ~n1420;
  assign n1422 = ~n1040 & ~n1421;
  assign n1423 = ~x96 & x224;
  assign n1424 = ~x95 & x223;
  assign n1425 = ~n1423 & ~n1424;
  assign n1426 = ~n1422 & n1425;
  assign n1427 = x97 & ~x225;
  assign n1428 = x96 & ~x224;
  assign n1429 = ~n1427 & ~n1428;
  assign n1430 = ~n1426 & n1429;
  assign n1431 = ~x97 & x225;
  assign n1432 = ~n1430 & ~n1431;
  assign n1433 = ~n1039 & ~n1432;
  assign n1434 = ~x99 & x227;
  assign n1435 = ~x98 & x226;
  assign n1436 = ~n1434 & ~n1435;
  assign n1437 = ~n1433 & n1436;
  assign n1438 = x100 & ~x228;
  assign n1439 = x99 & ~x227;
  assign n1440 = ~n1438 & ~n1439;
  assign n1441 = ~n1437 & n1440;
  assign n1442 = ~x101 & x229;
  assign n1443 = ~x100 & x228;
  assign n1444 = ~n1442 & ~n1443;
  assign n1445 = ~n1441 & n1444;
  assign n1446 = x101 & ~x229;
  assign n1447 = ~n1445 & ~n1446;
  assign n1448 = ~n1038 & ~n1447;
  assign n1449 = x103 & ~x231;
  assign n1450 = x102 & ~x230;
  assign n1451 = ~n1449 & ~n1450;
  assign n1452 = ~n1448 & n1451;
  assign n1453 = ~x104 & x232;
  assign n1454 = ~x103 & x231;
  assign n1455 = ~n1453 & ~n1454;
  assign n1456 = ~n1452 & n1455;
  assign n1457 = x105 & ~x233;
  assign n1458 = x104 & ~x232;
  assign n1459 = ~n1457 & ~n1458;
  assign n1460 = ~n1456 & n1459;
  assign n1461 = ~x105 & x233;
  assign n1462 = ~n1460 & ~n1461;
  assign n1463 = ~n1037 & ~n1462;
  assign n1464 = ~x107 & x235;
  assign n1465 = ~x106 & x234;
  assign n1466 = ~n1464 & ~n1465;
  assign n1467 = ~n1463 & n1466;
  assign n1468 = x108 & ~x236;
  assign n1469 = x107 & ~x235;
  assign n1470 = ~n1468 & ~n1469;
  assign n1471 = ~n1467 & n1470;
  assign n1472 = ~x109 & x237;
  assign n1473 = ~x108 & x236;
  assign n1474 = ~n1472 & ~n1473;
  assign n1475 = ~n1471 & n1474;
  assign n1476 = x109 & ~x237;
  assign n1477 = ~n1475 & ~n1476;
  assign n1478 = ~n1036 & ~n1477;
  assign n1479 = x111 & ~x239;
  assign n1480 = x110 & ~x238;
  assign n1481 = ~n1479 & ~n1480;
  assign n1482 = ~n1478 & n1481;
  assign n1483 = ~x112 & x240;
  assign n1484 = ~x111 & x239;
  assign n1485 = ~n1483 & ~n1484;
  assign n1486 = ~n1482 & n1485;
  assign n1487 = x113 & ~x241;
  assign n1488 = x112 & ~x240;
  assign n1489 = ~n1487 & ~n1488;
  assign n1490 = ~n1486 & n1489;
  assign n1491 = ~x113 & x241;
  assign n1492 = ~n1490 & ~n1491;
  assign n1493 = ~n1035 & ~n1492;
  assign n1494 = ~x115 & x243;
  assign n1495 = ~x114 & x242;
  assign n1496 = ~n1494 & ~n1495;
  assign n1497 = ~n1493 & n1496;
  assign n1498 = x116 & ~x244;
  assign n1499 = x115 & ~x243;
  assign n1500 = ~n1498 & ~n1499;
  assign n1501 = ~n1497 & n1500;
  assign n1502 = ~x116 & x244;
  assign n1503 = ~n1501 & ~n1502;
  assign n1504 = ~n1034 & ~n1503;
  assign n1505 = ~x118 & x246;
  assign n1506 = ~x117 & x245;
  assign n1507 = ~n1505 & ~n1506;
  assign n1508 = ~n1504 & n1507;
  assign n1509 = x119 & ~x247;
  assign n1510 = x118 & ~x246;
  assign n1511 = ~n1509 & ~n1510;
  assign n1512 = ~n1508 & n1511;
  assign n1513 = ~x119 & x247;
  assign n1514 = ~n1512 & ~n1513;
  assign n1515 = ~n1033 & ~n1514;
  assign n1516 = ~x121 & x249;
  assign n1517 = ~x120 & x248;
  assign n1518 = ~n1516 & ~n1517;
  assign n1519 = ~n1515 & n1518;
  assign n1520 = x121 & ~x249;
  assign n1521 = ~n1519 & ~n1520;
  assign n1522 = ~n1032 & ~n1521;
  assign n1523 = x123 & ~x251;
  assign n1524 = x122 & ~x250;
  assign n1525 = ~n1523 & ~n1524;
  assign n1526 = ~n1522 & n1525;
  assign n1527 = ~x125 & x253;
  assign n1528 = ~x126 & x254;
  assign n1529 = ~n1527 & ~n1528;
  assign n1530 = ~x123 & x251;
  assign n1531 = ~x124 & x252;
  assign n1532 = ~n1530 & ~n1531;
  assign n1533 = n1529 & n1532;
  assign n1534 = ~n1526 & n1533;
  assign n1535 = x125 & ~x253;
  assign n1536 = x124 & ~x252;
  assign n1537 = ~n1535 & ~n1536;
  assign n1538 = n1529 & ~n1537;
  assign n1539 = ~x127 & x255;
  assign n1540 = x126 & ~x254;
  assign n1541 = ~n1539 & ~n1540;
  assign n1542 = ~n1538 & n1541;
  assign n1543 = ~n1534 & n1542;
  assign n1544 = x127 & ~x255;
  assign n1545 = ~n1543 & ~n1544;
  assign n1546 = x250 ^ x122;
  assign n1547 = ~n1545 & n1546;
  assign n1548 = n1547 ^ x122;
  assign n1549 = n1031 & ~n1548;
  assign n1550 = x248 ^ x120;
  assign n1551 = ~n1545 & n1550;
  assign n1552 = n1551 ^ x120;
  assign n1553 = x504 ^ x376;
  assign n1554 = ~n1028 & n1553;
  assign n1555 = n1554 ^ x376;
  assign n1556 = n1552 & ~n1555;
  assign n1557 = x238 ^ x110;
  assign n1558 = ~n1545 & n1557;
  assign n1559 = n1558 ^ x110;
  assign n1560 = x494 ^ x366;
  assign n1561 = ~n1028 & n1560;
  assign n1562 = n1561 ^ x366;
  assign n1563 = ~n1559 & n1562;
  assign n1564 = x236 ^ x108;
  assign n1565 = ~n1545 & n1564;
  assign n1566 = n1565 ^ x108;
  assign n1567 = x492 ^ x364;
  assign n1568 = ~n1028 & n1567;
  assign n1569 = n1568 ^ x364;
  assign n1570 = n1566 & ~n1569;
  assign n1571 = x229 ^ x101;
  assign n1572 = ~n1545 & n1571;
  assign n1573 = n1572 ^ x101;
  assign n1574 = x485 ^ x357;
  assign n1575 = ~n1028 & n1574;
  assign n1576 = n1575 ^ x357;
  assign n1577 = ~n1573 & n1576;
  assign n1578 = x225 ^ x97;
  assign n1579 = ~n1545 & n1578;
  assign n1580 = n1579 ^ x97;
  assign n1581 = x481 ^ x353;
  assign n1582 = ~n1028 & n1581;
  assign n1583 = n1582 ^ x353;
  assign n1584 = n1580 & ~n1583;
  assign n1585 = x200 ^ x72;
  assign n1586 = ~n1545 & n1585;
  assign n1587 = n1586 ^ x72;
  assign n1588 = x456 ^ x328;
  assign n1589 = ~n1028 & n1588;
  assign n1590 = n1589 ^ x328;
  assign n1591 = ~n1587 & n1590;
  assign n1592 = x452 ^ x324;
  assign n1593 = ~n1028 & n1592;
  assign n1594 = n1593 ^ x324;
  assign n1595 = x196 ^ x68;
  assign n1596 = ~n1545 & n1595;
  assign n1597 = n1596 ^ x68;
  assign n1598 = ~n1594 & n1597;
  assign n1599 = x441 ^ x313;
  assign n1600 = ~n1028 & n1599;
  assign n1601 = n1600 ^ x313;
  assign n1602 = x185 ^ x57;
  assign n1603 = ~n1545 & n1602;
  assign n1604 = n1603 ^ x57;
  assign n1605 = ~n1601 & n1604;
  assign n1606 = x437 ^ x309;
  assign n1607 = ~n1028 & n1606;
  assign n1608 = n1607 ^ x309;
  assign n1609 = x181 ^ x53;
  assign n1610 = ~n1545 & n1609;
  assign n1611 = n1610 ^ x53;
  assign n1612 = n1608 & ~n1611;
  assign n1613 = x432 ^ x304;
  assign n1614 = ~n1028 & n1613;
  assign n1615 = n1614 ^ x304;
  assign n1616 = x176 ^ x48;
  assign n1617 = ~n1545 & n1616;
  assign n1618 = n1617 ^ x48;
  assign n1619 = n1615 & ~n1618;
  assign n1620 = x174 ^ x46;
  assign n1621 = ~n1545 & n1620;
  assign n1622 = n1621 ^ x46;
  assign n1623 = x430 ^ x302;
  assign n1624 = ~n1028 & n1623;
  assign n1625 = n1624 ^ x302;
  assign n1626 = n1622 & ~n1625;
  assign n1627 = x170 ^ x42;
  assign n1628 = ~n1545 & n1627;
  assign n1629 = n1628 ^ x42;
  assign n1630 = x426 ^ x298;
  assign n1631 = ~n1028 & n1630;
  assign n1632 = n1631 ^ x298;
  assign n1633 = ~n1629 & n1632;
  assign n1634 = x167 ^ x39;
  assign n1635 = ~n1545 & n1634;
  assign n1636 = n1635 ^ x39;
  assign n1637 = x423 ^ x295;
  assign n1638 = ~n1028 & n1637;
  assign n1639 = n1638 ^ x295;
  assign n1640 = ~n1636 & n1639;
  assign n1641 = x421 ^ x293;
  assign n1642 = ~n1028 & n1641;
  assign n1643 = n1642 ^ x293;
  assign n1644 = x165 ^ x37;
  assign n1645 = ~n1545 & n1644;
  assign n1646 = n1645 ^ x37;
  assign n1647 = ~n1643 & n1646;
  assign n1648 = x418 ^ x290;
  assign n1649 = ~n1028 & n1648;
  assign n1650 = n1649 ^ x290;
  assign n1651 = x162 ^ x34;
  assign n1652 = ~n1545 & n1651;
  assign n1653 = n1652 ^ x34;
  assign n1654 = ~n1650 & n1653;
  assign n1655 = x160 ^ x32;
  assign n1656 = ~n1545 & n1655;
  assign n1657 = n1656 ^ x32;
  assign n1658 = x416 ^ x288;
  assign n1659 = ~n1028 & n1658;
  assign n1660 = n1659 ^ x288;
  assign n1661 = ~n1657 & n1660;
  assign n1662 = x414 ^ x286;
  assign n1663 = ~n1028 & n1662;
  assign n1664 = n1663 ^ x286;
  assign n1665 = x158 ^ x30;
  assign n1666 = ~n1545 & n1665;
  assign n1667 = n1666 ^ x30;
  assign n1668 = ~n1664 & n1667;
  assign n1669 = x411 ^ x283;
  assign n1670 = ~n1028 & n1669;
  assign n1671 = n1670 ^ x283;
  assign n1672 = x155 ^ x27;
  assign n1673 = ~n1545 & n1672;
  assign n1674 = n1673 ^ x27;
  assign n1675 = ~n1671 & n1674;
  assign n1676 = x153 ^ x25;
  assign n1677 = ~n1545 & n1676;
  assign n1678 = n1677 ^ x25;
  assign n1679 = x409 ^ x281;
  assign n1680 = ~n1028 & n1679;
  assign n1681 = n1680 ^ x281;
  assign n1682 = ~n1678 & n1681;
  assign n1683 = x405 ^ x277;
  assign n1684 = ~n1028 & n1683;
  assign n1685 = n1684 ^ x277;
  assign n1686 = x149 ^ x21;
  assign n1687 = ~n1545 & n1686;
  assign n1688 = n1687 ^ x21;
  assign n1689 = ~n1685 & n1688;
  assign n1690 = x146 ^ x18;
  assign n1691 = ~n1545 & n1690;
  assign n1692 = n1691 ^ x18;
  assign n1693 = x402 ^ x274;
  assign n1694 = ~n1028 & n1693;
  assign n1695 = n1694 ^ x274;
  assign n1696 = n1692 & ~n1695;
  assign n1697 = x400 ^ x272;
  assign n1698 = ~n1028 & n1697;
  assign n1699 = n1698 ^ x272;
  assign n1700 = x144 ^ x16;
  assign n1701 = ~n1545 & n1700;
  assign n1702 = n1701 ^ x16;
  assign n1703 = n1699 & ~n1702;
  assign n1704 = x392 ^ x264;
  assign n1705 = ~n1028 & n1704;
  assign n1706 = n1705 ^ x264;
  assign n1707 = x136 ^ x8;
  assign n1708 = ~n1545 & n1707;
  assign n1709 = n1708 ^ x8;
  assign n1710 = ~n1706 & n1709;
  assign n1711 = x133 ^ x5;
  assign n1712 = ~n1545 & n1711;
  assign n1713 = n1712 ^ x5;
  assign n1714 = x389 ^ x261;
  assign n1715 = ~n1028 & n1714;
  assign n1716 = n1715 ^ x261;
  assign n1717 = n1713 & ~n1716;
  assign n1718 = x385 ^ x257;
  assign n1719 = ~n1028 & n1718;
  assign n1720 = n1719 ^ x257;
  assign n1721 = x129 ^ x1;
  assign n1722 = ~n1545 & n1721;
  assign n1723 = n1722 ^ x1;
  assign n1724 = n1720 & ~n1723;
  assign n1725 = x384 ^ x256;
  assign n1726 = ~n1028 & n1725;
  assign n1727 = n1726 ^ x256;
  assign n1728 = x128 ^ x0;
  assign n1729 = ~n1545 & n1728;
  assign n1730 = n1729 ^ x0;
  assign n1731 = ~n1727 & n1730;
  assign n1732 = ~n1724 & n1731;
  assign n1733 = x386 ^ x258;
  assign n1734 = ~n1028 & n1733;
  assign n1735 = n1734 ^ x258;
  assign n1736 = x130 ^ x2;
  assign n1737 = ~n1545 & n1736;
  assign n1738 = n1737 ^ x2;
  assign n1739 = ~n1735 & n1738;
  assign n1740 = ~n1720 & n1723;
  assign n1741 = ~n1739 & ~n1740;
  assign n1742 = ~n1732 & n1741;
  assign n1743 = n1735 & ~n1738;
  assign n1744 = x387 ^ x259;
  assign n1745 = ~n1028 & n1744;
  assign n1746 = n1745 ^ x259;
  assign n1747 = x131 ^ x3;
  assign n1748 = ~n1545 & n1747;
  assign n1749 = n1748 ^ x3;
  assign n1750 = n1746 & ~n1749;
  assign n1751 = ~n1743 & ~n1750;
  assign n1752 = ~n1742 & n1751;
  assign n1753 = ~n1746 & n1749;
  assign n1754 = x132 ^ x4;
  assign n1755 = ~n1545 & n1754;
  assign n1756 = n1755 ^ x4;
  assign n1757 = x388 ^ x260;
  assign n1758 = ~n1028 & n1757;
  assign n1759 = n1758 ^ x260;
  assign n1760 = n1756 & ~n1759;
  assign n1761 = ~n1753 & ~n1760;
  assign n1762 = ~n1752 & n1761;
  assign n1763 = ~n1756 & n1759;
  assign n1764 = ~n1762 & ~n1763;
  assign n1765 = ~n1717 & ~n1764;
  assign n1766 = ~n1713 & n1716;
  assign n1767 = x390 ^ x262;
  assign n1768 = ~n1028 & n1767;
  assign n1769 = n1768 ^ x262;
  assign n1770 = x134 ^ x6;
  assign n1771 = ~n1545 & n1770;
  assign n1772 = n1771 ^ x6;
  assign n1773 = n1769 & ~n1772;
  assign n1774 = ~n1766 & ~n1773;
  assign n1775 = ~n1765 & n1774;
  assign n1776 = ~n1769 & n1772;
  assign n1777 = x135 ^ x7;
  assign n1778 = ~n1545 & n1777;
  assign n1779 = n1778 ^ x7;
  assign n1780 = x391 ^ x263;
  assign n1781 = ~n1028 & n1780;
  assign n1782 = n1781 ^ x263;
  assign n1783 = n1779 & ~n1782;
  assign n1784 = ~n1776 & ~n1783;
  assign n1785 = ~n1775 & n1784;
  assign n1786 = ~n1779 & n1782;
  assign n1787 = ~n1785 & ~n1786;
  assign n1788 = ~n1710 & ~n1787;
  assign n1789 = n1706 & ~n1709;
  assign n1790 = x393 ^ x265;
  assign n1791 = ~n1028 & n1790;
  assign n1792 = n1791 ^ x265;
  assign n1793 = x137 ^ x9;
  assign n1794 = ~n1545 & n1793;
  assign n1795 = n1794 ^ x9;
  assign n1796 = n1792 & ~n1795;
  assign n1797 = ~n1789 & ~n1796;
  assign n1798 = ~n1788 & n1797;
  assign n1799 = ~n1792 & n1795;
  assign n1800 = x138 ^ x10;
  assign n1801 = ~n1545 & n1800;
  assign n1802 = n1801 ^ x10;
  assign n1803 = x394 ^ x266;
  assign n1804 = ~n1028 & n1803;
  assign n1805 = n1804 ^ x266;
  assign n1806 = n1802 & ~n1805;
  assign n1807 = ~n1799 & ~n1806;
  assign n1808 = ~n1798 & n1807;
  assign n1809 = ~n1802 & n1805;
  assign n1810 = x139 ^ x11;
  assign n1811 = ~n1545 & n1810;
  assign n1812 = n1811 ^ x11;
  assign n1813 = x395 ^ x267;
  assign n1814 = ~n1028 & n1813;
  assign n1815 = n1814 ^ x267;
  assign n1816 = ~n1812 & n1815;
  assign n1817 = ~n1809 & ~n1816;
  assign n1818 = ~n1808 & n1817;
  assign n1819 = n1812 & ~n1815;
  assign n1820 = x140 ^ x12;
  assign n1821 = ~n1545 & n1820;
  assign n1822 = n1821 ^ x12;
  assign n1823 = x396 ^ x268;
  assign n1824 = ~n1028 & n1823;
  assign n1825 = n1824 ^ x268;
  assign n1826 = n1822 & ~n1825;
  assign n1827 = ~n1819 & ~n1826;
  assign n1828 = ~n1818 & n1827;
  assign n1829 = ~n1822 & n1825;
  assign n1830 = x397 ^ x269;
  assign n1831 = ~n1028 & n1830;
  assign n1832 = n1831 ^ x269;
  assign n1833 = x141 ^ x13;
  assign n1834 = ~n1545 & n1833;
  assign n1835 = n1834 ^ x13;
  assign n1836 = n1832 & ~n1835;
  assign n1837 = ~n1829 & ~n1836;
  assign n1838 = ~n1828 & n1837;
  assign n1839 = ~n1832 & n1835;
  assign n1840 = x398 ^ x270;
  assign n1841 = ~n1028 & n1840;
  assign n1842 = n1841 ^ x270;
  assign n1843 = x142 ^ x14;
  assign n1844 = ~n1545 & n1843;
  assign n1845 = n1844 ^ x14;
  assign n1846 = ~n1842 & n1845;
  assign n1847 = ~n1839 & ~n1846;
  assign n1848 = ~n1838 & n1847;
  assign n1849 = x143 ^ x15;
  assign n1850 = ~n1545 & n1849;
  assign n1851 = n1850 ^ x15;
  assign n1852 = x399 ^ x271;
  assign n1853 = ~n1028 & n1852;
  assign n1854 = n1853 ^ x271;
  assign n1855 = ~n1851 & n1854;
  assign n1856 = n1842 & ~n1845;
  assign n1857 = ~n1855 & ~n1856;
  assign n1858 = ~n1848 & n1857;
  assign n1859 = n1851 & ~n1854;
  assign n1860 = ~n1858 & ~n1859;
  assign n1861 = ~n1703 & ~n1860;
  assign n1862 = ~n1699 & n1702;
  assign n1863 = x145 ^ x17;
  assign n1864 = ~n1545 & n1863;
  assign n1865 = n1864 ^ x17;
  assign n1866 = x401 ^ x273;
  assign n1867 = ~n1028 & n1866;
  assign n1868 = n1867 ^ x273;
  assign n1869 = n1865 & ~n1868;
  assign n1870 = ~n1862 & ~n1869;
  assign n1871 = ~n1861 & n1870;
  assign n1872 = ~n1865 & n1868;
  assign n1873 = ~n1871 & ~n1872;
  assign n1874 = ~n1696 & ~n1873;
  assign n1875 = ~n1692 & n1695;
  assign n1876 = x403 ^ x275;
  assign n1877 = ~n1028 & n1876;
  assign n1878 = n1877 ^ x275;
  assign n1879 = x147 ^ x19;
  assign n1880 = ~n1545 & n1879;
  assign n1881 = n1880 ^ x19;
  assign n1882 = n1878 & ~n1881;
  assign n1883 = ~n1875 & ~n1882;
  assign n1884 = ~n1874 & n1883;
  assign n1885 = ~n1878 & n1881;
  assign n1886 = x148 ^ x20;
  assign n1887 = ~n1545 & n1886;
  assign n1888 = n1887 ^ x20;
  assign n1889 = x404 ^ x276;
  assign n1890 = ~n1028 & n1889;
  assign n1891 = n1890 ^ x276;
  assign n1892 = n1888 & ~n1891;
  assign n1893 = ~n1885 & ~n1892;
  assign n1894 = ~n1884 & n1893;
  assign n1895 = ~n1888 & n1891;
  assign n1896 = ~n1894 & ~n1895;
  assign n1897 = ~n1689 & ~n1896;
  assign n1898 = n1685 & ~n1688;
  assign n1899 = x406 ^ x278;
  assign n1900 = ~n1028 & n1899;
  assign n1901 = n1900 ^ x278;
  assign n1902 = x150 ^ x22;
  assign n1903 = ~n1545 & n1902;
  assign n1904 = n1903 ^ x22;
  assign n1905 = n1901 & ~n1904;
  assign n1906 = ~n1898 & ~n1905;
  assign n1907 = ~n1897 & n1906;
  assign n1908 = ~n1901 & n1904;
  assign n1909 = x407 ^ x279;
  assign n1910 = ~n1028 & n1909;
  assign n1911 = n1910 ^ x279;
  assign n1912 = x151 ^ x23;
  assign n1913 = ~n1545 & n1912;
  assign n1914 = n1913 ^ x23;
  assign n1915 = ~n1911 & n1914;
  assign n1916 = ~n1908 & ~n1915;
  assign n1917 = ~n1907 & n1916;
  assign n1918 = n1911 & ~n1914;
  assign n1919 = x152 ^ x24;
  assign n1920 = ~n1545 & n1919;
  assign n1921 = n1920 ^ x24;
  assign n1922 = x408 ^ x280;
  assign n1923 = ~n1028 & n1922;
  assign n1924 = n1923 ^ x280;
  assign n1925 = ~n1921 & n1924;
  assign n1926 = ~n1918 & ~n1925;
  assign n1927 = ~n1917 & n1926;
  assign n1928 = n1921 & ~n1924;
  assign n1929 = ~n1927 & ~n1928;
  assign n1930 = ~n1682 & ~n1929;
  assign n1931 = x154 ^ x26;
  assign n1932 = ~n1545 & n1931;
  assign n1933 = n1932 ^ x26;
  assign n1934 = x410 ^ x282;
  assign n1935 = ~n1028 & n1934;
  assign n1936 = n1935 ^ x282;
  assign n1937 = n1933 & ~n1936;
  assign n1938 = n1678 & ~n1681;
  assign n1939 = ~n1937 & ~n1938;
  assign n1940 = ~n1930 & n1939;
  assign n1941 = ~n1933 & n1936;
  assign n1942 = ~n1940 & ~n1941;
  assign n1943 = ~n1675 & ~n1942;
  assign n1944 = n1671 & ~n1674;
  assign n1945 = x156 ^ x28;
  assign n1946 = ~n1545 & n1945;
  assign n1947 = n1946 ^ x28;
  assign n1948 = x412 ^ x284;
  assign n1949 = ~n1028 & n1948;
  assign n1950 = n1949 ^ x284;
  assign n1951 = ~n1947 & n1950;
  assign n1952 = ~n1944 & ~n1951;
  assign n1953 = ~n1943 & n1952;
  assign n1954 = n1947 & ~n1950;
  assign n1955 = x157 ^ x29;
  assign n1956 = ~n1545 & n1955;
  assign n1957 = n1956 ^ x29;
  assign n1958 = x413 ^ x285;
  assign n1959 = ~n1028 & n1958;
  assign n1960 = n1959 ^ x285;
  assign n1961 = n1957 & ~n1960;
  assign n1962 = ~n1954 & ~n1961;
  assign n1963 = ~n1953 & n1962;
  assign n1964 = ~n1957 & n1960;
  assign n1965 = ~n1963 & ~n1964;
  assign n1966 = ~n1668 & ~n1965;
  assign n1967 = n1664 & ~n1667;
  assign n1968 = x159 ^ x31;
  assign n1969 = ~n1545 & n1968;
  assign n1970 = n1969 ^ x31;
  assign n1971 = x415 ^ x287;
  assign n1972 = ~n1028 & n1971;
  assign n1973 = n1972 ^ x287;
  assign n1974 = ~n1970 & n1973;
  assign n1975 = ~n1967 & ~n1974;
  assign n1976 = ~n1966 & n1975;
  assign n1977 = n1970 & ~n1973;
  assign n1978 = ~n1976 & ~n1977;
  assign n1979 = ~n1661 & ~n1978;
  assign n1980 = x161 ^ x33;
  assign n1981 = ~n1545 & n1980;
  assign n1982 = n1981 ^ x33;
  assign n1983 = x417 ^ x289;
  assign n1984 = ~n1028 & n1983;
  assign n1985 = n1984 ^ x289;
  assign n1986 = n1982 & ~n1985;
  assign n1987 = n1657 & ~n1660;
  assign n1988 = ~n1986 & ~n1987;
  assign n1989 = ~n1979 & n1988;
  assign n1990 = ~n1982 & n1985;
  assign n1991 = ~n1989 & ~n1990;
  assign n1992 = ~n1654 & ~n1991;
  assign n1993 = n1650 & ~n1653;
  assign n1994 = x163 ^ x35;
  assign n1995 = ~n1545 & n1994;
  assign n1996 = n1995 ^ x35;
  assign n1997 = x419 ^ x291;
  assign n1998 = ~n1028 & n1997;
  assign n1999 = n1998 ^ x291;
  assign n2000 = ~n1996 & n1999;
  assign n2001 = ~n1993 & ~n2000;
  assign n2002 = ~n1992 & n2001;
  assign n2003 = n1996 & ~n1999;
  assign n2004 = x164 ^ x36;
  assign n2005 = ~n1545 & n2004;
  assign n2006 = n2005 ^ x36;
  assign n2007 = x420 ^ x292;
  assign n2008 = ~n1028 & n2007;
  assign n2009 = n2008 ^ x292;
  assign n2010 = n2006 & ~n2009;
  assign n2011 = ~n2003 & ~n2010;
  assign n2012 = ~n2002 & n2011;
  assign n2013 = ~n2006 & n2009;
  assign n2014 = ~n2012 & ~n2013;
  assign n2015 = ~n1647 & ~n2014;
  assign n2016 = n1643 & ~n1646;
  assign n2017 = x166 ^ x38;
  assign n2018 = ~n1545 & n2017;
  assign n2019 = n2018 ^ x38;
  assign n2020 = x422 ^ x294;
  assign n2021 = ~n1028 & n2020;
  assign n2022 = n2021 ^ x294;
  assign n2023 = ~n2019 & n2022;
  assign n2024 = ~n2016 & ~n2023;
  assign n2025 = ~n2015 & n2024;
  assign n2026 = n2019 & ~n2022;
  assign n2027 = ~n2025 & ~n2026;
  assign n2028 = ~n1640 & ~n2027;
  assign n2029 = n1636 & ~n1639;
  assign n2030 = x168 ^ x40;
  assign n2031 = ~n1545 & n2030;
  assign n2032 = n2031 ^ x40;
  assign n2033 = x424 ^ x296;
  assign n2034 = ~n1028 & n2033;
  assign n2035 = n2034 ^ x296;
  assign n2036 = n2032 & ~n2035;
  assign n2037 = ~n2029 & ~n2036;
  assign n2038 = ~n2028 & n2037;
  assign n2039 = ~n2032 & n2035;
  assign n2040 = x169 ^ x41;
  assign n2041 = ~n1545 & n2040;
  assign n2042 = n2041 ^ x41;
  assign n2043 = x425 ^ x297;
  assign n2044 = ~n1028 & n2043;
  assign n2045 = n2044 ^ x297;
  assign n2046 = ~n2042 & n2045;
  assign n2047 = ~n2039 & ~n2046;
  assign n2048 = ~n2038 & n2047;
  assign n2049 = n2042 & ~n2045;
  assign n2050 = ~n2048 & ~n2049;
  assign n2051 = ~n1633 & ~n2050;
  assign n2052 = n1629 & ~n1632;
  assign n2053 = x427 ^ x299;
  assign n2054 = ~n1028 & n2053;
  assign n2055 = n2054 ^ x299;
  assign n2056 = x171 ^ x43;
  assign n2057 = ~n1545 & n2056;
  assign n2058 = n2057 ^ x43;
  assign n2059 = ~n2055 & n2058;
  assign n2060 = ~n2052 & ~n2059;
  assign n2061 = ~n2051 & n2060;
  assign n2062 = n2055 & ~n2058;
  assign n2063 = x428 ^ x300;
  assign n2064 = ~n1028 & n2063;
  assign n2065 = n2064 ^ x300;
  assign n2066 = x172 ^ x44;
  assign n2067 = ~n1545 & n2066;
  assign n2068 = n2067 ^ x44;
  assign n2069 = n2065 & ~n2068;
  assign n2070 = ~n2062 & ~n2069;
  assign n2071 = ~n2061 & n2070;
  assign n2072 = ~n2065 & n2068;
  assign n2073 = x173 ^ x45;
  assign n2074 = ~n1545 & n2073;
  assign n2075 = n2074 ^ x45;
  assign n2076 = x429 ^ x301;
  assign n2077 = ~n1028 & n2076;
  assign n2078 = n2077 ^ x301;
  assign n2079 = n2075 & ~n2078;
  assign n2080 = ~n2072 & ~n2079;
  assign n2081 = ~n2071 & n2080;
  assign n2082 = ~n2075 & n2078;
  assign n2083 = ~n2081 & ~n2082;
  assign n2084 = ~n1626 & ~n2083;
  assign n2085 = ~n1622 & n1625;
  assign n2086 = x175 ^ x47;
  assign n2087 = ~n1545 & n2086;
  assign n2088 = n2087 ^ x47;
  assign n2089 = x431 ^ x303;
  assign n2090 = ~n1028 & n2089;
  assign n2091 = n2090 ^ x303;
  assign n2092 = ~n2088 & n2091;
  assign n2093 = ~n2085 & ~n2092;
  assign n2094 = ~n2084 & n2093;
  assign n2095 = n2088 & ~n2091;
  assign n2096 = ~n2094 & ~n2095;
  assign n2097 = ~n1619 & ~n2096;
  assign n2098 = ~n1615 & n1618;
  assign n2099 = x177 ^ x49;
  assign n2100 = ~n1545 & n2099;
  assign n2101 = n2100 ^ x49;
  assign n2102 = x433 ^ x305;
  assign n2103 = ~n1028 & n2102;
  assign n2104 = n2103 ^ x305;
  assign n2105 = n2101 & ~n2104;
  assign n2106 = ~n2098 & ~n2105;
  assign n2107 = ~n2097 & n2106;
  assign n2108 = ~n2101 & n2104;
  assign n2109 = x434 ^ x306;
  assign n2110 = ~n1028 & n2109;
  assign n2111 = n2110 ^ x306;
  assign n2112 = x178 ^ x50;
  assign n2113 = ~n1545 & n2112;
  assign n2114 = n2113 ^ x50;
  assign n2115 = n2111 & ~n2114;
  assign n2116 = ~n2108 & ~n2115;
  assign n2117 = ~n2107 & n2116;
  assign n2118 = ~n2111 & n2114;
  assign n2119 = x435 ^ x307;
  assign n2120 = ~n1028 & n2119;
  assign n2121 = n2120 ^ x307;
  assign n2122 = x179 ^ x51;
  assign n2123 = ~n1545 & n2122;
  assign n2124 = n2123 ^ x51;
  assign n2125 = ~n2121 & n2124;
  assign n2126 = ~n2118 & ~n2125;
  assign n2127 = ~n2117 & n2126;
  assign n2128 = x180 ^ x52;
  assign n2129 = ~n1545 & n2128;
  assign n2130 = n2129 ^ x52;
  assign n2131 = x436 ^ x308;
  assign n2132 = ~n1028 & n2131;
  assign n2133 = n2132 ^ x308;
  assign n2134 = ~n2130 & n2133;
  assign n2135 = n2121 & ~n2124;
  assign n2136 = ~n2134 & ~n2135;
  assign n2137 = ~n2127 & n2136;
  assign n2138 = n2130 & ~n2133;
  assign n2139 = ~n2137 & ~n2138;
  assign n2140 = ~n1612 & ~n2139;
  assign n2141 = ~n1608 & n1611;
  assign n2142 = x182 ^ x54;
  assign n2143 = ~n1545 & n2142;
  assign n2144 = n2143 ^ x54;
  assign n2145 = x438 ^ x310;
  assign n2146 = ~n1028 & n2145;
  assign n2147 = n2146 ^ x310;
  assign n2148 = n2144 & ~n2147;
  assign n2149 = ~n2141 & ~n2148;
  assign n2150 = ~n2140 & n2149;
  assign n2151 = ~n2144 & n2147;
  assign n2152 = x439 ^ x311;
  assign n2153 = ~n1028 & n2152;
  assign n2154 = n2153 ^ x311;
  assign n2155 = x183 ^ x55;
  assign n2156 = ~n1545 & n2155;
  assign n2157 = n2156 ^ x55;
  assign n2158 = n2154 & ~n2157;
  assign n2159 = ~n2151 & ~n2158;
  assign n2160 = ~n2150 & n2159;
  assign n2161 = x184 ^ x56;
  assign n2162 = ~n1545 & n2161;
  assign n2163 = n2162 ^ x56;
  assign n2164 = x440 ^ x312;
  assign n2165 = ~n1028 & n2164;
  assign n2166 = n2165 ^ x312;
  assign n2167 = n2163 & ~n2166;
  assign n2168 = ~n2154 & n2157;
  assign n2169 = ~n2167 & ~n2168;
  assign n2170 = ~n2160 & n2169;
  assign n2171 = ~n2163 & n2166;
  assign n2172 = ~n2170 & ~n2171;
  assign n2173 = ~n1605 & ~n2172;
  assign n2174 = n1601 & ~n1604;
  assign n2175 = x442 ^ x314;
  assign n2176 = ~n1028 & n2175;
  assign n2177 = n2176 ^ x314;
  assign n2178 = x186 ^ x58;
  assign n2179 = ~n1545 & n2178;
  assign n2180 = n2179 ^ x58;
  assign n2181 = n2177 & ~n2180;
  assign n2182 = ~n2174 & ~n2181;
  assign n2183 = ~n2173 & n2182;
  assign n2184 = ~n2177 & n2180;
  assign n2185 = x443 ^ x315;
  assign n2186 = ~n1028 & n2185;
  assign n2187 = n2186 ^ x315;
  assign n2188 = x187 ^ x59;
  assign n2189 = ~n1545 & n2188;
  assign n2190 = n2189 ^ x59;
  assign n2191 = ~n2187 & n2190;
  assign n2192 = ~n2184 & ~n2191;
  assign n2193 = ~n2183 & n2192;
  assign n2194 = n2187 & ~n2190;
  assign n2195 = x188 ^ x60;
  assign n2196 = ~n1545 & n2195;
  assign n2197 = n2196 ^ x60;
  assign n2198 = x444 ^ x316;
  assign n2199 = ~n1028 & n2198;
  assign n2200 = n2199 ^ x316;
  assign n2201 = ~n2197 & n2200;
  assign n2202 = ~n2194 & ~n2201;
  assign n2203 = ~n2193 & n2202;
  assign n2204 = n2197 & ~n2200;
  assign n2205 = x445 ^ x317;
  assign n2206 = ~n1028 & n2205;
  assign n2207 = n2206 ^ x317;
  assign n2208 = x189 ^ x61;
  assign n2209 = ~n1545 & n2208;
  assign n2210 = n2209 ^ x61;
  assign n2211 = ~n2207 & n2210;
  assign n2212 = ~n2204 & ~n2211;
  assign n2213 = ~n2203 & n2212;
  assign n2214 = n2207 & ~n2210;
  assign n2215 = x190 ^ x62;
  assign n2216 = ~n1545 & n2215;
  assign n2217 = n2216 ^ x62;
  assign n2218 = x446 ^ x318;
  assign n2219 = ~n1028 & n2218;
  assign n2220 = n2219 ^ x318;
  assign n2221 = ~n2217 & n2220;
  assign n2222 = ~n2214 & ~n2221;
  assign n2223 = ~n2213 & n2222;
  assign n2224 = n2217 & ~n2220;
  assign n2225 = x191 ^ x63;
  assign n2226 = ~n1545 & n2225;
  assign n2227 = n2226 ^ x63;
  assign n2228 = n780 & ~n1028;
  assign n2229 = n2228 ^ x319;
  assign n2230 = n2227 & ~n2229;
  assign n2231 = ~n2224 & ~n2230;
  assign n2232 = ~n2223 & n2231;
  assign n2233 = ~n2227 & n2229;
  assign n2234 = x192 ^ x64;
  assign n2235 = ~n1545 & n2234;
  assign n2236 = n2235 ^ x64;
  assign n2237 = x448 ^ x320;
  assign n2238 = ~n1028 & n2237;
  assign n2239 = n2238 ^ x320;
  assign n2240 = ~n2236 & n2239;
  assign n2241 = ~n2233 & ~n2240;
  assign n2242 = ~n2232 & n2241;
  assign n2243 = n2236 & ~n2239;
  assign n2244 = x193 ^ x65;
  assign n2245 = ~n1545 & n2244;
  assign n2246 = n2245 ^ x65;
  assign n2247 = x449 ^ x321;
  assign n2248 = ~n1028 & n2247;
  assign n2249 = n2248 ^ x321;
  assign n2250 = n2246 & ~n2249;
  assign n2251 = ~n2243 & ~n2250;
  assign n2252 = ~n2242 & n2251;
  assign n2253 = ~n2246 & n2249;
  assign n2254 = x194 ^ x66;
  assign n2255 = ~n1545 & n2254;
  assign n2256 = n2255 ^ x66;
  assign n2257 = x450 ^ x322;
  assign n2258 = ~n1028 & n2257;
  assign n2259 = n2258 ^ x322;
  assign n2260 = ~n2256 & n2259;
  assign n2261 = ~n2253 & ~n2260;
  assign n2262 = ~n2252 & n2261;
  assign n2263 = n2256 & ~n2259;
  assign n2264 = x195 ^ x67;
  assign n2265 = ~n1545 & n2264;
  assign n2266 = n2265 ^ x67;
  assign n2267 = x451 ^ x323;
  assign n2268 = ~n1028 & n2267;
  assign n2269 = n2268 ^ x323;
  assign n2270 = n2266 & ~n2269;
  assign n2271 = ~n2263 & ~n2270;
  assign n2272 = ~n2262 & n2271;
  assign n2273 = ~n2266 & n2269;
  assign n2274 = ~n2272 & ~n2273;
  assign n2275 = ~n1598 & ~n2274;
  assign n2276 = x197 ^ x69;
  assign n2277 = ~n1545 & n2276;
  assign n2278 = n2277 ^ x69;
  assign n2279 = x453 ^ x325;
  assign n2280 = ~n1028 & n2279;
  assign n2281 = n2280 ^ x325;
  assign n2282 = ~n2278 & n2281;
  assign n2283 = n1594 & ~n1597;
  assign n2284 = ~n2282 & ~n2283;
  assign n2285 = ~n2275 & n2284;
  assign n2286 = n2278 & ~n2281;
  assign n2287 = x198 ^ x70;
  assign n2288 = ~n1545 & n2287;
  assign n2289 = n2288 ^ x70;
  assign n2290 = x454 ^ x326;
  assign n2291 = ~n1028 & n2290;
  assign n2292 = n2291 ^ x326;
  assign n2293 = n2289 & ~n2292;
  assign n2294 = ~n2286 & ~n2293;
  assign n2295 = ~n2285 & n2294;
  assign n2296 = ~n2289 & n2292;
  assign n2297 = x199 ^ x71;
  assign n2298 = ~n1545 & n2297;
  assign n2299 = n2298 ^ x71;
  assign n2300 = x455 ^ x327;
  assign n2301 = ~n1028 & n2300;
  assign n2302 = n2301 ^ x327;
  assign n2303 = ~n2299 & n2302;
  assign n2304 = ~n2296 & ~n2303;
  assign n2305 = ~n2295 & n2304;
  assign n2306 = n2299 & ~n2302;
  assign n2307 = ~n2305 & ~n2306;
  assign n2308 = ~n1591 & ~n2307;
  assign n2309 = n1587 & ~n1590;
  assign n2310 = x457 ^ x329;
  assign n2311 = ~n1028 & n2310;
  assign n2312 = n2311 ^ x329;
  assign n2313 = x201 ^ x73;
  assign n2314 = ~n1545 & n2313;
  assign n2315 = n2314 ^ x73;
  assign n2316 = ~n2312 & n2315;
  assign n2317 = ~n2309 & ~n2316;
  assign n2318 = ~n2308 & n2317;
  assign n2319 = n2312 & ~n2315;
  assign n2320 = x202 ^ x74;
  assign n2321 = ~n1545 & n2320;
  assign n2322 = n2321 ^ x74;
  assign n2323 = x458 ^ x330;
  assign n2324 = ~n1028 & n2323;
  assign n2325 = n2324 ^ x330;
  assign n2326 = ~n2322 & n2325;
  assign n2327 = ~n2319 & ~n2326;
  assign n2328 = ~n2318 & n2327;
  assign n2329 = x459 ^ x331;
  assign n2330 = ~n1028 & n2329;
  assign n2331 = n2330 ^ x331;
  assign n2332 = x203 ^ x75;
  assign n2333 = ~n1545 & n2332;
  assign n2334 = n2333 ^ x75;
  assign n2335 = ~n2331 & n2334;
  assign n2336 = n2322 & ~n2325;
  assign n2337 = ~n2335 & ~n2336;
  assign n2338 = ~n2328 & n2337;
  assign n2339 = x204 ^ x76;
  assign n2340 = ~n1545 & n2339;
  assign n2341 = n2340 ^ x76;
  assign n2342 = x460 ^ x332;
  assign n2343 = ~n1028 & n2342;
  assign n2344 = n2343 ^ x332;
  assign n2345 = ~n2341 & n2344;
  assign n2346 = n2331 & ~n2334;
  assign n2347 = ~n2345 & ~n2346;
  assign n2348 = ~n2338 & n2347;
  assign n2349 = x461 ^ x333;
  assign n2350 = ~n1028 & n2349;
  assign n2351 = n2350 ^ x333;
  assign n2352 = x205 ^ x77;
  assign n2353 = ~n1545 & n2352;
  assign n2354 = n2353 ^ x77;
  assign n2355 = ~n2351 & n2354;
  assign n2356 = n2341 & ~n2344;
  assign n2357 = ~n2355 & ~n2356;
  assign n2358 = ~n2348 & n2357;
  assign n2359 = x462 ^ x334;
  assign n2360 = ~n1028 & n2359;
  assign n2361 = n2360 ^ x334;
  assign n2362 = x206 ^ x78;
  assign n2363 = ~n1545 & n2362;
  assign n2364 = n2363 ^ x78;
  assign n2365 = n2361 & ~n2364;
  assign n2366 = n2351 & ~n2354;
  assign n2367 = ~n2365 & ~n2366;
  assign n2368 = ~n2358 & n2367;
  assign n2369 = ~n2361 & n2364;
  assign n2370 = ~n2368 & ~n2369;
  assign n2371 = x207 ^ x79;
  assign n2372 = ~n1545 & n2371;
  assign n2373 = n2372 ^ x79;
  assign n2374 = x463 ^ x335;
  assign n2375 = ~n1028 & n2374;
  assign n2376 = n2375 ^ x335;
  assign n2377 = ~n2373 & n2376;
  assign n2378 = ~n2370 & ~n2377;
  assign n2379 = x208 ^ x80;
  assign n2380 = ~n1545 & n2379;
  assign n2381 = n2380 ^ x80;
  assign n2382 = x464 ^ x336;
  assign n2383 = ~n1028 & n2382;
  assign n2384 = n2383 ^ x336;
  assign n2385 = n2381 & ~n2384;
  assign n2386 = n2373 & ~n2376;
  assign n2387 = ~n2385 & ~n2386;
  assign n2388 = ~n2378 & n2387;
  assign n2389 = ~n2381 & n2384;
  assign n2390 = x209 ^ x81;
  assign n2391 = ~n1545 & n2390;
  assign n2392 = n2391 ^ x81;
  assign n2393 = x465 ^ x337;
  assign n2394 = ~n1028 & n2393;
  assign n2395 = n2394 ^ x337;
  assign n2396 = ~n2392 & n2395;
  assign n2397 = ~n2389 & ~n2396;
  assign n2398 = ~n2388 & n2397;
  assign n2399 = n2392 & ~n2395;
  assign n2400 = ~n2398 & ~n2399;
  assign n2401 = x466 ^ x338;
  assign n2402 = ~n1028 & n2401;
  assign n2403 = n2402 ^ x338;
  assign n2404 = x210 ^ x82;
  assign n2405 = ~n1545 & n2404;
  assign n2406 = n2405 ^ x82;
  assign n2407 = n2403 & ~n2406;
  assign n2408 = ~n2400 & ~n2407;
  assign n2409 = x211 ^ x83;
  assign n2410 = ~n1545 & n2409;
  assign n2411 = n2410 ^ x83;
  assign n2412 = x467 ^ x339;
  assign n2413 = ~n1028 & n2412;
  assign n2414 = n2413 ^ x339;
  assign n2415 = n2411 & ~n2414;
  assign n2416 = ~n2403 & n2406;
  assign n2417 = ~n2415 & ~n2416;
  assign n2418 = ~n2408 & n2417;
  assign n2419 = x212 ^ x84;
  assign n2420 = ~n1545 & n2419;
  assign n2421 = n2420 ^ x84;
  assign n2422 = x468 ^ x340;
  assign n2423 = ~n1028 & n2422;
  assign n2424 = n2423 ^ x340;
  assign n2425 = ~n2421 & n2424;
  assign n2426 = ~n2411 & n2414;
  assign n2427 = ~n2425 & ~n2426;
  assign n2428 = ~n2418 & n2427;
  assign n2429 = x213 ^ x85;
  assign n2430 = ~n1545 & n2429;
  assign n2431 = n2430 ^ x85;
  assign n2432 = x469 ^ x341;
  assign n2433 = ~n1028 & n2432;
  assign n2434 = n2433 ^ x341;
  assign n2435 = n2431 & ~n2434;
  assign n2436 = n2421 & ~n2424;
  assign n2437 = ~n2435 & ~n2436;
  assign n2438 = ~n2428 & n2437;
  assign n2439 = x470 ^ x342;
  assign n2440 = ~n1028 & n2439;
  assign n2441 = n2440 ^ x342;
  assign n2442 = x214 ^ x86;
  assign n2443 = ~n1545 & n2442;
  assign n2444 = n2443 ^ x86;
  assign n2445 = n2441 & ~n2444;
  assign n2446 = ~n2431 & n2434;
  assign n2447 = ~n2445 & ~n2446;
  assign n2448 = ~n2438 & n2447;
  assign n2449 = ~n2441 & n2444;
  assign n2450 = x215 ^ x87;
  assign n2451 = ~n1545 & n2450;
  assign n2452 = n2451 ^ x87;
  assign n2453 = x471 ^ x343;
  assign n2454 = ~n1028 & n2453;
  assign n2455 = n2454 ^ x343;
  assign n2456 = n2452 & ~n2455;
  assign n2457 = ~n2449 & ~n2456;
  assign n2458 = ~n2448 & n2457;
  assign n2459 = x472 ^ x344;
  assign n2460 = ~n1028 & n2459;
  assign n2461 = n2460 ^ x344;
  assign n2462 = x216 ^ x88;
  assign n2463 = ~n1545 & n2462;
  assign n2464 = n2463 ^ x88;
  assign n2465 = n2461 & ~n2464;
  assign n2466 = ~n2452 & n2455;
  assign n2467 = ~n2465 & ~n2466;
  assign n2468 = ~n2458 & n2467;
  assign n2469 = x473 ^ x345;
  assign n2470 = ~n1028 & n2469;
  assign n2471 = n2470 ^ x345;
  assign n2472 = x217 ^ x89;
  assign n2473 = ~n1545 & n2472;
  assign n2474 = n2473 ^ x89;
  assign n2475 = ~n2471 & n2474;
  assign n2476 = ~n2461 & n2464;
  assign n2477 = ~n2475 & ~n2476;
  assign n2478 = ~n2468 & n2477;
  assign n2479 = x474 ^ x346;
  assign n2480 = ~n1028 & n2479;
  assign n2481 = n2480 ^ x346;
  assign n2482 = x218 ^ x90;
  assign n2483 = ~n1545 & n2482;
  assign n2484 = n2483 ^ x90;
  assign n2485 = n2481 & ~n2484;
  assign n2486 = n2471 & ~n2474;
  assign n2487 = ~n2485 & ~n2486;
  assign n2488 = ~n2478 & n2487;
  assign n2489 = x219 ^ x91;
  assign n2490 = ~n1545 & n2489;
  assign n2491 = n2490 ^ x91;
  assign n2492 = x475 ^ x347;
  assign n2493 = ~n1028 & n2492;
  assign n2494 = n2493 ^ x347;
  assign n2495 = n2491 & ~n2494;
  assign n2496 = ~n2481 & n2484;
  assign n2497 = ~n2495 & ~n2496;
  assign n2498 = ~n2488 & n2497;
  assign n2499 = x476 ^ x348;
  assign n2500 = ~n1028 & n2499;
  assign n2501 = n2500 ^ x348;
  assign n2502 = x220 ^ x92;
  assign n2503 = ~n1545 & n2502;
  assign n2504 = n2503 ^ x92;
  assign n2505 = n2501 & ~n2504;
  assign n2506 = ~n2491 & n2494;
  assign n2507 = ~n2505 & ~n2506;
  assign n2508 = ~n2498 & n2507;
  assign n2509 = x477 ^ x349;
  assign n2510 = ~n1028 & n2509;
  assign n2511 = n2510 ^ x349;
  assign n2512 = x221 ^ x93;
  assign n2513 = ~n1545 & n2512;
  assign n2514 = n2513 ^ x93;
  assign n2515 = ~n2511 & n2514;
  assign n2516 = ~n2501 & n2504;
  assign n2517 = ~n2515 & ~n2516;
  assign n2518 = ~n2508 & n2517;
  assign n2519 = n2511 & ~n2514;
  assign n2520 = ~n2518 & ~n2519;
  assign n2521 = x478 ^ x350;
  assign n2522 = ~n1028 & n2521;
  assign n2523 = n2522 ^ x350;
  assign n2524 = x222 ^ x94;
  assign n2525 = ~n1545 & n2524;
  assign n2526 = n2525 ^ x94;
  assign n2527 = ~n2523 & n2526;
  assign n2528 = ~n2520 & ~n2527;
  assign n2529 = x479 ^ x351;
  assign n2530 = ~n1028 & n2529;
  assign n2531 = n2530 ^ x351;
  assign n2532 = x223 ^ x95;
  assign n2533 = ~n1545 & n2532;
  assign n2534 = n2533 ^ x95;
  assign n2535 = n2531 & ~n2534;
  assign n2536 = n2523 & ~n2526;
  assign n2537 = ~n2535 & ~n2536;
  assign n2538 = ~n2528 & n2537;
  assign n2539 = x224 ^ x96;
  assign n2540 = ~n1545 & n2539;
  assign n2541 = n2540 ^ x96;
  assign n2542 = x480 ^ x352;
  assign n2543 = ~n1028 & n2542;
  assign n2544 = n2543 ^ x352;
  assign n2545 = n2541 & ~n2544;
  assign n2546 = ~n2531 & n2534;
  assign n2547 = ~n2545 & ~n2546;
  assign n2548 = ~n2538 & n2547;
  assign n2549 = ~n1580 & n1583;
  assign n2550 = ~n2541 & n2544;
  assign n2551 = ~n2549 & ~n2550;
  assign n2552 = ~n2548 & n2551;
  assign n2553 = ~n1584 & ~n2552;
  assign n2554 = x482 ^ x354;
  assign n2555 = ~n1028 & n2554;
  assign n2556 = n2555 ^ x354;
  assign n2557 = x226 ^ x98;
  assign n2558 = ~n1545 & n2557;
  assign n2559 = n2558 ^ x98;
  assign n2560 = n2556 & ~n2559;
  assign n2561 = ~n2553 & ~n2560;
  assign n2562 = x483 ^ x355;
  assign n2563 = ~n1028 & n2562;
  assign n2564 = n2563 ^ x355;
  assign n2565 = x227 ^ x99;
  assign n2566 = ~n1545 & n2565;
  assign n2567 = n2566 ^ x99;
  assign n2568 = ~n2564 & n2567;
  assign n2569 = ~n2556 & n2559;
  assign n2570 = ~n2568 & ~n2569;
  assign n2571 = ~n2561 & n2570;
  assign n2572 = x228 ^ x100;
  assign n2573 = ~n1545 & n2572;
  assign n2574 = n2573 ^ x100;
  assign n2575 = x484 ^ x356;
  assign n2576 = ~n1028 & n2575;
  assign n2577 = n2576 ^ x356;
  assign n2578 = ~n2574 & n2577;
  assign n2579 = n2564 & ~n2567;
  assign n2580 = ~n2578 & ~n2579;
  assign n2581 = ~n2571 & n2580;
  assign n2582 = n1573 & ~n1576;
  assign n2583 = n2574 & ~n2577;
  assign n2584 = ~n2582 & ~n2583;
  assign n2585 = ~n2581 & n2584;
  assign n2586 = ~n1577 & ~n2585;
  assign n2587 = x486 ^ x358;
  assign n2588 = ~n1028 & n2587;
  assign n2589 = n2588 ^ x358;
  assign n2590 = x230 ^ x102;
  assign n2591 = ~n1545 & n2590;
  assign n2592 = n2591 ^ x102;
  assign n2593 = ~n2589 & n2592;
  assign n2594 = ~n2586 & ~n2593;
  assign n2595 = x487 ^ x359;
  assign n2596 = ~n1028 & n2595;
  assign n2597 = n2596 ^ x359;
  assign n2598 = x231 ^ x103;
  assign n2599 = ~n1545 & n2598;
  assign n2600 = n2599 ^ x103;
  assign n2601 = n2597 & ~n2600;
  assign n2602 = n2589 & ~n2592;
  assign n2603 = ~n2601 & ~n2602;
  assign n2604 = ~n2594 & n2603;
  assign n2605 = x232 ^ x104;
  assign n2606 = ~n1545 & n2605;
  assign n2607 = n2606 ^ x104;
  assign n2608 = x488 ^ x360;
  assign n2609 = ~n1028 & n2608;
  assign n2610 = n2609 ^ x360;
  assign n2611 = n2607 & ~n2610;
  assign n2612 = ~n2597 & n2600;
  assign n2613 = ~n2611 & ~n2612;
  assign n2614 = ~n2604 & n2613;
  assign n2615 = ~n2607 & n2610;
  assign n2616 = ~n2614 & ~n2615;
  assign n2617 = x489 ^ x361;
  assign n2618 = ~n1028 & n2617;
  assign n2619 = n2618 ^ x361;
  assign n2620 = x233 ^ x105;
  assign n2621 = ~n1545 & n2620;
  assign n2622 = n2621 ^ x105;
  assign n2623 = ~n2619 & n2622;
  assign n2624 = ~n2616 & ~n2623;
  assign n2625 = x490 ^ x362;
  assign n2626 = ~n1028 & n2625;
  assign n2627 = n2626 ^ x362;
  assign n2628 = x234 ^ x106;
  assign n2629 = ~n1545 & n2628;
  assign n2630 = n2629 ^ x106;
  assign n2631 = n2627 & ~n2630;
  assign n2632 = n2619 & ~n2622;
  assign n2633 = ~n2631 & ~n2632;
  assign n2634 = ~n2624 & n2633;
  assign n2635 = x491 ^ x363;
  assign n2636 = ~n1028 & n2635;
  assign n2637 = n2636 ^ x363;
  assign n2638 = x235 ^ x107;
  assign n2639 = ~n1545 & n2638;
  assign n2640 = n2639 ^ x107;
  assign n2641 = ~n2637 & n2640;
  assign n2642 = ~n2627 & n2630;
  assign n2643 = ~n2641 & ~n2642;
  assign n2644 = ~n2634 & n2643;
  assign n2645 = n2637 & ~n2640;
  assign n2646 = ~n2644 & ~n2645;
  assign n2647 = ~n1570 & ~n2646;
  assign n2648 = x237 ^ x109;
  assign n2649 = ~n1545 & n2648;
  assign n2650 = n2649 ^ x109;
  assign n2651 = x493 ^ x365;
  assign n2652 = ~n1028 & n2651;
  assign n2653 = n2652 ^ x365;
  assign n2654 = ~n2650 & n2653;
  assign n2655 = ~n1566 & n1569;
  assign n2656 = ~n2654 & ~n2655;
  assign n2657 = ~n2647 & n2656;
  assign n2658 = n1559 & ~n1562;
  assign n2659 = n2650 & ~n2653;
  assign n2660 = ~n2658 & ~n2659;
  assign n2661 = ~n2657 & n2660;
  assign n2662 = ~n1563 & ~n2661;
  assign n2663 = x495 ^ x367;
  assign n2664 = ~n1028 & n2663;
  assign n2665 = n2664 ^ x367;
  assign n2666 = x239 ^ x111;
  assign n2667 = ~n1545 & n2666;
  assign n2668 = n2667 ^ x111;
  assign n2669 = ~n2665 & n2668;
  assign n2670 = ~n2662 & ~n2669;
  assign n2671 = x496 ^ x368;
  assign n2672 = ~n1028 & n2671;
  assign n2673 = n2672 ^ x368;
  assign n2674 = x240 ^ x112;
  assign n2675 = ~n1545 & n2674;
  assign n2676 = n2675 ^ x112;
  assign n2677 = n2673 & ~n2676;
  assign n2678 = n2665 & ~n2668;
  assign n2679 = ~n2677 & ~n2678;
  assign n2680 = ~n2670 & n2679;
  assign n2681 = x241 ^ x113;
  assign n2682 = ~n1545 & n2681;
  assign n2683 = n2682 ^ x113;
  assign n2684 = x497 ^ x369;
  assign n2685 = ~n1028 & n2684;
  assign n2686 = n2685 ^ x369;
  assign n2687 = n2683 & ~n2686;
  assign n2688 = ~n2673 & n2676;
  assign n2689 = ~n2687 & ~n2688;
  assign n2690 = ~n2680 & n2689;
  assign n2691 = x498 ^ x370;
  assign n2692 = ~n1028 & n2691;
  assign n2693 = n2692 ^ x370;
  assign n2694 = x242 ^ x114;
  assign n2695 = ~n1545 & n2694;
  assign n2696 = n2695 ^ x114;
  assign n2697 = n2693 & ~n2696;
  assign n2698 = ~n2683 & n2686;
  assign n2699 = ~n2697 & ~n2698;
  assign n2700 = ~n2690 & n2699;
  assign n2701 = x499 ^ x371;
  assign n2702 = ~n1028 & n2701;
  assign n2703 = n2702 ^ x371;
  assign n2704 = x243 ^ x115;
  assign n2705 = ~n1545 & n2704;
  assign n2706 = n2705 ^ x115;
  assign n2707 = ~n2703 & n2706;
  assign n2708 = ~n2693 & n2696;
  assign n2709 = ~n2707 & ~n2708;
  assign n2710 = ~n2700 & n2709;
  assign n2711 = x244 ^ x116;
  assign n2712 = ~n1545 & n2711;
  assign n2713 = n2712 ^ x116;
  assign n2714 = x500 ^ x372;
  assign n2715 = ~n1028 & n2714;
  assign n2716 = n2715 ^ x372;
  assign n2717 = ~n2713 & n2716;
  assign n2718 = n2703 & ~n2706;
  assign n2719 = ~n2717 & ~n2718;
  assign n2720 = ~n2710 & n2719;
  assign n2721 = x245 ^ x117;
  assign n2722 = ~n1545 & n2721;
  assign n2723 = n2722 ^ x117;
  assign n2724 = x501 ^ x373;
  assign n2725 = ~n1028 & n2724;
  assign n2726 = n2725 ^ x373;
  assign n2727 = n2723 & ~n2726;
  assign n2728 = n2713 & ~n2716;
  assign n2729 = ~n2727 & ~n2728;
  assign n2730 = ~n2720 & n2729;
  assign n2731 = x502 ^ x374;
  assign n2732 = ~n1028 & n2731;
  assign n2733 = n2732 ^ x374;
  assign n2734 = x246 ^ x118;
  assign n2735 = ~n1545 & n2734;
  assign n2736 = n2735 ^ x118;
  assign n2737 = n2733 & ~n2736;
  assign n2738 = ~n2723 & n2726;
  assign n2739 = ~n2737 & ~n2738;
  assign n2740 = ~n2730 & n2739;
  assign n2741 = x503 ^ x375;
  assign n2742 = ~n1028 & n2741;
  assign n2743 = n2742 ^ x375;
  assign n2744 = x247 ^ x119;
  assign n2745 = ~n1545 & n2744;
  assign n2746 = n2745 ^ x119;
  assign n2747 = ~n2743 & n2746;
  assign n2748 = ~n2733 & n2736;
  assign n2749 = ~n2747 & ~n2748;
  assign n2750 = ~n2740 & n2749;
  assign n2751 = n2743 & ~n2746;
  assign n2752 = ~n2750 & ~n2751;
  assign n2753 = ~n1556 & ~n2752;
  assign n2754 = x249 ^ x121;
  assign n2755 = ~n1545 & n2754;
  assign n2756 = n2755 ^ x121;
  assign n2757 = x505 ^ x377;
  assign n2758 = ~n1028 & n2757;
  assign n2759 = n2758 ^ x377;
  assign n2760 = ~n2756 & n2759;
  assign n2761 = ~n1552 & n1555;
  assign n2762 = ~n2760 & ~n2761;
  assign n2763 = ~n2753 & n2762;
  assign n2764 = n2756 & ~n2759;
  assign n2765 = ~n1031 & n1548;
  assign n2766 = ~n2764 & ~n2765;
  assign n2767 = ~n2763 & n2766;
  assign n2768 = ~n1549 & ~n2767;
  assign n2769 = x507 ^ x379;
  assign n2770 = ~n1028 & n2769;
  assign n2771 = n2770 ^ x379;
  assign n2772 = x251 ^ x123;
  assign n2773 = ~n1545 & n2772;
  assign n2774 = n2773 ^ x123;
  assign n2775 = ~n2771 & n2774;
  assign n2776 = ~n2768 & ~n2775;
  assign n2777 = x508 ^ x380;
  assign n2778 = ~n1028 & n2777;
  assign n2779 = n2778 ^ x380;
  assign n2780 = x252 ^ x124;
  assign n2781 = ~n1545 & n2780;
  assign n2782 = n2781 ^ x124;
  assign n2783 = n2779 & ~n2782;
  assign n2784 = n2771 & ~n2774;
  assign n2785 = ~n2783 & ~n2784;
  assign n2786 = ~n2776 & n2785;
  assign n2787 = x253 ^ x125;
  assign n2788 = ~n1545 & n2787;
  assign n2789 = n2788 ^ x125;
  assign n2790 = x509 ^ x381;
  assign n2791 = ~n1028 & n2790;
  assign n2792 = n2791 ^ x381;
  assign n2793 = n2789 & ~n2792;
  assign n2794 = ~n2779 & n2782;
  assign n2795 = ~n2793 & ~n2794;
  assign n2796 = ~n2786 & n2795;
  assign n2797 = x510 ^ x382;
  assign n2798 = ~n1028 & n2797;
  assign n2799 = n2798 ^ x382;
  assign n2800 = x254 ^ x126;
  assign n2801 = ~n1545 & n2800;
  assign n2802 = n2801 ^ x126;
  assign n2803 = n2799 & ~n2802;
  assign n2804 = ~n2789 & n2792;
  assign n2805 = ~n2803 & ~n2804;
  assign n2806 = ~n2796 & n2805;
  assign n2807 = x127 & x255;
  assign n2808 = x383 & x511;
  assign n2809 = ~n2807 & n2808;
  assign n2810 = ~n2799 & n2802;
  assign n2811 = ~n2809 & ~n2810;
  assign n2812 = ~n2806 & n2811;
  assign n2813 = n2807 & ~n2808;
  assign n2814 = ~n2812 & ~n2813;
  assign n2815 = n1730 ^ n1727;
  assign n2816 = n2814 & n2815;
  assign n2817 = n2816 ^ n1727;
  assign n2818 = n1723 ^ n1720;
  assign n2819 = n2814 & n2818;
  assign n2820 = n2819 ^ n1720;
  assign n2821 = n1738 ^ n1735;
  assign n2822 = n2814 & n2821;
  assign n2823 = n2822 ^ n1735;
  assign n2824 = n1749 ^ n1746;
  assign n2825 = n2814 & n2824;
  assign n2826 = n2825 ^ n1746;
  assign n2827 = n1759 ^ n1756;
  assign n2828 = ~n2814 & n2827;
  assign n2829 = n2828 ^ n1756;
  assign n2830 = n1716 ^ n1713;
  assign n2831 = ~n2814 & n2830;
  assign n2832 = n2831 ^ n1713;
  assign n2833 = n1772 ^ n1769;
  assign n2834 = n2814 & n2833;
  assign n2835 = n2834 ^ n1769;
  assign n2836 = n1782 ^ n1779;
  assign n2837 = ~n2814 & n2836;
  assign n2838 = n2837 ^ n1779;
  assign n2839 = n1709 ^ n1706;
  assign n2840 = n2814 & n2839;
  assign n2841 = n2840 ^ n1706;
  assign n2842 = n1795 ^ n1792;
  assign n2843 = n2814 & n2842;
  assign n2844 = n2843 ^ n1792;
  assign n2845 = n1805 ^ n1802;
  assign n2846 = ~n2814 & n2845;
  assign n2847 = n2846 ^ n1802;
  assign n2848 = n1815 ^ n1812;
  assign n2849 = ~n2814 & n2848;
  assign n2850 = n2849 ^ n1812;
  assign n2851 = n1825 ^ n1822;
  assign n2852 = ~n2814 & n2851;
  assign n2853 = n2852 ^ n1822;
  assign n2854 = n1835 ^ n1832;
  assign n2855 = n2814 & n2854;
  assign n2856 = n2855 ^ n1832;
  assign n2857 = n1845 ^ n1842;
  assign n2858 = n2814 & n2857;
  assign n2859 = n2858 ^ n1842;
  assign n2860 = n1854 ^ n1851;
  assign n2861 = ~n2814 & n2860;
  assign n2862 = n2861 ^ n1851;
  assign n2863 = n1702 ^ n1699;
  assign n2864 = n2814 & n2863;
  assign n2865 = n2864 ^ n1699;
  assign n2866 = n1868 ^ n1865;
  assign n2867 = ~n2814 & n2866;
  assign n2868 = n2867 ^ n1865;
  assign n2869 = n1695 ^ n1692;
  assign n2870 = ~n2814 & n2869;
  assign n2871 = n2870 ^ n1692;
  assign n2872 = n1881 ^ n1878;
  assign n2873 = n2814 & n2872;
  assign n2874 = n2873 ^ n1878;
  assign n2875 = n1891 ^ n1888;
  assign n2876 = ~n2814 & n2875;
  assign n2877 = n2876 ^ n1888;
  assign n2878 = n1688 ^ n1685;
  assign n2879 = n2814 & n2878;
  assign n2880 = n2879 ^ n1685;
  assign n2881 = n1904 ^ n1901;
  assign n2882 = n2814 & n2881;
  assign n2883 = n2882 ^ n1901;
  assign n2884 = n1914 ^ n1911;
  assign n2885 = n2814 & n2884;
  assign n2886 = n2885 ^ n1911;
  assign n2887 = n1924 ^ n1921;
  assign n2888 = ~n2814 & n2887;
  assign n2889 = n2888 ^ n1921;
  assign n2890 = n1681 ^ n1678;
  assign n2891 = ~n2814 & n2890;
  assign n2892 = n2891 ^ n1678;
  assign n2893 = n1936 ^ n1933;
  assign n2894 = ~n2814 & n2893;
  assign n2895 = n2894 ^ n1933;
  assign n2896 = n1674 ^ n1671;
  assign n2897 = n2814 & n2896;
  assign n2898 = n2897 ^ n1671;
  assign n2899 = n1950 ^ n1947;
  assign n2900 = ~n2814 & n2899;
  assign n2901 = n2900 ^ n1947;
  assign n2902 = n1960 ^ n1957;
  assign n2903 = ~n2814 & n2902;
  assign n2904 = n2903 ^ n1957;
  assign n2905 = n1667 ^ n1664;
  assign n2906 = n2814 & n2905;
  assign n2907 = n2906 ^ n1664;
  assign n2908 = n1973 ^ n1970;
  assign n2909 = ~n2814 & n2908;
  assign n2910 = n2909 ^ n1970;
  assign n2911 = n1660 ^ n1657;
  assign n2912 = ~n2814 & n2911;
  assign n2913 = n2912 ^ n1657;
  assign n2914 = n1985 ^ n1982;
  assign n2915 = ~n2814 & n2914;
  assign n2916 = n2915 ^ n1982;
  assign n2917 = n1653 ^ n1650;
  assign n2918 = n2814 & n2917;
  assign n2919 = n2918 ^ n1650;
  assign n2920 = n1999 ^ n1996;
  assign n2921 = ~n2814 & n2920;
  assign n2922 = n2921 ^ n1996;
  assign n2923 = n2009 ^ n2006;
  assign n2924 = ~n2814 & n2923;
  assign n2925 = n2924 ^ n2006;
  assign n2926 = n1646 ^ n1643;
  assign n2927 = n2814 & n2926;
  assign n2928 = n2927 ^ n1643;
  assign n2929 = n2022 ^ n2019;
  assign n2930 = ~n2814 & n2929;
  assign n2931 = n2930 ^ n2019;
  assign n2932 = n1639 ^ n1636;
  assign n2933 = ~n2814 & n2932;
  assign n2934 = n2933 ^ n1636;
  assign n2935 = n2035 ^ n2032;
  assign n2936 = ~n2814 & n2935;
  assign n2937 = n2936 ^ n2032;
  assign n2938 = n2045 ^ n2042;
  assign n2939 = ~n2814 & n2938;
  assign n2940 = n2939 ^ n2042;
  assign n2941 = n1632 ^ n1629;
  assign n2942 = ~n2814 & n2941;
  assign n2943 = n2942 ^ n1629;
  assign n2944 = n2058 ^ n2055;
  assign n2945 = n2814 & n2944;
  assign n2946 = n2945 ^ n2055;
  assign n2947 = n2068 ^ n2065;
  assign n2948 = n2814 & n2947;
  assign n2949 = n2948 ^ n2065;
  assign n2950 = n2078 ^ n2075;
  assign n2951 = ~n2814 & n2950;
  assign n2952 = n2951 ^ n2075;
  assign n2953 = n1625 ^ n1622;
  assign n2954 = ~n2814 & n2953;
  assign n2955 = n2954 ^ n1622;
  assign n2956 = n2091 ^ n2088;
  assign n2957 = ~n2814 & n2956;
  assign n2958 = n2957 ^ n2088;
  assign n2959 = n1618 ^ n1615;
  assign n2960 = n2814 & n2959;
  assign n2961 = n2960 ^ n1615;
  assign n2962 = n2104 ^ n2101;
  assign n2963 = ~n2814 & n2962;
  assign n2964 = n2963 ^ n2101;
  assign n2965 = n2114 ^ n2111;
  assign n2966 = n2814 & n2965;
  assign n2967 = n2966 ^ n2111;
  assign n2968 = n2124 ^ n2121;
  assign n2969 = n2814 & n2968;
  assign n2970 = n2969 ^ n2121;
  assign n2971 = n2133 ^ n2130;
  assign n2972 = ~n2814 & n2971;
  assign n2973 = n2972 ^ n2130;
  assign n2974 = n1611 ^ n1608;
  assign n2975 = n2814 & n2974;
  assign n2976 = n2975 ^ n1608;
  assign n2977 = n2147 ^ n2144;
  assign n2978 = ~n2814 & n2977;
  assign n2979 = n2978 ^ n2144;
  assign n2980 = n2157 ^ n2154;
  assign n2981 = n2814 & n2980;
  assign n2982 = n2981 ^ n2154;
  assign n2983 = n2166 ^ n2163;
  assign n2984 = ~n2814 & n2983;
  assign n2985 = n2984 ^ n2163;
  assign n2986 = n1604 ^ n1601;
  assign n2987 = n2814 & n2986;
  assign n2988 = n2987 ^ n1601;
  assign n2989 = n2180 ^ n2177;
  assign n2990 = n2814 & n2989;
  assign n2991 = n2990 ^ n2177;
  assign n2992 = n2190 ^ n2187;
  assign n2993 = n2814 & n2992;
  assign n2994 = n2993 ^ n2187;
  assign n2995 = n2200 ^ n2197;
  assign n2996 = ~n2814 & n2995;
  assign n2997 = n2996 ^ n2197;
  assign n2998 = n2210 ^ n2207;
  assign n2999 = n2814 & n2998;
  assign n3000 = n2999 ^ n2207;
  assign n3001 = n2220 ^ n2217;
  assign n3002 = ~n2814 & n3001;
  assign n3003 = n3002 ^ n2217;
  assign n3004 = n2229 ^ n2227;
  assign n3005 = ~n2814 & n3004;
  assign n3006 = n3005 ^ n2227;
  assign n3007 = n2239 ^ n2236;
  assign n3008 = ~n2814 & n3007;
  assign n3009 = n3008 ^ n2236;
  assign n3010 = n2249 ^ n2246;
  assign n3011 = ~n2814 & n3010;
  assign n3012 = n3011 ^ n2246;
  assign n3013 = n2259 ^ n2256;
  assign n3014 = ~n2814 & n3013;
  assign n3015 = n3014 ^ n2256;
  assign n3016 = n2269 ^ n2266;
  assign n3017 = ~n2814 & n3016;
  assign n3018 = n3017 ^ n2266;
  assign n3019 = n1597 ^ n1594;
  assign n3020 = n2814 & n3019;
  assign n3021 = n3020 ^ n1594;
  assign n3022 = n2281 ^ n2278;
  assign n3023 = ~n2814 & n3022;
  assign n3024 = n3023 ^ n2278;
  assign n3025 = n2292 ^ n2289;
  assign n3026 = ~n2814 & n3025;
  assign n3027 = n3026 ^ n2289;
  assign n3028 = n2302 ^ n2299;
  assign n3029 = ~n2814 & n3028;
  assign n3030 = n3029 ^ n2299;
  assign n3031 = n1590 ^ n1587;
  assign n3032 = ~n2814 & n3031;
  assign n3033 = n3032 ^ n1587;
  assign n3034 = n2315 ^ n2312;
  assign n3035 = n2814 & n3034;
  assign n3036 = n3035 ^ n2312;
  assign n3037 = n2325 ^ n2322;
  assign n3038 = ~n2814 & n3037;
  assign n3039 = n3038 ^ n2322;
  assign n3040 = n2334 ^ n2331;
  assign n3041 = n2814 & n3040;
  assign n3042 = n3041 ^ n2331;
  assign n3043 = n2344 ^ n2341;
  assign n3044 = ~n2814 & n3043;
  assign n3045 = n3044 ^ n2341;
  assign n3046 = n2354 ^ n2351;
  assign n3047 = n2814 & n3046;
  assign n3048 = n3047 ^ n2351;
  assign n3049 = n2364 ^ n2361;
  assign n3050 = n2814 & n3049;
  assign n3051 = n3050 ^ n2361;
  assign n3052 = n2376 ^ n2373;
  assign n3053 = ~n2814 & n3052;
  assign n3054 = n3053 ^ n2373;
  assign n3055 = n2384 ^ n2381;
  assign n3056 = ~n2814 & n3055;
  assign n3057 = n3056 ^ n2381;
  assign n3058 = n2395 ^ n2392;
  assign n3059 = ~n2814 & n3058;
  assign n3060 = n3059 ^ n2392;
  assign n3061 = n2406 ^ n2403;
  assign n3062 = n2814 & n3061;
  assign n3063 = n3062 ^ n2403;
  assign n3064 = n2414 ^ n2411;
  assign n3065 = ~n2814 & n3064;
  assign n3066 = n3065 ^ n2411;
  assign n3067 = n2424 ^ n2421;
  assign n3068 = ~n2814 & n3067;
  assign n3069 = n3068 ^ n2421;
  assign n3070 = n2434 ^ n2431;
  assign n3071 = ~n2814 & n3070;
  assign n3072 = n3071 ^ n2431;
  assign n3073 = n2444 ^ n2441;
  assign n3074 = n2814 & n3073;
  assign n3075 = n3074 ^ n2441;
  assign n3076 = n2455 ^ n2452;
  assign n3077 = ~n2814 & n3076;
  assign n3078 = n3077 ^ n2452;
  assign n3079 = n2464 ^ n2461;
  assign n3080 = n2814 & n3079;
  assign n3081 = n3080 ^ n2461;
  assign n3082 = n2474 ^ n2471;
  assign n3083 = n2814 & n3082;
  assign n3084 = n3083 ^ n2471;
  assign n3085 = n2484 ^ n2481;
  assign n3086 = n2814 & n3085;
  assign n3087 = n3086 ^ n2481;
  assign n3088 = n2494 ^ n2491;
  assign n3089 = ~n2814 & n3088;
  assign n3090 = n3089 ^ n2491;
  assign n3091 = n2504 ^ n2501;
  assign n3092 = n2814 & n3091;
  assign n3093 = n3092 ^ n2501;
  assign n3094 = n2514 ^ n2511;
  assign n3095 = n2814 & n3094;
  assign n3096 = n3095 ^ n2511;
  assign n3097 = n2526 ^ n2523;
  assign n3098 = n2814 & n3097;
  assign n3099 = n3098 ^ n2523;
  assign n3100 = n2534 ^ n2531;
  assign n3101 = n2814 & n3100;
  assign n3102 = n3101 ^ n2531;
  assign n3103 = n2544 ^ n2541;
  assign n3104 = ~n2814 & n3103;
  assign n3105 = n3104 ^ n2541;
  assign n3106 = n1583 ^ n1580;
  assign n3107 = ~n2814 & n3106;
  assign n3108 = n3107 ^ n1580;
  assign n3109 = n2559 ^ n2556;
  assign n3110 = n2814 & n3109;
  assign n3111 = n3110 ^ n2556;
  assign n3112 = n2567 ^ n2564;
  assign n3113 = n2814 & n3112;
  assign n3114 = n3113 ^ n2564;
  assign n3115 = n2577 ^ n2574;
  assign n3116 = ~n2814 & n3115;
  assign n3117 = n3116 ^ n2574;
  assign n3118 = n1576 ^ n1573;
  assign n3119 = ~n2814 & n3118;
  assign n3120 = n3119 ^ n1573;
  assign n3121 = n2592 ^ n2589;
  assign n3122 = n2814 & n3121;
  assign n3123 = n3122 ^ n2589;
  assign n3124 = n2600 ^ n2597;
  assign n3125 = n2814 & n3124;
  assign n3126 = n3125 ^ n2597;
  assign n3127 = n2610 ^ n2607;
  assign n3128 = ~n2814 & n3127;
  assign n3129 = n3128 ^ n2607;
  assign n3130 = n2622 ^ n2619;
  assign n3131 = n2814 & n3130;
  assign n3132 = n3131 ^ n2619;
  assign n3133 = n2630 ^ n2627;
  assign n3134 = n2814 & n3133;
  assign n3135 = n3134 ^ n2627;
  assign n3136 = n2640 ^ n2637;
  assign n3137 = n2814 & n3136;
  assign n3138 = n3137 ^ n2637;
  assign n3139 = n1569 ^ n1566;
  assign n3140 = ~n2814 & n3139;
  assign n3141 = n3140 ^ n1566;
  assign n3142 = n2653 ^ n2650;
  assign n3143 = ~n2814 & n3142;
  assign n3144 = n3143 ^ n2650;
  assign n3145 = n1562 ^ n1559;
  assign n3146 = ~n2814 & n3145;
  assign n3147 = n3146 ^ n1559;
  assign n3148 = n2668 ^ n2665;
  assign n3149 = n2814 & n3148;
  assign n3150 = n3149 ^ n2665;
  assign n3151 = n2676 ^ n2673;
  assign n3152 = n2814 & n3151;
  assign n3153 = n3152 ^ n2673;
  assign n3154 = n2686 ^ n2683;
  assign n3155 = ~n2814 & n3154;
  assign n3156 = n3155 ^ n2683;
  assign n3157 = n2696 ^ n2693;
  assign n3158 = n2814 & n3157;
  assign n3159 = n3158 ^ n2693;
  assign n3160 = n2706 ^ n2703;
  assign n3161 = n2814 & n3160;
  assign n3162 = n3161 ^ n2703;
  assign n3163 = n2716 ^ n2713;
  assign n3164 = ~n2814 & n3163;
  assign n3165 = n3164 ^ n2713;
  assign n3166 = n2726 ^ n2723;
  assign n3167 = ~n2814 & n3166;
  assign n3168 = n3167 ^ n2723;
  assign n3169 = n2736 ^ n2733;
  assign n3170 = n2814 & n3169;
  assign n3171 = n3170 ^ n2733;
  assign n3172 = n2746 ^ n2743;
  assign n3173 = n2814 & n3172;
  assign n3174 = n3173 ^ n2743;
  assign n3175 = n1555 ^ n1552;
  assign n3176 = ~n2814 & n3175;
  assign n3177 = n3176 ^ n1552;
  assign n3178 = n2759 ^ n2756;
  assign n3179 = ~n2814 & n3178;
  assign n3180 = n3179 ^ n2756;
  assign n3181 = n1548 ^ n1031;
  assign n3182 = n2814 & n3181;
  assign n3183 = n3182 ^ n1031;
  assign n3184 = n2774 ^ n2771;
  assign n3185 = n2814 & n3184;
  assign n3186 = n3185 ^ n2771;
  assign n3187 = n2782 ^ n2779;
  assign n3188 = n2814 & n3187;
  assign n3189 = n3188 ^ n2779;
  assign n3190 = n2792 ^ n2789;
  assign n3191 = ~n2814 & n3190;
  assign n3192 = n3191 ^ n2789;
  assign n3193 = n2802 ^ n2799;
  assign n3194 = n2814 & n3193;
  assign n3195 = n3194 ^ n2799;
  assign n3196 = n2807 & n2808;
  assign n3197 = n1545 ^ n1028;
  assign n3198 = n2814 & n3197;
  assign n3199 = n3198 ^ n1028;
  assign y0 = n2817;
  assign y1 = n2820;
  assign y2 = n2823;
  assign y3 = n2826;
  assign y4 = n2829;
  assign y5 = n2832;
  assign y6 = n2835;
  assign y7 = n2838;
  assign y8 = n2841;
  assign y9 = n2844;
  assign y10 = n2847;
  assign y11 = n2850;
  assign y12 = n2853;
  assign y13 = n2856;
  assign y14 = n2859;
  assign y15 = n2862;
  assign y16 = n2865;
  assign y17 = n2868;
  assign y18 = n2871;
  assign y19 = n2874;
  assign y20 = n2877;
  assign y21 = n2880;
  assign y22 = n2883;
  assign y23 = n2886;
  assign y24 = n2889;
  assign y25 = n2892;
  assign y26 = n2895;
  assign y27 = n2898;
  assign y28 = n2901;
  assign y29 = n2904;
  assign y30 = n2907;
  assign y31 = n2910;
  assign y32 = n2913;
  assign y33 = n2916;
  assign y34 = n2919;
  assign y35 = n2922;
  assign y36 = n2925;
  assign y37 = n2928;
  assign y38 = n2931;
  assign y39 = n2934;
  assign y40 = n2937;
  assign y41 = n2940;
  assign y42 = n2943;
  assign y43 = n2946;
  assign y44 = n2949;
  assign y45 = n2952;
  assign y46 = n2955;
  assign y47 = n2958;
  assign y48 = n2961;
  assign y49 = n2964;
  assign y50 = n2967;
  assign y51 = n2970;
  assign y52 = n2973;
  assign y53 = n2976;
  assign y54 = n2979;
  assign y55 = n2982;
  assign y56 = n2985;
  assign y57 = n2988;
  assign y58 = n2991;
  assign y59 = n2994;
  assign y60 = n2997;
  assign y61 = n3000;
  assign y62 = n3003;
  assign y63 = n3006;
  assign y64 = n3009;
  assign y65 = n3012;
  assign y66 = n3015;
  assign y67 = n3018;
  assign y68 = n3021;
  assign y69 = n3024;
  assign y70 = n3027;
  assign y71 = n3030;
  assign y72 = n3033;
  assign y73 = n3036;
  assign y74 = n3039;
  assign y75 = n3042;
  assign y76 = n3045;
  assign y77 = n3048;
  assign y78 = n3051;
  assign y79 = n3054;
  assign y80 = n3057;
  assign y81 = n3060;
  assign y82 = n3063;
  assign y83 = n3066;
  assign y84 = n3069;
  assign y85 = n3072;
  assign y86 = n3075;
  assign y87 = n3078;
  assign y88 = n3081;
  assign y89 = n3084;
  assign y90 = n3087;
  assign y91 = n3090;
  assign y92 = n3093;
  assign y93 = n3096;
  assign y94 = n3099;
  assign y95 = n3102;
  assign y96 = n3105;
  assign y97 = n3108;
  assign y98 = n3111;
  assign y99 = n3114;
  assign y100 = n3117;
  assign y101 = n3120;
  assign y102 = n3123;
  assign y103 = n3126;
  assign y104 = n3129;
  assign y105 = n3132;
  assign y106 = n3135;
  assign y107 = n3138;
  assign y108 = n3141;
  assign y109 = n3144;
  assign y110 = n3147;
  assign y111 = n3150;
  assign y112 = n3153;
  assign y113 = n3156;
  assign y114 = n3159;
  assign y115 = n3162;
  assign y116 = n3165;
  assign y117 = n3168;
  assign y118 = n3171;
  assign y119 = n3174;
  assign y120 = n3177;
  assign y121 = n3180;
  assign y122 = n3183;
  assign y123 = n3186;
  assign y124 = n3189;
  assign y125 = n3192;
  assign y126 = n3195;
  assign y127 = n3196;
  assign y128 = ~n3199;
  assign y129 = ~n2814;
endmodule
