module top(n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437);
  input n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63;
  output n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437;
  wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373;
  assign n12261 = n51 ^ n50;
  assign n12205 = n41 ^ n40;
  assign n12225 = n49 ^ n48;
  assign n12307 = n60 ^ n59;
  assign n12280 = n62 ^ n61;
  assign n12276 = n35 ^ n34;
  assign n12287 = n56 ^ n55;
  assign n12309 = n50 ^ n49;
  assign n12305 = n58 ^ n57;
  assign n12292 = n40 ^ n39;
  assign n12202 = n39 ^ n38;
  assign n12176 = n57 ^ n56;
  assign n12291 = n36 ^ n35;
  assign n12302 = n38 ^ n37;
  assign n12223 = n37 ^ n36;
  assign n12286 = n52 ^ n51;
  assign n12258 = n45 ^ n44;
  assign n12299 = n34 ^ n33;
  assign n12301 = n46 ^ n45;
  assign n12214 = n43 ^ n42;
  assign n12279 = n44 ^ n43;
  assign n12238 = n47 ^ n46;
  assign n12229 = n59 ^ n58;
  assign n12297 = n48 ^ n47;
  assign n12200 = n55 ^ n54;
  assign n12283 = n54 ^ n53;
  assign n12192 = n62 ^ n63;
  assign n12312 = n42 ^ n41;
  assign n12271 = n53 ^ n52;
  assign n12254 = n61 ^ n60;
  assign n5209 = n63 & n5;
  assign n12349 = n0 & n58;
  assign n6057 = n63 & n21;
  assign n6158 = n63 & n25;
  assign n12367 = n0 & n34;
  assign n12372 = n0 & n40;
  assign n12364 = n0 & n60;
  assign n6423 = n63 & n26;
  assign n6227 = n63 & n15;
  assign n6425 = n63 & n18;
  assign n12369 = n0 & n42;
  assign n6273 = n63 & n14;
  assign n6404 = n63 & n3;
  assign n6221 = n63 & n8;
  assign n12368 = n0 & n52;
  assign n12350 = n0 & n56;
  assign n5138 = n63 & n29;
  assign n10228 = n63 & n0;
  assign n12373 = n0 & n36;
  assign n6144 = n63 & n22;
  assign n5082 = n63 & n16;
  assign n12361 = n0 & n54;
  assign n5052 = n63 & n10;
  assign n5299 = n63 & n2;
  assign n12356 = n0 & n38;
  assign n5068 = n63 & n9;
  assign n6118 = n63 & n17;
  assign n6050 = n30 & n63;
  assign n5163 = n63 & n27;
  assign n5249 = n63 & n23;
  assign n6304 = n63 & n24;
  assign n5277 = n63 & n12;
  assign n12347 = n0 & n44;
  assign n5173 = n63 & n6;
  assign n12374 = n32 & n0;
  assign n6247 = n63 & n7;
  assign n6149 = n63 & n11;
  assign n6204 = n63 & n28;
  assign n5175 = n63 & n20;
  assign n12365 = n0 & n62;
  assign n12362 = n0 & n48;
  assign n5028 = n63 & n1;
  assign n12363 = n0 & n46;
  assign n6358 = n63 & n13;
  assign n12348 = n0 & n50;
  assign n12327 = n32 & n33;
  assign n6384 = n63 & n4;
  assign n6315 = n63 & n19;
  assign n10997 = ~n26;
  assign n10965 = ~n18;
  assign n10949 = ~n13;
  assign n11344 = ~n55;
  assign n12355 = ~n54;
  assign n11000 = ~n25;
  assign n12370 = ~n38;
  assign n9939 = ~n31;
  assign n10996 = ~n23;
  assign n11332 = ~n59;
  assign n7004 = ~n33;
  assign n12359 = ~n52;
  assign n11004 = ~n7;
  assign n11129 = ~n41;
  assign n11593 = ~n57;
  assign n12343 = ~n56;
  assign n12354 = ~n62;
  assign n11337 = ~n51;
  assign n10992 = ~n28;
  assign n10962 = ~n20;
  assign n11340 = ~n47;
  assign n10957 = ~n9;
  assign n11342 = ~n35;
  assign n10990 = ~n2;
  assign n10954 = ~n4;
  assign n10971 = ~n12;
  assign n12371 = ~n44;
  assign n10988 = ~n19;
  assign n11739 = ~n53;
  assign n11898 = ~n61;
  assign n11007 = ~n0;
  assign n10973 = ~n1;
  assign n10994 = ~n16;
  assign n10952 = ~n6;
  assign n12345 = ~n32;
  assign n10999 = ~n3;
  assign n12353 = ~n48;
  assign n10979 = ~n5;
  assign n12366 = ~n46;
  assign n11005 = ~n17;
  assign n11137 = ~n39;
  assign n10981 = ~n11;
  assign n10961 = ~n29;
  assign n12346 = ~n34;
  assign n12352 = ~n60;
  assign n10977 = ~n30;
  assign n10959 = ~n22;
  assign n11166 = ~n43;
  assign n10974 = ~n10;
  assign n11003 = ~n15;
  assign n11320 = ~n63;
  assign n12344 = ~n58;
  assign n11327 = ~n49;
  assign n10989 = ~n21;
  assign n12357 = ~n40;
  assign n12358 = ~n42;
  assign n10972 = ~n14;
  assign n12351 = ~n36;
  assign n10966 = ~n27;
  assign n11104 = ~n45;
  assign n10963 = ~n24;
  assign n11329 = ~n37;
  assign n10969 = ~n8;
  assign n12360 = ~n50;
  assign n6082 = n12279 & n0;
  assign n12152 = n11320 & n12280;
  assign n6340 = n12283 & n0;
  assign n12149 = n12286 & n53;
  assign n12133 = n11593 & n12287;
  assign n6360 = n12291 & n0;
  assign n12131 = n11129 & n12292;
  assign n12128 = n12297 & n49;
  assign n12157 = n12287 & n57;
  assign n6282 = n12287 & n0;
  assign n12155 = n12279 & n45;
  assign n12138 = n12299 & n35;
  assign n12150 = n11340 & n12301;
  assign n9706 = n12299 & n0;
  assign n12147 = n11137 & n12302;
  assign n12139 = n11344 & n12283;
  assign n12129 = n12305 & n59;
  assign n12143 = n12307 & n61;
  assign n12151 = n12309 & n51;
  assign n12130 = n11104 & n12279;
  assign n9670 = n12301 & n0;
  assign n12134 = n11166 & n12312;
  assign n9676 = n12297 & n0;
  assign n9674 = n12309 & n0;
  assign n12148 = n12283 & n55;
  assign n9672 = n12286 & n0;
  assign n12136 = n12292 & n41;
  assign n12127 = n12312 & n43;
  assign n6260 = n12305 & n0;
  assign n12156 = n11329 & n12291;
  assign n12154 = n12280 & n63;
  assign n6092 = n12312 & n0;
  assign n9188 = n12292 & n0;
  assign n12140 = n11739 & n12286;
  assign n12158 = n11898 & n12307;
  assign n12145 = n12302 & n39;
  assign n12142 = n11337 & n12309;
  assign n9684 = n12302 & n0;
  assign n12137 = n12301 & n47;
  assign n12144 = n12291 & n37;
  assign n6192 = n12307 & n0;
  assign n12126 = n11327 & n12297;
  assign n12153 = n11332 & n12305;
  assign n9704 = n12280 & n0;
  assign n12146 = n11342 & n12299;
  assign n12316 = n10971 & n12327;
  assign n12199 = ~n12283;
  assign n12320 = n10973 & n12327;
  assign n12323 = n10999 & n12327;
  assign n12253 = ~n12307;
  assign n12293 = n10997 & n12327;
  assign n12300 = n10992 & n12327;
  assign n12311 = n10966 & n12327;
  assign n12322 = n9939 & n12327;
  assign n12318 = n10954 & n12327;
  assign n12237 = ~n12301;
  assign n12285 = n10965 & n12327;
  assign n12213 = ~n12312;
  assign n12288 = n10961 & n12327;
  assign n12275 = ~n12299;
  assign n12298 = n10994 & n12327;
  assign n12306 = n11000 & n12327;
  assign n12317 = n10979 & n12327;
  assign n12321 = n10972 & n12327;
  assign n12313 = n11004 & n12327;
  assign n12257 = ~n12279;
  assign n12175 = ~n12287;
  assign n12324 = n10949 & n12327;
  assign n12303 = n11005 & n12327;
  assign n12304 = n10959 & n12327;
  assign n12260 = ~n12309;
  assign n12296 = n10969 & n12327;
  assign n12228 = ~n12305;
  assign n12201 = ~n12302;
  assign n12315 = n10977 & n12327;
  assign n12289 = n11003 & n12327;
  assign n12326 = n10952 & n12327;
  assign n11081 = ~n12280;
  assign n12281 = n10963 & n12327;
  assign n12290 = n10981 & n12327;
  assign n12270 = ~n12286;
  assign n12222 = ~n12291;
  assign n12282 = n10962 & n12327;
  assign n12319 = n10988 & n12327;
  assign n12204 = ~n12292;
  assign n12314 = n10996 & n12327;
  assign n12310 = n10974 & n12327;
  assign n12308 = n10989 & n12327;
  assign n12325 = n10990 & n12327;
  assign n12294 = n10957 & n12327;
  assign n12224 = ~n12297;
  assign n12338 = n11007 & n12343;
  assign n6992 = ~n6404;
  assign n12328 = n11007 & n12344;
  assign n6704 = ~n6204;
  assign n12278 = n12345 & n33;
  assign n6708 = ~n6384;
  assign n6976 = ~n5173;
  assign n6961 = ~n6057;
  assign n12337 = n11007 & n12346;
  assign n11097 = ~n12347;
  assign n11095 = ~n12348;
  assign n11085 = ~n12349;
  assign n11077 = ~n12350;
  assign n12330 = n11007 & n12351;
  assign n7974 = ~n5163;
  assign n6967 = ~n5175;
  assign n12329 = n11007 & n12352;
  assign n6990 = ~n5082;
  assign n12341 = n11007 & n12353;
  assign n12339 = n11007 & n12354;
  assign n12334 = n11007 & n12355;
  assign n6988 = ~n5277;
  assign n8006 = ~n5138;
  assign n6700 = ~n6050;
  assign n6711 = ~n6144;
  assign n6957 = ~n5068;
  assign n6968 = ~n6247;
  assign n6962 = ~n6227;
  assign n6999 = ~n6425;
  assign n6972 = ~n6273;
  assign n11093 = ~n12356;
  assign n12332 = n11007 & n12357;
  assign n12333 = n11007 & n12358;
  assign n6995 = ~n6118;
  assign n12340 = n11007 & n12359;
  assign n12331 = n11007 & n12360;
  assign n11083 = ~n12361;
  assign n6958 = ~n6304;
  assign n11091 = ~n12362;
  assign n6996 = ~n6149;
  assign n12295 = ~n12374;
  assign n11099 = ~n12363;
  assign n6975 = ~n5249;
  assign n11089 = ~n12364;
  assign n6983 = ~n6358;
  assign n6997 = ~n5299;
  assign n11075 = ~n12365;
  assign n12336 = n11007 & n12366;
  assign n6956 = ~n6221;
  assign n7000 = ~n5028;
  assign n11087 = ~n12367;
  assign n11334 = ~n12327;
  assign n11065 = ~n10228;
  assign n6984 = ~n5209;
  assign n11073 = ~n12368;
  assign n11079 = ~n12369;
  assign n12284 = n7004 & n32;
  assign n12335 = n11007 & n12370;
  assign n12342 = n11007 & n12371;
  assign n6966 = ~n6423;
  assign n7002 = ~n5052;
  assign n6977 = ~n6315;
  assign n11101 = ~n12372;
  assign n6981 = ~n6158;
  assign n11071 = ~n12373;
  assign n12008 = n12126 & n22;
  assign n11267 = n12127 & n10962;
  assign n11642 = n12128 & n11000;
  assign n11844 = n12129 & n10974;
  assign n11758 = n12130 & n14;
  assign n11541 = n12131 & n16;
  assign n12123 = n12133 & n15;
  assign n11955 = n12128 & n10977;
  assign n11111 = n12134 & n10;
  assign n11372 = n12129 & n10997;
  assign n12066 = n12134 & n21;
  assign n11250 = n12136 & n10961;
  assign n12094 = n12128 & n10959;
  assign n11275 = n12137 & n10999;
  assign n11614 = n12137 & n10981;
  assign n11221 = n12138 & n11005;
  assign n11852 = n12139 & n20;
  assign n11851 = n12140 & n30;
  assign n11820 = n12134 & n12;
  assign n11443 = n12130 & n10;
  assign n12043 = n12142 & n23;
  assign n11144 = n12143 & n10969;
  assign n11814 = n12134 & n28;
  assign n11829 = n12140 & n11;
  assign n11170 = n12133 & n9;
  assign n11429 = n12144 & n10962;
  assign n11364 = n12143 & n10989;
  assign n11556 = n12145 & n10959;
  assign n11230 = n12146 & n21;
  assign n11300 = n12129 & n10973;
  assign n11188 = n12147 & n5;
  assign n11617 = n12145 & n11000;
  assign n11621 = n12137 & n10957;
  assign n11168 = n12126 & n17;
  assign n11784 = n12148 & n10996;
  assign n11653 = n12130 & n17;
  assign n11173 = n12148 & n11005;
  assign n11591 = n12149 & n10990;
  assign n11962 = n12147 & n7;
  assign n11688 = n12150 & n20;
  assign n11366 = n12151 & n10965;
  assign n11394 = n12145 & n10979;
  assign n11505 = n12138 & n10977;
  assign n11874 = n12126 & n16;
  assign n11384 = n12147 & n26;
  assign n11590 = n12144 & n10952;
  assign n11791 = n12134 & n8;
  assign n11859 = n12152 & n3;
  assign n11728 = n12152 & n18;
  assign n11607 = n12128 & n10963;
  assign n11873 = n12153 & n15;
  assign n12020 = n12154 & n10977;
  assign n12067 = n12143 & n11005;
  assign n11440 = n12131 & n5;
  assign n11523 = n12126 & n5;
  assign n11139 = n12127 & n10959;
  assign n11322 = n12140 & n18;
  assign n11245 = n12149 & n9939;
  assign n11474 = n12146 & n24;
  assign n11839 = n12133 & n30;
  assign n11495 = n12128 & n10992;
  assign n11298 = n12150 & n11;
  assign n11836 = n12150 & n12;
  assign n12049 = n12140 & n20;
  assign n11268 = n12149 & n10954;
  assign n12064 = n12127 & n9939;
  assign n11572 = n12130 & n6;
  assign n11175 = n12136 & n10949;
  assign n12116 = n12140 & n6;
  assign n11378 = n12154 & n11000;
  assign n11449 = n12155 & n10992;
  assign n11684 = n12156 & n18;
  assign n11731 = n12133 & n25;
  assign n11659 = n12147 & n22;
  assign n11757 = n12156 & n19;
  assign n11244 = n12150 & n27;
  assign n11206 = n12154 & n10979;
  assign n11783 = n12152 & n24;
  assign n11813 = n12139 & n4;
  assign n11373 = n12157 & n10971;
  assign n12039 = n12156 & n2;
  assign n11317 = n12136 & n9939;
  assign n11468 = n12154 & n11005;
  assign n12080 = n12155 & n10952;
  assign n11521 = n12148 & n10959;
  assign n11699 = n12133 & n18;
  assign n11908 = n12126 & n21;
  assign n11557 = n12143 & n10966;
  assign n11507 = n12155 & n10972;
  assign n11509 = n12145 & n10954;
  assign n11216 = n12155 & n9939;
  assign n11877 = n12143 & n10972;
  assign n11239 = n12152 & n23;
  assign n11626 = n12157 & n10962;
  assign n12061 = n12155 & n10962;
  assign n11876 = n12146 & n11;
  assign n11123 = n12127 & n10966;
  assign n11426 = n12138 & n10972;
  assign n11675 = n12156 & n7;
  assign n12095 = n12147 & n18;
  assign n11549 = n12157 & n10972;
  assign n11819 = n12139 & n31;
  assign n11946 = n12139 & n22;
  assign n11790 = n12134 & n23;
  assign n11938 = n12147 & n9;
  assign n11910 = n12131 & n21;
  assign n11589 = n12129 & n10949;
  assign n11855 = n12134 & n9;
  assign n11539 = n12151 & n10996;
  assign n11700 = n12134 & n30;
  assign n11587 = n12145 & n10949;
  assign n11148 = n12151 & n10994;
  assign n11548 = n12142 & n25;
  assign n11542 = n12154 & n10969;
  assign n11424 = n12129 & n10963;
  assign n11463 = n12149 & n10992;
  assign n11948 = n12145 & n10996;
  assign n11725 = n12126 & n30;
  assign n11446 = n12144 & n10949;
  assign n11260 = n12151 & n10992;
  assign n11132 = n12153 & n10;
  assign n11550 = n12136 & n10959;
  assign n11297 = n12134 & n20;
  assign n11183 = n12151 & n11004;
  assign n12074 = n12143 & n10974;
  assign n11179 = n12152 & n17;
  assign n11568 = n12146 & n25;
  assign n11409 = n12137 & n10977;
  assign n11402 = n12155 & n10994;
  assign n11125 = n12137 & n10965;
  assign n11433 = n12149 & n10972;
  assign n11309 = n12130 & n2;
  assign n11160 = n12151 & n10954;
  assign n11525 = n12153 & n21;
  assign n11737 = n12140 & n31;
  assign n11365 = n12155 & n11005;
  assign n11760 = n12154 & n10961;
  assign n11276 = n12138 & n10971;
  assign n11871 = n12139 & n30;
  assign n11734 = n12142 & n11;
  assign n11743 = n12126 & n2;
  assign n11376 = n12137 & n10972;
  assign n11395 = n12137 & n10988;
  assign n11520 = n12140 & n12;
  assign n11857 = n12134 & n5;
  assign n11296 = n12148 & n10961;
  assign n11255 = n12147 & n14;
  assign n11278 = n12143 & n10992;
  assign n11214 = n12138 & n10961;
  assign n11696 = n12131 & n14;
  assign n11517 = n12158 & n11;
  assign n11577 = n12145 & n10965;
  assign n11455 = n12145 & n10990;
  assign n11360 = n12149 & n11004;
  assign n11800 = n12130 & n24;
  assign n11545 = n12151 & n10989;
  assign n11664 = n12156 & n23;
  assign n11996 = n12150 & n16;
  assign n11532 = n12151 & n10997;
  assign n11131 = n12146 & n14;
  assign n11724 = n12158 & n22;
  assign n11697 = n12147 & n15;
  assign n11442 = n12149 & n10996;
  assign n11182 = n12127 & n10992;
  assign n11315 = n12152 & n25;
  assign n11226 = n12157 & n10959;
  assign n11115 = n12144 & n11003;
  assign n12065 = n12142 & n17;
  assign n12016 = n12152 & n16;
  assign n12019 = n12142 & n6;
  assign n11211 = n12126 & n15;
  assign n11686 = n12150 & n15;
  assign n11515 = n12151 & n10973;
  assign n11894 = n12146 & n18;
  assign n12120 = n12139 & n2;
  assign n11405 = n12145 & n10997;
  assign n11708 = n12150 & n2;
  assign n11253 = n12140 & n22;
  assign n11205 = n12142 & n14;
  assign n11674 = n12130 & n18;
  assign n11143 = n12136 & n10996;
  assign n11914 = n12148 & n10979;
  assign n11552 = n12137 & n10954;
  assign n11909 = n12138 & n10974;
  assign n11679 = n12148 & n10974;
  assign n11622 = n12131 & n23;
  assign n11251 = n12142 & n5;
  assign n11274 = n12129 & n10971;
  assign n12115 = n12140 & n9;
  assign n11325 = n12142 & n21;
  assign n11146 = n12157 & n9939;
  assign n11834 = n12153 & n18;
  assign n12068 = n12156 & n22;
  assign n12050 = n12150 & n26;
  assign n12119 = n12134 & n7;
  assign n11238 = n12157 & n10973;
  assign n11768 = n12133 & n31;
  assign n11511 = n12129 & n10957;
  assign n11887 = n12148 & n10962;
  assign n11553 = n12136 & n10963;
  assign n12104 = n12157 & n11005;
  assign n11693 = n12156 & n27;
  assign n11625 = n12152 & n26;
  assign n11733 = n12149 & n10971;
  assign n12057 = n12138 & n10966;
  assign n11282 = n12138 & n11003;
  assign n11262 = n12127 & n10989;
  assign n11258 = n12146 & n7;
  assign n11257 = n12136 & n10954;
  assign n11281 = n12138 & n10994;
  assign n11907 = n12149 & n11005;
  assign n11504 = n12145 & n11004;
  assign n11611 = n12136 & n10973;
  assign n11573 = n12130 & n21;
  assign n11538 = n12129 & n10989;
  assign n11242 = n12146 & n8;
  assign n11945 = n12152 & n5;
  assign n11904 = n12151 & n9939;
  assign n11736 = n12126 & n13;
  assign n11303 = n12131 & n11;
  assign n11499 = n12130 & n3;
  assign n11727 = n12146 & n28;
  assign n11831 = n12158 & n19;
  assign n11285 = n12128 & n9939;
  assign n11286 = n12156 & n15;
  assign n11514 = n12129 & n11000;
  assign n11940 = n12127 & n11005;
  assign n11729 = n12142 & n24;
  assign n11492 = n12144 & n10994;
  assign n11135 = n12144 & n10981;
  assign n12075 = n12148 & n10965;
  assign n11761 = n12158 & n2;
  assign n11218 = n12133 & n14;
  assign n12055 = n12150 & n7;
  assign n11690 = n12158 & n7;
  assign n11406 = n12129 & n10979;
  assign n11830 = n12150 & n22;
  assign n11155 = n12147 & n4;
  assign n11269 = n12140 & n16;
  assign n11991 = n12153 & n31;
  assign n12078 = n12142 & n31;
  assign n11646 = n12142 & n27;
  assign n12005 = n12149 & n10974;
  assign n11954 = n12149 & n10969;
  assign n11763 = n12147 & n19;
  assign n11689 = n12140 & n4;
  assign n11191 = n12136 & n10990;
  assign n11601 = n12145 & n10969;
  assign n11987 = n12146 & n26;
  assign n11338 = n12144 & n10990;
  assign n11256 = n12130 & n30;
  assign n11990 = n12147 & n13;
  assign n11762 = n12128 & n10969;
  assign n11796 = n12158 & n13;
  assign n11892 = n12142 & n29;
  assign n11585 = n12142 & n15;
  assign n11751 = n12152 & n11;
  assign n11321 = n12146 & n22;
  assign n11837 = n12156 & n13;
  assign n11672 = n12130 & n31;
  assign n11326 = n12145 & n10972;
  assign n12017 = n12138 & n10981;
  assign n11362 = n12148 & n10972;
  assign n11217 = n12139 & n6;
  assign n11973 = n12139 & n27;
  assign n11164 = n12158 & n10;
  assign n11172 = n12146 & n13;
  assign n11287 = n12153 & n12;
  assign n12030 = n12130 & n27;
  assign n11512 = n12137 & n10952;
  assign n11403 = n12137 & n11004;
  assign n11192 = n12137 & n10966;
  assign n11236 = n12144 & n10996;
  assign n11219 = n12151 & n10979;
  assign n11252 = n12129 & n10992;
  assign n11534 = n12136 & n10994;
  assign n11158 = n12154 & n10989;
  assign n11655 = n12139 & n17;
  assign n11543 = n12151 & n10990;
  assign n11469 = n12136 & n10965;
  assign n11289 = n12152 & n15;
  assign n11259 = n12157 & n10952;
  assign n12097 = n12152 & n29;
  assign n11723 = n12147 & n21;
  assign n11698 = n12158 & n1;
  assign n11412 = n12136 & n10997;
  assign n11201 = n12153 & n11;
  assign n11311 = n12144 & n10965;
  assign n11869 = n12154 & n10965;
  assign n11453 = n12140 & n5;
  assign n11858 = n12133 & n3;
  assign n11209 = n12137 & n11000;
  assign n11397 = n12129 & n10977;
  assign n11234 = n12156 & n16;
  assign n11126 = n12140 & n24;
  assign n11650 = n12143 & n9939;
  assign n11475 = n12149 & n10963;
  assign n11110 = n12156 & n12;
  assign n11107 = n12143 & n10971;
  assign n11220 = n12130 & n28;
  assign n11306 = n12147 & n6;
  assign n11254 = n12137 & n11005;
  assign n11213 = n12136 & n10969;
  assign n11263 = n12150 & n4;
  assign n12087 = n12136 & n10989;
  assign n11330 = n12157 & n10979;
  assign n11243 = n12143 & n11000;
  assign n12112 = n12146 & n31;
  assign n11464 = n12155 & n10999;
  assign n11392 = n12138 & n10957;
  assign n11826 = n12139 & n3;
  assign n11578 = n12148 & n10981;
  assign n11452 = n12154 & n10997;
  assign n12109 = n12139 & n18;
  assign n11307 = n12142 & n28;
  assign n11189 = n12148 & n10963;
  assign n11456 = n12155 & n10961;
  assign n11726 = n12133 & n29;
  assign n11524 = n12138 & n10962;
  assign n11347 = n12150 & n17;
  assign n11695 = n12131 & n30;
  assign n11312 = n12147 & n31;
  assign n11775 = n12156 & n8;
  assign n12096 = n12129 & n10959;
  assign n11756 = n12133 & n21;
  assign n12018 = n12133 & n1;
  assign n11603 = n12154 & n10988;
  assign n11290 = n12150 & n9;
  assign n11627 = n12155 & n11004;
  assign n11853 = n12130 & n25;
  assign n11151 = n12137 & n10996;
  assign n11140 = n12153 & n2;
  assign n11116 = n12146 & n1;
  assign n11416 = n12129 & n10969;
  assign n11640 = n12128 & n10957;
  assign n11157 = n12146 & n2;
  assign n11414 = n12136 & n10979;
  assign n11197 = n12155 & n10981;
  assign n12007 = n12137 & n10989;
  assign n11235 = n12143 & n10988;
  assign n11974 = n12134 & n17;
  assign n11842 = n12153 & n9;
  assign n11594 = n12144 & n10972;
  assign n11313 = n12136 & n11005;
  assign n11202 = n12129 & n10988;
  assign n11380 = n12145 & n10994;
  assign n11988 = n12126 & n14;
  assign n11497 = n12144 & n10973;
  assign n11795 = n12150 & n13;
  assign n12077 = n12140 & n13;
  assign n11413 = n12137 & n10961;
  assign n11215 = n12128 & n10972;
  assign n11984 = n12149 & n10957;
  assign n11639 = n12158 & n23;
  assign n11371 = n12128 & n10997;
  assign n11367 = n12144 & n10966;
  assign n11706 = n12150 & n24;
  assign n11812 = n12142 & n1;
  assign n11998 = n12144 & n10974;
  assign n11546 = n12143 & n10962;
  assign n11224 = n12144 & n10954;
  assign n11162 = n12154 & n10990;
  assign n11863 = n12147 & n23;
  assign n11310 = n12153 & n22;
  assign n11799 = n12158 & n12;
  assign n11802 = n12156 & n30;
  assign n11906 = n12143 & n10949;
  assign n11559 = n12149 & n10962;
  assign n11266 = n12142 & n18;
  assign n11122 = n12146 & n12;
  assign n11533 = n12144 & n10969;
  assign n11584 = n12144 & n10988;
  assign n11501 = n12128 & n10965;
  assign n12047 = n12134 & n16;
  assign n11379 = n12127 & n11000;
  assign n12003 = n12153 & n17;
  assign n11561 = n12157 & n10988;
  assign n11425 = n12137 & n11003;
  assign n11658 = n12133 & n28;
  assign n11357 = n12138 & n10989;
  assign n11503 = n12128 & n11005;
  assign n11701 = n12158 & n4;
  assign n11391 = n12138 & n10979;
  assign n11323 = n12131 & n28;
  assign n11133 = n12144 & n10997;
  assign n11500 = n12145 & n10963;
  assign n11393 = n12156 & n24;
  assign n11754 = n12150 & n5;
  assign n11953 = n12144 & n10977;
  assign n11558 = n12128 & n10962;
  assign n11370 = n12142 & n9;
  assign n11119 = n12142 & n4;
  assign n11588 = n12154 & n10994;
  assign n12121 = n12134 & n19;
  assign n11891 = n12131 & n20;
  assign n11369 = n12129 & n10962;
  assign n11823 = n12139 & n24;
  assign n11510 = n12150 & n19;
  assign n11964 = n12138 & n10990;
  assign n11586 = n12128 & n10999;
  assign n11537 = n12127 & n10974;
  assign n11161 = n12156 & n17;
  assign n11461 = n12153 & n13;
  assign n12070 = n12146 & n4;
  assign n11608 = n12157 & n10963;
  assign n11732 = n12140 & n3;
  assign n11454 = n12154 & n10959;
  assign n11579 = n12144 & n10999;
  assign n11536 = n12151 & n10962;
  assign n11193 = n12144 & n10961;
  assign n11609 = n12153 & n23;
  assign n11294 = n12151 & n10999;
  assign n11551 = n12146 & n17;
  assign n11632 = n12139 & n23;
  assign n11417 = n12139 & n25;
  assign n11544 = n12131 & n19;
  assign n11363 = n12150 & n29;
  assign n11470 = n12146 & n5;
  assign n11445 = n12145 & n10989;
  assign n11194 = n12136 & n10957;
  assign n11227 = n12157 & n10961;
  assign n11660 = n12150 & n6;
  assign n12032 = n12148 & n10990;
  assign n11527 = n12156 & n4;
  assign n11434 = n12144 & n11005;
  assign n11195 = n12152 & n19;
  assign n11522 = n12126 & n10;
  assign n11261 = n12151 & n10963;
  assign n11481 = n12155 & n11000;
  assign n11595 = n12126 & n9;
  assign n11498 = n12154 & n10974;
  assign n11518 = n12128 & n10949;
  assign n12045 = n12147 & n12;
  assign n11437 = n12136 & n10977;
  assign n11368 = n12145 & n10966;
  assign n11422 = n12137 & n10979;
  assign n11399 = n12155 & n10989;
  assign n11401 = n12138 & n10996;
  assign n11827 = n12131 & n15;
  assign n11979 = n12131 & n9;
  assign n11432 = n12131 & n17;
  assign n11661 = n12137 & n10959;
  assign n12084 = n12157 & n10957;
  assign n11506 = n12128 & n10966;
  assign n11305 = n12158 & n5;
  assign n12114 = n12133 & n17;
  assign n11335 = n12153 & n26;
  assign n11516 = n12127 & n10977;
  assign n11770 = n12142 & n19;
  assign n11759 = n12134 & n25;
  assign n11508 = n12143 & n10965;
  assign n11411 = n12137 & n10992;
  assign n11937 = n12152 & n14;
  assign n11845 = n12142 & n7;
  assign n11847 = n12152 & n13;
  assign n11436 = n12157 & n10997;
  assign n11676 = n12142 & n2;
  assign n11109 = n12134 & n11;
  assign n11581 = n12147 & n27;
  assign n11890 = n12130 & n5;
  assign n11124 = n12140 & n23;
  assign n11375 = n12145 & n10957;
  assign n12124 = n12158 & n17;
  assign n11237 = n12146 & n16;
  assign n11153 = n12129 & n11003;
  assign n11540 = n12149 & n10965;
  assign n11624 = n12154 & n10992;
  assign n11324 = n12127 & n10988;
  assign n11560 = n12145 & n10999;
  assign n11654 = n12152 & n21;
  assign n11496 = n12144 & n10979;
  assign n11410 = n12147 & n8;
  assign n11471 = n12155 & n10959;
  assign n11273 = n12148 & n9939;
  assign n11566 = n12147 & n2;
  assign n11969 = n12150 & n21;
  assign n11896 = n12126 & n28;
  assign n11473 = n12143 & n10977;
  assign n11883 = n12139 & n13;
  assign n11833 = n12158 & n28;
  assign n11576 = n12136 & n10981;
  assign n12004 = n12158 & n9;
  assign n11668 = n12156 & n5;
  assign n11482 = n12133 & n5;
  assign n12072 = n12157 & n11004;
  assign n11600 = n12129 & n10972;
  assign n11912 = n12131 & n1;
  assign n11704 = n12130 & n29;
  assign n11240 = n12152 & n20;
  assign n11295 = n12127 & n10973;
  assign n11620 = n12139 & n16;
  assign n11478 = n12127 & n10999;
  assign n11163 = n12140 & n26;
  assign n11400 = n12152 & n31;
  assign n11806 = n12154 & n11003;
  assign n11941 = n12148 & n11003;
  assign n11749 = n12131 & n3;
  assign n11707 = n12146 & n15;
  assign n11604 = n12151 & n11005;
  assign n11810 = n12139 & n29;
  assign n12076 = n12156 & n10;
  assign n11486 = n12157 & n10977;
  assign n11702 = n12139 & n10;
  assign n11174 = n12140 & n7;
  assign n11304 = n12140 & n21;
  assign n11292 = n12136 & n11003;
  assign n11662 = n12134 & n3;
  assign n11476 = n12148 & n10997;
  assign n11742 = n12140 & n17;
  assign n11747 = n12152 & n27;
  assign n11288 = n12134 & n26;
  assign n11899 = n12154 & n10999;
  assign n11994 = n12156 & n29;
  assign n11299 = n12142 & n16;
  assign n11861 = n12147 & n17;
  assign n11169 = n12149 & n10949;
  assign n11901 = n12157 & n11003;
  assign n11615 = n12130 & n13;
  assign n11744 = n12145 & n10971;
  assign n12105 = n12129 & n10954;
  assign n12090 = n12153 & n14;
  assign n12111 = n12158 & n8;
  assign n12086 = n12151 & n11003;
  assign n12046 = n12149 & n10979;
  assign n12083 = n12131 & n12;
  assign n12052 = n12154 & n10952;
  assign n12073 = n12126 & n7;
  assign n11815 = n12139 & n9;
  assign n11716 = n12146 & n29;
  assign n11293 = n12143 & n10957;
  assign n11134 = n12137 & n10949;
  assign n11479 = n12157 & n10974;
  assign n11316 = n12131 & n2;
  assign n11712 = n12139 & n11;
  assign n11149 = n12138 & n9939;
  assign n11777 = n12133 & n24;
  assign n12071 = n12158 & n14;
  assign n11888 = n12133 & n6;
  assign n11222 = n12153 & n16;
  assign n11967 = n12129 & n10961;
  assign n11748 = n12147 & n3;
  assign n11547 = n12153 & n20;
  assign n11489 = n12155 & n10957;
  assign n11862 = n12134 & n14;
  assign n11767 = n12136 & n10992;
  assign n12092 = n12134 & n18;
  assign n11447 = n12151 & n10959;
  assign n11975 = n12130 & n9;
  assign n11792 = n12139 & n26;
  assign n11786 = n12131 & n6;
  assign n11860 = n12142 & n13;
  assign n11381 = n12154 & n10973;
  assign n11203 = n12138 & n10952;
  assign n11746 = n12153 & n6;
  assign n11241 = n12138 & n10997;
  assign n11633 = n12158 & n30;
  assign n11911 = n12148 & n10988;
  assign n11352 = n12145 & n10961;
  assign n11687 = n12131 & n4;
  assign n12048 = n12136 & n10952;
  assign n11893 = n12155 & n10990;
  assign n11494 = n12151 & n10952;
  assign n11878 = n12147 & n20;
  assign n12091 = n12130 & n19;
  assign n11919 = n12128 & n10990;
  assign n11223 = n12126 & n3;
  assign n11816 = n12150 & n23;
  assign n11772 = n12127 & n10965;
  assign n11936 = n12140 & n8;
  assign n11270 = n12157 & n10969;
  assign n11480 = n12146 & n30;
  assign n11952 = n12133 & n27;
  assign n11526 = n12127 & n10954;
  assign n11854 = n12150 & n1;
  assign n11619 = n12153 & n4;
  assign n11850 = n12144 & n11000;
  assign n12028 = n12130 & n7;
  assign n12015 = n12139 & n8;
  assign n11670 = n12133 & n12;
  assign n11458 = n12154 & n10954;
  assign n11374 = n12151 & n10974;
  assign n11868 = n12142 & n8;
  assign n11355 = n12154 & n10971;
  assign n11118 = n12126 & n19;
  assign n11711 = n12133 & n2;
  assign n11648 = n12145 & n9939;
  assign n11947 = n12140 & n27;
  assign n11565 = n12149 & n10959;
  assign n11450 = n12151 & n10961;
  assign n11567 = n12144 & n10963;
  assign n11444 = n12157 & n10965;
  assign n11483 = n12157 & n10996;
  assign n11407 = n12136 & n10999;
  assign n11198 = n12133 & n4;
  assign n11824 = n12131 & n25;
  assign n11881 = n12158 & n24;
  assign n11821 = n12153 & n30;
  assign n11848 = n12145 & n10981;
  assign n11752 = n12134 & n24;
  assign n12103 = n12158 & n25;
  assign n11977 = n12152 & n10;
  assign n11832 = n12139 & n5;
  assign n11184 = n12127 & n10994;
  assign n12056 = n12126 & n23;
  assign n11685 = n12139 & n15;
  assign n11875 = n12131 & n31;
  assign n11818 = n12153 & n19;
  assign n11142 = n12139 & n7;
  assign n11843 = n12142 & n20;
  assign n11838 = n12142 & n3;
  assign n11755 = n12146 & n27;
  assign n11319 = n12144 & n9939;
  assign n11117 = n12152 & n30;
  assign n11985 = n12153 & n3;
  assign n12100 = n12148 & n10971;
  assign n11905 = n12156 & n6;
  assign n11872 = n12138 & n10973;
  assign n11448 = n12143 & n10973;
  assign n12088 = n12131 & n27;
  assign n11356 = n12151 & n10977;
  assign n11663 = n12133 & n8;
  assign n11435 = n12127 & n10969;
  assign n11694 = n12146 & n9;
  assign n11472 = n12143 & n10996;
  assign n12079 = n12153 & n7;
  assign n12006 = n12151 & n10972;
  assign n11531 = n12146 & n10;
  assign n11420 = n12155 & n10965;
  assign n11308 = n12130 & n20;
  assign n11502 = n12154 & n10963;
  assign n11864 = n12153 & n5;
  assign n11913 = n12142 & n30;
  assign n11835 = n12140 & n28;
  assign n11741 = n12131 & n26;
  assign n11788 = n12150 & n28;
  assign n11519 = n12128 & n10979;
  assign n11804 = n12150 & n10;
  assign n11709 = n12152 & n1;
  assign n11377 = n12151 & n10969;
  assign n11284 = n12143 & n10963;
  assign n11703 = n12133 & n11;
  assign n11636 = n12157 & n10966;
  assign n11383 = n12158 & n31;
  assign n11886 = n12127 & n10997;
  assign n11950 = n12129 & n10952;
  assign n12037 = n12134 & n13;
  assign n11419 = n12154 & n10962;
  assign n11459 = n12136 & n10966;
  assign n11999 = n12126 & n4;
  assign n11885 = n12153 & n25;
  assign n11580 = n12151 & n10981;
  assign n11102 = n12149 & n10999;
  assign n11943 = n12133 & n16;
  assign n12038 = n12148 & n10992;
  assign n11225 = n12150 & n8;
  assign n11785 = n12127 & n10996;
  assign n11171 = n12137 & n10963;
  assign n11154 = n12139 & n21;
  assign n12027 = n12156 & n26;
  assign n11388 = n12137 & n10997;
  assign n11822 = n12134 & n22;
  assign n11961 = n12129 & n11005;
  assign n11265 = n12128 & n10952;
  assign n11605 = n12157 & n10992;
  assign n11349 = n12143 & n10999;
  assign n11248 = n12129 & n9939;
  assign n11972 = n12133 & n19;
  assign n11966 = n12144 & n10989;
  assign n11740 = n12147 & n24;
  assign n11981 = n12131 & n7;
  assign n11196 = n12128 & n10974;
  assign n11797 = n12147 & n30;
  assign n11635 = n12157 & n10990;
  assign n11616 = n12129 & n10990;
  assign n11466 = n12155 & n11003;
  assign n11493 = n12134 & n4;
  assign n11722 = n12131 & n13;
  assign n11465 = n12131 & n8;
  assign n11773 = n12130 & n11;
  assign n11264 = n12156 & n28;
  assign n11673 = n12126 & n1;
  assign n11867 = n12158 & n26;
  assign n11487 = n12155 & n10974;
  assign n12041 = n12147 & n28;
  assign n11598 = n12128 & n11004;
  assign n11421 = n12127 & n11003;
  assign n11127 = n12148 & n10973;
  assign n11968 = n12133 & n20;
  assign n11575 = n12127 & n10957;
  assign n11922 = n12126 & n20;
  assign n11825 = n12138 & n10965;
  assign n11346 = n12128 & n10981;
  assign n11150 = n12145 & n10988;
  assign n11884 = n12126 & n25;
  assign n11717 = n12150 & n25;
  assign n11345 = n12156 & n14;
  assign n11918 = n12145 & n11005;
  assign n11618 = n12134 & n15;
  assign n11880 = n12130 & n16;
  assign n11112 = n12137 & n10969;
  assign n12001 = n12153 & n1;
  assign n11986 = n12158 & n21;
  assign n11190 = n12149 & n11000;
  assign n11408 = n12149 & n10961;
  assign n11715 = n12146 & n23;
  assign n12035 = n12136 & n10974;
  assign n11634 = n12155 & n10988;
  assign n11631 = n12137 & n10971;
  assign n11491 = n12151 & n10949;
  assign n11900 = n12144 & n10992;
  assign n11389 = n12154 & n10957;
  assign n12034 = n12129 & n10996;
  assign n11978 = n12158 & n27;
  assign n11571 = n12154 & n10981;
  assign n11204 = n12129 & n11004;
  assign n11460 = n12149 & n10977;
  assign n11720 = n12152 & n4;
  assign n11993 = n12149 & n10989;
  assign n11530 = n12155 & n10979;
  assign n12051 = n12129 & n10999;
  assign n11705 = n12133 & n22;
  assign n12014 = n12158 & n18;
  assign n11207 = n12136 & n10971;
  assign n11680 = n12140 & n10;
  assign n11613 = n12148 & n10966;
  assign n11710 = n12152 & n28;
  assign n11682 = n12134 & n6;
  assign n12113 = n12145 & n10973;
  assign n11669 = n12126 & n8;
  assign n12042 = n12150 & n3;
  assign n11529 = n12128 & n10961;
  assign n11415 = n12128 & n10996;
  assign n12029 = n12126 & n24;
  assign n11348 = n12155 & n10971;
  assign n11354 = n12145 & n10952;
  assign n11927 = n12126 & n31;
  assign n11771 = n12140 & n25;
  assign n11730 = n12154 & n10966;
  assign n11778 = n12148 & n11000;
  assign n11879 = n12139 & n12;
  assign n11849 = n12140 & n19;
  assign n11959 = n12144 & n10959;
  assign n11467 = n12143 & n10990;
  assign n11485 = n12145 & n11003;
  assign n11353 = n12155 & n10973;
  assign n11957 = n12148 & n10994;
  assign n11457 = n12143 & n11004;
  assign n12040 = n12128 & n10971;
  assign n11939 = n12129 & n10994;
  assign n11513 = n12136 & n11004;
  assign n11130 = n12146 & n19;
  assign n11870 = n12138 & n10963;
  assign n12033 = n12144 & n11004;
  assign n11178 = n12133 & n26;
  assign n11246 = n12131 & n10;
  assign n11187 = n12137 & n10973;
  assign n11314 = n12143 & n10981;
  assign n11120 = n12127 & n10981;
  assign n11965 = n12158 & n29;
  assign n11441 = n12149 & n10973;
  assign n11484 = n12149 & n11003;
  assign n11105 = n12155 & n10963;
  assign n11681 = n12138 & n11004;
  assign n11992 = n12145 & n10977;
  assign n11606 = n12149 & n10952;
  assign n11971 = n12128 & n10954;
  assign n11902 = n12148 & n10957;
  assign n12025 = n12138 & n10969;
  assign n12118 = n12130 & n4;
  assign n11358 = n12148 & n10977;
  assign n11995 = n12143 & n10997;
  assign n11846 = n12158 & n3;
  assign n12023 = n12128 & n10989;
  assign n12069 = n12137 & n10994;
  assign n11638 = n12157 & n10989;
  assign n11769 = n12133 & n7;
  assign n12098 = n12146 & n6;
  assign n11721 = n12131 & n22;
  assign n11477 = n12151 & n11000;
  assign n11649 = n12137 & n9939;
  assign n12110 = n12136 & n10972;
  assign n11623 = n12138 & n10949;
  assign n11641 = n12157 & n10949;
  assign n12024 = n12154 & n11004;
  assign n11942 = n12143 & n11003;
  assign n11789 = n12139 & n1;
  assign n11350 = n12136 & n10962;
  assign n11210 = n12148 & n10999;
  assign n11718 = n12152 & n22;
  assign n11283 = n12155 & n10966;
  assign n12053 = n12136 & n10988;
  assign n11361 = n12157 & n10954;
  assign n12009 = n12157 & n10999;
  assign n11776 = n12151 & n10971;
  assign n11980 = n12140 & n2;
  assign n12054 = n12157 & n11000;
  assign n11351 = n12154 & n10972;
  assign n11811 = n12126 & n27;
  assign n12085 = n12153 & n28;
  assign n11949 = n12128 & n11003;
  assign n11989 = n12131 & n24;
  assign n11803 = n12150 & n14;
  assign n11610 = n12129 & n10965;
  assign n11753 = n12140 & n15;
  assign n11960 = n12139 & n28;
  assign n12060 = n12140 & n1;
  assign n12031 = n12134 & n1;
  assign n11780 = n12126 & n11;
  assign n12122 = n12150 & n18;
  assign n11180 = n12139 & n19;
  assign n11793 = n12156 & n20;
  assign n11882 = n12127 & n11004;
  assign n11841 = n12156 & n31;
  assign n11554 = n12127 & n10972;
  assign n11774 = n12156 & n11;
  assign n11612 = n12152 & n12;
  assign n11387 = n12144 & n10957;
  assign n11764 = n12148 & n10969;
  assign n11856 = n12130 & n23;
  assign n11199 = n12156 & n1;
  assign n11766 = n12126 & n6;
  assign n11535 = n12130 & n12;
  assign n11106 = n12127 & n10961;
  assign n11944 = n12147 & n1;
  assign n11569 = n12145 & n10962;
  assign n11599 = n12155 & n10977;
  assign n12011 = n12151 & n10957;
  assign n11794 = n12158 & n16;
  assign n12093 = n12131 & n18;
  assign n11765 = n12157 & n10994;
  assign n11186 = n12127 & n10949;
  assign n12022 = n12151 & n10966;
  assign n11108 = n12139 & n14;
  assign n11145 = n12150 & n31;
  assign n11817 = n12156 & n9;
  assign n11597 = n12137 & n10974;
  assign n11563 = n12137 & n10990;
  assign n12010 = n12149 & n10966;
  assign n11382 = n12138 & n10954;
  assign n12106 = n12155 & n10949;
  assign n12117 = n12147 & n16;
  assign n11805 = n12147 & n10;
  assign n12012 = n12133 & n10;
  assign n11398 = n12145 & n10974;
  assign n11665 = n12143 & n10959;
  assign n11958 = n12134 & n2;
  assign n11963 = n12130 & n8;
  assign n12082 = n12148 & n11004;
  assign n11596 = n12133 & n23;
  assign n11828 = n12158 & n20;
  assign n12044 = n12153 & n24;
  assign n11247 = n12127 & n10971;
  assign n11840 = n12152 & n7;
  assign n11562 = n12148 & n10952;
  assign n11396 = n12128 & n10994;
  assign n11630 = n12143 & n10961;
  assign n11779 = n12153 & n27;
  assign n12013 = n12148 & n10954;
  assign n11667 = n12131 & n29;
  assign n11570 = n12143 & n10994;
  assign n11976 = n12149 & n10988;
  assign n11951 = n12144 & n10971;
  assign n11647 = n12148 & n10989;
  assign n12026 = n12150 & n30;
  assign n11318 = n12148 & n10949;
  assign n11147 = n12142 & n10;
  assign n11678 = n12138 & n10992;
  assign n11956 = n12153 & n8;
  assign n11208 = n12152 & n8;
  assign n11564 = n12157 & n10981;
  assign n11666 = n12130 & n22;
  assign n11277 = n12126 & n29;
  assign n11787 = n12134 & n31;
  assign n11359 = n12149 & n10997;
  assign n11645 = n12138 & n10988;
  assign n11637 = n12154 & n10996;
  assign n11121 = n12147 & n11;
  assign n11185 = n12127 & n10952;
  assign n11801 = n12152 & n2;
  assign n12062 = n12142 & n26;
  assign n11671 = n12134 & n29;
  assign n11970 = n12128 & n10973;
  assign n11291 = n12128 & n10988;
  assign n11677 = n12156 & n25;
  assign n11782 = n12133 & n13;
  assign n11735 = n12142 & n22;
  assign n11781 = n12155 & n10996;
  assign n11915 = n12130 & n26;
  assign n11719 = n12142 & n12;
  assign n12021 = n12134 & n27;
  assign n11897 = n12126 & n12;
  assign n11683 = n12126 & n18;
  assign n11423 = n12143 & n10954;
  assign n12036 = n12153 & n29;
  assign n12099 = n12154 & n10949;
  assign n12000 = n12155 & n10954;
  assign n11583 = n12129 & n10966;
  assign n11997 = n12140 & n14;
  assign n12002 = n12151 & n10988;
  assign n11602 = n12138 & n11000;
  assign n11903 = n12152 & n6;
  assign n12081 = n12130 & n1;
  assign n11451 = n12145 & n10992;
  assign n11574 = n12149 & n10994;
  assign n12125 = n12126 & n26;
  assign n11745 = n12146 & n3;
  assign n11231 = n12136 & n11000;
  assign n11488 = n12156 & n21;
  assign n11404 = n12158 & n15;
  assign n11528 = n12129 & n10981;
  assign n11555 = n12155 & n10997;
  assign n12063 = n12138 & n10959;
  assign n11798 = n12130 & n15;
  assign n11582 = n12143 & n10952;
  assign n11462 = n12156 & n3;
  assign n11390 = n12149 & n10981;
  assign n11249 = n12158 & n6;
  assign n11200 = n12147 & n29;
  assign n11181 = n12127 & n10963;
  assign n11152 = n12137 & n10962;
  assign n11159 = n12146 & n20;
  assign n11418 = n12127 & n10990;
  assign n12089 = n12147 & n25;
  assign n11212 = n12155 & n10969;
  assign n11141 = n12154 & n9939;
  assign n11490 = n12127 & n10979;
  assign n11167 = n12138 & n10999;
  assign n11809 = n12152 & n9;
  assign n11895 = n12140 & n29;
  assign n11750 = n12143 & n10979;
  assign n9950 = ~n9706;
  assign n11592 = n12175 & n12176;
  assign n6994 = ~n6092;
  assign n7041 = ~n12127;
  assign n9944 = ~n9674;
  assign n7049 = ~n12143;
  assign n7010 = ~n12128;
  assign n11138 = n11081 & n12192;
  assign n7053 = ~n12137;
  assign n7047 = ~n12157;
  assign n9941 = ~n6360;
  assign n9946 = ~n9670;
  assign n11343 = n12199 & n12200;
  assign n11136 = n12201 & n12202;
  assign n6970 = ~n6192;
  assign n11128 = n12204 & n12205;
  assign n7027 = ~n12155;
  assign n9945 = ~n9188;
  assign n7057 = ~n12151;
  assign n7043 = ~n12129;
  assign n11165 = n12213 & n12214;
  assign n7045 = ~n12136;
  assign n7059 = ~n12148;
  assign n6974 = ~n6260;
  assign n11328 = n12222 & n12223;
  assign n11156 = n12224 & n12225;
  assign n11331 = n12228 & n12229;
  assign n7055 = ~n12145;
  assign n11339 = n12237 & n12238;
  assign n6982 = ~n6282;
  assign n9943 = ~n9672;
  assign n7003 = ~n6082;
  assign n11889 = n12253 & n12254;
  assign n7061 = ~n12144;
  assign n11103 = n12257 & n12258;
  assign n9948 = ~n9704;
  assign n7073 = ~n12138;
  assign n6986 = ~n6340;
  assign n11336 = n12260 & n12261;
  assign n11738 = n12270 & n12271;
  assign n7051 = ~n12149;
  assign n9947 = ~n9676;
  assign n11341 = n12275 & n12276;
  assign n9942 = ~n9684;
  assign n7039 = ~n12154;
  assign n12216 = n12278 & n11004;
  assign n11644 = ~n12281;
  assign n11233 = ~n12282;
  assign n12232 = n12284 & n11;
  assign n11917 = ~n12285;
  assign n12184 = n12278 & n10988;
  assign n12227 = n12284 & n31;
  assign n12172 = n12284 & n24;
  assign n11386 = ~n12288;
  assign n12102 = ~n12289;
  assign n11714 = ~n12290;
  assign n12195 = n12278 & n10969;
  assign n11229 = ~n12293;
  assign n12191 = n12278 & n10952;
  assign n12180 = n12278 & n10997;
  assign n11692 = ~n12294;
  assign n12188 = n12278 & n10954;
  assign n12197 = n12284 & n21;
  assign n7971 = n12295 & n33;
  assign n11657 = ~n12296;
  assign n11114 = ~n12298;
  assign n12181 = n12278 & n10962;
  assign n11431 = ~n12300;
  assign n12173 = n12284 & n3;
  assign n12269 = n12278 & n10959;
  assign n12171 = n12284 & n16;
  assign n12268 = n12284 & n20;
  assign n11629 = ~n12303;
  assign n11302 = ~n12304;
  assign n11439 = ~n12306;
  assign n12198 = n12278 & n10994;
  assign n12242 = n12284 & n6;
  assign n12193 = n12278 & n11007;
  assign n12190 = n12284 & n23;
  assign n12178 = n12284 & n1;
  assign n12183 = n12278 & n10966;
  assign n12220 = n12284 & n8;
  assign n11866 = ~n12308;
  assign n12255 = n12278 & n11003;
  assign n12249 = n12278 & n10974;
  assign n12196 = n12284 & n18;
  assign n11280 = ~n12310;
  assign n12259 = n12278 & n10971;
  assign n12262 = n12278 & n11000;
  assign n12186 = n12284 & n22;
  assign n12108 = ~n12311;
  assign n12174 = n12278 & n10977;
  assign n12248 = n12284 & n14;
  assign n12210 = n12284 & n17;
  assign n12236 = n12278 & n10999;
  assign n11808 = ~n12313;
  assign n12217 = n12278 & n10979;
  assign n12177 = n12284 & n9;
  assign n12211 = n12284 & n2;
  assign n12274 = n12278 & n10973;
  assign n12189 = n12278 & n10996;
  assign n12256 = n12284 & n26;
  assign n12218 = n12278 & n9939;
  assign n11428 = ~n12314;
  assign n11933 = ~n12315;
  assign n12240 = n12284 & n12;
  assign n12277 = n12284 & n5;
  assign n12215 = n12284 & n4;
  assign n12273 = n12278 & n11005;
  assign n11926 = ~n12316;
  assign n12187 = n12278 & n10989;
  assign n12239 = n12278 & n10965;
  assign n12219 = n12278 & n10963;
  assign n12209 = n12284 & n15;
  assign n12233 = n12284 & n19;
  assign n11983 = ~n12317;
  assign n12251 = n12284 & n29;
  assign n11652 = ~n12318;
  assign n12247 = n12284 & n13;
  assign n12208 = n12284 & n28;
  assign n12185 = n12284 & n27;
  assign n12212 = n12284 & n25;
  assign n12194 = n12278 & n10990;
  assign n11929 = ~n12319;
  assign n11931 = ~n12320;
  assign n12244 = n12278 & n10981;
  assign n11924 = ~n12321;
  assign n12267 = n12278 & n10972;
  assign n12252 = n12278 & n10957;
  assign n11272 = ~n12322;
  assign n12264 = n12278 & n10961;
  assign n11935 = ~n12323;
  assign n12263 = n12284 & n30;
  assign n12243 = n12284 & n7;
  assign n11177 = ~n12324;
  assign n12265 = n12278 & n10992;
  assign n11921 = ~n12325;
  assign n12059 = ~n12326;
  assign n12241 = n12278 & n10949;
  assign n12234 = n12284 & n10;
  assign n12182 = ~n12328;
  assign n12221 = ~n12329;
  assign n12266 = ~n12330;
  assign n12245 = ~n12331;
  assign n12203 = ~n12332;
  assign n12246 = ~n12333;
  assign n12235 = ~n12334;
  assign n12207 = ~n12335;
  assign n12272 = ~n12336;
  assign n12206 = ~n12337;
  assign n12231 = ~n12338;
  assign n12179 = ~n12339;
  assign n12226 = ~n12340;
  assign n12250 = ~n12341;
  assign n12230 = ~n12342;
  assign n8106 = ~n11102;
  assign n11006 = n11103 & n11104;
  assign n9144 = ~n11105;
  assign n8430 = ~n11106;
  assign n8164 = ~n11107;
  assign n8888 = ~n11108;
  assign n9192 = ~n11109;
  assign n9506 = ~n11110;
  assign n9342 = ~n11111;
  assign n9146 = ~n11112;
  assign n8504 = ~n11115;
  assign n9934 = ~n11116;
  assign n8838 = ~n11117;
  assign n9646 = ~n11118;
  assign n8122 = ~n11119;
  assign n9186 = ~n11120;
  assign n9440 = ~n11121;
  assign n9570 = ~n11122;
  assign n8878 = ~n11123;
  assign n9422 = ~n11124;
  assign n8966 = ~n11125;
  assign n8344 = ~n11126;
  assign n9044 = ~n11127;
  assign n10958 = n11128 & n11129;
  assign n9178 = ~n11130;
  assign n8800 = ~n11131;
  assign n9058 = ~n11132;
  assign n8210 = ~n11133;
  assign n8482 = ~n11134;
  assign n9556 = ~n11135;
  assign n10964 = n11136 & n11137;
  assign n10968 = n11138 & n63;
  assign n9370 = ~n11139;
  assign n8548 = ~n11140;
  assign n9668 = ~n11141;
  assign n8284 = ~n11142;
  assign n9080 = ~n11143;
  assign n9062 = ~n11144;
  assign n8884 = ~n11145;
  assign n8936 = ~n11146;
  assign n9838 = ~n11147;
  assign n9514 = ~n11148;
  assign n8252 = ~n11149;
  assign n8822 = ~n11150;
  assign n8840 = ~n11151;
  assign n9666 = ~n11152;
  assign n8130 = ~n11153;
  assign n9438 = ~n11154;
  assign n8094 = ~n11155;
  assign n10967 = n11156 & n49;
  assign n8008 = ~n11157;
  assign n8982 = ~n11158;
  assign n9098 = ~n11159;
  assign n9806 = ~n11160;
  assign n9184 = ~n11161;
  assign n9180 = ~n11162;
  assign n8572 = ~n11163;
  assign n8624 = ~n11164;
  assign n10995 = n11165 & n11166;
  assign n9002 = ~n11167;
  assign n9644 = ~n11168;
  assign n9614 = ~n11169;
  assign n9078 = ~n11170;
  assign n8338 = ~n11171;
  assign n9892 = ~n11172;
  assign n8422 = ~n11173;
  assign n8510 = ~n11174;
  assign n9018 = ~n11175;
  assign n8984 = ~n11178;
  assign n8416 = ~n11179;
  assign n8184 = ~n11180;
  assign n9520 = ~n11181;
  assign n8756 = ~n11182;
  assign n9540 = ~n11183;
  assign n8714 = ~n11184;
  assign n8318 = ~n11185;
  assign n8634 = ~n11186;
  assign n9736 = ~n11187;
  assign n9660 = ~n11188;
  assign n8642 = ~n11189;
  assign n8810 = ~n11190;
  assign n9068 = ~n11191;
  assign n8162 = ~n11192;
  assign n8042 = ~n11193;
  assign n9456 = ~n11194;
  assign n8490 = ~n11195;
  assign n9546 = ~n11196;
  assign n8198 = ~n11197;
  assign n9236 = ~n11198;
  assign n9920 = ~n11199;
  assign n9372 = ~n11200;
  assign n8852 = ~n11201;
  assign n8828 = ~n11202;
  assign n8972 = ~n11203;
  assign n9896 = ~n11204;
  assign n9010 = ~n11205;
  assign n9444 = ~n11206;
  assign n9300 = ~n11207;
  assign n8976 = ~n11208;
  assign n8402 = ~n11209;
  assign n9174 = ~n11210;
  assign n9828 = ~n11211;
  assign n8512 = ~n11212;
  assign n9526 = ~n11213;
  assign n9844 = ~n11214;
  assign n8148 = ~n11215;
  assign n8304 = ~n11216;
  assign n8594 = ~n11217;
  assign n8560 = ~n11218;
  assign n8248 = ~n11219;
  assign n8282 = ~n11220;
  assign n9722 = ~n11221;
  assign n9864 = ~n11222;
  assign n9326 = ~n11223;
  assign n9286 = ~n11224;
  assign n8072 = ~n11225;
  assign n8696 = ~n11226;
  assign n9904 = ~n11227;
  assign n9022 = ~n11230;
  assign n9602 = ~n11231;
  assign n9492 = ~n11234;
  assign n8376 = ~n11235;
  assign n8342 = ~n11236;
  assign n9388 = ~n11237;
  assign n8736 = ~n11238;
  assign n8120 = ~n11239;
  assign n9136 = ~n11240;
  assign n8516 = ~n11241;
  assign n9744 = ~n11242;
  assign n8458 = ~n11243;
  assign n8076 = ~n11244;
  assign n8812 = ~n11245;
  assign n9402 = ~n11246;
  assign n9108 = ~n11247;
  assign n9268 = ~n11248;
  assign n9780 = ~n11249;
  assign n8916 = ~n11250;
  assign n8160 = ~n11251;
  assign n9544 = ~n11252;
  assign n9028 = ~n11253;
  assign n9430 = ~n11254;
  assign n9294 = ~n11255;
  assign n9620 = ~n11256;
  assign n9416 = ~n11257;
  assign n9760 = ~n11258;
  assign n8226 = ~n11259;
  assign n8686 = ~n11260;
  assign n9880 = ~n11261;
  assign n8424 = ~n11262;
  assign n9380 = ~n11263;
  assign n8078 = ~n11264;
  assign n9152 = ~n11265;
  assign n9410 = ~n11266;
  assign n8214 = ~n11267;
  assign n8086 = ~n11268;
  assign n9138 = ~n11269;
  assign n9932 = ~n11270;
  assign n8462 = ~n11273;
  assign n8978 = ~n11274;
  assign n8636 = ~n11275;
  assign n8054 = ~n11276;
  assign n9656 = ~n11277;
  assign n8530 = ~n11278;
  assign n8240 = ~n11281;
  assign n9454 = ~n11282;
  assign n9338 = ~n11283;
  assign n8374 = ~n11284;
  assign n8328 = ~n11285;
  assign n8762 = ~n11286;
  assign n8546 = ~n11287;
  assign n9822 = ~n11288;
  assign n8970 = ~n11289;
  assign n9056 = ~n11290;
  assign n9304 = ~n11291;
  assign n8398 = ~n11292;
  assign n8790 = ~n11293;
  assign n9198 = ~n11294;
  assign n9730 = ~n11295;
  assign n8744 = ~n11296;
  assign n8218 = ~n11297;
  assign n9412 = ~n11298;
  assign n9494 = ~n11299;
  assign n9848 = ~n11300;
  assign n9332 = ~n11303;
  assign n8386 = ~n11304;
  assign n9890 = ~n11305;
  assign n8826 = ~n11306;
  assign n8690 = ~n11307;
  assign n9598 = ~n11308;
  assign n9306 = ~n11309;
  assign n8208 = ~n11310;
  assign n8154 = ~n11311;
  assign n8876 = ~n11312;
  assign n8844 = ~n11313;
  assign n8680 = ~n11314;
  assign n8740 = ~n11315;
  assign n9752 = ~n11316;
  assign n8656 = ~n11317;
  assign n9280 = ~n11318;
  assign n9360 = ~n11319;
  assign n10991 = n11138 & n11320;
  assign n8944 = ~n11321;
  assign n9020 = ~n11322;
  assign n9084 = ~n11323;
  assign n8320 = ~n11324;
  assign n8772 = ~n11325;
  assign n8898 = ~n11326;
  assign n11014 = n11156 & n11327;
  assign n10955 = n11328 & n11329;
  assign n8288 = ~n11330;
  assign n11013 = n11331 & n11332;
  assign n8348 = ~n11335;
  assign n10947 = n11336 & n11337;
  assign n8394 = ~n11338;
  assign n11001 = n11339 & n11340;
  assign n10946 = n11341 & n11342;
  assign n11012 = n11343 & n11344;
  assign n9408 = ~n11345;
  assign n8486 = ~n11346;
  assign n8492 = ~n11347;
  assign n10987 = n11103 & n45;
  assign n8404 = ~n11348;
  assign n9816 = ~n11349;
  assign n8564 = ~n11350;
  assign n9308 = ~n11351;
  assign n8998 = ~n11352;
  assign n8346 = ~n11353;
  assign n8262 = ~n11354;
  assign n9794 = ~n11355;
  assign n9810 = ~n11356;
  assign n8644 = ~n11357;
  assign n8286 = ~n11358;
  assign n8568 = ~n11359;
  assign n8508 = ~n11360;
  assign n9228 = ~n11361;
  assign n9552 = ~n11362;
  assign n9382 = ~n11363;
  assign n9586 = ~n11364;
  assign n8298 = ~n11365;
  assign n9710 = ~n11366;
  assign n8802 = ~n11367;
  assign n9624 = ~n11368;
  assign n9076 = ~n11369;
  assign n8500 = ~n11370;
  assign n8432 = ~n11371;
  assign n9640 = ~n11372;
  assign n9072 = ~n11373;
  assign n9906 = ~n11374;
  assign n9214 = ~n11375;
  assign n8554 = ~n11376;
  assign n8750 = ~n11377;
  assign n8694 = ~n11378;
  assign n9290 = ~n11379;
  assign n9014 = ~n11380;
  assign n8506 = ~n11381;
  assign n9832 = ~n11382;
  assign n8052 = ~n11383;
  assign n9912 = ~n11384;
  assign n9158 = ~n11387;
  assign n8046 = ~n11388;
  assign n8688 = ~n11389;
  assign n9424 = ~n11390;
  assign n9176 = ~n11391;
  assign n8080 = ~n11392;
  assign n8542 = ~n11393;
  assign n8912 = ~n11394;
  assign n9588 = ~n11395;
  assign n8088 = ~n11396;
  assign n9200 = ~n11397;
  assign n9522 = ~n11398;
  assign n9719 = ~n11399;
  assign n9066 = ~n11400;
  assign n9168 = ~n11401;
  assign n8534 = ~n11402;
  assign n8712 = ~n11403;
  assign n9368 = ~n11404;
  assign n8020 = ~n11405;
  assign n8022 = ~n11406;
  assign n8666 = ~n11407;
  assign n9384 = ~n11408;
  assign n8332 = ~n11409;
  assign n8792 = ~n11410;
  assign n8062 = ~n11411;
  assign n9448 = ~n11412;
  assign n9378 = ~n11413;
  assign n9568 = ~n11414;
  assign n9762 = ~n11415;
  assign n9040 = ~n11416;
  assign n8396 = ~n11417;
  assign n9572 = ~n11418;
  assign n9530 = ~n11419;
  assign n8232 = ~n11420;
  assign n9130 = ~n11421;
  assign n9536 = ~n11422;
  assign n8384 = ~n11423;
  assign n8428 = ~n11424;
  assign n8370 = ~n11425;
  assign n8360 = ~n11426;
  assign n8954 = ~n11429;
  assign n8846 = ~n11432;
  assign n9490 = ~n11433;
  assign n9182 = ~n11434;
  assign n8056 = ~n11435;
  assign n9566 = ~n11436;
  assign n8266 = ~n11437;
  assign n8782 = ~n11440;
  assign n9204 = ~n11441;
  assign n9914 = ~n11442;
  assign n9114 = ~n11443;
  assign n8068 = ~n11444;
  assign n8206 = ~n11445;
  assign n8116 = ~n11446;
  assign n8532 = ~n11447;
  assign n8246 = ~n11448;
  assign n8748 = ~n11449;
  assign n8892 = ~n11450;
  assign n8420 = ~n11451;
  assign n9594 = ~n11452;
  assign n8774 = ~n11453;
  assign n8468 = ~n11454;
  assign n9212 = ~n11455;
  assign n8118 = ~n11456;
  assign n8950 = ~n11457;
  assign n8896 = ~n11458;
  assign n9270 = ~n11459;
  assign n9434 = ~n11460;
  assign n8454 = ~n11461;
  assign n9034 = ~n11462;
  assign n9662 = ~n11463;
  assign n10976 = n11339 & n47;
  assign n9574 = ~n11464;
  assign n8222 = ~n11465;
  assign n8692 = ~n11466;
  assign n8356 = ~n11467;
  assign n8408 = ~n11468;
  assign n8734 = ~n11469;
  assign n8778 = ~n11470;
  assign n9202 = ~n11471;
  assign n9486 = ~n11472;
  assign n8280 = ~n11473;
  assign n8698 = ~n11474;
  assign n8658 = ~n11475;
  assign n9748 = ~n11476;
  assign n9466 = ~n11477;
  assign n9788 = ~n11478;
  assign n8250 = ~n11479;
  assign n9782 = ~n11480;
  assign n8890 = ~n11481;
  assign n8292 = ~n11482;
  assign n8260 = ~n11483;
  assign n8496 = ~n11484;
  assign n9148 = ~n11485;
  assign n10978 = n11343 & n55;
  assign n9278 = ~n11486;
  assign n9112 = ~n11487;
  assign n8866 = ~n11488;
  assign n8710 = ~n11489;
  assign n9714 = ~n11490;
  assign n9862 = ~n11491;
  assign n9724 = ~n11492;
  assign n9582 = ~n11493;
  assign n8930 = ~n11494;
  assign n8932 = ~n11495;
  assign n9774 = ~n11496;
  assign n9260 = ~n11497;
  assign n8064 = ~n11498;
  assign n9842 = ~n11499;
  assign n8578 = ~n11500;
  assign n9504 = ~n11501;
  assign n9580 = ~n11502;
  assign n9094 = ~n11503;
  assign n8036 = ~n11504;
  assign n9778 = ~n11505;
  assign n9502 = ~n11506;
  assign n8798 = ~n11507;
  assign n8582 = ~n11508;
  assign n8788 = ~n11509;
  assign n9652 = ~n11510;
  assign n9396 = ~n11511;
  assign n9248 = ~n11512;
  assign n8662 = ~n11513;
  assign n8716 = ~n11514;
  assign n8770 = ~n11515;
  assign n8256 = ~n11516;
  assign n8682 = ~n11517;
  assign n8324 = ~n11518;
  assign n9222 = ~n11519;
  assign n8040 = ~n11520;
  assign n9142 = ~n11521;
  assign n8732 = ~n11522;
  assign n9244 = ~n11523;
  assign n9528 = ~n11524;
  assign n8388 = ~n11525;
  assign n9622 = ~n11526;
  assign n9804 = ~n11527;
  assign n8850 = ~n11528;
  assign n8938 = ~n11529;
  assign n9756 = ~n11530;
  assign n9638 = ~n11531;
  assign n9190 = ~n11532;
  assign n9654 = ~n11533;
  assign n8924 = ~n11534;
  assign n9016 = ~n11535;
  assign n8814 = ~n11536;
  assign n8908 = ~n11537;
  assign n8540 = ~n11538;
  assign n8098 = ~n11539;
  assign n8586 = ~n11540;
  assign n8928 = ~n11541;
  assign n8768 = ~n11542;
  assign n8378 = ~n11543;
  assign n8494 = ~n11544;
  assign n8470 = ~n11545;
  assign n8176 = ~n11546;
  assign n8676 = ~n11547;
  assign n9472 = ~n11548;
  assign n8558 = ~n11549;
  assign n8182 = ~n11550;
  assign n9330 = ~n11551;
  assign n9446 = ~n11552;
  assign n8618 = ~n11553;
  assign n8964 = ~n11554;
  assign n8574 = ~n11555;
  assign n8728 = ~n11556;
  assign n8988 = ~n11557;
  assign n9052 = ~n11558;
  assign n8628 = ~n11559;
  assign n9576 = ~n11560;
  assign n9420 = ~n11561;
  assign n8592 = ~n11562;
  assign n8446 = ~n11563;
  assign n9354 = ~n11564;
  assign n9166 = ~n11565;
  assign n9784 = ~n11566;
  assign n9860 = ~n11567;
  assign n8476 = ~n11568;
  assign n8704 = ~n11569;
  assign n8060 = ~n11570;
  assign n8110 = ~n11571;
  assign n9432 = ~n11572;
  assign n9856 = ~n11573;
  assign n9134 = ~n11574;
  assign n8242 = ~n11575;
  assign n9808 = ~n11576;
  assign n10975 = n11136 & n39;
  assign n8946 = ~n11577;
  assign n9866 = ~n11578;
  assign n9814 = ~n11579;
  assign n9632 = ~n11580;
  assign n8808 = ~n11581;
  assign n9534 = ~n11582;
  assign n9878 = ~n11583;
  assign n9048 = ~n11584;
  assign n8034 = ~n11585;
  assign n8904 = ~n11586;
  assign n9812 = ~n11587;
  assign n8596 = ~n11588;
  assign n8448 = ~n11589;
  assign n8460 = ~n11590;
  assign n9802 = ~n11591;
  assign n11002 = n11592 & n11593;
  assign n9406 = ~n11594;
  assign n8836 = ~n11595;
  assign n8268 = ~n11596;
  assign n9096 = ~n11597;
  assign n8058 = ~n11598;
  assign n9612 = ~n11599;
  assign n8312 = ~n11600;
  assign n9746 = ~n11601;
  assign n8474 = ~n11602;
  assign n8664 = ~n11603;
  assign n8352 = ~n11604;
  assign n8438 = ~n11605;
  assign n8742 = ~n11606;
  assign n8296 = ~n11607;
  assign n8974 = ~n11608;
  assign n9374 = ~n11609;
  assign n9876 = ~n11610;
  assign n9086 = ~n11611;
  assign n9800 = ~n11612;
  assign n9242 = ~n11613;
  assign n8440 = ~n11614;
  assign n8870 = ~n11615;
  assign n8544 = ~n11616;
  assign n9852 = ~n11617;
  assign n8858 = ~n11618;
  assign n8238 = ~n11619;
  assign n9436 = ~n11620;
  assign n9288 = ~n11621;
  assign n9840 = ~n11622;
  assign n8090 = ~n11623;
  assign n9462 = ~n11624;
  assign n10980 = n11336 & n51;
  assign n8216 = ~n11625;
  assign n9350 = ~n11626;
  assign n9314 = ~n11627;
  assign n9036 = ~n11630;
  assign n9634 = ~n11631;
  assign n8150 = ~n11632;
  assign n8400 = ~n11633;
  assign n9728 = ~n11634;
  assign n8722 = ~n11635;
  assign n8856 = ~n11636;
  assign n9364 = ~n11637;
  assign n9070 = ~n11638;
  assign n8958 = ~n11639;
  assign n8832 = ~n11640;
  assign n8910 = ~n11641;
  assign n9334 = ~n11642;
  assign n9194 = ~n11645;
  assign n8622 = ~n11646;
  assign n8274 = ~n11647;
  assign n8872 = ~n11648;
  assign n10993 = n11341 & n35;
  assign n8882 = ~n11649;
  assign n8254 = ~n11650;
  assign n8302 = ~n11653;
  assign n8990 = ~n11654;
  assign n10948 = n11328 & n37;
  assign n8426 = ~n11655;
  assign n9132 = ~n11658;
  assign n8514 = ~n11659;
  assign n9250 = ~n11660;
  assign n9090 = ~n11661;
  assign n9608 = ~n11662;
  assign n9922 = ~n11663;
  assign n8230 = ~n11664;
  assign n9442 = ~n11665;
  assign n9488 = ~n11666;
  assign n8922 = ~n11667;
  assign n9772 = ~n11668;
  assign n8766 = ~n11669;
  assign n9282 = ~n11670;
  assign n8436 = ~n11671;
  assign n9336 = ~n11672;
  assign n9584 = ~n11673;
  assign n8234 = ~n11674;
  assign n9790 = ~n11675;
  assign n9296 = ~n11676;
  assign n8316 = ~n11677;
  assign n8134 = ~n11678;
  assign n8012 = ~n11679;
  assign n8202 = ~n11680;
  assign n9758 = ~n11681;
  assign n9512 = ~n11682;
  assign n9510 = ~n11683;
  assign n9106 = ~n11684;
  assign n8906 = ~n11685;
  assign n8372 = ~n11686;
  assign n9630 = ~n11687;
  assign n9358 = ~n11688;
  assign n8940 = ~n11689;
  assign n9392 = ~n11690;
  assign n9160 = ~n11693;
  assign n8026 = ~n11694;
  assign n8520 = ~n11695;
  assign n9140 = ~n11696;
  assign n9226 = ~n11697;
  assign n8412 = ~n11698;
  assign n9592 = ~n11699;
  assign n8264 = ~n11700;
  assign n8684 = ~n11701;
  assign n8044 = ~n11702;
  assign n8994 = ~n11703;
  assign n8126 = ~n11704;
  assign n8702 = ~n11705;
  assign n8552 = ~n11706;
  assign n8172 = ~n11707;
  assign n9518 = ~n11708;
  assign n9928 = ~n11709;
  assign n8502 = ~n11710;
  assign n8724 = ~n11711;
  assign n9894 = ~n11712;
  assign n8806 = ~n11715;
  assign n9846 = ~n11716;
  assign n8410 = ~n11717;
  assign n8480 = ~n11718;
  assign n8192 = ~n11719;
  assign n9542 = ~n11720;
  assign n8186 = ~n11721;
  assign n9196 = ~n11722;
  assign n8178 = ~n11723;
  assign n9650 = ~n11724;
  assign n8632 = ~n11725;
  assign n8392 = ~n11726;
  assign n8136 = ~n11727;
  assign n8674 = ~n11728;
  assign n9776 = ~n11729;
  assign n9550 = ~n11730;
  assign n9648 = ~n11731;
  assign n9032 = ~n11732;
  assign n8050 = ~n11733;
  assign n8340 = ~n11734;
  assign n8066 = ~n11735;
  assign n8326 = ~n11736;
  assign n8830 = ~n11737;
  assign n10986 = n11738 & n11739;
  assign n8142 = ~n11740;
  assign n9450 = ~n11741;
  assign n9102 = ~n11742;
  assign n8926 = ~n11743;
  assign n9006 = ~n11744;
  assign n8082 = ~n11745;
  assign n9768 = ~n11746;
  assign n8900 = ~n11747;
  assign n9764 = ~n11748;
  assign n9664 = ~n11749;
  assign n8010 = ~n11750;
  assign n8114 = ~n11751;
  assign n9524 = ~n11752;
  assign n9272 = ~n11753;
  assign n9322 = ~n11754;
  assign n8364 = ~n11755;
  assign n9232 = ~n11756;
  assign n9042 = ~n11757;
  assign n8804 = ~n11758;
  assign n9578 = ~n11759;
  assign n8048 = ~n11760;
  assign n8358 = ~n11761;
  assign n8918 = ~n11762;
  assign n10956 = n11592 & n57;
  assign n8824 = ~n11763;
  assign n9124 = ~n11764;
  assign n8630 = ~n11765;
  assign n9154 = ~n11766;
  assign n9082 = ~n11767;
  assign n9292 = ~n11768;
  assign n8784 = ~n11769;
  assign n8886 = ~n11770;
  assign n8818 = ~n11771;
  assign n9100 = ~n11772;
  assign n8224 = ~n11773;
  assign n9900 = ~n11774;
  assign n9858 = ~n11775;
  assign n8190 = ~n11776;
  assign n8466 = ~n11777;
  assign n8638 = ~n11778;
  assign n9884 = ~n11779;
  assign n8488 = ~n11780;
  assign n9376 = ~n11781;
  assign n8362 = ~n11782;
  assign n9390 = ~n11783;
  assign n9302 = ~n11784;
  assign n9264 = ~n11785;
  assign n9590 = ~n11786;
  assign n8158 = ~n11787;
  assign n8914 = ~n11788;
  assign n9046 = ~n11789;
  assign n8786 = ~n11790;
  assign n9712 = ~n11791;
  assign n10970 = n11165 & n43;
  assign n9740 = ~n11792;
  assign n8956 = ~n11793;
  assign n8128 = ~n11794;
  assign n8484 = ~n11795;
  assign n8140 = ~n11796;
  assign n9118 = ~n11797;
  assign n8272 = ~n11798;
  assign n8290 = ~n11799;
  assign n9150 = ~n11800;
  assign n8102 = ~n11801;
  assign n9458 = ~n11802;
  assign n8556 = ~n11803;
  assign n8700 = ~n11804;
  assign n8294 = ~n11805;
  assign n9246 = ~n11806;
  assign n8590 = ~n11809;
  assign n8754 = ~n11810;
  assign n9508 = ~n11811;
  assign n8478 = ~n11812;
  assign n9726 = ~n11813;
  assign n8760 = ~n11814;
  assign n9792 = ~n11815;
  assign n8842 = ~n11816;
  assign n9604 = ~n11817;
  assign n8708 = ~n11818;
  assign n8096 = ~n11819;
  assign n9468 = ~n11820;
  assign n9754 = ~n11821;
  assign n8074 = ~n11822;
  assign n8650 = ~n11823;
  assign n9606 = ~n11824;
  assign n8168 = ~n11825;
  assign n8854 = ~n11826;
  assign n8354 = ~n11827;
  assign n8180 = ~n11828;
  assign n9868 = ~n11829;
  assign n8196 = ~n11830;
  assign n8382 = ~n11831;
  assign n8608 = ~n11832;
  assign n8550 = ~n11833;
  assign n9216 = ~n11834;
  assign n9210 = ~n11835;
  assign n8730 = ~n11836;
  assign n9538 = ~n11837;
  assign n8780 = ~n11838;
  assign n9274 = ~n11839;
  assign n9012 = ~n11840;
  assign n9262 = ~n11841;
  assign n8874 = ~n11842;
  assign n8820 = ~n11843;
  assign n9126 = ~n11844;
  assign n8758 = ~n11845;
  assign n9818 = ~n11846;
  assign n9394 = ~n11847;
  assign n9328 = ~n11848;
  assign n9924 = ~n11849;
  assign n8992 = ~n11850;
  assign n9554 = ~n11851;
  assign n9836 = ~n11852;
  assign n8894 = ~n11853;
  assign n9548 = ~n11854;
  assign n8980 = ~n11855;
  assign n8084 = ~n11856;
  assign n9564 = ~n11857;
  assign n8418 = ~n11858;
  assign n9824 = ~n11859;
  assign n8670 = ~n11860;
  assign n9474 = ~n11861;
  assign n8968 = ~n11862;
  assign n8368 = ~n11863;
  assign n9930 = ~n11864;
  assign n9346 = ~n11867;
  assign n8752 = ~n11868;
  assign n8028 = ~n11869;
  assign n8276 = ~n11870;
  assign n8310 = ~n11871;
  assign n9886 = ~n11872;
  assign n8132 = ~n11873;
  assign n9208 = ~n11874;
  assign n8660 = ~n11875;
  assign n8450 = ~n11876;
  assign n9898 = ~n11877;
  assign n8706 = ~n11878;
  assign n9476 = ~n11879;
  assign n8536 = ~n11880;
  assign n8390 = ~n11881;
  assign n9480 = ~n11882;
  assign n9284 = ~n11883;
  assign n8212 = ~n11884;
  assign n8720 = ~n11885;
  assign n9122 = ~n11886;
  assign n9830 = ~n11887;
  assign n8228 = ~n11888;
  assign n10960 = n11889 & n61;
  assign n9478 = ~n11890;
  assign n8566 = ~n11891;
  assign n8794 = ~n11892;
  assign n9310 = ~n11893;
  assign n9258 = ~n11894;
  assign n9464 = ~n11895;
  assign n9164 = ~n11896;
  assign n8562 = ~n11897;
  assign n10998 = n11889 & n11898;
  assign n8816 = ~n11899;
  assign n8442 = ~n11900;
  assign n8952 = ~n11901;
  assign n8018 = ~n11902;
  assign n9234 = ~n11903;
  assign n9220 = ~n11904;
  assign n9750 = ~n11905;
  assign n8138 = ~n11906;
  assign n9218 = ~n11907;
  assign n9000 = ~n11908;
  assign n9693 = ~n11909;
  assign n8336 = ~n11910;
  assign n9596 = ~n11911;
  assign n10951 = n11738 & n53;
  assign n9938 = ~n11912;
  assign n9074 = ~n11913;
  assign n8606 = ~n11914;
  assign n8580 = ~n11915;
  assign n9414 = ~n11918;
  assign n9004 = ~n11919;
  assign n9054 = ~n11922;
  assign n9626 = ~n11927;
  assign n8528 = ~n11936;
  assign n9240 = ~n11937;
  assign n9060 = ~n11938;
  assign n9658 = ~n11939;
  assign n8598 = ~n11940;
  assign n8902 = ~n11941;
  assign n9366 = ~n11942;
  assign n9266 = ~n11943;
  assign n10953 = n11128 & n41;
  assign n9820 = ~n11944;
  assign n8244 = ~n11945;
  assign n9156 = ~n11946;
  assign n9224 = ~n11947;
  assign n8366 = ~n11948;
  assign n9826 = ~n11949;
  assign n9766 = ~n11950;
  assign n9902 = ~n11951;
  assign n8860 = ~n11952;
  assign n8576 = ~n11953;
  assign n9742 = ~n11954;
  assign n8626 = ~n11955;
  assign n9498 = ~n11956;
  assign n8570 = ~n11957;
  assign n8124 = ~n11958;
  assign n9734 = ~n11959;
  assign n8156 = ~n11960;
  assign n9452 = ~n11961;
  assign n8032 = ~n11962;
  assign n9344 = ~n11963;
  assign n8472 = ~n11964;
  assign n9872 = ~n11965;
  assign n8864 = ~n11966;
  assign n9516 = ~n11967;
  assign n9356 = ~n11968;
  assign n9404 = ~n11969;
  assign n8038 = ~n11970;
  assign n9252 = ~n11971;
  assign n9024 = ~n11972;
  assign n9256 = ~n11973;
  assign n8602 = ~n11974;
  assign n8640 = ~n11975;
  assign n8414 = ~n11976;
  assign n8434 = ~n11977;
  assign n9030 = ~n11978;
  assign n8584 = ~n11979;
  assign n9120 = ~n11980;
  assign n9882 = ~n11981;
  assign n8306 = ~n11984;
  assign n8406 = ~n11985;
  assign n9418 = ~n11986;
  assign n8518 = ~n11987;
  assign n8380 = ~n11988;
  assign n9910 = ~n11989;
  assign n9320 = ~n11990;
  assign n9532 = ~n11991;
  assign n9116 = ~n11992;
  assign n8270 = ~n11993;
  assign n9636 = ~n11994;
  assign n9340 = ~n11995;
  assign n8146 = ~n11996;
  assign n9642 = ~n11997;
  assign n9316 = ~n11998;
  assign n9254 = ~n11999;
  assign n9026 = ~n12000;
  assign n8070 = ~n12001;
  assign n8738 = ~n12002;
  assign n9460 = ~n12003;
  assign n8834 = ~n12004;
  assign n8200 = ~n12005;
  assign n8278 = ~n12006;
  assign n9400 = ~n12007;
  assign n10950 = n11331 & n59;
  assign n8616 = ~n12008;
  assign n8610 = ~n12009;
  assign n8350 = ~n12010;
  assign n8498 = ~n12011;
  assign n9496 = ~n12012;
  assign n8718 = ~n12013;
  assign n9038 = ~n12014;
  assign n8220 = ~n12015;
  assign n8604 = ~n12016;
  assign n8092 = ~n12017;
  assign n8862 = ~n12018;
  assign n8934 = ~n12019;
  assign n8648 = ~n12020;
  assign n8880 = ~n12021;
  assign n9936 = ~n12022;
  assign n8996 = ~n12023;
  assign n9008 = ~n12024;
  assign n8016 = ~n12025;
  assign n9092 = ~n12026;
  assign n9170 = ~n12027;
  assign n9362 = ~n12028;
  assign n8300 = ~n12029;
  assign n8652 = ~n12030;
  assign n8464 = ~n12031;
  assign n8960 = ~n12032;
  assign n8764 = ~n12033;
  assign n8174 = ~n12034;
  assign n9172 = ~n12035;
  assign n8668 = ~n12036;
  assign n9088 = ~n12037;
  assign n9470 = ~n12038;
  assign n9850 = ~n12039;
  assign n8522 = ~n12040;
  assign n9738 = ~n12041;
  assign n8678 = ~n12042;
  assign n8104 = ~n12043;
  assign n9500 = ~n12044;
  assign n9398 = ~n12045;
  assign n8776 = ~n12046;
  assign n9870 = ~n12047;
  assign n9558 = ~n12048;
  assign n9918 = ~n12049;
  assign n8014 = ~n12050;
  assign n8654 = ~n12051;
  assign n9600 = ~n12052;
  assign n9770 = ~n12053;
  assign n9318 = ~n12054;
  assign n8646 = ~n12055;
  assign n8672 = ~n12056;
  assign n9238 = ~n12057;
  assign n9206 = ~n12060;
  assign n9908 = ~n12061;
  assign n9128 = ~n12062;
  assign n8942 = ~n12063;
  assign n8152 = ~n12064;
  assign n9298 = ~n12065;
  assign n8108 = ~n12066;
  assign n8848 = ~n12067;
  assign n8796 = ~n12068;
  assign n8144 = ~n12069;
  assign n9834 = ~n12070;
  assign n9786 = ~n12071;
  assign n9796 = ~n12072;
  assign n9050 = ~n12073;
  assign n8620 = ~n12074;
  assign n8456 = ~n12075;
  assign n8030 = ~n12076;
  assign n9616 = ~n12077;
  assign n9230 = ~n12078;
  assign n9732 = ~n12079;
  assign n9874 = ~n12080;
  assign n9428 = ~n12081;
  assign n8166 = ~n12082;
  assign n9560 = ~n12083;
  assign n8170 = ~n12084;
  assign n9562 = ~n12085;
  assign n9610 = ~n12086;
  assign n8330 = ~n12087;
  assign n8612 = ~n12088;
  assign n9926 = ~n12089;
  assign n8314 = ~n12090;
  assign n9618 = ~n12091;
  assign n8588 = ~n12092;
  assign n9484 = ~n12093;
  assign n8614 = ~n12094;
  assign n8948 = ~n12095;
  assign n8204 = ~n12096;
  assign n8100 = ~n12097;
  assign n9798 = ~n12098;
  assign n9386 = ~n12099;
  assign n8538 = ~n12100;
  assign n9324 = ~n12103;
  assign n8188 = ~n12104;
  assign n8726 = ~n12105;
  assign n8868 = ~n12106;
  assign n9888 = ~n12109;
  assign n9854 = ~n12110;
  assign n8024 = ~n12111;
  assign n9426 = ~n12112;
  assign n9162 = ~n12113;
  assign n8194 = ~n12114;
  assign n8308 = ~n12115;
  assign n8746 = ~n12116;
  assign n9104 = ~n12117;
  assign n8334 = ~n12118;
  assign n9482 = ~n12119;
  assign n8962 = ~n12120;
  assign n8322 = ~n12121;
  assign n8524 = ~n12122;
  assign n8444 = ~n12123;
  assign n9276 = ~n12124;
  assign n8986 = ~n12125;
  assign n11080 = ~n11138;
  assign n11020 = ~n12171;
  assign n11058 = ~n12172;
  assign n11011 = ~n12173;
  assign n11271 = ~n12174;
  assign n11009 = ~n12177;
  assign n11052 = ~n12178;
  assign n12141 = n12179 & n61;
  assign n12107 = ~n12180;
  assign n11865 = ~n12181;
  assign n12162 = n12182 & n57;
  assign n11430 = ~n12183;
  assign n11232 = ~n12184;
  assign n10985 = ~n12185;
  assign n11067 = ~n12186;
  assign n11301 = ~n12187;
  assign n11982 = ~n12188;
  assign n11643 = ~n12189;
  assign n11022 = ~n12190;
  assign n11807 = ~n12191;
  assign n11930 = ~n12193;
  assign n11934 = ~n12194;
  assign n11691 = ~n12195;
  assign n11026 = ~n12196;
  assign n10983 = ~n12197;
  assign n11628 = ~n12198;
  assign n12135 = n12203 & n39;
  assign n12168 = n12206 & n33;
  assign n12165 = n12207 & n37;
  assign n11024 = ~n12208;
  assign n11062 = ~n12209;
  assign n11056 = ~n12210;
  assign n11016 = ~n12211;
  assign n11034 = ~n12212;
  assign n11018 = ~n12215;
  assign n11656 = ~n12216;
  assign n12058 = ~n12217;
  assign n11333 = ~n12218;
  assign n11438 = ~n12219;
  assign n11054 = ~n12220;
  assign n12132 = n12221 & n59;
  assign n12160 = n12226 & n51;
  assign n11046 = ~n12227;
  assign n12161 = n12230 & n43;
  assign n12164 = n12231 & n55;
  assign n11032 = ~n12232;
  assign n11048 = ~n12233;
  assign n11050 = ~n12234;
  assign n12159 = n12235 & n53;
  assign n11651 = ~n12236;
  assign n11928 = ~n12239;
  assign n11038 = ~n12240;
  assign n11923 = ~n12241;
  assign n11064 = ~n12242;
  assign n11069 = ~n12243;
  assign n11925 = ~n12244;
  assign n12166 = n12245 & n49;
  assign n12167 = n12246 & n41;
  assign n11028 = ~n12247;
  assign n11040 = ~n12248;
  assign n11713 = ~n12249;
  assign n12170 = n12250 & n47;
  assign n11036 = ~n12251;
  assign n11279 = ~n12252;
  assign n11113 = ~n12255;
  assign n11044 = ~n12256;
  assign n11176 = ~n12259;
  assign n11228 = ~n12262;
  assign n11030 = ~n12263;
  assign n11932 = ~n12264;
  assign n11385 = ~n12265;
  assign n12163 = n12266 & n35;
  assign n12101 = ~n12267;
  assign n11042 = ~n12268;
  assign n11427 = ~n12269;
  assign n12169 = n12272 & n45;
  assign n11916 = ~n12273;
  assign n11920 = ~n12274;
  assign n11060 = ~n12277;
  assign n10507 = n10946 & n2;
  assign n10469 = n10947 & n10;
  assign n10334 = n10948 & n10949;
  assign n10410 = n10950 & n9939;
  assign n10361 = n10951 & n10952;
  assign n10405 = n10953 & n10954;
  assign n10862 = n10955 & n16;
  assign n10117 = n10956 & n10957;
  assign n10511 = n10958 & n22;
  assign n10509 = n10947 & n13;
  assign n10699 = n10958 & n2;
  assign n10860 = n10947 & n30;
  assign n10404 = n10948 & n10959;
  assign n10399 = n10960 & n10961;
  assign n10401 = n10953 & n10962;
  assign n10261 = n10953 & n10963;
  assign n10260 = n10950 & n10959;
  assign n10595 = n10964 & n11;
  assign n10508 = n10955 & n9;
  assign n10400 = n10950 & n10965;
  assign n10396 = n10951 & n10954;
  assign n10398 = n10950 & n10966;
  assign n10259 = n10967 & n10952;
  assign n10257 = n10968 & n10969;
  assign n10258 = n10970 & n10971;
  assign n10678 = n10964 & n19;
  assign n10254 = n10968 & n10972;
  assign n10393 = n10956 & n10973;
  assign n10247 = n10956 & n10974;
  assign n10255 = n10975 & n10971;
  assign n10394 = n10976 & n10977;
  assign n10253 = n10978 & n10979;
  assign n10252 = n10968 & n10952;
  assign n10390 = n10980 & n10974;
  assign n10251 = n10967 & n10981;
  assign n10249 = n10980 & n10963;
  assign n10388 = n10968 & n10963;
  assign n10387 = n10970 & n10981;
  assign n10350 = n10951 & n10949;
  assign n10385 = n10968 & n10979;
  assign n10606 = n10986 & n22;
  assign n10246 = n10970 & n10949;
  assign n10245 = n10970 & n10973;
  assign n10383 = n10948 & n10969;
  assign n10242 = n10987 & n10952;
  assign n10380 = n10960 & n10988;
  assign n10501 = n10986 & n0;
  assign n10243 = n10975 & n10954;
  assign n10706 = n10946 & n22;
  assign n10591 = n10964 & n20;
  assign n10239 = n10968 & n10962;
  assign n10241 = n10951 & n10989;
  assign n10378 = n10967 & n10957;
  assign n10374 = n10950 & n10971;
  assign n10377 = n10950 & n10979;
  assign n10375 = n10975 & n10990;
  assign n10493 = n10946 & n31;
  assign n10750 = n10991 & n24;
  assign n10372 = n10948 & n10954;
  assign n10370 = n10976 & n10992;
  assign n10369 = n10953 & n10990;
  assign n10365 = n10968 & n10977;
  assign n10367 = n10956 & n10977;
  assign n10368 = n10993 & n10994;
  assign n10871 = n10995 & n5;
  assign n10024 = n10956 & n10969;
  assign n10366 = n10976 & n10954;
  assign n10492 = n10955 & n0;
  assign n10364 = n10950 & n10996;
  assign n10204 = n10951 & n10963;
  assign n10363 = n10987 & n10997;
  assign n9960 = n10975 & n10994;
  assign n10362 = n10980 & n10952;
  assign n10705 = n10964 & n9;
  assign n10470 = n10995 & n22;
  assign n10830 = n10998 & n20;
  assign n10357 = n10948 & n10971;
  assign n10359 = n10976 & n10988;
  assign n10360 = n10978 & n10966;
  assign n10583 = n10998 & n13;
  assign n10389 = n10951 & n10999;
  assign n10582 = n10946 & n0;
  assign n10843 = n10946 & n12;
  assign n9961 = n10995 & n18;
  assign n10581 = n10955 & n24;
  assign n10578 = n10964 & n16;
  assign n10240 = n10980 & n10989;
  assign n10486 = n10998 & n5;
  assign n10352 = n10956 & n11000;
  assign n10686 = n11001 & n11;
  assign n10902 = n10946 & n25;
  assign n10483 = n11002 & n11;
  assign n10225 = n10987 & n10963;
  assign n10348 = n10987 & n10979;
  assign n10795 = n10998 & n9;
  assign n10238 = n10987 & n10988;
  assign n10237 = n10967 & n10971;
  assign n10235 = n10950 & n10963;
  assign n10233 = n10987 & n10990;
  assign n10343 = n10951 & n10959;
  assign n10234 = n10967 & n10992;
  assign n10231 = n10978 & n10981;
  assign n10347 = n10967 & n11003;
  assign n10477 = n10964 & n5;
  assign n10761 = n10995 & n2;
  assign n10230 = n10993 & n10957;
  assign n10226 = n10980 & n10997;
  assign n9962 = n10998 & n7;
  assign n10222 = n10980 & n10969;
  assign n10224 = n10968 & n11004;
  assign n10339 = n10968 & n10996;
  assign n10471 = n10991 & n21;
  assign n10223 = n10960 & n10972;
  assign n10221 = n10951 & n10977;
  assign n10336 = n10993 & n10961;
  assign n10220 = n10970 & n10997;
  assign n10219 = n10987 & n10992;
  assign n10340 = n10967 & n11005;
  assign n10472 = n11006 & n2;
  assign n10018 = n10960 & n10992;
  assign n9966 = n10964 & n22;
  assign n10703 = n11006 & n11;
  assign n10021 = n10967 & n10990;
  assign n10425 = n10975 & n11007;
  assign n10485 = n11001 & n29;
  assign n10356 = n10967 & n10994;
  assign n10016 = n10968 & n10973;
  assign n10291 = n10993 & n11005;
  assign n9952 = n10986 & n29;
  assign n10579 = n10986 & n8;
  assign n10337 = n10960 & n10962;
  assign n10338 = n10948 & n10992;
  assign n10019 = n10976 & n10996;
  assign n10087 = n10960 & n10997;
  assign n10482 = n10955 & n2;
  assign n10845 = n10995 & n8;
  assign n10857 = n10947 & n6;
  assign n10011 = n10980 & n10988;
  assign n10332 = n10976 & n11000;
  assign n10711 = n10991 & n7;
  assign n10510 = n11001 & n4;
  assign n10333 = n10953 & n10957;
  assign n10759 = n10995 & n14;
  assign n10700 = n10986 & n21;
  assign n10466 = n11006 & n8;
  assign n10012 = n10960 & n10963;
  assign n10467 = n11012 & n3;
  assign n10358 = n10980 & n11005;
  assign n10008 = n10987 & n10994;
  assign n10774 = n11001 & n8;
  assign n10152 = n10953 & n10988;
  assign n10574 = n11012 & n0;
  assign n10696 = n11013 & n18;
  assign n10020 = n10960 & n10999;
  assign n10858 = n11014 & n25;
  assign n10694 = n10955 & n11;
  assign n10602 = n10998 & n23;
  assign n10476 = n10958 & n25;
  assign n10524 = n10991 & n8;
  assign n10473 = n11013 & n29;
  assign n10603 = n10991 & n4;
  assign n9974 = n10968 & n10954;
  assign n9978 = n10978 & n10961;
  assign n9980 = n10975 & n10952;
  assign n9982 = n10950 & n10952;
  assign n9983 = n10948 & n10979;
  assign n9985 = n10951 & n10996;
  assign n9996 = n10978 & n10994;
  assign n9988 = n10948 & n10972;
  assign n9990 = n10980 & n10996;
  assign n10847 = n10991 & n14;
  assign n9993 = n10953 & n10965;
  assign n9995 = n10978 & n10999;
  assign n10000 = n10967 & n10972;
  assign n9998 = n10953 & n10981;
  assign n9999 = n10956 & n11003;
  assign n10001 = n10976 & n10949;
  assign n10002 = n10993 & n10992;
  assign n10114 = n10975 & n10961;
  assign n10487 = n10995 & n15;
  assign n10855 = n11006 & n6;
  assign n10010 = n10956 & n10996;
  assign n10013 = n10993 & n10990;
  assign n10014 = n10948 & n11004;
  assign n10022 = n10956 & n10954;
  assign n10846 = n11014 & n4;
  assign n10015 = n10950 & n10961;
  assign n10027 = n10975 & n11000;
  assign n10033 = n10960 & n10981;
  assign n10034 = n10980 & n10994;
  assign n9997 = n10950 & n10957;
  assign n10040 = n10976 & n10973;
  assign n10575 = n11013 & n13;
  assign n9991 = n10953 & n10952;
  assign n10045 = n10960 & n10979;
  assign n10046 = n10987 & n10972;
  assign n10048 = n10968 & n10974;
  assign n10049 = n10968 & n10990;
  assign n10704 = n10995 & n9;
  assign n10051 = n10960 & n11004;
  assign n10052 = n10975 & n10963;
  assign n10525 = n10947 & n17;
  assign n10057 = n10950 & n10972;
  assign n9994 = n10956 & n10952;
  assign n10063 = n10975 & n10999;
  assign n10064 = n10950 & n10994;
  assign n10023 = n10987 & n10973;
  assign n10069 = n10953 & n10989;
  assign n10072 = n10978 & n11004;
  assign n10074 = n10956 & n10979;
  assign n10075 = n10953 & n10966;
  assign n10077 = n10950 & n10999;
  assign n10080 = n10970 & n10961;
  assign n10082 = n10978 & n10952;
  assign n10086 = n10970 & n10965;
  assign n10267 = n10964 & n6;
  assign n10088 = n10967 & n10977;
  assign n10488 = n10995 & n11;
  assign n10094 = n10975 & n10959;
  assign n9992 = n10993 & n10989;
  assign n10097 = n10948 & n10981;
  assign n10100 = n10960 & n10965;
  assign n10218 = n10967 & n10959;
  assign n10101 = n10980 & n10954;
  assign n10605 = n10986 & n18;
  assign n10106 = n10975 & n10997;
  assign n10107 = n10956 & n10988;
  assign n10119 = n10956 & n10966;
  assign n10120 = n10978 & n10974;
  assign n10121 = n10976 & n11004;
  assign n10122 = n10960 & n10949;
  assign n10115 = n10967 & n10999;
  assign n10128 = n10978 & n10959;
  assign n10130 = n10976 & n11005;
  assign n10131 = n10976 & n10971;
  assign n10133 = n10968 & n10965;
  assign n9989 = n10975 & n11004;
  assign n10135 = n10978 & n11005;
  assign n10136 = n10987 & n10954;
  assign n10137 = n10978 & n10957;
  assign n10138 = n10960 & n10969;
  assign n10140 = n10970 & n10954;
  assign n10762 = n11013 & n15;
  assign n10712 = n10947 & n23;
  assign n10144 = n10948 & n10988;
  assign n10576 = n10998 & n11;
  assign n10145 = n10970 & n10952;
  assign n10211 = n10950 & n10981;
  assign n10147 = n10980 & n10957;
  assign n10149 = n10956 & n10965;
  assign n10123 = n10950 & n10973;
  assign n10151 = n10956 & n10949;
  assign n10153 = n10978 & n11003;
  assign n10155 = n10976 & n10952;
  assign n9987 = n10960 & n10966;
  assign n10216 = n10951 & n10974;
  assign n10157 = n10956 & n10999;
  assign n10160 = n10960 & n10990;
  assign n10163 = n10967 & n10989;
  assign n9976 = n10960 & n10989;
  assign n10165 = n10980 & n10949;
  assign n10167 = n10967 & n10961;
  assign n10170 = n10950 & n10992;
  assign n10174 = n10956 & n10994;
  assign n10176 = n10980 & n10966;
  assign n10179 = n10967 & n11004;
  assign n10580 = n11014 & n20;
  assign n9986 = n10993 & n10971;
  assign n10181 = n10967 & n11000;
  assign n10185 = n10970 & n10972;
  assign n10186 = n10993 & n10954;
  assign n10191 = n10960 & n10954;
  assign n10763 = n10995 & n26;
  assign n10197 = n10993 & n10949;
  assign n10198 = n10980 & n10990;
  assign n9984 = n10953 & n10973;
  assign n10127 = n10978 & n11000;
  assign n10202 = n10987 & n10959;
  assign n10203 = n10970 & n10990;
  assign n10210 = n10968 & n10992;
  assign n10341 = n10960 & n11003;
  assign n10205 = n10976 & n10963;
  assign n10207 = n10960 & n10994;
  assign n10215 = n10948 & n10962;
  assign n10213 = n10970 & n10999;
  assign n10214 = n10956 & n10997;
  assign n10118 = n10978 & n10949;
  assign n10126 = n10968 & n10966;
  assign n10335 = n10987 & n10949;
  assign n10125 = n10956 & n11005;
  assign n10232 = n10956 & n10971;
  assign n10212 = n10987 & n10981;
  assign n10236 = n10960 & n10959;
  assign n10124 = n10951 & n11003;
  assign n9981 = n10978 & n10962;
  assign n10248 = n10993 & n10962;
  assign n10209 = n10978 & n10990;
  assign n9979 = n10953 & n11004;
  assign n10208 = n10950 & n10974;
  assign n10263 = n10956 & n10961;
  assign n10264 = n10953 & n10999;
  assign n10342 = n10948 & n10990;
  assign n9977 = n10976 & n10981;
  assign n10206 = n10975 & n10965;
  assign n10474 = n11012 & n8;
  assign n9975 = n10970 & n11004;
  assign n10281 = n10978 & n10977;
  assign n10283 = n10948 & n10997;
  assign n10109 = n10951 & n10973;
  assign n10549 = n10964 & n27;
  assign n10545 = n10975 & n10974;
  assign n10331 = n10970 & n10992;
  assign n10292 = n10967 & n10954;
  assign n10293 = n10948 & n10977;
  assign n9958 = n10953 & n10971;
  assign n10297 = n10951 & n10971;
  assign n10116 = n10956 & n10972;
  assign n10312 = n10975 & n10969;
  assign n10113 = n10960 & n11000;
  assign n10201 = n10960 & n10974;
  assign n10112 = n10948 & n10952;
  assign n10200 = n10993 & n10959;
  assign n10842 = n10958 & n4;
  assign n10111 = n10956 & n10992;
  assign n10199 = n10953 & n10997;
  assign n10110 = n10968 & n10989;
  assign n10754 = n11002 & n28;
  assign n10003 = n10948 & n10973;
  assign n10108 = n10968 & n10994;
  assign n10196 = n10987 & n10961;
  assign n10850 = n10964 & n0;
  assign n10861 = n10986 & n3;
  assign n10701 = n11014 & n8;
  assign n10379 = n10993 & n10952;
  assign n10841 = n11006 & n21;
  assign n10105 = n10993 & n11003;
  assign n10104 = n10950 & n11004;
  assign n10189 = n10970 & n10994;
  assign n10395 = n10967 & n10969;
  assign n10103 = n10953 & n11003;
  assign n10344 = n10970 & n10974;
  assign n10190 = n10993 & n10974;
  assign n10102 = n10987 & n10977;
  assign n10187 = n10980 & n10979;
  assign n10093 = n10967 & n10949;
  assign n10838 = n11002 & n29;
  assign n10559 = n11006 & n27;
  assign n10188 = n10970 & n10966;
  assign n10424 = n10968 & n11007;
  assign n10229 = n10993 & n11004;
  assign n10430 = n10967 & n11007;
  assign n10099 = n10960 & n10996;
  assign n10432 = n10980 & n11007;
  assign n10436 = n10978 & n11007;
  assign n10437 = n10970 & n10969;
  assign n10837 = n11014 & n10;
  assign n10183 = n10960 & n10977;
  assign n10562 = n10955 & n25;
  assign n10445 = n10964 & n8;
  assign n10447 = n10986 & n15;
  assign n10835 = n11002 & n25;
  assign n10449 = n10955 & n29;
  assign n10184 = n10951 & n10979;
  assign n10453 = n11012 & n11;
  assign n10096 = n10976 & n10989;
  assign n10457 = n11012 & n12;
  assign n10182 = n10953 & n11005;
  assign n10461 = n10946 & n17;
  assign n10463 = n10958 & n18;
  assign n10095 = n10968 & n10957;
  assign n10464 = n11002 & n15;
  assign n10475 = n10968 & n11003;
  assign n10468 = n10998 & n15;
  assign n10345 = n10978 & n10997;
  assign n10497 = n10968 & n10961;
  assign n10090 = n10950 & n11000;
  assign n10478 = n11013 & n21;
  assign n10834 = n10998 & n31;
  assign n10480 = n10998 & n24;
  assign n10484 = n10964 & n3;
  assign n10092 = n10993 & n10997;
  assign n10698 = n10955 & n4;
  assign n10490 = n10951 & n10992;
  assign n10495 = n10946 & n11;
  assign n10180 = n10975 & n10981;
  assign n10091 = n10953 & n10949;
  assign n10481 = n10980 & n11003;
  assign n10177 = n10948 & n10957;
  assign n10505 = n10958 & n12;
  assign n10465 = n10946 & n3;
  assign n10849 = n10995 & n24;
  assign n10351 = n10956 & n11004;
  assign n10178 = n10951 & n10961;
  assign n10515 = n10970 & n10979;
  assign n10175 = n10993 & n10966;
  assign n10532 = n10998 & n3;
  assign n10523 = n10958 & n31;
  assign n10089 = n10970 & n10977;
  assign n10572 = n10986 & n20;
  assign n10851 = n11002 & n27;
  assign n10534 = n10991 & n10;
  assign n10533 = n10970 & n10959;
  assign n10538 = n10958 & n15;
  assign n10682 = n10948 & n10963;
  assign n10586 = n11014 & n30;
  assign n10541 = n10964 & n29;
  assign n10173 = n10950 & n10988;
  assign n10462 = n11006 & n16;
  assign n10571 = n10995 & n29;
  assign n10713 = n10986 & n4;
  assign n10547 = n11014 & n24;
  assign n10004 = n10980 & n10961;
  assign n10553 = n11001 & n30;
  assign n10349 = n10980 & n10981;
  assign n10564 = n11012 & n7;
  assign n10330 = n10968 & n10971;
  assign n10573 = n10991 & n13;
  assign n9959 = n11001 & n19;
  assign n10005 = n10967 & n10979;
  assign n10577 = n10991 & n6;
  assign n10692 = n10998 & n18;
  assign n10585 = n11006 & n19;
  assign n10570 = n10958 & n14;
  assign n10596 = n10946 & n6;
  assign n10760 = n10998 & n16;
  assign n10568 = n11013 & n1;
  assign n10328 = n10968 & n10959;
  assign n10608 = n10947 & n26;
  assign n10691 = n11002 & n23;
  assign n10624 = n10947 & n28;
  assign n10628 = n11013 & n26;
  assign n10569 = n10947 & n18;
  assign n10632 = n10946 & n15;
  assign n10639 = n10947 & n7;
  assign n10327 = n10987 & n10957;
  assign n10636 = n10947 & n0;
  assign n10689 = n11012 & n19;
  assign n10690 = n11013 & n30;
  assign n10455 = n11014 & n9;
  assign n10460 = n10998 & n30;
  assign n10757 = n11006 & n10;
  assign n10656 = n10955 & n18;
  assign n10459 = n11013 & n24;
  assign n10688 = n11013 & n9;
  assign n10663 = n11001 & n2;
  assign n10479 = n10964 & n31;
  assign n10491 = n11012 & n30;
  assign n10671 = n10958 & n20;
  assign n10673 = n11013 & n19;
  assign n10674 = n11002 & n18;
  assign n10687 = n11014 & n17;
  assign n10567 = n10986 & n31;
  assign n10755 = n10958 & n27;
  assign n10326 = n10976 & n10999;
  assign n10458 = n10947 & n14;
  assign n10831 = n11001 & n17;
  assign n10695 = n10995 & n4;
  assign n10134 = n10956 & n10990;
  assign n10268 = n10976 & n10961;
  assign n10566 = n10958 & n23;
  assign n10565 = n11014 & n12;
  assign n10587 = n10998 & n29;
  assign n10717 = n11012 & n2;
  assign n10325 = n10948 & n10999;
  assign n10413 = n10951 & n9939;
  assign n10729 = n11002 & n7;
  assign n10323 = n10978 & n10971;
  assign n10733 = n11001 & n28;
  assign n10456 = n11001 & n27;
  assign n10744 = n11012 & n27;
  assign n10685 = n10946 & n1;
  assign n10584 = n11012 & n29;
  assign n10752 = n10947 & n16;
  assign n10756 = n10958 & n1;
  assign n10563 = n10995 & n19;
  assign n10764 = n10958 & n5;
  assign n10324 = n10948 & n11003;
  assign n10780 = n11013 & n17;
  assign n10792 = n10998 & n25;
  assign n10797 = n10964 & n17;
  assign n10801 = n10998 & n6;
  assign n10561 = n10946 & n8;
  assign n10807 = n10998 & n14;
  assign n10129 = n10993 & n10963;
  assign n10817 = n10995 & n1;
  assign n10821 = n10946 & n5;
  assign n10454 = n10955 & n14;
  assign n10444 = n10995 & n0;
  assign n10829 = n10991 & n19;
  assign n10833 = n10947 & n11;
  assign n10322 = n10951 & n10969;
  assign n10836 = n11012 & n22;
  assign n10840 = n10991 & n11;
  assign n10844 = n11014 & n18;
  assign n10494 = n10991 & n12;
  assign n10848 = n10986 & n5;
  assign n10852 = n11006 & n13;
  assign n10856 = n11012 & n25;
  assign n10217 = n10987 & n10971;
  assign n10513 = n10947 & n1;
  assign n10868 = n10995 & n16;
  assign n10872 = n11013 & n5;
  assign n10874 = n11013 & n27;
  assign n10876 = n10998 & n4;
  assign n10880 = n11001 & n22;
  assign n10321 = n10993 & n10981;
  assign n10017 = n10968 & n11005;
  assign n10270 = n10948 & n11005;
  assign n10028 = n10951 & n10988;
  assign n10888 = n10995 & n31;
  assign n10891 = n10955 & n12;
  assign n10892 = n11002 & n1;
  assign n10896 = n11002 & n17;
  assign n10898 = n11012 & n10;
  assign n10859 = n10946 & n28;
  assign n10681 = n10995 & n21;
  assign n10827 = n10986 & n23;
  assign n10814 = n10947 & n9;
  assign n10823 = n11001 & n13;
  assign n10589 = n10998 & n1;
  assign n10753 = n11002 & n3;
  assign n10828 = n11001 & n10;
  assign n10683 = n10986 & n12;
  assign n10452 = n11001 & n1;
  assign n10751 = n10991 & n2;
  assign n10899 = n10995 & n12;
  assign n10526 = n11001 & n7;
  assign n10320 = n10951 & n10957;
  assign n10244 = n10978 & n10992;
  assign n10680 = n11014 & n11;
  assign n10714 = n10991 & n31;
  assign n10029 = n10987 & n10962;
  assign n10826 = n11013 & n7;
  assign n10450 = n10946 & n23;
  assign n10502 = n11001 & n16;
  assign n10451 = n11006 & n3;
  assign n10294 = n10948 & n10961;
  assign n10825 = n10986 & n28;
  assign n10679 = n11006 & n12;
  assign n10903 = n10955 & n26;
  assign n10824 = n10946 & n13;
  assign n10609 = n11012 & n16;
  assign n10697 = n10995 & n13;
  assign n10945 = n10976 & n10974;
  assign n10298 = n10953 & n10972;
  assign n10250 = n10951 & n10990;
  assign n10715 = n11013 & n10;
  assign n10295 = n10978 & n10989;
  assign n10139 = n10976 & n10966;
  assign n10897 = n10947 & n8;
  assign n10384 = n10975 & n10957;
  assign n10822 = n11002 & n14;
  assign n10610 = n10991 & n17;
  assign n10448 = n11014 & n26;
  assign n10716 = n10947 & n25;
  assign n10296 = n10953 & n10959;
  assign n10677 = n10955 & n23;
  assign n10030 = n10970 & n10962;
  assign n10749 = n11002 & n20;
  assign n10819 = n10958 & n17;
  assign n10611 = n10995 & n28;
  assign n10820 = n11002 & n12;
  assign n10676 = n10995 & n25;
  assign n10748 = n11014 & n19;
  assign n10895 = n10958 & n19;
  assign n10528 = n10946 & n16;
  assign n10272 = n10960 & n10952;
  assign n10854 = n10958 & n10;
  assign n10894 = n10964 & n12;
  assign n10775 = n10986 & n26;
  assign n10446 = n11014 & n15;
  assign n10527 = n10991 & n22;
  assign n10273 = n10980 & n11000;
  assign n10597 = n10995 & n6;
  assign n10818 = n11006 & n22;
  assign n10675 = n11006 & n14;
  assign n10031 = n10987 & n10965;
  assign n10607 = n10964 & n26;
  assign n10141 = n10978 & n10973;
  assign n10718 = n11002 & n10;
  assign n10893 = n10998 & n21;
  assign n10746 = n10955 & n28;
  assign n10906 = n10975 & n10989;
  assign n10416 = n10976 & n9939;
  assign n10085 = n10967 & n10966;
  assign n10907 = n10998 & n10;
  assign n10776 = n11006 & n31;
  assign n10271 = n10976 & n10972;
  assign n10747 = n10991 & n26;
  assign n10613 = n10955 & n3;
  assign n10719 = n11002 & n0;
  assign n10816 = n11001 & n31;
  assign n10439 = n10970 & n11007;
  assign n10275 = n10967 & n10962;
  assign n10560 = n11002 & n16;
  assign n10084 = n10967 & n10996;
  assign n10142 = n10980 & n10962;
  assign n10143 = n10975 & n10949;
  assign n10614 = n10991 & n5;
  assign n10503 = n11002 & n4;
  assign n10172 = n10980 & n10965;
  assign n10009 = n10948 & n10974;
  assign n10319 = n10987 & n11004;
  assign n10720 = n10986 & n10;
  assign n10299 = n10970 & n10963;
  assign n10672 = n11014 & n22;
  assign n10815 = n10986 & n19;
  assign n10615 = n10986 & n2;
  assign n10409 = n10967 & n9939;
  assign n10813 = n11013 & n4;
  assign n10274 = n10968 & n10988;
  assign n10318 = n10970 & n10957;
  assign n10866 = n10955 & n21;
  assign n10832 = n10955 & n6;
  assign n10276 = n10980 & n10971;
  assign n10670 = n10991 & n23;
  assign n10721 = n10955 & n13;
  assign n10668 = n10964 & n14;
  assign n10707 = n10958 & n8;
  assign n10890 = n10964 & n7;
  assign n10805 = n11002 & n6;
  assign n10035 = n10950 & n10954;
  assign n10864 = n10964 & n10;
  assign n10779 = n10947 & n2;
  assign n10669 = n11014 & n0;
  assign n10653 = n10955 & n22;
  assign n10353 = n10975 & n11003;
  assign n10742 = n10998 & n2;
  assign n10504 = n10995 & n23;
  assign n10770 = n11014 & n5;
  assign n10867 = n10986 & n7;
  assign n10667 = n10991 & n18;
  assign n10666 = n11012 & n23;
  assign n10265 = n10956 & n10962;
  assign n10558 = n10998 & n19;
  assign n10777 = n10995 & n3;
  assign n10434 = n10956 & n11007;
  assign n10557 = n11001 & n15;
  assign n10037 = n10975 & n10966;
  assign n10556 = n11006 & n7;
  assign n10743 = n10955 & n27;
  assign n10812 = n10991 & n20;
  assign n10617 = n11014 & n23;
  assign n10811 = n11013 & n6;
  assign n10665 = n11006 & n26;
  assign n10664 = n11001 & n20;
  assign n10301 = n10980 & n10973;
  assign n10772 = n11001 & n21;
  assign n9955 = n10964 & n25;
  assign n10278 = n10993 & n10979;
  assign n10723 = n10998 & n22;
  assign n10006 = n10976 & n10965;
  assign n10912 = n11002 & n19;
  assign n10660 = n11006 & n18;
  assign n10662 = n11001 & n25;
  assign n10427 = n10987 & n11007;
  assign n10810 = n10991 & n30;
  assign n10661 = n11006 & n4;
  assign n10391 = n10980 & n10972;
  assign n10910 = n10946 & n20;
  assign n10039 = n10993 & n10999;
  assign n10496 = n11012 & n31;
  assign n10279 = n10993 & n10965;
  assign n10038 = n10987 & n10969;
  assign n10392 = n10976 & n10959;
  assign n10741 = n11013 & n25;
  assign n10590 = n11012 & n24;
  assign n10913 = n10991 & n1;
  assign n10280 = n10950 & n10949;
  assign n10555 = n11012 & n18;
  assign n10809 = n11012 & n15;
  assign n10659 = n11013 & n28;
  assign n10282 = n10978 & n10988;
  assign n10914 = n10987 & n11003;
  assign n10554 = n11001 & n26;
  assign n10808 = n10986 & n9;
  assign n10738 = n11012 & n5;
  assign n10658 = n11014 & n1;
  assign n10171 = n10953 & n10977;
  assign n10657 = n10958 & n0;
  assign n10740 = n11001 & n0;
  assign n10915 = n11001 & n3;
  assign n10169 = n10950 & n10977;
  assign n10588 = n11002 & n22;
  assign n10506 = n11002 & n21;
  assign n10654 = n11013 & n0;
  assign n10739 = n11002 & n5;
  assign n10655 = n10991 & n9;
  assign n10806 = n10946 & n19;
  assign n10489 = n11012 & n14;
  assign n10737 = n10955 & n1;
  assign n10917 = n10991 & n15;
  assign n10168 = n10967 & n10973;
  assign n10552 = n10995 & n30;
  assign n10652 = n11002 & n2;
  assign n10443 = n10947 & n5;
  assign n10791 = n11014 & n3;
  assign n10373 = n10951 & n11004;
  assign n10420 = n10968 & n9939;
  assign n10422 = n10978 & n9939;
  assign n10651 = n11012 & n4;
  assign n10498 = n10958 & n11;
  assign n10803 = n10955 & n15;
  assign n10804 = n11014 & n28;
  assign n10419 = n10987 & n9939;
  assign n10736 = n11006 & n17;
  assign n10693 = n10964 & n28;
  assign n10516 = n11002 & n9;
  assign n10650 = n10958 & n3;
  assign n10256 = n10948 & n10965;
  assign n10551 = n10946 & n18;
  assign n10592 = n11014 & n29;
  assign n10734 = n10998 & n28;
  assign n10649 = n10986 & n17;
  assign n10800 = n10964 & n13;
  assign n10647 = n10946 & n14;
  assign n10517 = n10947 & n12;
  assign n10550 = n11014 & n13;
  assign n10802 = n11014 & n7;
  assign n10708 = n10986 & n24;
  assign n10376 = n10993 & n10969;
  assign n10735 = n11002 & n30;
  assign n10921 = n10993 & n10973;
  assign n10648 = n11001 & n9;
  assign n10041 = n10976 & n10990;
  assign n10499 = n10986 & n25;
  assign n10166 = n10968 & n10999;
  assign n10645 = n11002 & n26;
  assign n10514 = n10955 & n30;
  assign n10397 = n10953 & n10979;
  assign n10548 = n10958 & n13;
  assign n10598 = n10964 & n4;
  assign n10599 = n10946 & n4;
  assign n10646 = n10958 & n28;
  assign n10593 = n11001 & n14;
  assign n10918 = n10991 & n29;
  assign n10919 = n10986 & n11;
  assign n10889 = n10955 & n8;
  assign n10709 = n11002 & n8;
  assign n10923 = n11012 & n28;
  assign n9965 = n10964 & n23;
  assign n10643 = n11002 & n13;
  assign n10885 = n10998 & n0;
  assign n10773 = n11012 & n13;
  assign n10641 = n11013 & n20;
  assign n10042 = n10980 & n10999;
  assign n10766 = n11001 & n24;
  assign n10644 = n11006 & n24;
  assign n10518 = n10998 & n8;
  assign n10799 = n10986 & n14;
  assign n10386 = n10950 & n10969;
  assign n10798 = n10955 & n31;
  assign n10887 = n10964 & n24;
  assign n10600 = n11013 & n31;
  assign n10724 = n11013 & n3;
  assign n10500 = n11013 & n16;
  assign n10886 = n11006 & n1;
  assign n10285 = n10975 & n10972;
  assign n10642 = n11001 & n23;
  assign n10778 = n11006 & n5;
  assign n10043 = n10978 & n10972;
  assign n10796 = n10947 & n3;
  assign n10863 = n10958 & n16;
  assign n10881 = n11006 & n0;
  assign n10036 = n10967 & n10997;
  assign n10794 = n10964 & n2;
  assign n9954 = n10947 & n4;
  assign n10640 = n10991 & n27;
  assign n10884 = n11012 & n21;
  assign n10044 = n10993 & n10977;
  assign n10793 = n11013 & n11;
  assign n10638 = n10986 & n1;
  assign n10883 = n10958 & n24;
  assign n10882 = n10995 & n10;
  assign n10286 = n10980 & n10977;
  assign n10637 = n10998 & n27;
  assign n10879 = n10995 & n7;
  assign n10875 = n10946 & n9;
  assign n10870 = n10955 & n10;
  assign n10635 = n10955 & n7;
  assign n10873 = n11013 & n8;
  assign n10877 = n11002 & n24;
  assign n10930 = n10950 & n10962;
  assign n10302 = n10951 & n11005;
  assign n10790 = n11001 & n5;
  assign n10634 = n11001 & n6;
  assign n10428 = n10951 & n11007;
  assign n10789 = n11006 & n25;
  assign n10878 = n11013 & n23;
  assign n10633 = n10947 & n15;
  assign n10853 = n10958 & n7;
  assign n10788 = n10995 & n20;
  assign n10284 = n10993 & n10988;
  assign n10402 = n10950 & n10990;
  assign n10047 = n10968 & n10997;
  assign n10418 = n10993 & n9939;
  assign n10629 = n10964 & n18;
  assign n10631 = n10986 & n6;
  assign n10787 = n10964 & n15;
  assign n10442 = n10991 & n16;
  assign n10544 = n10958 & n26;
  assign n10618 = n11013 & n12;
  assign n10403 = n10950 & n11003;
  assign n10262 = n10970 & n11003;
  assign n10732 = n10946 & n21;
  assign n10931 = n10967 & n10988;
  assign n10546 = n10998 & n12;
  assign n10905 = n11006 & n30;
  assign n10083 = n10970 & n10996;
  assign n10288 = n10967 & n10965;
  assign n10630 = n11012 & n1;
  assign n10079 = n10975 & n10962;
  assign n10317 = n10968 & n10981;
  assign n10927 = n10975 & n10992;
  assign n10316 = n10951 & n10997;
  assign n10441 = n10991 & n0;
  assign n10381 = n10948 & n10994;
  assign n10933 = n11014 & n6;
  assign n10932 = n10951 & n10962;
  assign n10287 = n10978 & n10996;
  assign n10616 = n11014 & n27;
  assign n10758 = n10958 & n30;
  assign n10627 = n10998 & n17;
  assign n10543 = n11013 & n14;
  assign n10601 = n10958 & n9;
  assign n10081 = n10956 & n10959;
  assign n10440 = n11006 & n23;
  assign n10304 = n10948 & n11000;
  assign n10154 = n10951 & n11000;
  assign n10519 = n10958 & n29;
  assign n10934 = n10978 & n10963;
  assign n10542 = n11002 & n31;
  assign n10731 = n10947 & n31;
  assign n10423 = n10953 & n9939;
  assign n10539 = n10955 & n17;
  assign n10305 = n10987 & n10996;
  assign n10540 = n11006 & n15;
  assign n10786 = n10946 & n26;
  assign n10745 = n10998 & n26;
  assign n10785 = n11014 & n16;
  assign n10730 = n10995 & n17;
  assign n10306 = n10967 & n10963;
  assign n10078 = n10980 & n10992;
  assign n10626 = n11001 & n12;
  assign n10050 = n10948 & n10989;
  assign n10315 = n10951 & n10994;
  assign n10407 = n10978 & n10969;
  assign n10771 = n10986 & n16;
  assign n10937 = n10960 & n10973;
  assign n10938 = n10955 & n5;
  assign n10429 = n10948 & n11007;
  assign n10438 = n10953 & n11007;
  assign n10625 = n10947 & n20;
  assign n10722 = n10964 & n30;
  assign n10941 = n10987 & n11000;
  assign n10053 = n10950 & n10997;
  assign n10411 = n10948 & n9939;
  assign n10314 = n10975 & n11005;
  assign n10619 = n10995 & n27;
  assign n10431 = n10960 & n11007;
  assign n10065 = n10987 & n10974;
  assign n10623 = n10946 & n24;
  assign n10728 = n10946 & n10;
  assign n10289 = n10980 & n11004;
  assign n10936 = n11014 & n21;
  assign n10536 = n10955 & n19;
  assign n10300 = n10953 & n10992;
  assign n10727 = n10991 & n25;
  assign n10537 = n10946 & n29;
  assign n10621 = n11014 & n31;
  assign n10622 = n10986 & n27;
  assign n10277 = n10987 & n10989;
  assign n10408 = n10987 & n10999;
  assign n10308 = n10956 & n10963;
  assign n10781 = n11014 & n14;
  assign n10784 = n10946 & n7;
  assign n10620 = n10946 & n30;
  assign n10310 = n10980 & n10959;
  assign n9953 = n10986 & n30;
  assign n10156 = n10975 & n10977;
  assign n10783 = n10964 & n1;
  assign n10520 = n11012 & n17;
  assign n10726 = n10964 & n21;
  assign n10869 = n10958 & n6;
  assign n10939 = n10950 & n10989;
  assign n10782 = n10947 & n24;
  assign n10007 = n10950 & n11005;
  assign n10309 = n10951 & n10966;
  assign n10076 = n10987 & n11005;
  assign n10433 = n10950 & n11007;
  assign n10535 = n10991 & n28;
  assign n10313 = n10976 & n10969;
  assign n10073 = n10993 & n10996;
  assign n10725 = n11006 & n28;
  assign n10522 = n10947 & n21;
  assign n10531 = n11013 & n22;
  assign n10435 = n10976 & n11007;
  assign n10311 = n10953 & n10974;
  assign n9964 = n11006 & n29;
  assign n10940 = n10960 & n10957;
  assign n10594 = n10947 & n27;
  assign n10512 = n11001 & n18;
  assign n10164 = n10976 & n10979;
  assign n10071 = n10970 & n10988;
  assign n10070 = n10968 & n11000;
  assign n10426 = n10993 & n11007;
  assign n10161 = n10978 & n10954;
  assign n10066 = n10987 & n10966;
  assign n10068 = n10956 & n10989;
  assign n10132 = n10993 & n11000;
  assign n10059 = n10975 & n10988;
  assign n9956 = n11012 & n20;
  assign n10060 = n10975 & n10996;
  assign n10061 = n10976 & n11003;
  assign n10062 = n10976 & n10997;
  assign n10159 = n10960 & n11005;
  assign n10158 = n10953 & n10969;
  assign n10354 = n10953 & n11000;
  assign n10303 = n10951 & n10972;
  assign n10058 = n10970 & n11000;
  assign n10926 = n10947 & n22;
  assign n10710 = n10947 & n19;
  assign n10529 = n11012 & n9;
  assign n10612 = n10986 & n13;
  assign n10067 = n10978 & n10965;
  assign n10162 = n10960 & n10971;
  assign n10530 = n11006 & n20;
  assign n10765 = n11012 & n26;
  assign n10521 = n11012 & n6;
  assign n10604 = n11013 & n2;
  assign n10056 = n10993 & n10972;
  assign n10290 = n10968 & n10949;
  assign n10055 = n10951 & n10981;
  assign n10054 = n10975 & n10973;
  assign n10421 = n10970 & n9939;
  assign n10025 = n10951 & n10965;
  assign n10150 = n10948 & n10996;
  assign n10148 = n10975 & n10979;
  assign n10146 = n10953 & n10961;
  assign n10193 = n10970 & n10989;
  assign n10032 = n10948 & n10966;
  assign n10417 = n10975 & n9939;
  assign n10769 = n10946 & n27;
  assign n10943 = n10976 & n10957;
  assign n10684 = n10955 & n20;
  assign n10414 = n10960 & n9939;
  assign n10192 = n10953 & n10996;
  assign n10768 = n11006 & n9;
  assign n10865 = n10991 & n3;
  assign n10839 = n10958 & n21;
  assign n10194 = n10953 & n10994;
  assign n10415 = n10980 & n9939;
  assign n10944 = n10967 & n10974;
  assign n10269 = n10970 & n11005;
  assign n10195 = n10976 & n10962;
  assign n10767 = n10947 & n29;
  assign n10412 = n10956 & n9939;
  assign n10026 = n10976 & n10994;
  assign n10266 = n10956 & n10981;
  assign n10702 = n11014 & n2;
  assign n9940 = n11080 & n11081;
  assign n10382 = ~n10976;
  assign n10355 = ~n10975;
  assign n10346 = ~n10948;
  assign n9968 = ~n10951;
  assign n9967 = ~n10993;
  assign n10307 = ~n10970;
  assign n9970 = ~n10987;
  assign n9969 = ~n10953;
  assign n10329 = ~n10960;
  assign n9971 = ~n10967;
  assign n9973 = ~n10978;
  assign n9972 = ~n10956;
  assign n10406 = ~n10950;
  assign n10371 = ~n10980;
  assign n11019 = n11113 & n11114;
  assign n11027 = n11176 & n11177;
  assign n11043 = n11228 & n11229;
  assign n11041 = n11232 & n11233;
  assign n11045 = n11271 & n11272;
  assign n11049 = n11279 & n11280;
  assign n11066 = n11301 & n11302;
  assign n10900 = n11333 & n11334;
  assign n11035 = n11385 & n11386;
  assign n11021 = n11427 & n11428;
  assign n11023 = n11430 & n11431;
  assign n11033 = n11438 & n11439;
  assign n11055 = n11628 & n11629;
  assign n11057 = n11643 & n11644;
  assign n11017 = n11651 & n11652;
  assign n11053 = n11656 & n11657;
  assign n11008 = n11691 & n11692;
  assign n11031 = n11713 & n11714;
  assign n11068 = n11807 & n11808;
  assign n10982 = n11865 & n11866;
  assign n11025 = n11916 & n11917;
  assign n11015 = n11920 & n11921;
  assign n11039 = n11923 & n11924;
  assign n11037 = n11925 & n11926;
  assign n11047 = n11928 & n11929;
  assign n11051 = n11930 & n11931;
  assign n11029 = n11932 & n11933;
  assign n11010 = n11934 & n11935;
  assign n11059 = n11982 & n11983;
  assign n11063 = n12058 & n12059;
  assign n11061 = n12101 & n12102;
  assign n10984 = n12107 & n12108;
  assign n11088 = ~n12132;
  assign n11100 = ~n12135;
  assign n11074 = ~n12141;
  assign n11082 = ~n12159;
  assign n11072 = ~n12160;
  assign n11096 = ~n12161;
  assign n11084 = ~n12162;
  assign n11070 = ~n12163;
  assign n11076 = ~n12164;
  assign n11092 = ~n12165;
  assign n11094 = ~n12166;
  assign n11078 = ~n12167;
  assign n11086 = ~n12168;
  assign n11098 = ~n12169;
  assign n11090 = ~n12170;
  assign n8004 = n9939 ^ n9940;
  assign n9553 = ~n9952;
  assign n8829 = ~n9953;
  assign n8159 = ~n9954;
  assign n9911 = ~n9955;
  assign n9437 = ~n9956;
  assign n9017 = ~n9958;
  assign n9357 = ~n9959;
  assign n9413 = ~n9960;
  assign n8321 = ~n9961;
  assign n8023 = ~n9962;
  assign n9619 = ~n9964;
  assign n8141 = ~n9965;
  assign n8367 = ~n9966;
  assign n6406 = n9967 & n7073;
  assign n6198 = n9968 & n7051;
  assign n6160 = n9969 & n7045;
  assign n6352 = n9970 & n7027;
  assign n6252 = n9971 & n7010;
  assign n6166 = n9972 & n7047;
  assign n6320 = n9973 & n7059;
  assign n9443 = ~n9974;
  assign n8055 = ~n9975;
  assign n9441 = ~n9976;
  assign n9633 = ~n9977;
  assign n8285 = ~n9978;
  assign n9525 = ~n9979;
  assign n8035 = ~n9980;
  assign n8273 = ~n9981;
  assign n9895 = ~n9982;
  assign n8459 = ~n9983;
  assign n9067 = ~n9984;
  assign n8657 = ~n9985;
  assign n8089 = ~n9986;
  assign n8529 = ~n9987;
  assign n8503 = ~n9988;
  assign n9745 = ~n9989;
  assign n9879 = ~n9990;
  assign n8661 = ~n9991;
  assign n8941 = ~n9992;
  assign n9769 = ~n9993;
  assign n9795 = ~n9994;
  assign n8717 = ~n9995;
  assign n8421 = ~n9996;
  assign n9125 = ~n9997;
  assign n9299 = ~n9998;
  assign n8629 = ~n9999;
  assign n9825 = ~n10000;
  assign n8553 = ~n10001;
  assign n9843 = ~n10002;
  assign n8393 = ~n10003;
  assign n9809 = ~n10004;
  assign n9151 = ~n10005;
  assign n9587 = ~n10006;
  assign n9875 = ~n10007;
  assign n8297 = ~n10008;
  assign n9555 = ~n10009;
  assign n8973 = ~n10010;
  assign n8813 = ~n10011;
  assign n8457 = ~n10012;
  assign n9001 = ~n10013;
  assign n9653 = ~n10014;
  assign n9199 = ~n10015;
  assign n9179 = ~n10016;
  assign n8027 = ~n10017;
  assign n9035 = ~n10018;
  assign n8337 = ~n10019;
  assign n8383 = ~n10020;
  assign n8903 = ~n10021;
  assign n8287 = ~n10022;
  assign n9309 = ~n10023;
  assign n8169 = ~n10024;
  assign n8413 = ~n10025;
  assign n9429 = ~n10026;
  assign n8019 = ~n10027;
  assign n8627 = ~n10028;
  assign n9718 = ~n10029;
  assign n8423 = ~n10030;
  assign n9727 = ~n10031;
  assign n8441 = ~n10032;
  assign n8163 = ~n10033;
  assign n8351 = ~n10034;
  assign n8021 = ~n10035;
  assign n9501 = ~n10036;
  assign n8419 = ~n10037;
  assign n8709 = ~n10038;
  assign n9831 = ~n10039;
  assign n8445 = ~n10040;
  assign n8635 = ~n10041;
  assign n9805 = ~n10042;
  assign n8901 = ~n10043;
  assign n8251 = ~n10044;
  assign n9533 = ~n10045;
  assign n8691 = ~n10046;
  assign n9549 = ~n10047;
  assign n8109 = ~n10048;
  assign n8815 = ~n10049;
  assign n9733 = ~n10050;
  assign n9061 = ~n10051;
  assign n9851 = ~n10052;
  assign n9877 = ~n10053;
  assign n9211 = ~n10054;
  assign n8049 = ~n10055;
  assign n9453 = ~n10056;
  assign n8129 = ~n10057;
  assign n9121 = ~n10058;
  assign n8703 = ~n10059;
  assign n8577 = ~n10060;
  assign n8143 = ~n10061;
  assign n8161 = ~n10062;
  assign n8787 = ~n10063;
  assign n9451 = ~n10064;
  assign n8197 = ~n10065;
  assign n8747 = ~n10066;
  assign n9595 = ~n10067;
  assign n8695 = ~n10068;
  assign n8181 = ~n10069;
  assign n9593 = ~n10070;
  assign n8213 = ~n10071;
  assign n9123 = ~n10072;
  assign n8275 = ~n10073;
  assign n8225 = ~n10074;
  assign n9081 = ~n10075;
  assign n8231 = ~n10076;
  assign n8725 = ~n10077;
  assign n8891 = ~n10078;
  assign n8205 = ~n10079;
  assign n8255 = ~n10080;
  assign n8259 = ~n10081;
  assign n8165 = ~n10082;
  assign n9519 = ~n10083;
  assign n8295 = ~n10084;
  assign n8931 = ~n10085;
  assign n8319 = ~n10086;
  assign n8987 = ~n10087;
  assign n8327 = ~n10088;
  assign n8151 = ~n10089;
  assign n9639 = ~n10090;
  assign n9853 = ~n10091;
  assign n9237 = ~n10092;
  assign n8147 = ~n10093;
  assign n8365 = ~n10094;
  assign n8063 = ~n10095;
  assign n9089 = ~n10096;
  assign n9901 = ~n10097;
  assign n8373 = ~n10099;
  assign n8375 = ~n10100;
  assign n8247 = ~n10101;
  assign n8303 = ~n10102;
  assign n8923 = ~n10103;
  assign n9039 = ~n10104;
  assign n8239 = ~n10105;
  assign n9623 = ~n10106;
  assign n9349 = ~n10107;
  assign n8407 = ~n10108;
  assign n9801 = ~n10109;
  assign n8467 = ~n10110;
  assign n9903 = ~n10111;
  assign n8763 = ~n10112;
  assign n9339 = ~n10113;
  assign n9115 = ~n10114;
  assign n9251 = ~n10115;
  assign n8951 = ~n10116;
  assign n8249 = ~n10117;
  assign n9551 = ~n10118;
  assign n8437 = ~n10119;
  assign n9865 = ~n10120;
  assign n9145 = ~n10121;
  assign n9897 = ~n10122;
  assign n8543 = ~n10123;
  assign n9133 = ~n10124;
  assign n8067 = ~n10125;
  assign n9461 = ~n10126;
  assign n9747 = ~n10127;
  assign n9301 = ~n10128;
  assign n8473 = ~n10129;
  assign n8965 = ~n10130;
  assign n8481 = ~n10131;
  assign n8515 = ~n10132;
  assign n8663 = ~n10133;
  assign n8609 = ~n10134;
  assign n8455 = ~n10135;
  assign n9755 = ~n10136;
  assign n8011 = ~n10137;
  assign n8789 = ~n10138;
  assign n8061 = ~n10139;
  assign n9713 = ~n10140;
  assign n8959 = ~n10141;
  assign n8469 = ~n10142;
  assign n8897 = ~n10143;
  assign n8953 = ~n10144;
  assign n9479 = ~n10145;
  assign n8265 = ~n10146;
  assign n9905 = ~n10147;
  assign n8261 = ~n10148;
  assign n9419 = ~n10149;
  assign n9859 = ~n10150;
  assign n8557 = ~n10151;
  assign n8563 = ~n10152;
  assign n8569 = ~n10153;
  assign n8567 = ~n10154;
  assign n8711 = ~n10155;
  assign n8871 = ~n10156;
  assign n9227 = ~n10157;
  assign n9455 = ~n10158;
  assign n8581 = ~n10159;
  assign n9815 = ~n10160;
  assign n8605 = ~n10161;
  assign n8137 = ~n10162;
  assign n8613 = ~n10163;
  assign n9247 = ~n10164;
  assign n8277 = ~n10165;
  assign n8895 = ~n10166;
  assign n8625 = ~n10167;
  assign n9003 = ~n10168;
  assign n9267 = ~n10169;
  assign n9515 = ~n10170;
  assign n8655 = ~n10171;
  assign n8737 = ~n10172;
  assign n9075 = ~n10173;
  assign n8187 = ~n10174;
  assign n8133 = ~n10175;
  assign n8685 = ~n10176;
  assign n9315 = ~n10177;
  assign n9433 = ~n10178;
  assign n8917 = ~n10179;
  assign n9005 = ~n10180;
  assign n8431 = ~n10181;
  assign n8733 = ~n10182;
  assign n8253 = ~n10183;
  assign n8741 = ~n10184;
  assign n9129 = ~n10185;
  assign n9175 = ~n10186;
  assign n8929 = ~n10187;
  assign n8755 = ~n10188;
  assign n8597 = ~n10189;
  assign n8091 = ~n10190;
  assign n8009 = ~n10191;
  assign n8617 = ~n10192;
  assign n9369 = ~n10193;
  assign n8843 = ~n10194;
  assign n9399 = ~n10195;
  assign n9611 = ~n10196;
  assign n8359 = ~n10197;
  assign n9197 = ~n10198;
  assign n9269 = ~n10199;
  assign n9167 = ~n10200;
  assign n8679 = ~n10201;
  assign n9375 = ~n10202;
  assign n9787 = ~n10203;
  assign n8809 = ~n10204;
  assign n8401 = ~n10205;
  assign n8821 = ~n10206;
  assign n8847 = ~n10207;
  assign n8849 = ~n10208;
  assign n9173 = ~n10209;
  assign n8047 = ~n10210;
  assign n8977 = ~n10211;
  assign n8403 = ~n10212;
  assign n9621 = ~n10213;
  assign n8855 = ~n10214;
  assign n8863 = ~n10215;
  assign n9423 = ~n10216;
  assign n8867 = ~n10217;
  assign n9761 = ~n10218;
  assign n8117 = ~n10219;
  assign n8877 = ~n10220;
  assign n8811 = ~n10221;
  assign n8497 = ~n10222;
  assign n9365 = ~n10223;
  assign n8767 = ~n10224;
  assign n8889 = ~n10225;
  assign n9935 = ~n10226;
  assign n8015 = ~n10229;
  assign n9692 = ~n10230;
  assign n8537 = ~n10231;
  assign n8909 = ~n10232;
  assign n9573 = ~n10233;
  assign n8937 = ~n10234;
  assign n8715 = ~n10235;
  assign n9485 = ~n10236;
  assign n8323 = ~n10237;
  assign n9907 = ~n10238;
  assign n8981 = ~n10239;
  assign n8531 = ~n10240;
  assign n9165 = ~n10241;
  assign n9313 = ~n10242;
  assign n8911 = ~n10243;
  assign n8743 = ~n10244;
  assign n9571 = ~n10245;
  assign n8963 = ~n10246;
  assign n9353 = ~n10247;
  assign n8643 = ~n10248;
  assign n9465 = ~n10249;
  assign n8105 = ~n10250;
  assign n8521 = ~n10251;
  assign n9007 = ~n10252;
  assign n8591 = ~n10253;
  assign n9245 = ~n10254;
  assign n9811 = ~n10255;
  assign n9047 = ~n10256;
  assign n8687 = ~n10257;
  assign n8633 = ~n10258;
  assign n8057 = ~n10259;
  assign n8173 = ~n10260;
  assign n9601 = ~n10261;
  assign n8713 = ~n10262;
  assign n9277 = ~n10263;
  assign n9415 = ~n10264;
  assign n9069 = ~n10265;
  assign n9071 = ~n10266;
  assign n8031 = ~n10267;
  assign n8331 = ~n10268;
  assign n9099 = ~n10269;
  assign n8153 = ~n10270;
  assign n8369 = ~n10271;
  assign n8949 = ~n10272;
  assign n9189 = ~n10273;
  assign n9529 = ~n10274;
  assign n8995 = ~n10275;
  assign n9861 = ~n10276;
  assign n9201 = ~n10277;
  assign n8971 = ~n10278;
  assign n9193 = ~n10279;
  assign n8311 = ~n10280;
  assign n8461 = ~n10281;
  assign n9829 = ~n10282;
  assign n8801 = ~n10283;
  assign n9527 = ~n10284;
  assign n9147 = ~n10285;
  assign n9219 = ~n10286;
  assign n8641 = ~n10287;
  assign n9303 = ~n10288;
  assign n8749 = ~n10289;
  assign n9307 = ~n10290;
  assign n8167 = ~n10291;
  assign n9221 = ~n10292;
  assign n9359 = ~n10293;
  assign n8575 = ~n10294;
  assign n9141 = ~n10295;
  assign n9079 = ~n10296;
  assign n9613 = ~n10297;
  assign n8397 = ~n10298;
  assign n9289 = ~n10299;
  assign n8915 = ~n10300;
  assign n8377 = ~n10301;
  assign n8585 = ~n10302;
  assign n8495 = ~n10303;
  assign n8209 = ~n10304;
  assign n9143 = ~n10305;
  assign n9333 = ~n10306;
  assign n6346 = n10307 & n7041;
  assign n9317 = ~n10308;
  assign n9661 = ~n10309;
  assign n8097 = ~n10310;
  assign n9807 = ~n10311;
  assign n9213 = ~n10312;
  assign n9287 = ~n10313;
  assign n8945 = ~n10314;
  assign n9217 = ~n10315;
  assign n8349 = ~n10316;
  assign n9793 = ~n10317;
  assign n8907 = ~n10318;
  assign n8511 = ~n10319;
  assign n8199 = ~n10320;
  assign n8053 = ~n10321;
  assign n8305 = ~n10322;
  assign n9279 = ~n10323;
  assign n9723 = ~n10324;
  assign n9285 = ~n10325;
  assign n9445 = ~n10326;
  assign n9111 = ~n10327;
  assign n9363 = ~n10328;
  assign n6270 = n10329 & n7049;
  assign n9385 = ~n10330;
  assign n8429 = ~n10331;
  assign n8045 = ~n10332;
  assign n9171 = ~n10333;
  assign n9405 = ~n10334;
  assign n8797 = ~n10335;
  assign n9777 = ~n10336;
  assign n9585 = ~n10337;
  assign n8041 = ~n10338;
  assign n9579 = ~n10339;
  assign n9503 = ~n10340;
  assign n8059 = ~n10341;
  assign n9813 = ~n10342;
  assign n9913 = ~n10343;
  assign n9185 = ~n10344;
  assign n9241 = ~n10345;
  assign n6428 = n10346 & n7061;
  assign n8087 = ~n10347;
  assign n9873 = ~n10348;
  assign n8189 = ~n10349;
  assign n9489 = ~n10350;
  assign n9931 = ~n10351;
  assign n9565 = ~n10352;
  assign n9013 = ~n10353;
  assign n9447 = ~n10354;
  assign n6236 = n10355 & n7055;
  assign n9093 = ~n10356;
  assign n8115 = ~n10357;
  assign n9709 = ~n10358;
  assign n9665 = ~n10359;
  assign n9469 = ~n10360;
  assign n8507 = ~n10361;
  assign n9539 = ~n10362;
  assign n9337 = ~n10363;
  assign n8427 = ~n10364;
  assign n9667 = ~n10365;
  assign n9535 = ~n10366;
  assign n8935 = ~n10367;
  assign n9721 = ~n10368;
  assign n8665 = ~n10369;
  assign n9377 = ~n10370;
  assign n6308 = n10371 & n7057;
  assign n9773 = ~n10372;
  assign n9741 = ~n10373;
  assign n8447 = ~n10374;
  assign n9575 = ~n10375;
  assign n8079 = ~n10376;
  assign n9765 = ~n10377;
  assign n9545 = ~n10378;
  assign n9757 = ~n10379;
  assign n8175 = ~n10380;
  assign n9181 = ~n10381;
  assign n6242 = n10382 & n7053;
  assign n9157 = ~n10383;
  assign n9521 = ~n10384;
  assign n9599 = ~n10385;
  assign n9395 = ~n10386;
  assign n9107 = ~n10387;
  assign n8693 = ~n10388;
  assign n8085 = ~n10389;
  assign n9631 = ~n10390;
  assign n9609 = ~n10391;
  assign n8839 = ~n10392;
  assign n8721 = ~n10393;
  assign n8881 = ~n10394;
  assign n8831 = ~n10395;
  assign n8775 = ~n10396;
  assign n9557 = ~n10397;
  assign n9543 = ~n10398;
  assign n8279 = ~n10399;
  assign n8827 = ~n10400;
  assign n8329 = ~n10401;
  assign n8653 = ~n10402;
  assign n9657 = ~n10403;
  assign n8341 = ~n10404;
  assign n9567 = ~n10405;
  assign n6294 = n10406 & n7043;
  assign n8017 = ~n10407;
  assign n9025 = ~n10408;
  assign n9916 = ~n10409;
  assign n9348 = ~n10410;
  assign n9110 = ~n10411;
  assign n8112 = ~n10412;
  assign n8236 = ~n10413;
  assign n8258 = ~n10414;
  assign n8920 = ~n10415;
  assign n8526 = ~n10416;
  assign n8600 = ~n10417;
  assign n9352 = ~n10418;
  assign n9064 = ~n10419;
  assign n9716 = ~n10420;
  assign n9628 = ~n10421;
  assign n9312 = ~n10422;
  assign n8452 = ~n10423;
  assign n8505 = ~n10424;
  assign n9161 = ~n10425;
  assign n9885 = ~n10426;
  assign n8345 = ~n10427;
  assign n9203 = ~n10428;
  assign n9259 = ~n10429;
  assign n8037 = ~n10430;
  assign n8245 = ~n10431;
  assign n8769 = ~n10432;
  assign n9847 = ~n10433;
  assign n8735 = ~n10434;
  assign n9735 = ~n10435;
  assign n9043 = ~n10436;
  assign n8241 = ~n10437;
  assign n9085 = ~n10438;
  assign n9729 = ~n10439;
  assign n9149 = ~n10440;
  assign n9927 = ~n10441;
  assign n8415 = ~n10442;
  assign n8933 = ~n10443;
  assign n8463 = ~n10444;
  assign n9059 = ~n10445;
  assign n9207 = ~n10446;
  assign n9137 = ~n10447;
  assign n9507 = ~n10448;
  assign n9457 = ~n10449;
  assign n8697 = ~n10450;
  assign n8333 = ~n10451;
  assign n9517 = ~n10452;
  assign n9475 = ~n10453;
  assign n8761 = ~n10454;
  assign n8731 = ~n10455;
  assign n8913 = ~n10456;
  assign n9283 = ~n10457;
  assign n8033 = ~n10458;
  assign n8719 = ~n10459;
  assign n8051 = ~n10460;
  assign n9257 = ~n10461;
  assign n8301 = ~n10462;
  assign n8493 = ~n10463;
  assign n9265 = ~n10464;
  assign n9833 = ~n10465;
  assign n8639 = ~n10466;
  assign n9725 = ~n10467;
  assign n8127 = ~n10468;
  assign n8339 = ~n10469;
  assign n8785 = ~n10470;
  assign n8479 = ~n10471;
  assign n9841 = ~n10472;
  assign n9753 = ~n10473;
  assign n9791 = ~n10474;
  assign n8595 = ~n10475;
  assign n9449 = ~n10476;
  assign n8825 = ~n10477;
  assign n8207 = ~n10478;
  assign n8599 = ~n10479;
  assign n9323 = ~n10480;
  assign n9513 = ~n10481;
  assign n9033 = ~n10482;
  assign n9281 = ~n10483;
  assign n8093 = ~n10484;
  assign n9091 = ~n10485;
  assign n9779 = ~n10486;
  assign n9869 = ~n10487;
  assign n9467 = ~n10488;
  assign n8905 = ~n10489;
  assign n9383 = ~n10490;
  assign n8095 = ~n10491;
  assign n9919 = ~n10492;
  assign n9351 = ~n10493;
  assign n9393 = ~n10494;
  assign n9569 = ~n10495;
  assign n9311 = ~n10496;
  assign n8647 = ~n10497;
  assign n9559 = ~n10498;
  assign n8571 = ~n10499;
  assign n9459 = ~n10500;
  assign n9205 = ~n10501;
  assign n8491 = ~n10502;
  assign n8291 = ~n10503;
  assign n9523 = ~n10504;
  assign n9195 = ~n10505;
  assign n8701 = ~n10506;
  assign n8081 = ~n10507;
  assign n8029 = ~n10508;
  assign n9009 = ~n10509;
  assign n9321 = ~n10510;
  assign n9839 = ~n10511;
  assign n9651 = ~n10512;
  assign n9295 = ~n10513;
  assign n9261 = ~n10514;
  assign n8317 = ~n10515;
  assign n9495 = ~n10516;
  assign n8669 = ~n10517;
  assign n8833 = ~n10518;
  assign n8519 = ~n10519;
  assign n9887 = ~n10520;
  assign n8283 = ~n10521;
  assign n8065 = ~n10522;
  assign n8451 = ~n10523;
  assign n8589 = ~n10524;
  assign n9409 = ~n10525;
  assign n8071 = ~n10526;
  assign n8119 = ~n10527;
  assign n9329 = ~n10528;
  assign n8043 = ~n10529;
  assign n9855 = ~n10530;
  assign n9373 = ~n10531;
  assign n8683 = ~n10532;
  assign n9263 = ~n10533;
  assign n8113 = ~n10534;
  assign n8099 = ~n10535;
  assign n8955 = ~n10536;
  assign n9781 = ~n10537;
  assign n8927 = ~n10538;
  assign n9105 = ~n10539;
  assign n8535 = ~n10540;
  assign n9117 = ~n10541;
  assign n8111 = ~n10542;
  assign n8131 = ~n10543;
  assign n8611 = ~n10544;
  assign n9327 = ~n10545;
  assign n8139 = ~n10546;
  assign n8211 = ~n10547;
  assign n9139 = ~n10548;
  assign n9737 = ~n10549;
  assign n8379 = ~n10550;
  assign n9177 = ~n10551;
  assign n8157 = ~n10552;
  assign n8883 = ~n10553;
  assign n8075 = ~n10554;
  assign n8183 = ~n10555;
  assign n9343 = ~n10556;
  assign n8145 = ~n10557;
  assign n8179 = ~n10558;
  assign n8281 = ~n10559;
  assign n8193 = ~n10560;
  assign n8025 = ~n10561;
  assign n9169 = ~n10562;
  assign n8217 = ~n10563;
  assign n8219 = ~n10564;
  assign n8325 = ~n10565;
  assign n9909 = ~n10566;
  assign n8235 = ~n10567;
  assign n8547 = ~n10568;
  assign n8885 = ~n10569;
  assign n8353 = ~n10570;
  assign n8263 = ~n10571;
  assign n8385 = ~n10572;
  assign n9239 = ~n10573;
  assign n9045 = ~n10574;
  assign n8313 = ~n10575;
  assign n8289 = ~n10576;
  assign n9011 = ~n10577;
  assign n9473 = ~n10578;
  assign n8307 = ~n10579;
  assign n8999 = ~n10580;
  assign n8315 = ~n10581;
  assign n9933 = ~n10582;
  assign n9785 = ~n10583;
  assign n8309 = ~n10584;
  assign n9597 = ~n10585;
  assign n9625 = ~n10586;
  assign n8399 = ~n10587;
  assign n8267 = ~n10588;
  assign n8357 = ~n10589;
  assign n8395 = ~n10590;
  assign n8177 = ~n10591;
  assign n8631 = ~n10592;
  assign n8371 = ~n10593;
  assign n8689 = ~n10594;
  assign n9397 = ~n10595;
  assign n9759 = ~n10596;
  assign n9481 = ~n10597;
  assign n9659 = ~n10598;
  assign n8777 = ~n10599;
  assign n9347 = ~n10600;
  assign n9401 = ~n10601;
  assign n8389 = ~n10602;
  assign n8243 = ~n10603;
  assign n8405 = ~n10604;
  assign n9923 = ~n10605;
  assign n9421 = ~n10606;
  assign n8807 = ~n10607;
  assign n8621 = ~n10608;
  assign n8425 = ~n10609;
  assign n8673 = ~n10610;
  assign n8435 = ~n10611;
  assign n9641 = ~n10612;
  assign n9803 = ~n10613;
  assign n9233 = ~n10614;
  assign n9031 = ~n10615;
  assign n9163 = ~n10616;
  assign n8299 = ~n10617;
  assign n8453 = ~n10618;
  assign n8759 = ~n10619;
  assign n9425 = ~n10620;
  assign n9915 = ~n10621;
  assign n9209 = ~n10622;
  assign n8475 = ~n10623;
  assign n8793 = ~n10624;
  assign n8771 = ~n10625;
  assign n8483 = ~n10626;
  assign n9037 = ~n10627;
  assign n9883 = ~n10628;
  assign n8823 = ~n10629;
  assign n8961 = ~n10630;
  assign n8509 = ~n10631;
  assign n9387 = ~n10632;
  assign n9493 = ~n10633;
  assign n8645 = ~n10634;
  assign n9857 = ~n10635;
  assign n8477 = ~n10636;
  assign n8549 = ~n10637;
  assign n9119 = ~n10638;
  assign n8751 = ~n10639;
  assign n8501 = ~n10640;
  assign n8387 = ~n10641;
  assign n8551 = ~n10642;
  assign n8559 = ~n10643;
  assign n8893 = ~n10644;
  assign n8859 = ~n10645;
  assign n8921 = ~n10646;
  assign n8171 = ~n10647;
  assign n8699 = ~n10648;
  assign n9019 = ~n10649;
  assign n9629 = ~n10650;
  assign n8607 = ~n10651;
  assign n8417 = ~n10652;
  assign n8229 = ~n10653;
  assign n8069 = ~n10654;
  assign n8433 = ~n10655;
  assign n9041 = ~n10656;
  assign n9937 = ~n10657;
  assign n8925 = ~n10658;
  assign n8667 = ~n10659;
  assign n9617 = ~n10660;
  assign n9477 = ~n10661;
  assign n8013 = ~n10662;
  assign n8677 = ~n10663;
  assign n9403 = ~n10664;
  assign n8651 = ~n10665;
  assign n8649 = ~n10666;
  assign n8489 = ~n10667;
  assign n9225 = ~n10668;
  assign n9583 = ~n10669;
  assign n9389 = ~n10670;
  assign n8335 = ~n10671;
  assign n8671 = ~n10672;
  assign n8675 = ~n10673;
  assign n9023 = ~n10674;
  assign n8271 = ~n10675;
  assign n9821 = ~n10676;
  assign n8541 = ~n10677;
  assign n8705 = ~n10678;
  assign n8869 = ~n10679;
  assign n8561 = ~n10680;
  assign n8073 = ~n10681;
  assign n8991 = ~n10682;
  assign n9615 = ~n10683;
  assign n8865 = ~n10684;
  assign n8007 = ~n10685;
  assign n8729 = ~n10686;
  assign n9509 = ~n10687;
  assign n9057 = ~n10688;
  assign n9835 = ~n10689;
  assign n9531 = ~n10690;
  assign n8465 = ~n10691;
  assign n8381 = ~n10692;
  assign n9371 = ~n10693;
  assign n9505 = ~n10694;
  assign n9563 = ~n10695;
  assign n8707 = ~n10696;
  assign n8967 = ~n10697;
  assign n9771 = ~n10698;
  assign n9663 = ~n10699;
  assign n9027 = ~n10700;
  assign n8835 = ~n10701;
  assign n9325 = ~n10702;
  assign n9015 = ~n10703;
  assign n9341 = ~n10704;
  assign n8293 = ~n10705;
  assign n8805 = ~n10706;
  assign n8583 = ~n10707;
  assign n8817 = ~n10708;
  assign n9077 = ~n10709;
  assign n8819 = ~n10710;
  assign n8975 = ~n10711;
  assign n9775 = ~n10712;
  assign n8773 = ~n10713;
  assign n9715 = ~n10714;
  assign n8851 = ~n10715;
  assign n9127 = ~n10716;
  assign n8853 = ~n10717;
  assign n8993 = ~n10718;
  assign n8861 = ~n10719;
  assign n9867 = ~n10720;
  assign n9407 = ~n10721;
  assign n8875 = ~n10722;
  assign n8957 = ~n10723;
  assign n8237 = ~n10724;
  assign n8125 = ~n10725;
  assign n8513 = ~n10726;
  assign n8215 = ~n10727;
  assign n8449 = ~n10728;
  assign n9921 = ~n10729;
  assign n8587 = ~n10730;
  assign n8919 = ~n10731;
  assign n8943 = ~n10732;
  assign n9381 = ~n10733;
  assign n9871 = ~n10734;
  assign n9291 = ~n10735;
  assign n8233 = ~n10736;
  assign n9849 = ~n10737;
  assign n8593 = ~n10738;
  assign n8227 = ~n10739;
  assign n9547 = ~n10740;
  assign n8347 = ~n10741;
  assign n9817 = ~n10742;
  assign n8077 = ~n10743;
  assign n8155 = ~n10744;
  assign n9029 = ~n10745;
  assign n9635 = ~n10746;
  assign n8899 = ~n10747;
  assign n9053 = ~n10748;
  assign n9231 = ~n10749;
  assign n8739 = ~n10750;
  assign n9823 = ~n10751;
  assign n9297 = ~n10752;
  assign n9235 = ~n10753;
  assign n8391 = ~n10754;
  assign n9083 = ~n10755;
  assign n9751 = ~n10756;
  assign n8223 = ~n10757;
  assign n8659 = ~n10758;
  assign n8857 = ~n10759;
  assign n9275 = ~n10760;
  assign n9607 = ~n10761;
  assign n9863 = ~n10762;
  assign n8879 = ~n10763;
  assign n9589 = ~n10764;
  assign n9255 = ~n10765;
  assign n8409 = ~n10766;
  assign n9073 = ~n10767;
  assign n9113 = ~n10768;
  assign n8135 = ~n10769;
  assign n9153 = ~n10770;
  assign n9101 = ~n10771;
  assign n8195 = ~n10772;
  assign n8887 = ~n10773;
  assign n9055 = ~n10774;
  assign n9223 = ~n10775;
  assign n9063 = ~n10776;
  assign n9581 = ~n10777;
  assign n9431 = ~n10778;
  assign n8779 = ~n10779;
  assign n9215 = ~n10780;
  assign n9827 = ~n10781;
  assign n9471 = ~n10782;
  assign n9783 = ~n10783;
  assign n9743 = ~n10784;
  assign n9643 = ~n10785;
  assign n8363 = ~n10786;
  assign n9103 = ~n10787;
  assign n8107 = ~n10788;
  assign n8579 = ~n10789;
  assign n9249 = ~n10790;
  assign n9253 = ~n10791;
  assign n9345 = ~n10792;
  assign n8545 = ~n10793;
  assign n9763 = ~n10794;
  assign n8623 = ~n10795;
  assign n8121 = ~n10796;
  assign n8947 = ~n10797;
  assign n9109 = ~n10798;
  assign n9271 = ~n10799;
  assign n9293 = ~n10800;
  assign n9391 = ~n10801;
  assign n8765 = ~n10802;
  assign n9491 = ~n10803;
  assign n9655 = ~n10804;
  assign n8783 = ~n10805;
  assign n9097 = ~n10806;
  assign n9367 = ~n10807;
  assign n8201 = ~n10808;
  assign n9435 = ~n10809;
  assign n9065 = ~n10810;
  assign n9731 = ~n10811;
  assign n8989 = ~n10812;
  assign n9929 = ~n10813;
  assign n9837 = ~n10814;
  assign n9917 = ~n10815;
  assign n8525 = ~n10816;
  assign n8123 = ~n10817;
  assign n8083 = ~n10818;
  assign n9483 = ~n10819;
  assign n8361 = ~n10820;
  assign n9797 = ~n10821;
  assign n8443 = ~n10822;
  assign n8555 = ~n10823;
  assign n8799 = ~n10824;
  assign n9463 = ~n10825;
  assign n9497 = ~n10826;
  assign n8343 = ~n10827;
  assign n9411 = ~n10828;
  assign n9135 = ~n10829;
  assign n9417 = ~n10830;
  assign n8523 = ~n10831;
  assign n9789 = ~n10832;
  assign n8191 = ~n10833;
  assign n8257 = ~n10834;
  assign n8983 = ~n10835;
  assign n8149 = ~n10836;
  assign n8487 = ~n10837;
  assign n9273 = ~n10838;
  assign n8185 = ~n10839;
  assign n9799 = ~n10840;
  assign n9487 = ~n10841;
  assign n8781 = ~n10842;
  assign n9891 = ~n10843;
  assign n9645 = ~n10844;
  assign n8979 = ~n10845;
  assign n9243 = ~n10846;
  assign n8969 = ~n10847;
  assign n8745 = ~n10848;
  assign n9577 = ~n10849;
  assign n9819 = ~n10850;
  assign n9131 = ~n10851;
  assign n8803 = ~n10852;
  assign n8221 = ~n10853;
  assign n9331 = ~n10854;
  assign n9361 = ~n10855;
  assign n9739 = ~n10856;
  assign n8757 = ~n10857;
  assign n8985 = ~n10858;
  assign n9845 = ~n10859;
  assign n9229 = ~n10860;
  assign n8939 = ~n10861;
  assign n9183 = ~n10862;
  assign n8845 = ~n10863;
  assign n9439 = ~n10864;
  assign n9541 = ~n10865;
  assign n8795 = ~n10866;
  assign n8527 = ~n10867;
  assign n8601 = ~n10868;
  assign n9881 = ~n10869;
  assign n9899 = ~n10870;
  assign n9511 = ~n10871;
  assign n9767 = ~n10872;
  assign n8873 = ~n10873;
  assign n9561 = ~n10874;
  assign n9637 = ~n10875;
  assign n9889 = ~n10876;
  assign n9647 = ~n10877;
  assign n9499 = ~n10878;
  assign n9711 = ~n10879;
  assign n8841 = ~n10880;
  assign n9427 = ~n10881;
  assign n9191 = ~n10882;
  assign n9605 = ~n10883;
  assign n9155 = ~n10884;
  assign n8411 = ~n10885;
  assign n9305 = ~n10886;
  assign n9925 = ~n10887;
  assign n9627 = ~n10888;
  assign n9603 = ~n10889;
  assign n8791 = ~n10890;
  assign n9537 = ~n10891;
  assign n8723 = ~n10892;
  assign n9649 = ~n10893;
  assign n9319 = ~n10894;
  assign n8565 = ~n10895;
  assign n9591 = ~n10896;
  assign n8499 = ~n10897;
  assign n9893 = ~n10898;
  assign n9087 = ~n10899;
  assign n6064 = n10228 ^ n10900;
  assign n8517 = ~n10902;
  assign n9159 = ~n10903;
  assign n9335 = ~n10905;
  assign n8727 = ~n10906;
  assign n8681 = ~n10907;
  assign n9021 = ~n10910;
  assign n9355 = ~n10912;
  assign n8101 = ~n10913;
  assign n8533 = ~n10914;
  assign n9379 = ~n10915;
  assign n8603 = ~n10917;
  assign n8837 = ~n10918;
  assign n8039 = ~n10919;
  assign n8471 = ~n10921;
  assign n8753 = ~n10923;
  assign n8103 = ~n10926;
  assign n8997 = ~n10927;
  assign n8539 = ~n10930;
  assign n9051 = ~n10931;
  assign n8269 = ~n10932;
  assign n9049 = ~n10933;
  assign n8637 = ~n10934;
  assign n8615 = ~n10936;
  assign n8355 = ~n10937;
  assign n9749 = ~n10938;
  assign n8203 = ~n10939;
  assign n8619 = ~n10940;
  assign n8573 = ~n10941;
  assign n9095 = ~n10943;
  assign n8485 = ~n10944;
  assign n8439 = ~n10945;
  assign n6368 = n10982 & n10983;
  assign n6232 = n10984 & n10985;
  assign n5004 = n11008 & n11009;
  assign n7978 = n11010 & n11011;
  assign n9949 = n11015 & n11016;
  assign n5132 = n11017 & n11018;
  assign n9675 = n11019 & n11020;
  assign n6326 = n11021 & n11022;
  assign n5088 = n11023 & n11024;
  assign n9673 = n11025 & n11026;
  assign n7988 = n11027 & n11028;
  assign n9717 = n11029 & n11030;
  assign n4996 = n11031 & n11032;
  assign n6278 = n11033 & n11034;
  assign n7984 = n11035 & n11036;
  assign n6332 = n11037 & n11038;
  assign n9669 = n11039 & n11040;
  assign n9671 = n11041 & n11042;
  assign n5142 = n11043 & n11044;
  assign n7982 = n11045 & n11046;
  assign n7986 = n11047 & n11048;
  assign n6244 = n11049 & n11050;
  assign n9963 = n11051 & n11052;
  assign n9187 = n11053 & n11054;
  assign n7999 = n11055 & n11056;
  assign n5187 = n11057 & n11058;
  assign n8003 = n11059 & n11060;
  assign n8001 = n11061 & n11062;
  assign n9720 = n11063 & n11064;
  assign n10901 = n10900 & n11065;
  assign n5219 = n11066 & n11067;
  assign n7980 = n11068 & n11069;
  assign n10922 = n11070 & n11071;
  assign n10942 = n11072 & n11073;
  assign n10908 = n11074 & n11075;
  assign n10911 = n11076 & n11077;
  assign n10929 = n11078 & n11079;
  assign n10925 = n11082 & n11083;
  assign n10904 = n11084 & n11085;
  assign n10916 = n11086 & n11087;
  assign n9957 = n11088 & n11089;
  assign n10935 = n11090 & n11091;
  assign n10928 = n11092 & n11093;
  assign n10924 = n11094 & n11095;
  assign n10227 = ~n10900;
  assign n10920 = n11096 & n11097;
  assign n10909 = n11098 & n11099;
  assign n10098 = n11100 & n11101;
  assign n6954 = n8004 & n63;
  assign n7112 = n8007 & n8008;
  assign n7121 = n8009 & n8010;
  assign n7129 = n8011 & n8012;
  assign n7168 = n8013 & n8014;
  assign n7255 = n8015 & n8016;
  assign n7123 = n8017 & n8018;
  assign n7141 = n8019 & n8020;
  assign n7125 = n8021 & n8022;
  assign n7664 = n8023 & n8024;
  assign n7952 = n8025 & n8026;
  assign n7103 = n8027 & n8028;
  assign n7742 = n8029 & n8030;
  assign n7356 = n8031 & n8032;
  assign n7350 = n8033 & n8034;
  assign n7357 = n8035 & n8036;
  assign n7119 = n8037 & n8038;
  assign n7164 = n8039 & n8040;
  assign n7945 = n8041 & n8042;
  assign n7128 = n8043 & n8044;
  assign n7169 = n8045 & n8046;
  assign n7139 = n8047 & n8048;
  assign n7165 = n8049 & n8050;
  assign n7920 = n8051 & n8052;
  assign n7349 = n8053 & n8054;
  assign n7185 = n8055 & n8056;
  assign n7133 = n8057 & n8058;
  assign n7709 = n8059 & n8060;
  assign n7939 = n8061 & n8062;
  assign n7155 = n8063 & n8064;
  assign n7160 = n8065 & n8066;
  assign n7581 = n8067 & n8068;
  assign n7450 = n8069 & n8070;
  assign n7700 = n8071 & n8072;
  assign n7162 = n8073 & n8074;
  assign n7210 = n8075 & n8076;
  assign n7150 = n8077 & n8078;
  assign n7953 = n8079 & n8080;
  assign n7108 = n8081 & n8082;
  assign n7796 = n8083 & n8084;
  assign n7615 = n8085 & n8086;
  assign n7531 = n8087 & n8088;
  assign n7515 = n8089 & n8090;
  assign n7663 = n8091 & n8092;
  assign n7748 = n8093 & n8094;
  assign n7092 = n8095 & n8096;
  assign n7175 = n8097 & n8098;
  assign n7138 = n8099 & n8100;
  assign n7130 = n8101 & n8102;
  assign n7174 = n8103 & n8104;
  assign n7179 = n8105 & n8106;
  assign n7470 = n8107 & n8108;
  assign n7181 = n8109 & n8110;
  assign n7046 = n8111 & n8112;
  assign n7180 = n8113 & n8114;
  assign n7843 = n8115 & n8116;
  assign n7183 = n8117 & n8118;
  assign n7468 = n8119 & n8120;
  assign n7194 = n8121 & n8122;
  assign n7936 = n8123 & n8124;
  assign n7182 = n8125 & n8126;
  assign n7708 = n8127 & n8128;
  assign n7189 = n8129 & n8130;
  assign n7188 = n8131 & n8132;
  assign n7191 = n8133 & n8134;
  assign n7190 = n8135 & n8136;
  assign n7193 = n8137 & n8138;
  assign n7192 = n8139 & n8140;
  assign n7196 = n8141 & n8142;
  assign n7201 = n8143 & n8144;
  assign n7200 = n8145 & n8146;
  assign n7205 = n8147 & n8148;
  assign n7684 = n8149 & n8150;
  assign n7207 = n8151 & n8152;
  assign n7307 = n8153 & n8154;
  assign n7950 = n8155 & n8156;
  assign n7206 = n8157 & n8158;
  assign n7642 = n8159 & n8160;
  assign n7211 = n8161 & n8162;
  assign n7265 = n8163 & n8164;
  assign n7267 = n8165 & n8166;
  assign n7741 = n8167 & n8168;
  assign n7965 = n8169 & n8170;
  assign n7482 = n8171 & n8172;
  assign n7177 = n8173 & n8174;
  assign n7217 = n8175 & n8176;
  assign n7362 = n8177 & n8178;
  assign n7216 = n8179 & n8180;
  assign n7229 = n8181 & n8182;
  assign n7224 = n8183 & n8184;
  assign n7228 = n8185 & n8186;
  assign n7227 = n8187 & n8188;
  assign n7231 = n8189 & n8190;
  assign n7230 = n8191 & n8192;
  assign n7226 = n8193 & n8194;
  assign n7678 = n8195 & n8196;
  assign n7681 = n8197 & n8198;
  assign n7235 = n8199 & n8200;
  assign n7234 = n8201 & n8202;
  assign n7233 = n8203 & n8204;
  assign n7363 = n8205 & n8206;
  assign n7232 = n8207 & n8208;
  assign n7239 = n8209 & n8210;
  assign n7236 = n8211 & n8212;
  assign n7241 = n8213 & n8214;
  assign n7212 = n8215 & n8216;
  assign n7240 = n8217 & n8218;
  assign n7242 = n8219 & n8220;
  assign n7882 = n8221 & n8222;
  assign n7680 = n8223 & n8224;
  assign n7245 = n8225 & n8226;
  assign n7244 = n8227 & n8228;
  assign n7446 = n8229 & n8230;
  assign n7247 = n8231 & n8232;
  assign n7246 = n8233 & n8234;
  assign n7050 = n8235 & n8236;
  assign n7252 = n8237 & n8238;
  assign n7439 = n8239 & n8240;
  assign n7759 = n8241 & n8242;
  assign n7830 = n8243 & n8244;
  assign n7323 = n8245 & n8246;
  assign n7643 = n8247 & n8248;
  assign n7857 = n8249 & n8250;
  assign n7929 = n8251 & n8252;
  assign n7921 = n8253 & n8254;
  assign n7257 = n8255 & n8256;
  assign n7048 = n8257 & n8258;
  assign n7259 = n8259 & n8260;
  assign n7943 = n8261 & n8262;
  assign n7256 = n8263 & n8264;
  assign n7383 = n8265 & n8266;
  assign n7258 = n8267 & n8268;
  assign n7261 = n8269 & n8270;
  assign n7486 = n8271 & n8272;
  assign n7823 = n8273 & n8274;
  assign n7489 = n8275 & n8276;
  assign n7713 = n8277 & n8278;
  assign n7263 = n8279 & n8280;
  assign n7126 = n8281 & n8282;
  assign n7266 = n8283 & n8284;
  assign n7199 = n8285 & n8286;
  assign n7269 = n8287 & n8288;
  assign n7264 = n8289 & n8290;
  assign n7268 = n8291 & n8292;
  assign n7880 = n8293 & n8294;
  assign n7271 = n8295 & n8296;
  assign n7273 = n8297 & n8298;
  assign n7270 = n8299 & n8300;
  assign n7272 = n8301 & n8302;
  assign n7651 = n8303 & n8304;
  assign n7275 = n8305 & n8306;
  assign n7274 = n8307 & n8308;
  assign n7198 = n8309 & n8310;
  assign n7277 = n8311 & n8312;
  assign n7276 = n8313 & n8314;
  assign n7278 = n8315 & n8316;
  assign n7871 = n8317 & n8318;
  assign n7281 = n8319 & n8320;
  assign n7280 = n8321 & n8322;
  assign n7285 = n8323 & n8324;
  assign n7284 = n8325 & n8326;
  assign n7283 = n8327 & n8328;
  assign n7289 = n8329 & n8330;
  assign n7675 = n8331 & n8332;
  assign n7186 = n8333 & n8334;
  assign n7288 = n8335 & n8336;
  assign n7401 = n8337 & n8338;
  assign n7290 = n8339 & n8340;
  assign n7447 = n8341 & n8342;
  assign n7728 = n8343 & n8344;
  assign n7969 = n8345 & n8346;
  assign n7286 = n8347 & n8348;
  assign n7293 = n8349 & n8350;
  assign n7099 = n8351 & n8352;
  assign n7314 = n8353 & n8354;
  assign n7295 = n8355 & n8356;
  assign n7294 = n8357 & n8358;
  assign n7865 = n8359 & n8360;
  assign n7592 = n8361 & n8362;
  assign n7296 = n8363 & n8364;
  assign n7299 = n8365 & n8366;
  assign n7298 = n8367 & n8368;
  assign n7301 = n8369 & n8370;
  assign n7300 = n8371 & n8372;
  assign n7303 = n8373 & n8374;
  assign n7305 = n8375 & n8376;
  assign n7755 = n8377 & n8378;
  assign n7204 = n8379 & n8380;
  assign n7304 = n8381 & n8382;
  assign n7407 = n8383 & n8384;
  assign n7260 = n8385 & n8386;
  assign n7396 = n8387 & n8388;
  assign n7302 = n8389 & n8390;
  assign n7586 = n8391 & n8392;
  assign n7107 = n8393 & n8394;
  assign n7480 = n8395 & n8396;
  assign n7315 = n8397 & n8398;
  assign n7262 = n8399 & n8400;
  assign n7319 = n8401 & n8402;
  assign n7641 = n8403 & n8404;
  assign n7316 = n8405 & n8406;
  assign n7321 = n8407 & n8408;
  assign n7318 = n8409 & n8410;
  assign n7322 = n8411 & n8412;
  assign n7325 = n8413 & n8414;
  assign n7320 = n8415 & n8416;
  assign n7222 = n8417 & n8418;
  assign n7313 = n8419 & n8420;
  assign n7327 = n8421 & n8422;
  assign n7471 = n8423 & n8424;
  assign n7326 = n8425 & n8426;
  assign n7855 = n8427 & n8428;
  assign n7333 = n8429 & n8430;
  assign n7673 = n8431 & n8432;
  assign n7154 = n8433 & n8434;
  assign n7332 = n8435 & n8436;
  assign n7339 = n8437 & n8438;
  assign n7541 = n8439 & n8440;
  assign n7151 = n8441 & n8442;
  assign n7340 = n8443 & n8444;
  assign n7877 = n8445 & n8446;
  assign n7345 = n8447 & n8448;
  assign n7662 = n8449 & n8450;
  assign n7044 = n8451 & n8452;
  assign n7344 = n8453 & n8454;
  assign n7035 = n8455 & n8456;
  assign n7077 = n8457 & n8458;
  assign n7347 = n8459 & n8460;
  assign n7093 = n8461 & n8462;
  assign n7166 = n8463 & n8464;
  assign n7156 = n8465 & n8466;
  assign n7359 = n8467 & n8468;
  assign n7377 = n8469 & n8470;
  assign n7113 = n8471 & n8472;
  assign n7361 = n8473 & n8474;
  assign n7360 = n8475 & n8476;
  assign n7774 = n8477 & n8478;
  assign n7358 = n8479 & n8480;
  assign n7365 = n8481 & n8482;
  assign n7364 = n8483 & n8484;
  assign n7367 = n8485 & n8486;
  assign n7366 = n8487 & n8488;
  assign n7782 = n8489 & n8490;
  assign n7820 = n8491 & n8492;
  assign n7368 = n8493 & n8494;
  assign n7753 = n8495 & n8496;
  assign n7371 = n8497 & n8498;
  assign n7370 = n8499 & n8500;
  assign n7330 = n8501 & n8502;
  assign n7029 = n8503 & n8504;
  assign n7343 = n8505 & n8506;
  assign n7373 = n8507 & n8508;
  assign n7372 = n8509 & n8510;
  assign n7781 = n8511 & n8512;
  assign n7378 = n8513 & n8514;
  assign n7381 = n8515 & n8516;
  assign n7380 = n8517 & n8518;
  assign n7382 = n8519 & n8520;
  assign n7413 = n8521 & n8522;
  assign n7136 = n8523 & n8524;
  assign n7052 = n8525 & n8526;
  assign n7388 = n8527 & n8528;
  assign n7385 = n8529 & n8530;
  assign n7161 = n8531 & n8532;
  assign n7393 = n8533 & n8534;
  assign n7392 = n8535 & n8536;
  assign n7785 = n8537 & n8538;
  assign n7397 = n8539 & n8540;
  assign n7398 = n8541 & n8542;
  assign n7403 = n8543 & n8544;
  assign n7394 = n8545 & n8546;
  assign n7402 = n8547 & n8548;
  assign n7384 = n8549 & n8550;
  assign n7400 = n8551 & n8552;
  assign n7409 = n8553 & n8554;
  assign n7408 = n8555 & n8556;
  assign n7411 = n8557 & n8558;
  assign n7410 = n8559 & n8560;
  assign n7412 = n8561 & n8562;
  assign n7415 = n8563 & n8564;
  assign n7414 = n8565 & n8566;
  assign n7417 = n8567 & n8568;
  assign n7419 = n8569 & n8570;
  assign n7416 = n8571 & n8572;
  assign n7421 = n8573 & n8574;
  assign n7839 = n8575 & n8576;
  assign n7197 = n8577 & n8578;
  assign n7420 = n8579 & n8580;
  assign n7423 = n8581 & n8582;
  assign n7840 = n8583 & n8584;
  assign n7429 = n8585 & n8586;
  assign n7430 = n8587 & n8588;
  assign n7484 = n8589 & n8590;
  assign n7433 = n8591 & n8592;
  assign n7432 = n8593 & n8594;
  assign n7435 = n8595 & n8596;
  assign n7441 = n8597 & n8598;
  assign n7054 = n8599 & n8600;
  assign n7440 = n8601 & n8602;
  assign n7434 = n8603 & n8604;
  assign n7443 = n8605 & n8606;
  assign n7442 = n8607 & n8608;
  assign n7223 = n8609 & n8610;
  assign n7070 = n8611 & n8612;
  assign n7445 = n8613 & n8614;
  assign n7444 = n8615 & n8616;
  assign n7014 = n8617 & n8618;
  assign n7453 = n8619 & n8620;
  assign n7686 = n8621 & n8622;
  assign n7452 = n8623 & n8624;
  assign n7455 = n8625 & n8626;
  assign n7767 = n8627 & n8628;
  assign n7143 = n8629 & n8630;
  assign n7454 = n8631 & n8632;
  assign n7677 = n8633 & n8634;
  assign n7153 = n8635 & n8636;
  assign n7481 = n8637 & n8638;
  assign n7504 = n8639 & n8640;
  assign n7849 = n8641 & n8642;
  assign n7337 = n8643 & n8644;
  assign n7566 = n8645 & n8646;
  assign n7427 = n8647 & n8648;
  assign n7848 = n8649 & n8650;
  assign n7460 = n8651 & n8652;
  assign n7317 = n8653 & n8654;
  assign n7463 = n8655 & n8656;
  assign n7729 = n8657 & n8658;
  assign n7462 = n8659 & n8660;
  assign n7477 = n8661 & n8662;
  assign n7783 = n8663 & n8664;
  assign n7963 = n8665 & n8666;
  assign n7456 = n8667 & n8668;
  assign n7110 = n8669 & n8670;
  assign n7466 = n8671 & n8672;
  assign n7102 = n8673 & n8674;
  assign n7464 = n8675 & n8676;
  assign n7152 = n8677 & n8678;
  assign n7473 = n8679 & n8680;
  assign n7472 = n8681 & n8682;
  assign n7406 = n8683 & n8684;
  assign n7479 = n8685 & n8686;
  assign n7485 = n8687 & n8688;
  assign n7478 = n8689 & n8690;
  assign n7487 = n8691 & n8692;
  assign n7495 = n8693 & n8694;
  assign n7311 = n8695 & n8696;
  assign n7488 = n8697 & n8698;
  assign n7644 = n8699 & n8700;
  assign n7310 = n8701 & n8702;
  assign n7491 = n8703 & n8704;
  assign n7490 = n8705 & n8706;
  assign n7542 = n8707 & n8708;
  assign n7505 = n8709 & n8710;
  assign n7567 = n8711 & n8712;
  assign n7497 = n8713 & n8714;
  assign n7499 = n8715 & n8716;
  assign n7087 = n8717 & n8718;
  assign n7498 = n8719 & n8720;
  assign n7501 = n8721 & n8722;
  assign n7500 = n8723 & n8724;
  assign n7253 = n8725 & n8726;
  assign n7379 = n8727 & n8728;
  assign n7930 = n8729 & n8730;
  assign n7502 = n8731 & n8732;
  assign n7507 = n8733 & n8734;
  assign n7569 = n8735 & n8736;
  assign n7583 = n8737 & n8738;
  assign n7494 = n8739 & n8740;
  assign n7511 = n8741 & n8742;
  assign n7509 = n8743 & n8744;
  assign n7510 = n8745 & n8746;
  assign n7127 = n8747 & n8748;
  assign n7513 = n8749 & n8750;
  assign n7512 = n8751 & n8752;
  assign n7508 = n8753 & n8754;
  assign n7517 = n8755 & n8756;
  assign n7892 = n8757 & n8758;
  assign n7516 = n8759 & n8760;
  assign n7028 = n8761 & n8762;
  assign n7020 = n8763 & n8764;
  assign n7600 = n8765 & n8766;
  assign n7519 = n8767 & n8768;
  assign n7775 = n8769 & n8770;
  assign n7376 = n8771 & n8772;
  assign n7606 = n8773 & n8774;
  assign n7607 = n8775 & n8776;
  assign n7616 = n8777 & n8778;
  assign n7724 = n8779 & n8780;
  assign n7730 = n8781 & n8782;
  assign n7080 = n8783 & n8784;
  assign n7948 = n8785 & n8786;
  assign n7749 = n8787 & n8788;
  assign n7545 = n8789 & n8790;
  assign n7202 = n8791 & n8792;
  assign n7248 = n8793 & n8794;
  assign n7522 = n8795 & n8796;
  assign n7525 = n8797 & n8798;
  assign n7864 = n8799 & n8800;
  assign n7115 = n8801 & n8802;
  assign n7524 = n8803 & n8804;
  assign n7528 = n8805 & n8806;
  assign n7926 = n8807 & n8808;
  assign n7533 = n8809 & n8810;
  assign n7535 = n8811 & n8812;
  assign n7537 = n8813 & n8814;
  assign n7405 = n8815 & n8816;
  assign n7532 = n8817 & n8818;
  assign n7536 = n8819 & n8820;
  assign n7539 = n8821 & n8822;
  assign n7538 = n8823 & n8824;
  assign n7942 = n8825 & n8826;
  assign n7543 = n8827 & n8828;
  assign n7534 = n8829 & n8830;
  assign n7549 = n8831 & n8832;
  assign n7544 = n8833 & n8834;
  assign n7548 = n8835 & n8836;
  assign n7426 = n8837 & n8838;
  assign n7547 = n8839 & n8840;
  assign n7546 = n8841 & n8842;
  assign n7553 = n8843 & n8844;
  assign n7552 = n8845 & n8846;
  assign n7555 = n8847 & n8848;
  assign n7557 = n8849 & n8850;
  assign n7556 = n8851 & n8852;
  assign n7560 = n8853 & n8854;
  assign n7559 = n8855 & n8856;
  assign n7562 = n8857 & n8858;
  assign n7558 = n8859 & n8860;
  assign n7568 = n8861 & n8862;
  assign n7571 = n8863 & n8864;
  assign n7570 = n8865 & n8866;
  assign n7575 = n8867 & n8868;
  assign n7574 = n8869 & n8870;
  assign n7573 = n8871 & n8872;
  assign n7808 = n8873 & n8874;
  assign n7572 = n8875 & n8876;
  assign n7159 = n8877 & n8878;
  assign n7158 = n8879 & n8880;
  assign n7579 = n8881 & n8882;
  assign n7578 = n8883 & n8884;
  assign n7582 = n8885 & n8886;
  assign n7966 = n8887 & n8888;
  assign n7565 = n8889 & n8890;
  assign n7249 = n8891 & n8892;
  assign n7564 = n8893 & n8894;
  assign n7375 = n8895 & n8896;
  assign n7018 = n8897 & n8898;
  assign n7448 = n8899 & n8900;
  assign n7589 = n8901 & n8902;
  assign n7771 = n8903 & n8904;
  assign n7588 = n8905 & n8906;
  assign n7779 = n8907 & n8908;
  assign n7593 = n8909 & n8910;
  assign n7959 = n8911 & n8912;
  assign n7938 = n8913 & n8914;
  assign n7599 = n8915 & n8916;
  assign n7601 = n8917 & n8918;
  assign n7056 = n8919 & n8920;
  assign n7598 = n8921 & n8922;
  assign n7603 = n8923 & n8924;
  assign n7802 = n8925 & n8926;
  assign n7602 = n8927 & n8928;
  assign n7609 = n8929 & n8930;
  assign n7707 = n8931 & n8932;
  assign n7608 = n8933 & n8934;
  assign n7597 = n8935 & n8936;
  assign n7613 = n8937 & n8938;
  assign n7614 = n8939 & n8940;
  assign n7623 = n8941 & n8942;
  assign n7622 = n8943 & n8944;
  assign n7625 = n8945 & n8946;
  assign n7624 = n8947 & n8948;
  assign n7807 = n8949 & n8950;
  assign n7341 = n8951 & n8952;
  assign n7735 = n8953 & n8954;
  assign n7734 = n8955 & n8956;
  assign n7604 = n8957 & n8958;
  assign n7629 = n8959 & n8960;
  assign n7628 = n8961 & n8962;
  assign n7631 = n8963 & n8964;
  assign n7137 = n8965 & n8966;
  assign n7630 = n8967 & n8968;
  assign n7626 = n8969 & n8970;
  assign n7083 = n8971 & n8972;
  assign n7157 = n8973 & n8974;
  assign n7518 = n8975 & n8976;
  assign n7395 = n8977 & n8978;
  assign n7758 = n8979 & n8980;
  assign n7633 = n8981 & n8982;
  assign n7898 = n8983 & n8984;
  assign n7672 = n8985 & n8986;
  assign n7639 = n8987 & n8988;
  assign n7632 = n8989 & n8990;
  assign n7279 = n8991 & n8992;
  assign n7798 = n8993 & n8994;
  assign n7635 = n8995 & n8996;
  assign n7683 = n8997 & n8998;
  assign n7634 = n8999 & n9000;
  assign n7109 = n9001 & n9002;
  assign n7803 = n9003 & n9004;
  assign n7811 = n9005 & n9006;
  assign n7637 = n9007 & n9008;
  assign n7712 = n9009 & n9010;
  assign n7636 = n9011 & n9012;
  assign n7689 = n9013 & n9014;
  assign n7640 = n9015 & n9016;
  assign n7723 = n9017 & n9018;
  assign n7428 = n9019 & n9020;
  assign n7336 = n9021 & n9022;
  assign n7832 = n9023 & n9024;
  assign n7187 = n9025 & n9026;
  assign n7900 = n9027 & n9028;
  assign n7638 = n9029 & n9030;
  assign n7178 = n9031 & n9032;
  assign n7218 = n9033 & n9034;
  assign n7747 = n9035 & n9036;
  assign n7422 = n9037 & n9038;
  assign n7861 = n9039 & n9040;
  assign n7648 = n9041 & n9042;
  assign n7653 = n9043 & n9044;
  assign n7652 = n9045 & n9046;
  assign n7649 = n9047 & n9048;
  assign n7132 = n9049 & n9050;
  assign n7657 = n9051 & n9052;
  assign n7656 = n9053 & n9054;
  assign n7658 = n9055 & n9056;
  assign n7660 = n9057 & n9058;
  assign n7890 = n9059 & n9060;
  assign n7665 = n9061 & n9062;
  assign n7026 = n9063 & n9064;
  assign n7768 = n9065 & n9066;
  assign n7033 = n9067 & n9068;
  assign n7667 = n9069 & n9070;
  assign n7905 = n9071 & n9072;
  assign n7720 = n9073 & n9074;
  assign n7465 = n9075 & n9076;
  assign n7964 = n9077 & n9078;
  assign n7147 = n9079 & n9080;
  assign n7671 = n9081 & n9082;
  assign n7670 = n9083 & n9084;
  assign n7025 = n9085 & n9086;
  assign n7676 = n9087 & n9088;
  assign n7679 = n9089 & n9090;
  assign n7674 = n9091 & n9092;
  assign n7933 = n9093 & n9094;
  assign n7645 = n9095 & n9096;
  assign n7874 = n9097 & n9098;
  assign n7431 = n9099 & n9100;
  assign n7584 = n9101 & n9102;
  assign n7688 = n9103 & n9104;
  assign n7306 = n9105 & n9106;
  assign n7693 = n9107 & n9108;
  assign n7060 = n9109 & n9110;
  assign n7751 = n9111 & n9112;
  assign n7750 = n9113 & n9114;
  assign n7521 = n9115 & n9116;
  assign n7520 = n9117 & n9118;
  assign n7694 = n9119 & n9120;
  assign n7309 = n9121 & n9122;
  assign n7243 = n9123 & n9124;
  assign n7661 = n9125 & n9126;
  assign n7716 = n9127 & n9128;
  assign n7563 = n9129 & n9130;
  assign n7338 = n9131 & n9132;
  assign n7493 = n9133 & n9134;
  assign n7956 = n9135 & n9136;
  assign n7492 = n9137 & n9138;
  assign n7698 = n9139 & n9140;
  assign n7697 = n9141 & n9142;
  assign n7703 = n9143 & n9144;
  assign n7701 = n9145 & n9146;
  assign n7691 = n9147 & n9148;
  assign n7702 = n9149 & n9150;
  assign n7705 = n9151 & n9152;
  assign n7704 = n9153 & n9154;
  assign n7696 = n9155 & n9156;
  assign n7917 = n9157 & n9158;
  assign n7114 = n9159 & n9160;
  assign n7091 = n9161 & n9162;
  assign n7706 = n9163 & n9164;
  assign n7901 = n9165 & n9166;
  assign n7529 = n9167 & n9168;
  assign n7238 = n9169 & n9170;
  assign n7815 = n9171 & n9172;
  assign n7561 = n9173 & n9174;
  assign n7617 = n9175 & n9176;
  assign n7710 = n9177 & n9178;
  assign n7131 = n9179 & n9180;
  assign n7715 = n9181 & n9182;
  assign n7714 = n9183 & n9184;
  assign n7719 = n9185 & n9186;
  assign n6070 = n9187 ^ n9188;
  assign n7717 = n9189 & n9190;
  assign n7718 = n9191 & n9192;
  assign n7711 = n9193 & n9194;
  assign n7722 = n9195 & n9196;
  assign n7725 = n9197 & n9198;
  assign n7031 = n9199 & n9200;
  assign n7851 = n9201 & n9202;
  assign n7459 = n9203 & n9204;
  assign n7458 = n9205 & n9206;
  assign n7530 = n9207 & n9208;
  assign n7960 = n9209 & n9210;
  assign n7063 = n9211 & n9212;
  assign n7891 = n9213 & n9214;
  assign n7066 = n9215 & n9216;
  assign n7585 = n9217 & n9218;
  assign n7941 = n9219 & n9220;
  assign n7761 = n9221 & n9222;
  assign n7292 = n9223 & n9224;
  assign n7690 = n9225 & n9226;
  assign n7425 = n9227 & n9228;
  assign n7940 = n9229 & n9230;
  assign n7666 = n9231 & n9232;
  assign n7732 = n9233 & n9234;
  assign n7424 = n9235 & n9236;
  assign n7297 = n9237 & n9238;
  assign n7858 = n9239 & n9240;
  assign n7391 = n9241 & n9242;
  assign n7760 = n9243 & n9244;
  assign n7627 = n9245 & n9246;
  assign n7887 = n9247 & n9248;
  assign n7886 = n9249 & n9250;
  assign n7737 = n9251 & n9252;
  assign n7736 = n9253 & n9254;
  assign n7390 = n9255 & n9256;
  assign n7740 = n9257 & n9258;
  assign n7621 = n9259 & n9260;
  assign n7902 = n9261 & n9262;
  assign n7949 = n9263 & n9264;
  assign n7142 = n9265 & n9266;
  assign n7777 = n9267 & n9268;
  assign n7071 = n9269 & n9270;
  assign n7752 = n9271 & n9272;
  assign n7738 = n9273 & n9274;
  assign n7554 = n9275 & n9276;
  assign n7739 = n9277 & n9278;
  assign n7251 = n9279 & n9280;
  assign n7904 = n9281 & n9282;
  assign n7250 = n9283 & n9284;
  assign n7085 = n9285 & n9286;
  assign n7659 = n9287 & n9288;
  assign n7215 = n9289 & n9290;
  assign n7596 = n9291 & n9292;
  assign n7017 = n9293 & n9294;
  assign n7754 = n9295 & n9296;
  assign n7098 = n9297 & n9298;
  assign n7757 = n9299 & n9300;
  assign n7685 = n9301 & n9302;
  assign n7791 = n9303 & n9304;
  assign n7924 = n9305 & n9306;
  assign n7859 = n9307 & n9308;
  assign n7925 = n9309 & n9310;
  assign n7058 = n9311 & n9312;
  assign n7763 = n9313 & n9314;
  assign n7743 = n9315 & n9316;
  assign n7527 = n9317 & n9318;
  assign n7576 = n9319 & n9320;
  assign n7764 = n9321 & n9322;
  assign n7076 = n9323 & n9324;
  assign n7770 = n9325 & n9326;
  assign n7827 = n9327 & n9328;
  assign n7912 = n9329 & n9330;
  assign n7170 = n9331 & n9332;
  assign n7237 = n9333 & n9334;
  assign n7650 = n9335 & n9336;
  assign n7461 = n9337 & n9338;
  assign n7773 = n9339 & n9340;
  assign n7778 = n9341 & n9342;
  assign n7780 = n9343 & n9344;
  assign n7772 = n9345 & n9346;
  assign n7042 = n9347 & n9348;
  assign n7787 = n9349 & n9350;
  assign n7072 = n9351 & n9352;
  assign n7799 = n9353 & n9354;
  assign n7786 = n9355 & n9356;
  assign n7884 = n9357 & n9358;
  assign n7903 = n9359 & n9360;
  assign n7762 = n9361 & n9362;
  assign n7469 = n9363 & n9364;
  assign n7793 = n9365 & n9366;
  assign n7792 = n9367 & n9368;
  assign n7163 = n9369 & n9370;
  assign n7682 = n9371 & n9372;
  assign n7176 = n9373 & n9374;
  assign n7797 = n9375 & n9376;
  assign n7805 = n9377 & n9378;
  assign n7800 = n9379 & n9380;
  assign n7804 = n9381 & n9382;
  assign n7145 = n9383 & n9384;
  assign n7813 = n9385 & n9386;
  assign n7438 = n9387 & n9388;
  assign n7220 = n9389 & n9390;
  assign n7806 = n9391 & n9392;
  assign n7812 = n9393 & n9394;
  assign n7809 = n9395 & n9396;
  assign n7810 = n9397 & n9398;
  assign n7149 = n9399 & n9400;
  assign n7814 = n9401 & n9402;
  assign n7148 = n9403 & n9404;
  assign n7817 = n9405 & n9406;
  assign n7816 = n9407 & n9408;
  assign n7910 = n9409 & n9410;
  assign n7540 = n9411 & n9412;
  assign n7655 = n9413 & n9414;
  assign n7935 = n9415 & n9416;
  assign n7896 = n9417 & n9418;
  assign n7833 = n9419 & n9420;
  assign n7354 = n9421 & n9422;
  assign n7135 = n9423 & n9424;
  assign n7928 = n9425 & n9426;
  assign n7968 = n9427 & n9428;
  assign n7821 = n9429 & n9430;
  assign n7824 = n9431 & n9432;
  assign n7647 = n9433 & n9434;
  assign n7418 = n9435 & n9436;
  assign n7822 = n9437 & n9438;
  assign n7826 = n9439 & n9440;
  assign n7829 = n9441 & n9442;
  assign n7831 = n9443 & n9444;
  assign n7801 = n9445 & n9446;
  assign n7835 = n9447 & n9448;
  assign n7834 = n9449 & n9450;
  assign n7837 = n9451 & n9452;
  assign n7483 = n9453 & n9454;
  assign n7841 = n9455 & n9456;
  assign n7838 = n9457 & n9458;
  assign n7836 = n9459 & n9460;
  assign n7331 = n9461 & n9462;
  assign n7144 = n9463 & n9464;
  assign n7853 = n9465 & n9466;
  assign n7692 = n9467 & n9468;
  assign n7951 = n9469 & n9470;
  assign n7852 = n9471 & n9472;
  assign n7654 = n9473 & n9474;
  assign n7784 = n9475 & n9476;
  assign n7844 = n9477 & n9478;
  assign n7847 = n9479 & n9480;
  assign n7846 = n9481 & n9482;
  assign n7506 = n9483 & n9484;
  assign n7605 = n9485 & n9486;
  assign n7850 = n9487 & n9488;
  assign n7863 = n9489 & n9490;
  assign n7908 = n9491 & n9492;
  assign n7872 = n9493 & n9494;
  assign n7856 = n9495 & n9496;
  assign n7860 = n9497 & n9498;
  assign n7854 = n9499 & n9500;
  assign n7867 = n9501 & n9502;
  assign n7012 = n9503 & n9504;
  assign n7868 = n9505 & n9506;
  assign n7866 = n9507 & n9508;
  assign n7011 = n9509 & n9510;
  assign n7870 = n9511 & n9512;
  assign n7873 = n9513 & n9514;
  assign n7457 = n9515 & n9516;
  assign n7876 = n9517 & n9518;
  assign n7879 = n9519 & n9520;
  assign n7881 = n9521 & n9522;
  assign n7878 = n9523 & n9524;
  assign n7883 = n9525 & n9526;
  assign n7875 = n9527 & n9528;
  assign n7957 = n9529 & n9530;
  assign n7776 = n9531 & n9532;
  assign n7551 = n9533 & n9534;
  assign n7765 = n9535 & n9536;
  assign n7842 = n9537 & n9538;
  assign n7893 = n9539 & n9540;
  assign n7374 = n9541 & n9542;
  assign n7745 = n9543 & n9544;
  assign n7503 = n9545 & n9546;
  assign n7888 = n9547 & n9548;
  assign n7449 = n9549 & n9550;
  assign n7967 = n9551 & n9552;
  assign n7646 = n9553 & n9554;
  assign n7895 = n9555 & n9556;
  assign n7907 = n9557 & n9558;
  assign n7756 = n9559 & n9560;
  assign n7744 = n9561 & n9562;
  assign n7788 = n9563 & n9564;
  assign n7899 = n9565 & n9566;
  assign n7731 = n9567 & n9568;
  assign n7348 = n9569 & n9570;
  assign n7937 = n9571 & n9572;
  assign n7795 = n9573 & n9574;
  assign n7037 = n9575 & n9576;
  assign n7214 = n9577 & n9578;
  assign n7221 = n9579 & n9580;
  assign n7818 = n9581 & n9582;
  assign n7118 = n9583 & n9584;
  assign n7897 = n9585 & n9586;
  assign n7173 = n9587 & n9588;
  assign n7906 = n9589 & n9590;
  assign n7580 = n9591 & n9592;
  assign n7213 = n9593 & n9594;
  assign n7225 = n9595 & n9596;
  assign n7328 = n9597 & n9598;
  assign n7733 = n9599 & n9600;
  assign n7915 = n9601 & n9602;
  assign n7916 = n9603 & n9604;
  assign n7914 = n9605 & n9606;
  assign n7918 = n9607 & n9608;
  assign n7351 = n9609 & n9610;
  assign n7611 = n9611 & n9612;
  assign n7923 = n9613 & n9614;
  assign n7922 = n9615 & n9616;
  assign n7668 = n9617 & n9618;
  assign n7610 = n9619 & n9620;
  assign n7819 = n9621 & n9622;
  assign n7927 = n9623 & n9624;
  assign n7282 = n9625 & n9626;
  assign n7040 = n9627 & n9628;
  assign n7934 = n9629 & n9630;
  assign n7291 = n9631 & n9632;
  assign n7931 = n9633 & n9634;
  assign n7944 = n9635 & n9636;
  assign n7946 = n9637 & n9638;
  assign n7287 = n9639 & n9640;
  assign n7862 = n9641 & n9642;
  assign n7932 = n9643 & n9644;
  assign n7790 = n9645 & n9646;
  assign n7526 = n9647 & n9648;
  assign n7828 = n9649 & n9650;
  assign n7172 = n9651 & n9652;
  assign n7727 = n9653 & n9654;
  assign n7612 = n9655 & n9656;
  assign n7955 = n9657 & n9658;
  assign n7958 = n9659 & n9660;
  assign n7961 = n9661 & n9662;
  assign n7962 = n9663 & n9664;
  assign n7885 = n9665 & n9666;
  assign n7769 = n9667 & n9668;
  assign n7976 = n6294 & n5163;
  assign n6078 = n9669 ^ n9670;
  assign n6072 = n9671 ^ n9672;
  assign n6074 = n9673 ^ n9674;
  assign n6076 = n9675 ^ n9676;
  assign n7947 = n9692 & n9693;
  assign n7911 = n9709 & n9710;
  assign n7184 = n9711 & n9712;
  assign n7789 = n9713 & n9714;
  assign n7038 = n9715 & n9716;
  assign n6068 = n9717 ^ n9704;
  assign n7209 = n9718 & n9719;
  assign n6066 = n9720 ^ n9684;
  assign n7975 = n6270 & n5138;
  assign n7913 = n9721 & n9722;
  assign n7909 = n9723 & n9724;
  assign n7086 = n9725 & n9726;
  assign n7669 = n9727 & n9728;
  assign n7167 = n9729 & n9730;
  assign n7334 = n9731 & n9732;
  assign n7523 = n9733 & n9734;
  assign n7889 = n9735 & n9736;
  assign n7312 = n9737 & n9738;
  assign n7474 = n9739 & n9740;
  assign n7389 = n9741 & n9742;
  assign n7254 = n9743 & n9744;
  assign n7203 = n9745 & n9746;
  assign n7475 = n9747 & n9748;
  assign n7346 = n9749 & n9750;
  assign n7032 = n9751 & n9752;
  assign n7030 = n9753 & n9754;
  assign n7845 = n9755 & n9756;
  assign n7016 = n9757 & n9758;
  assign n7015 = n9759 & n9760;
  assign n7467 = n9761 & n9762;
  assign n7036 = n9763 & n9764;
  assign n7065 = n9765 & n9766;
  assign n7064 = n9767 & n9768;
  assign n7369 = n9769 & n9770;
  assign n7436 = n9771 & n9772;
  assign n7437 = n9773 & n9774;
  assign n7116 = n9775 & n9776;
  assign n7023 = n9777 & n9778;
  assign n7550 = n9779 & n9780;
  assign n7022 = n9781 & n9782;
  assign n7062 = n9783 & n9784;
  assign n7074 = n9785 & n9786;
  assign n7919 = n9787 & n9788;
  assign n7019 = n9789 & n9790;
  assign n7122 = n9791 & n9792;
  assign n7079 = n9793 & n9794;
  assign n7081 = n9795 & n9796;
  assign n7082 = n9797 & n9798;
  assign n7078 = n9799 & n9800;
  assign n7695 = n9801 & n9802;
  assign n7084 = n9803 & n9804;
  assign n7195 = n9805 & n9806;
  assign n7171 = n9807 & n9808;
  assign n7721 = n9809 & n9810;
  assign n7577 = n9811 & n9812;
  assign n7219 = n9813 & n9814;
  assign n7089 = n9815 & n9816;
  assign n7088 = n9817 & n9818;
  assign n7090 = n9819 & n9820;
  assign n7308 = n9821 & n9822;
  assign n7404 = n9823 & n9824;
  assign n7595 = n9825 & n9826;
  assign n7594 = n9827 & n9828;
  assign n7095 = n9829 & n9830;
  assign n7097 = n9831 & n9832;
  assign n7096 = n9833 & n9834;
  assign n7094 = n9835 & n9836;
  assign n7386 = n9837 & n9838;
  assign n7146 = n9839 & n9840;
  assign n7794 = n9841 & n9842;
  assign n7101 = n9843 & n9844;
  assign n7100 = n9845 & n9846;
  assign n7451 = n9847 & n9848;
  assign n7106 = n9849 & n9850;
  assign n7105 = n9851 & n9852;
  assign n7699 = n9853 & n9854;
  assign n7208 = n9855 & n9856;
  assign n7726 = n9857 & n9858;
  assign n7399 = n9859 & n9860;
  assign n7111 = n9861 & n9862;
  assign n7954 = n9863 & n9864;
  assign n7069 = n9865 & n9866;
  assign n7134 = n9867 & n9868;
  assign n7496 = n9869 & n9870;
  assign n7746 = n9871 & n9872;
  assign n7825 = n9873 & n9874;
  assign n7067 = n9875 & n9876;
  assign n7619 = n9877 & n9878;
  assign n7117 = n9879 & n9880;
  assign n7476 = n9881 & n9882;
  assign n7618 = n9883 & n9884;
  assign n7353 = n9885 & n9886;
  assign n7034 = n9887 & n9888;
  assign n7120 = n9889 & n9890;
  assign n7514 = n9891 & n9892;
  assign n7068 = n9893 & n9894;
  assign n7335 = n9895 & n9896;
  assign n7075 = n9897 & n9898;
  assign n7894 = n9899 & n9900;
  assign n7869 = n9901 & n9902;
  assign n7587 = n9903 & n9904;
  assign n7387 = n9905 & n9906;
  assign n7329 = n9907 & n9908;
  assign n7013 = n9909 & n9910;
  assign n7140 = n9911 & n9912;
  assign n7355 = n9913 & n9914;
  assign n7009 = n9915 & n9916;
  assign n7766 = n9917 & n9918;
  assign n7620 = n9919 & n9920;
  assign n7590 = n9921 & n9922;
  assign n7324 = n9923 & n9924;
  assign n7104 = n9925 & n9926;
  assign n7342 = n9927 & n9928;
  assign n7124 = n9929 & n9930;
  assign n7591 = n9931 & n9932;
  assign n7352 = n9933 & n9934;
  assign n7687 = n9935 & n9936;
  assign n7024 = n9937 & n9938;
  assign n9679 = n5132 & n9941;
  assign n9680 = n9720 & n9942;
  assign n9687 = n9671 & n9943;
  assign n6991 = ~n6406;
  assign n7973 = ~n6294;
  assign n6971 = ~n6198;
  assign n6959 = ~n6160;
  assign n6965 = ~n6242;
  assign n6980 = ~n6352;
  assign n6973 = ~n6236;
  assign n6985 = ~n6428;
  assign n6989 = ~n6252;
  assign n8005 = ~n6270;
  assign n6998 = ~n6166;
  assign n6969 = ~n6320;
  assign n6960 = ~n6346;
  assign n6979 = ~n6308;
  assign n9694 = n9673 & n9944;
  assign n9689 = n9187 & n9945;
  assign n9685 = n9669 & n9946;
  assign n9700 = n9675 & n9947;
  assign n9702 = n9717 & n9948;
  assign n9678 = n9949 & n9950;
  assign n7983 = n9957 & n61;
  assign n7972 = ~n9963;
  assign n6093 = n10098 & n41;
  assign n6572 = ~n6278;
  assign n9681 = ~n7984;
  assign n9695 = ~n9669;
  assign n9951 = n10227 & n10228;
  assign n6544 = ~n6232;
  assign n9690 = ~n7982;
  assign n9701 = ~n9187;
  assign n9688 = ~n7986;
  assign n9696 = ~n8003;
  assign n6466 = ~n10901;
  assign n6616 = ~n6368;
  assign n6444 = ~n6244;
  assign n6534 = ~n5088;
  assign n9698 = ~n9675;
  assign n6582 = ~n5187;
  assign n6560 = ~n5142;
  assign n9697 = ~n9671;
  assign n6676 = ~n6332;
  assign n9703 = ~n9717;
  assign n6686 = ~n4996;
  assign n6594 = ~n6326;
  assign n9707 = ~n9673;
  assign n9686 = ~n7999;
  assign n9705 = ~n9949;
  assign n9683 = ~n9720;
  assign n9708 = ~n7980;
  assign n6606 = ~n5219;
  assign n9677 = ~n5132;
  assign n9691 = ~n8001;
  assign n9682 = ~n7978;
  assign n6446 = ~n5004;
  assign n9699 = ~n7988;
  assign n6219 = n10904 & n59;
  assign n7981 = n10908 & n63;
  assign n8000 = n10909 & n47;
  assign n6267 = n10911 & n57;
  assign n7977 = n10916 & n35;
  assign n7987 = n10920 & n45;
  assign n8002 = n10922 & n37;
  assign n7985 = n10924 & n51;
  assign n6311 = n10925 & n55;
  assign n7979 = n10928 & n39;
  assign n6211 = n10929 & n43;
  assign n7998 = n10935 & n49;
  assign n6343 = n10942 & n53;
  assign n3202 = n6954 ^ n6700;
  assign n3890 = n7009 & n7010;
  assign n6380 = n7011 & n7012;
  assign n6421 = n7013 & n7014;
  assign n6094 = n7015 & n7016;
  assign n6071 = n7017 & n7018;
  assign n6129 = n7019 & n7020;
  assign n6063 = n7022 & n7023;
  assign n6347 = n7024 & n7025;
  assign n6408 = n7026 & n7027;
  assign n6418 = n7028 & n7029;
  assign n4967 = n7030 & n7031;
  assign n6243 = n7032 & n7033;
  assign n6223 = n7034 & n7035;
  assign n6348 = n7036 & n7037;
  assign n6051 = n7038 & n7039;
  assign n6146 = n7040 & n7041;
  assign n4139 = n7042 & n7043;
  assign n6230 = n7044 & n7045;
  assign n5189 = n7046 & n7047;
  assign n4174 = n7048 & n7049;
  assign n4136 = n7050 & n7051;
  assign n3894 = n7052 & n7053;
  assign n6296 = n7054 & n7055;
  assign n6054 = n7056 & n7057;
  assign n5038 = n7058 & n7059;
  assign n3896 = n7060 & n7061;
  assign n6069 = n7062 & n7063;
  assign n6140 = n7064 & n7065;
  assign n6411 = n7066 & n7067;
  assign n5020 = n7068 & n7069;
  assign n5273 = n7070 & n7071;
  assign n6049 = n7072 & n7073;
  assign n6179 = n7074 & n7075;
  assign n6193 = n7076 & n7077;
  assign n5016 = n7078 & n7079;
  assign n5058 = n7080 & n7081;
  assign n6114 = n7082 & n7083;
  assign n6113 = n7084 & n7085;
  assign n6265 = n7086 & n7087;
  assign n5046 = n7088 & n7089;
  assign n6098 = n7090 & n7091;
  assign n6197 = n7092 & n7093;
  assign n6106 = n7094 & n7095;
  assign n6065 = n7096 & n7097;
  assign n5269 = n7098 & n7099;
  assign n6134 = n7100 & n7101;
  assign n6187 = n7102 & n7103;
  assign n6133 = n7104 & n7105;
  assign n6090 = n7106 & n7107;
  assign n6102 = n7108 & n7109;
  assign n6156 = n7110 & n7111;
  assign n6359 = n7112 & n7113;
  assign n5060 = n7114 & n7115;
  assign n6180 = n7116 & n7117;
  assign n5285 = n7118 & n7119;
  assign n6062 = n7120 & n7121;
  assign n6153 = n7122 & n7123;
  assign n6135 = n7124 & n7125;
  assign n6222 = n7126 & n7127;
  assign n6126 = n7128 & n7129;
  assign n6141 = n7130 & n7131;
  assign n5203 = n7132 & n7133;
  assign n6155 = n7134 & n7135;
  assign n5050 = n7136 & n7137;
  assign n6058 = n7138 & n7139;
  assign n6142 = n7140 & n7141;
  assign n5108 = n7142 & n7143;
  assign n6285 = n7144 & n7145;
  assign n5042 = n7146 & n7147;
  assign n6415 = n7148 & n7149;
  assign n6151 = n7150 & n7151;
  assign n6389 = n7152 & n7153;
  assign n5112 = n7154 & n7155;
  assign n6186 = n7156 & n7157;
  assign n5205 = n7158 & n7159;
  assign n6229 = n7160 & n7161;
  assign n5022 = n7162 & n7163;
  assign n6152 = n7164 & n7165;
  assign n6130 = n7166 & n7167;
  assign n6224 = n7168 & n7169;
  assign n5253 = n7170 & n7171;
  assign n6122 = n7172 & n7173;
  assign n6172 = n7174 & n7175;
  assign n6286 = n7176 & n7177;
  assign n5199 = n7178 & n7179;
  assign n6171 = n7180 & n7181;
  assign n5064 = n7182 & n7183;
  assign n5257 = n7184 & n7185;
  assign n5263 = n7186 & n7187;
  assign n6162 = n7188 & n7189;
  assign n6067 = n7190 & n7191;
  assign n6161 = n7192 & n7193;
  assign n6355 = n7194 & n7195;
  assign n6176 = n7196 & n7197;
  assign n6290 = n7198 & n7199;
  assign n6175 = n7200 & n7201;
  assign n6430 = n7202 & n7203;
  assign n5074 = n7204 & n7205;
  assign n6159 = n7206 & n7207;
  assign n6119 = n7208 & n7209;
  assign n5062 = n7210 & n7211;
  assign n6303 = n7212 & n7213;
  assign n6420 = n7214 & n7215;
  assign n6184 = n7216 & n7217;
  assign n5010 = n7218 & n7219;
  assign n6127 = n7220 & n7221;
  assign n6238 = n7222 & n7223;
  assign n6164 = n7224 & n7225;
  assign n6163 = n7226 & n7227;
  assign n6178 = n7228 & n7229;
  assign n6177 = n7230 & n7231;
  assign n6183 = n7232 & n7233;
  assign n5076 = n7234 & n7235;
  assign n5066 = n7236 & n7237;
  assign n6170 = n7238 & n7239;
  assign n6169 = n7240 & n7241;
  assign n5070 = n7242 & n7243;
  assign n6174 = n7244 & n7245;
  assign n6173 = n7246 & n7247;
  assign n6228 = n7248 & n7249;
  assign n5281 = n7250 & n7251;
  assign n5072 = n7252 & n7253;
  assign n6091 = n7254 & n7255;
  assign n3892 = n7256 & n7257;
  assign n5114 = n7258 & n7259;
  assign n6055 = n7260 & n7261;
  assign n6424 = n7262 & n7263;
  assign n5110 = n7264 & n7265;
  assign n6214 = n7266 & n7267;
  assign n6213 = n7268 & n7269;
  assign n6226 = n7270 & n7271;
  assign n5100 = n7272 & n7273;
  assign n6210 = n7274 & n7275;
  assign n6225 = n7276 & n7277;
  assign n6209 = n7278 & n7279;
  assign n5098 = n7280 & n7281;
  assign n6241 = n7282 & n7283;
  assign n6216 = n7284 & n7285;
  assign n6289 = n7286 & n7287;
  assign n6215 = n7288 & n7289;
  assign n5102 = n7290 & n7291;
  assign n5124 = n7292 & n7293;
  assign n6208 = n7294 & n7295;
  assign n6202 = n7296 & n7297;
  assign n6201 = n7298 & n7299;
  assign n5094 = n7300 & n7301;
  assign n5177 = n7302 & n7303;
  assign n6246 = n7304 & n7305;
  assign n6338 = n7306 & n7307;
  assign n6409 = n7308 & n7309;
  assign n6317 = n7310 & n7311;
  assign n5305 = n7312 & n7313;
  assign n6324 = n7314 & n7315;
  assign n6182 = n7316 & n7317;
  assign n5126 = n7318 & n7319;
  assign n6245 = n7320 & n7321;
  assign n6181 = n7322 & n7323;
  assign n6240 = n7324 & n7325;
  assign n6239 = n7326 & n7327;
  assign n5291 = n7328 & n7329;
  assign n5265 = n7330 & n7331;
  assign n5134 = n7332 & n7333;
  assign n5024 = n7334 & n7335;
  assign n6312 = n7336 & n7337;
  assign n6302 = n7338 & n7339;
  assign n6254 = n7340 & n7341;
  assign n5044 = n7342 & n7343;
  assign n6253 = n7344 & n7345;
  assign n5002 = n7346 & n7347;
  assign n6077 = n7348 & n7349;
  assign n6123 = n7350 & n7351;
  assign n7005 = n7352 & n7353;
  assign n6150 = n7354 & n7355;
  assign n6381 = n7356 & n7357;
  assign n6301 = n7358 & n7359;
  assign n6220 = n7360 & n7361;
  assign n6234 = n7362 & n7363;
  assign n6233 = n7364 & n7365;
  assign n5118 = n7366 & n7367;
  assign n6256 = n7368 & n7369;
  assign n6255 = n7370 & n7371;
  assign n5136 = n7372 & n7373;
  assign n4992 = n7374 & n7375;
  assign n6248 = n7376 & n7377;
  assign n5086 = n7378 & n7379;
  assign n6191 = n7380 & n7381;
  assign n4963 = n7382 & n7383;
  assign n6059 = n7384 & n7385;
  assign n6196 = n7386 & n7387;
  assign n6195 = n7388 & n7389;
  assign n5034 = n7390 & n7391;
  assign n5092 = n7392 & n7393;
  assign n5185 = n7394 & n7395;
  assign n6056 = n7396 & n7397;
  assign n6200 = n7398 & n7399;
  assign n6300 = n7400 & n7401;
  assign n6199 = n7402 & n7403;
  assign n6121 = n7404 & n7405;
  assign n6139 = n7406 & n7407;
  assign n6206 = n7408 & n7409;
  assign n6299 = n7410 & n7411;
  assign n6205 = n7412 & n7413;
  assign n5096 = n7414 & n7415;
  assign n6280 = n7416 & n7417;
  assign n5171 = n7418 & n7419;
  assign n6292 = n7420 & n7421;
  assign n6279 = n7422 & n7423;
  assign n5104 = n7424 & n7425;
  assign n6203 = n7426 & n7427;
  assign n6291 = n7428 & n7429;
  assign n6218 = n7430 & n7431;
  assign n6217 = n7432 & n7433;
  assign n5169 = n7434 & n7435;
  assign n4941 = n7436 & n7437;
  assign n5259 = n7438 & n7439;
  assign n6231 = n7440 & n7441;
  assign n5116 = n7442 & n7443;
  assign n6295 = n7444 & n7445;
  assign n6237 = n7446 & n7447;
  assign n5056 = n7448 & n7449;
  assign n5120 = n7450 & n7451;
  assign n5179 = n7452 & n7453;
  assign n6274 = n7454 & n7455;
  assign n6386 = n7456 & n7457;
  assign n5237 = n7458 & n7459;
  assign n5122 = n7460 & n7461;
  assign n6235 = n7462 & n7463;
  assign n5197 = n7464 & n7465;
  assign n6250 = n7466 & n7467;
  assign n5084 = n7468 & n7469;
  assign n6154 = n7470 & n7471;
  assign n6249 = n7472 & n7473;
  assign n6188 = n7474 & n7475;
  assign n6322 = n7476 & n7477;
  assign n6318 = n7478 & n7479;
  assign n5128 = n7480 & n7481;
  assign n6086 = n7482 & n7483;
  assign n5130 = n7484 & n7485;
  assign n5140 = n7486 & n7487;
  assign n6259 = n7488 & n7489;
  assign n5144 = n7490 & n7491;
  assign n6400 = n7492 & n7493;
  assign n6385 = n7494 & n7495;
  assign n6266 = n7496 & n7497;
  assign n6316 = n7498 & n7499;
  assign n5150 = n7500 & n7501;
  assign n6261 = n7502 & n7503;
  assign n5255 = n7504 & n7505;
  assign n5148 = n7506 & n7507;
  assign n5195 = n7508 & n7509;
  assign n6258 = n7510 & n7511;
  assign n6257 = n7512 & n7513;
  assign n6306 = n7514 & n7515;
  assign n6168 = n7516 & n7517;
  assign n6167 = n7518 & n7519;
  assign n6410 = n7520 & n7521;
  assign n6264 = n7522 & n7523;
  assign n6263 = n7524 & n7525;
  assign n5036 = n7526 & n7527;
  assign n6268 = n7528 & n7529;
  assign n6422 = n7530 & n7531;
  assign n5225 = n7532 & n7533;
  assign n6307 = n7534 & n7535;
  assign n6052 = n7536 & n7537;
  assign n6138 = n7538 & n7539;
  assign n6137 = n7540 & n7541;
  assign n6354 = n7542 & n7543;
  assign n5207 = n7544 & n7545;
  assign n6334 = n7546 & n7547;
  assign n5159 = n7548 & n7549;
  assign n6084 = n7550 & n7551;
  assign n6276 = n7552 & n7553;
  assign n6353 = n7554 & n7555;
  assign n6333 = n7556 & n7557;
  assign n5261 = n7558 & n7559;
  assign n5165 = n7560 & n7561;
  assign n6277 = n7562 & n7563;
  assign n5193 = n7564 & n7565;
  assign n6371 = n7566 & n7567;
  assign n6272 = n7568 & n7569;
  assign n6271 = n7570 & n7571;
  assign n6427 = n7572 & n7573;
  assign n5157 = n7574 & n7575;
  assign n6362 = n7576 & n7577;
  assign n6351 = n7578 & n7579;
  assign n6147 = n7580 & n7581;
  assign n6314 = n7582 & n7583;
  assign n6313 = n7584 & n7585;
  assign n6194 = n7586 & n7587;
  assign n6342 = n7588 & n7589;
  assign n6125 = n7590 & n7591;
  assign n6341 = n7592 & n7593;
  assign n6131 = n7594 & n7595;
  assign n6319 = n7596 & n7597;
  assign n5217 = n7598 & n7599;
  assign n6189 = n7600 & n7601;
  assign n5183 = n7602 & n7603;
  assign n6350 = n7604 & n7605;
  assign n5161 = n7606 & n7607;
  assign n6298 = n7608 & n7609;
  assign n3888 = n7610 & n7611;
  assign n5227 = n7612 & n7613;
  assign n6297 = n7614 & n7615;
  assign n6097 = n7616 & n7617;
  assign n5090 = n7618 & n7619;
  assign n6101 = n7620 & n7621;
  assign n6281 = n7622 & n7623;
  assign n5181 = n7624 & n7625;
  assign n6357 = n7626 & n7627;
  assign n6309 = n7628 & n7629;
  assign n5191 = n7630 & n7631;
  assign n6349 = n7632 & n7633;
  assign n6336 = n7634 & n7635;
  assign n6335 = n7636 & n7637;
  assign n5040 = n7638 & n7639;
  assign n5321 = n7640 & n7641;
  assign n6323 = n7642 & n7643;
  assign n6190 = n7644 & n7645;
  assign n6426 = n7646 & n7647;
  assign n6325 = n7648 & n7649;
  assign n6345 = n7650 & n7651;
  assign n5201 = n7652 & n7653;
  assign n6330 = n7654 & n7655;
  assign n5231 = n7656 & n7657;
  assign n6329 = n7658 & n7659;
  assign n6364 = n7660 & n7661;
  assign n6382 = n7662 & n7663;
  assign n6363 = n7664 & n7665;
  assign n6378 = n7666 & n7667;
  assign n6136 = n7668 & n7669;
  assign n6365 = n7670 & n7671;
  assign n6148 = n7672 & n7673;
  assign n4974 = n7674 & n7675;
  assign n6284 = n7676 & n7677;
  assign n5233 = n7678 & n7679;
  assign n6283 = n7680 & n7681;
  assign n6328 = n7682 & n7683;
  assign n6377 = n7684 & n7685;
  assign n5223 = n7686 & n7687;
  assign n5215 = n7688 & n7689;
  assign n6372 = n7690 & n7691;
  assign n6337 = n7692 & n7693;
  assign n6356 = n7694 & n7695;
  assign n5271 = n7696 & n7697;
  assign n5213 = n7698 & n7699;
  assign n6108 = n7700 & n7701;
  assign n6399 = n7702 & n7703;
  assign n6107 = n7704 & n7705;
  assign n6407 = n7706 & n7707;
  assign n5275 = n7708 & n7709;
  assign n6344 = n7710 & n7711;
  assign n4994 = n7712 & n7713;
  assign n6367 = n7714 & n7715;
  assign n6412 = n7716 & n7717;
  assign n5221 = n7718 & n7719;
  assign n6185 = n7720 & n7721;
  assign n6370 = n7722 & n7723;
  assign n6369 = n7724 & n7725;
  assign n5319 = n7726 & n7727;
  assign n6414 = n7728 & n7729;
  assign n5297 = n7730 & n7731;
  assign n6383 = n7732 & n7733;
  assign n6310 = n7734 & n7735;
  assign n6103 = n7736 & n7737;
  assign n3898 = n7738 & n7739;
  assign n5030 = n7740 & n7741;
  assign n5293 = n7742 & n7743;
  assign n6143 = n7744 & n7745;
  assign n6157 = n7746 & n7747;
  assign n5000 = n7748 & n7749;
  assign n5211 = n7750 & n7751;
  assign n6419 = n7752 & n7753;
  assign n6374 = n7754 & n7755;
  assign n6373 = n7756 & n7757;
  assign n6417 = n7758 & n7759;
  assign n5239 = n7760 & n7761;
  assign n5245 = n7762 & n7763;
  assign n6361 = n7764 & n7765;
  assign n5106 = n7766 & n7767;
  assign n6269 = n7768 & n7769;
  assign n5247 = n7770 & n7771;
  assign n6128 = n7772 & n7773;
  assign n6387 = n7774 & n7775;
  assign n6165 = n7776 & n7777;
  assign n6376 = n7778 & n7779;
  assign n6375 = n7780 & n7781;
  assign n6117 = n7782 & n7783;
  assign n6115 = n7784 & n7785;
  assign n6060 = n7786 & n7787;
  assign n5167 = n7788 & n7789;
  assign n6403 = n7790 & n7791;
  assign n6096 = n7792 & n7793;
  assign n6079 = n7794 & n7795;
  assign n6327 = n7796 & n7797;
  assign n5146 = n7798 & n7799;
  assign n6394 = n7800 & n7801;
  assign n6393 = n7802 & n7803;
  assign n5008 = n7804 & n7805;
  assign n5279 = n7806 & n7807;
  assign n6416 = n7808 & n7809;
  assign n6073 = n7810 & n7811;
  assign n6095 = n7812 & n7813;
  assign n6392 = n7814 & n7815;
  assign n6391 = n7816 & n7817;
  assign n6431 = n7818 & n7819;
  assign n6132 = n7820 & n7821;
  assign n5006 = n7822 & n7823;
  assign n6396 = n7824 & n7825;
  assign n6390 = n7826 & n7827;
  assign n5251 = n7828 & n7829;
  assign n6061 = n7830 & n7831;
  assign n6100 = n7832 & n7833;
  assign n6398 = n7834 & n7835;
  assign n6099 = n7836 & n7837;
  assign n6397 = n7838 & n7839;
  assign n6085 = n7840 & n7841;
  assign n5229 = n7842 & n7843;
  assign n6440 = n7844 & n7845;
  assign n6439 = n7846 & n7847;
  assign n5155 = n7848 & n7849;
  assign n6438 = n7850 & n7851;
  assign n5014 = n7852 & n7853;
  assign n6433 = n7854 & n7855;
  assign n6437 = n7856 & n7857;
  assign n6413 = n7858 & n7859;
  assign n5303 = n7860 & n7861;
  assign n6116 = n7862 & n7863;
  assign n6075 = n7864 & n7865;
  assign n5012 = n7866 & n7867;
  assign n6402 = n7868 & n7869;
  assign n6401 = n7870 & n7871;
  assign n6379 = n7872 & n7873;
  assign n6339 = n7874 & n7875;
  assign n6288 = n7876 & n7877;
  assign n5078 = n7878 & n7879;
  assign n6287 = n7880 & n7881;
  assign n5267 = n7882 & n7883;
  assign n6083 = n7884 & n7885;
  assign n6104 = n7886 & n7887;
  assign n6305 = n7888 & n7889;
  assign n5283 = n7890 & n7891;
  assign n6275 = n7892 & n7893;
  assign n6321 = n7894 & n7895;
  assign n4998 = n7896 & n7897;
  assign n5287 = n7898 & n7899;
  assign n6105 = n7900 & n7901;
  assign n6405 = n7902 & n7903;
  assign n6366 = n7904 & n7905;
  assign n6429 = n7906 & n7907;
  assign n5289 = n7908 & n7909;
  assign n5243 = n7910 & n7911;
  assign n6388 = n7912 & n7913;
  assign n6124 = n7914 & n7915;
  assign n6436 = n7916 & n7917;
  assign n6435 = n7918 & n7919;
  assign n6293 = n7920 & n7921;
  assign n5026 = n7922 & n7923;
  assign n6432 = n7924 & n7925;
  assign n5032 = n7926 & n7927;
  assign n6110 = n7928 & n7929;
  assign n6262 = n7930 & n7931;
  assign n6109 = n7932 & n7933;
  assign n6331 = n7934 & n7935;
  assign n4990 = n7936 & n7937;
  assign n6145 = n7938 & n7939;
  assign n6251 = n7940 & n7941;
  assign n4988 = n7942 & n7943;
  assign n6112 = n7944 & n7945;
  assign n6081 = n7946 & n7947;
  assign n6111 = n7948 & n7949;
  assign n6434 = n7950 & n7951;
  assign n6212 = n7952 & n7953;
  assign n5054 = n7954 & n7955;
  assign n6053 = n7956 & n7957;
  assign n6088 = n7958 & n7959;
  assign n5080 = n7960 & n7961;
  assign n6087 = n7962 & n7963;
  assign n6120 = n7964 & n7965;
  assign n5235 = n7966 & n7967;
  assign n5301 = n7968 & n7969;
  assign n12375 = n7971 ^ n7972;
  assign n7021 = n7973 & n7974;
  assign n5362 = ~n7975;
  assign n5458 = ~n7976;
  assign n7006 = n7977 ^ n7978;
  assign n4431 = n7979 ^ n7980;
  assign n4435 = n7981 ^ n7982;
  assign n4983 = n7983 ^ n7984;
  assign n4349 = n7985 ^ n7986;
  assign n3906 = n7987 ^ n7988;
  assign n4987 = n7998 ^ n7999;
  assign n6080 = n8000 ^ n8001;
  assign n4979 = n8002 ^ n8003;
  assign n7970 = n8005 & n8006;
  assign n7989 = n9677 & n6360;
  assign n6048 = n7972 & n7971;
  assign n7008 = ~n9678;
  assign n6462 = ~n9679;
  assign n6458 = ~n9680;
  assign n6207 = n9681 & n7983;
  assign n4946 = n9682 & n7977;
  assign n7993 = n9683 & n9684;
  assign n6670 = ~n9685;
  assign n6395 = n9686 & n7998;
  assign n6628 = ~n9687;
  assign n5241 = n9688 & n7985;
  assign n6452 = ~n9689;
  assign n5048 = n9690 & n7981;
  assign n4006 = n9691 & n8000;
  assign n6646 = ~n9694;
  assign n7995 = n9695 & n9670;
  assign n6089 = n9696 & n8002;
  assign n7996 = n9697 & n9672;
  assign n7994 = n9698 & n9676;
  assign n5295 = n9699 & n7987;
  assign n6658 = ~n9700;
  assign n7992 = n9701 & n9188;
  assign n6484 = ~n9702;
  assign n7991 = n9703 & n9704;
  assign n7997 = n9705 & n9706;
  assign n7990 = n9707 & n9674;
  assign n5018 = n9708 & n7979;
  assign n5348 = ~n9951;
  assign n3928 = n33 ^ n6049;
  assign n4429 = n6050 ^ n6051;
  assign n3916 = n6052 ^ n4963;
  assign n3902 = n6053 ^ n6054;
  assign n3908 = n6055 ^ n3892;
  assign n3912 = n6056 ^ n3894;
  assign n3914 = n6057 ^ n4136;
  assign n3920 = n6058 ^ n4139;
  assign n3922 = n6059 ^ n4967;
  assign n3930 = n6060 ^ n4974;
  assign n3932 = n6061 ^ n6049;
  assign n4433 = n33 ^ n6062;
  assign n3296 = n6063 ^ n6064;
  assign n4977 = n6065 ^ n6066;
  assign n4427 = n6067 ^ n6068;
  assign n3904 = n6069 ^ n6070;
  assign n4516 = n6071 ^ n6072;
  assign n3243 = n6073 ^ n6074;
  assign n4523 = n6075 ^ n6076;
  assign n3326 = n6077 ^ n6078;
  assign n4437 = n6079 ^ n6080;
  assign n4989 = n6081 ^ n6082;
  assign n4993 = n6083 ^ n6084;
  assign n5230 = n6085 ^ n6086;
  assign n4997 = n6087 ^ n6088;
  assign n4976 = n6089 ^ n6090;
  assign n5001 = n6091 ^ n6092;
  assign n5154 = n6093 ^ n6094;
  assign n5009 = n6095 ^ n6096;
  assign n5011 = n6097 ^ n6098;
  assign n5015 = n6099 ^ n6100;
  assign n4978 = n6101 ^ n6102;
  assign n5031 = n6103 ^ n6104;
  assign n4965 = n6105 ^ n6106;
  assign n5214 = n6107 ^ n6108;
  assign n5033 = n6109 ^ n6110;
  assign n5021 = n6111 ^ n6112;
  assign n5019 = n6113 ^ n6114;
  assign n5306 = n6115 ^ n6116;
  assign n5037 = n6117 ^ n6118;
  assign n5025 = n6119 ^ n6120;
  assign n5029 = n6121 ^ n6122;
  assign n5027 = n6123 ^ n6124;
  assign n5292 = n6125 ^ n6126;
  assign n5039 = n6127 ^ n6128;
  assign n4980 = n6129 ^ n6130;
  assign n5043 = n6131 ^ n6132;
  assign n5045 = n6133 ^ n6134;
  assign n5047 = n6135 ^ n6136;
  assign n5160 = n6137 ^ n6138;
  assign n5049 = n6139 ^ n6140;
  assign n5051 = n6141 ^ n6142;
  assign n4968 = n6143 ^ n6144;
  assign n5053 = n6145 ^ n6146;
  assign n5055 = n6147 ^ n6148;
  assign n5007 = n6149 ^ n6150;
  assign n5023 = n6151 ^ n6152;
  assign n5059 = n6153 ^ n6154;
  assign n5061 = n6155 ^ n6156;
  assign n4966 = n6157 ^ n6158;
  assign n5063 = n6159 ^ n6160;
  assign n5065 = n6161 ^ n6162;
  assign n5067 = n6163 ^ n6164;
  assign n5057 = n6165 ^ n6166;
  assign n5174 = n6167 ^ n6168;
  assign n5071 = n6169 ^ n6170;
  assign n5069 = n6171 ^ n6172;
  assign n5073 = n6173 ^ n6174;
  assign n5075 = n6175 ^ n6176;
  assign n5077 = n6177 ^ n6178;
  assign n5017 = n6179 ^ n6180;
  assign n4982 = n6181 ^ n6182;
  assign n4969 = n6183 ^ n6184;
  assign n5081 = n6185 ^ n6186;
  assign n5083 = n6187 ^ n6188;
  assign n5184 = n6189 ^ n6190;
  assign n5087 = n6191 ^ n6192;
  assign n5085 = n6193 ^ n6194;
  assign n5089 = n6195 ^ n6196;
  assign n5091 = n6197 ^ n6198;
  assign n5093 = n6199 ^ n6200;
  assign n5095 = n6201 ^ n6202;
  assign n4970 = n6203 ^ n6204;
  assign n5097 = n6205 ^ n6206;
  assign n3910 = n6207 ^ n6208;
  assign n5099 = n6209 ^ n6210;
  assign n4981 = n6211 ^ n6212;
  assign n5101 = n6213 ^ n6214;
  assign n5103 = n6215 ^ n6216;
  assign n5105 = n6217 ^ n6218;
  assign n5141 = n6219 ^ n6220;
  assign n5107 = n6221 ^ n6222;
  assign n5109 = n6223 ^ n6224;
  assign n5111 = n6225 ^ n6226;
  assign n5115 = n6227 ^ n6228;
  assign n5113 = n6229 ^ n6230;
  assign n5117 = n6231 ^ n6232;
  assign n5119 = n6233 ^ n6234;
  assign n5123 = n6235 ^ n6236;
  assign n5121 = n6237 ^ n6238;
  assign n5127 = n6239 ^ n6240;
  assign n5125 = n6241 ^ n6242;
  assign n5003 = n6243 ^ n6244;
  assign n5129 = n6245 ^ n6246;
  assign n4964 = n6247 ^ n6248;
  assign n5131 = n6249 ^ n6250;
  assign n5035 = n6251 ^ n6252;
  assign n5135 = n6253 ^ n6254;
  assign n5137 = n6255 ^ n6256;
  assign n5143 = n6257 ^ n6258;
  assign n5145 = n6259 ^ n6260;
  assign n5149 = n6261 ^ n6262;
  assign n5153 = n6263 ^ n6264;
  assign n5151 = n6265 ^ n6266;
  assign n3918 = n6267 ^ n6268;
  assign n5139 = n6269 ^ n6270;
  assign n5158 = n6271 ^ n6272;
  assign n5156 = n6273 ^ n6274;
  assign n5162 = n6275 ^ n6276;
  assign n5166 = n6277 ^ n6278;
  assign n5170 = n6279 ^ n6280;
  assign n5182 = n6281 ^ n6282;
  assign n4984 = n6283 ^ n6284;
  assign n4999 = n6285 ^ n6286;
  assign n5268 = n6287 ^ n6288;
  assign n5178 = n6289 ^ n6290;
  assign n5172 = n6291 ^ n6292;
  assign n5164 = n6293 ^ n6294;
  assign n5180 = n6295 ^ n6296;
  assign n5188 = n6297 ^ n6298;
  assign n5186 = n6299 ^ n6300;
  assign n5176 = n6301 ^ n6302;
  assign n5190 = n6303 ^ n6304;
  assign n5284 = n6305 ^ n6306;
  assign n5262 = n6307 ^ n6308;
  assign n5192 = n6309 ^ n6310;
  assign n4985 = n6311 ^ n6312;
  assign n5194 = n6313 ^ n6314;
  assign n5196 = n6315 ^ n6316;
  assign n5198 = n6317 ^ n6318;
  assign n5041 = n6319 ^ n6320;
  assign n5168 = n6321 ^ n6322;
  assign n5200 = n6323 ^ n6324;
  assign n5202 = n6325 ^ n6326;
  assign n5147 = n6327 ^ n6328;
  assign n5204 = n6329 ^ n6330;
  assign n4991 = n6331 ^ n6332;
  assign n5208 = n6333 ^ n6334;
  assign n5210 = n6335 ^ n6336;
  assign n5212 = n6337 ^ n6338;
  assign n5216 = n6339 ^ n6340;
  assign n5218 = n6341 ^ n6342;
  assign n5256 = n6343 ^ n6344;
  assign n5013 = n6345 ^ n6346;
  assign n5005 = n6347 ^ n6348;
  assign n4971 = n6349 ^ n6350;
  assign n5224 = n6351 ^ n6352;
  assign n5226 = n6353 ^ n6354;
  assign n5220 = n6355 ^ n6356;
  assign n5228 = n6357 ^ n6358;
  assign n5133 = n6359 ^ n6360;
  assign n5248 = n6361 ^ n6362;
  assign n5232 = n6363 ^ n6364;
  assign n5234 = n6365 ^ n6366;
  assign n5222 = n6367 ^ n6368;
  assign n5238 = n6369 ^ n6370;
  assign n5240 = n6371 ^ n6372;
  assign n5290 = n6373 ^ n6374;
  assign n5242 = n6375 ^ n6376;
  assign n4973 = n6377 ^ n6378;
  assign n5079 = n6379 ^ n6380;
  assign n5298 = n6381 ^ n6382;
  assign n4975 = n6383 ^ n6384;
  assign n5250 = n6385 ^ n6386;
  assign n5254 = n6387 ^ n6388;
  assign n5286 = n6389 ^ n6390;
  assign n5258 = n6391 ^ n6392;
  assign n5260 = n6393 ^ n6394;
  assign n3926 = n6395 ^ n6396;
  assign n5300 = n6397 ^ n6398;
  assign n5236 = n6399 ^ n6400;
  assign n5264 = n6401 ^ n6402;
  assign n5270 = n6403 ^ n6404;
  assign n5274 = n6405 ^ n6406;
  assign n5272 = n6407 ^ n6408;
  assign n5244 = n6409 ^ n6410;
  assign n5276 = n6411 ^ n6412;
  assign n5278 = n6413 ^ n6414;
  assign n5280 = n6415 ^ n6416;
  assign n5246 = n6417 ^ n6418;
  assign n5282 = n6419 ^ n6420;
  assign n4995 = n6421 ^ n6422;
  assign n5266 = n6423 ^ n6424;
  assign n5288 = n6425 ^ n6426;
  assign n5206 = n6427 ^ n6428;
  assign n5294 = n6429 ^ n6430;
  assign n5296 = n6431 ^ n6432;
  assign n5252 = n6433 ^ n6434;
  assign n5302 = n6435 ^ n6436;
  assign n5304 = n6437 ^ n6438;
  assign n4986 = n6439 ^ n6440;
  assign n6720 = n6222 & n6956;
  assign n6722 = n6172 & n6957;
  assign n6724 = n5189 & n6958;
  assign n6725 = n6159 & n6959;
  assign n6729 = n5012 & n6960;
  assign n6730 = n4136 & n6961;
  assign n6731 = n6228 & n6962;
  assign n6737 = n6241 & n6965;
  assign n6741 = n6424 & n6966;
  assign n6746 = n6302 & n6967;
  assign n6749 = n6248 & n6968;
  assign n6750 = n6319 & n6969;
  assign n6752 = n6191 & n6970;
  assign n6754 = n6197 & n6971;
  assign n6757 = n6274 & n6972;
  assign n6758 = n5122 & n6973;
  assign n6760 = n6259 & n6974;
  assign n6762 = n6386 & n6975;
  assign n6763 = n6168 & n6976;
  assign n6764 = n6316 & n6977;
  assign n6772 = n6307 & n6979;
  assign n6773 = n6351 & n6980;
  assign n6775 = n4967 & n6981;
  assign n6777 = n6281 & n6982;
  assign n6778 = n5227 & n6983;
  assign n6779 = n6336 & n6984;
  assign n6780 = n6427 & n6985;
  assign n6783 = n6339 & n6986;
  assign n6790 = n6414 & n6988;
  assign n6791 = n6251 & n6989;
  assign n6792 = n6188 & n6990;
  assign n6793 = n6405 & n6991;
  assign n6796 = n5269 & n6992;
  assign n6800 = n6091 & n6994;
  assign n6802 = n5036 & n6995;
  assign n6808 = n6150 & n6996;
  assign n6810 = n6398 & n6997;
  assign n6811 = n6165 & n6998;
  assign n6814 = n6426 & n6999;
  assign n6815 = n6122 & n7000;
  assign n6818 = n6146 & n7002;
  assign n6819 = n4988 & n7003;
  assign n6822 = n6062 & n7004;
  assign n6823 = n6049 & n7004;
  assign n6824 = n6185 & n6186;
  assign n6825 = n6119 & n6120;
  assign n6826 = n6223 & n6224;
  assign n6827 = n6098 & n5010;
  assign n6828 = n5002 & n6244;
  assign n6829 = n6435 & n6436;
  assign n6830 = n3896 & n6384;
  assign n6831 = n6153 & n6154;
  assign n6832 = n6135 & n6136;
  assign n6833 = n6133 & n6134;
  assign n6834 = n6102 & n4979;
  assign n6835 = n6155 & n6156;
  assign n6836 = n7005 & n7006;
  assign n6837 = n6189 & n6190;
  assign n6838 = n6125 & n6126;
  assign n6839 = n5050 & n6142;
  assign n6840 = n6193 & n6194;
  assign n6841 = n6229 & n6230;
  assign n6842 = n6337 & n6338;
  assign n6843 = n6416 & n5279;
  assign n6844 = n6162 & n5064;
  assign n6845 = n6051 & n6050;
  assign n6846 = n6175 & n6176;
  assign n6847 = n6058 & n4139;
  assign n6848 = n6177 & n6178;
  assign n6849 = n6163 & n6164;
  assign n6850 = n6169 & n6170;
  assign n6851 = n6173 & n6174;
  assign n6852 = n3892 & n6055;
  assign n6853 = n6213 & n6214;
  assign n6854 = n6226 & n5110;
  assign n6855 = n6209 & n6210;
  assign n6856 = n6215 & n6216;
  assign n6857 = n6201 & n6202;
  assign n6858 = n6289 & n6290;
  assign n6859 = n6182 & n4983;
  assign n6860 = n5128 & n6246;
  assign n6861 = n6240 & n5126;
  assign n6862 = n6421 & n6422;
  assign n6863 = n6254 & n5134;
  assign n6864 = n6348 & n5004;
  assign n6865 = n6233 & n6234;
  assign n6866 = n4174 & n6204;
  assign n6867 = n6061 & n6049;
  assign n6868 = n6255 & n6256;
  assign n6869 = n3894 & n6056;
  assign n6870 = n6300 & n5185;
  assign n6871 = n6205 & n6206;
  assign n6872 = n6196 & n5088;
  assign n6873 = n6292 & n5171;
  assign n6874 = n6218 & n5104;
  assign n6875 = n6231 & n6232;
  assign n6876 = n6279 & n6280;
  assign n6877 = n6237 & n6238;
  assign n6878 = n6295 & n6296;
  assign n6879 = n6129 & n6130;
  assign n6880 = n6249 & n6250;
  assign n6881 = n6318 & n5197;
  assign n6882 = n6199 & n6200;
  assign n6883 = n6261 & n6262;
  assign n6884 = n6258 & n5142;
  assign n6885 = n6179 & n6180;
  assign n6886 = n6305 & n6306;
  assign n6887 = n6263 & n6264;
  assign n6888 = n6137 & n6138;
  assign n6889 = n6276 & n5161;
  assign n6890 = n6334 & n5207;
  assign n6891 = n5165 & n6278;
  assign n6892 = n6354 & n5225;
  assign n6893 = n6271 & n6272;
  assign n6894 = n6287 & n6288;
  assign n6895 = n6313 & n6314;
  assign n6896 = n6341 & n6342;
  assign n6897 = n6111 & n6112;
  assign n6898 = n6298 & n5187;
  assign n6899 = n6356 & n5219;
  assign n6900 = n6309 & n6310;
  assign n6901 = n6054 & n6350;
  assign n6902 = n6323 & n6324;
  assign n6903 = n6325 & n6326;
  assign n6904 = n6330 & n5203;
  assign n6905 = n6364 & n5231;
  assign n6906 = n6151 & n6152;
  assign n6907 = n6283 & n6284;
  assign n6908 = n4974 & n6378;
  assign n6909 = n6409 & n6410;
  assign n6910 = n6108 & n5213;
  assign n6911 = n6399 & n6400;
  assign n6912 = n5271 & n6408;
  assign n6913 = n6088 & n4996;
  assign n6914 = n6367 & n6368;
  assign n6915 = n6369 & n6370;
  assign n6916 = n6412 & n5275;
  assign n6917 = n6372 & n5239;
  assign n6918 = n6103 & n6104;
  assign n6919 = n6420 & n5281;
  assign n6920 = n6373 & n6374;
  assign n6921 = n6417 & n6418;
  assign n6922 = n6361 & n6362;
  assign n6923 = n6079 & n6080;
  assign n6924 = n6327 & n6328;
  assign n6925 = n6393 & n6394;
  assign n6926 = n5008 & n6096;
  assign n6927 = n6128 & n5038;
  assign n6928 = n6285 & n6286;
  assign n6929 = n6390 & n5285;
  assign n6930 = n6085 & n6086;
  assign n6931 = n6099 & n6100;
  assign n6932 = n6440 & n4987;
  assign n6933 = n6115 & n6116;
  assign n6934 = n6131 & n6132;
  assign n6935 = n6381 & n6382;
  assign n6936 = n6437 & n6438;
  assign n6937 = n6401 & n6402;
  assign n6938 = n3898 & n6144;
  assign n6939 = n6379 & n6380;
  assign n6940 = n6083 & n6084;
  assign n6941 = n6321 & n6322;
  assign n6942 = n6430 & n5293;
  assign n6943 = n6433 & n6434;
  assign n6944 = n6365 & n6366;
  assign n6945 = n6123 & n6124;
  assign n6946 = n6110 & n5032;
  assign n6947 = n6331 & n6332;
  assign n6948 = n6391 & n6392;
  assign n6949 = n6265 & n6266;
  assign n6950 = n6147 & n6148;
  assign n6951 = n6387 & n6388;
  assign n5741 = ~n6411;
  assign n6821 = ~n4967;
  assign n6586 = ~n6418;
  assign n6713 = ~n6094;
  assign n6627 = ~n6071;
  assign n6445 = ~n6348;
  assign n5753 = ~n5273;
  assign n5529 = ~n6347;
  assign n6608 = ~n6408;
  assign n5527 = ~n6243;
  assign n6804 = ~n6140;
  assign n6455 = ~n6223;
  assign n6699 = ~n6051;
  assign n6817 = ~n6146;
  assign n4346 = ~n4139;
  assign n6472 = ~n6230;
  assign n6742 = ~n5189;
  assign n3728 = ~n4174;
  assign n4347 = ~n4136;
  assign n4348 = ~n3894;
  assign n6542 = ~n6296;
  assign n4972 = ~n6054;
  assign n6626 = ~n5038;
  assign n4122 = ~n3896;
  assign n6465 = ~n6063;
  assign n5557 = ~n6187;
  assign n6599 = ~n6421;
  assign n6441 = ~n6129;
  assign n6709 = ~n6049;
  assign n5817 = ~n5301;
  assign n4126 = ~n3890;
  assign n6449 = ~n6179;
  assign n6463 = ~n6193;
  assign n5533 = ~n5016;
  assign n5535 = ~n5058;
  assign n6715 = ~n6114;
  assign n5537 = ~n6113;
  assign n6553 = ~n6265;
  assign n5539 = ~n5046;
  assign n6487 = ~n6098;
  assign n6714 = ~n6197;
  assign n6716 = ~n6106;
  assign n6457 = ~n6065;
  assign n6794 = ~n5269;
  assign n6520 = ~n6134;
  assign n6519 = ~n6133;
  assign n6717 = ~n6090;
  assign n6693 = ~n6102;
  assign n6468 = ~n6156;
  assign n6461 = ~n6359;
  assign n5551 = ~n5060;
  assign n6450 = ~n6180;
  assign n6650 = ~n5285;
  assign n6719 = ~n6062;
  assign n6453 = ~n6153;
  assign n6469 = ~n6135;
  assign n6806 = ~n6222;
  assign n6478 = ~n6126;
  assign n5561 = ~n6141;
  assign n6596 = ~n5203;
  assign n6467 = ~n6155;
  assign n6475 = ~n5050;
  assign n6451 = ~n6069;
  assign n6701 = ~n6058;
  assign n6476 = ~n6142;
  assign n5671 = ~n5108;
  assign n6447 = ~n6285;
  assign n5545 = ~n5042;
  assign n5775 = ~n6415;
  assign n6479 = ~n6151;
  assign n5789 = ~n6389;
  assign n5567 = ~n5112;
  assign n6678 = ~n6186;
  assign n5687 = ~n5205;
  assign n6471 = ~n6229;
  assign n5565 = ~n5022;
  assign n6480 = ~n6152;
  assign n6442 = ~n6130;
  assign n6456 = ~n6224;
  assign n5765 = ~n5253;
  assign n6738 = ~n6122;
  assign n5773 = ~n5259;
  assign n6744 = ~n6172;
  assign n6448 = ~n6286;
  assign n5711 = ~n5199;
  assign n5569 = ~n6171;
  assign n6482 = ~n5064;
  assign n5779 = ~n5257;
  assign n5803 = ~n5263;
  assign n6481 = ~n6162;
  assign n6483 = ~n6067;
  assign n5571 = ~n6161;
  assign n5725 = ~n6355;
  assign n6486 = ~n6176;
  assign n6498 = ~n6290;
  assign n6485 = ~n6175;
  assign n6671 = ~n6430;
  assign n5575 = ~n5074;
  assign n6723 = ~n6159;
  assign n6687 = ~n6119;
  assign n5577 = ~n5062;
  assign n5573 = ~n6303;
  assign n6623 = ~n6420;
  assign n6726 = ~n6184;
  assign n6488 = ~n5010;
  assign n5783 = ~n6127;
  assign n6546 = ~n6238;
  assign n6490 = ~n6164;
  assign n6489 = ~n6163;
  assign n6492 = ~n6178;
  assign n6491 = ~n6177;
  assign n5367 = ~n6183;
  assign n5579 = ~n5076;
  assign n5581 = ~n5066;
  assign n6494 = ~n6170;
  assign n6493 = ~n6169;
  assign n5583 = ~n5070;
  assign n6496 = ~n6174;
  assign n6495 = ~n6173;
  assign n6660 = ~n6380;
  assign n6728 = ~n6228;
  assign n6624 = ~n5281;
  assign n5585 = ~n5072;
  assign n6781 = ~n6091;
  assign n4345 = ~n3892;
  assign n5587 = ~n5114;
  assign n6702 = ~n6055;
  assign n6727 = ~n6424;
  assign n6500 = ~n5110;
  assign n6502 = ~n6214;
  assign n6501 = ~n6213;
  assign n6499 = ~n6226;
  assign n5589 = ~n5100;
  assign n6504 = ~n6210;
  assign n5591 = ~n6225;
  assign n6503 = ~n6209;
  assign n5593 = ~n5098;
  assign n6732 = ~n6241;
  assign n6506 = ~n6216;
  assign n6497 = ~n6289;
  assign n6505 = ~n6215;
  assign n5595 = ~n5102;
  assign n5597 = ~n5124;
  assign n6734 = ~n6208;
  assign n6510 = ~n6202;
  assign n6509 = ~n6201;
  assign n5599 = ~n5094;
  assign n5601 = ~n5177;
  assign n6514 = ~n6246;
  assign n6508 = ~n6338;
  assign n6555 = ~n6409;
  assign n5653 = ~n6317;
  assign n5799 = ~n5305;
  assign n6590 = ~n6324;
  assign n6691 = ~n6182;
  assign n6516 = ~n5126;
  assign n5605 = ~n6245;
  assign n5607 = ~n6181;
  assign n6515 = ~n6240;
  assign n5609 = ~n6239;
  assign n5563 = ~n5291;
  assign n5603 = ~n5265;
  assign n6518 = ~n5134;
  assign n5523 = ~n5024;
  assign n6766 = ~n6312;
  assign n6739 = ~n6302;
  assign n6517 = ~n6254;
  assign n5559 = ~n5044;
  assign n5613 = ~n6253;
  assign n6443 = ~n5002;
  assign n6669 = ~n6077;
  assign n6587 = ~n6123;
  assign n6695 = ~n7005;
  assign n6805 = ~n6150;
  assign n6637 = ~n6381;
  assign n5615 = ~n6301;
  assign n6743 = ~n6220;
  assign n6522 = ~n6234;
  assign n6521 = ~n6233;
  assign n5617 = ~n5118;
  assign n6524 = ~n6256;
  assign n6523 = ~n6255;
  assign n5619 = ~n5136;
  assign n5665 = ~n4992;
  assign n6747 = ~n6248;
  assign n5625 = ~n5086;
  assign n6751 = ~n6191;
  assign n5841 = ~n4963;
  assign n6748 = ~n6059;
  assign n6533 = ~n6196;
  assign n5627 = ~n6195;
  assign n5749 = ~n5034;
  assign n5633 = ~n5092;
  assign n6526 = ~n5185;
  assign n6703 = ~n6056;
  assign n6540 = ~n6200;
  assign n6525 = ~n6300;
  assign n6539 = ~n6199;
  assign n5727 = ~n6121;
  assign n5611 = ~n6139;
  assign n6528 = ~n6206;
  assign n5621 = ~n6299;
  assign n6527 = ~n6205;
  assign n5623 = ~n5096;
  assign n6530 = ~n6280;
  assign n6532 = ~n5171;
  assign n6531 = ~n6292;
  assign n6529 = ~n6279;
  assign n6538 = ~n5104;
  assign n5429 = ~n6203;
  assign n5629 = ~n6291;
  assign n6537 = ~n6218;
  assign n5631 = ~n6217;
  assign n5635 = ~n5169;
  assign n4441 = ~n4941;
  assign n6543 = ~n6231;
  assign n5637 = ~n5116;
  assign n6541 = ~n6295;
  assign n6545 = ~n6237;
  assign n5787 = ~n5056;
  assign n5639 = ~n5120;
  assign n5641 = ~n5179;
  assign n6755 = ~n6274;
  assign n6753 = ~n6386;
  assign n5743 = ~n5237;
  assign n6756 = ~n5122;
  assign n5647 = ~n6235;
  assign n6548 = ~n5197;
  assign n6552 = ~n6250;
  assign n5699 = ~n5084;
  assign n6454 = ~n6154;
  assign n6551 = ~n6249;
  assign n6712 = ~n6188;
  assign n6536 = ~n6322;
  assign n6547 = ~n6318;
  assign n6513 = ~n5128;
  assign n6652 = ~n6086;
  assign n5649 = ~n5130;
  assign n5310 = ~n5140;
  assign n6733 = ~n6259;
  assign n5655 = ~n5144;
  assign n6610 = ~n6400;
  assign n5651 = ~n6385;
  assign n6554 = ~n6266;
  assign n6759 = ~n6316;
  assign n5657 = ~n5150;
  assign n6557 = ~n6261;
  assign n5314 = ~n5255;
  assign n5659 = ~n5148;
  assign n5661 = ~n5195;
  assign n6559 = ~n6258;
  assign n5663 = ~n6257;
  assign n6666 = ~n6306;
  assign n6761 = ~n6168;
  assign n5667 = ~n6167;
  assign n6556 = ~n6410;
  assign n6562 = ~n6264;
  assign n6561 = ~n6263;
  assign n6795 = ~n5036;
  assign n6767 = ~n6268;
  assign n6600 = ~n6422;
  assign n6564 = ~n5225;
  assign n6745 = ~n6307;
  assign n6768 = ~n6052;
  assign n6566 = ~n6138;
  assign n6565 = ~n6137;
  assign n6563 = ~n6354;
  assign n6568 = ~n5207;
  assign n6567 = ~n6334;
  assign n5675 = ~n5159;
  assign n6664 = ~n6084;
  assign n6569 = ~n6276;
  assign n5673 = ~n6353;
  assign n5677 = ~n6333;
  assign n5683 = ~n5261;
  assign n6571 = ~n5165;
  assign n5681 = ~n6277;
  assign n5689 = ~n5193;
  assign n5745 = ~n6371;
  assign n6574 = ~n6272;
  assign n6573 = ~n6271;
  assign n6770 = ~n6427;
  assign n5685 = ~n5157;
  assign n6632 = ~n6362;
  assign n6771 = ~n6351;
  assign n6681 = ~n6147;
  assign n6576 = ~n6314;
  assign n6575 = ~n6313;
  assign n6464 = ~n6194;
  assign n6578 = ~n6342;
  assign n6477 = ~n6125;
  assign n6577 = ~n6341;
  assign n6549 = ~n6131;
  assign n6769 = ~n6319;
  assign n5691 = ~n5217;
  assign n6579 = ~n6189;
  assign n5833 = ~n5020;
  assign n5693 = ~n5183;
  assign n6705 = ~n6350;
  assign n6570 = ~n5161;
  assign n6581 = ~n6298;
  assign n4124 = ~n3888;
  assign n6774 = ~n5227;
  assign n5695 = ~n6297;
  assign n5543 = ~n6097;
  assign n5549 = ~n5090;
  assign n5547 = ~n6101;
  assign n6776 = ~n6281;
  assign n5701 = ~n5181;
  assign n5697 = ~n6357;
  assign n6583 = ~n6309;
  assign n5703 = ~n5191;
  assign n5705 = ~n6349;
  assign n6812 = ~n6336;
  assign n5709 = ~n6335;
  assign n5707 = ~n5040;
  assign n5843 = ~n5321;
  assign n6589 = ~n6323;
  assign n6580 = ~n6190;
  assign n6813 = ~n6426;
  assign n6593 = ~n6325;
  assign n5805 = ~n6345;
  assign n5713 = ~n5201;
  assign n6595 = ~n6330;
  assign n6598 = ~n5231;
  assign n5715 = ~n6329;
  assign n6597 = ~n6364;
  assign n6638 = ~n6382;
  assign n5717 = ~n6363;
  assign n6707 = ~n6378;
  assign n6470 = ~n6136;
  assign n6601 = ~n6365;
  assign n6682 = ~n6148;
  assign n6706 = ~n4974;
  assign n6604 = ~n6284;
  assign n5719 = ~n5233;
  assign n6603 = ~n6283;
  assign n6640 = ~n6328;
  assign n5831 = ~n6377;
  assign n5735 = ~n5223;
  assign n5721 = ~n5215;
  assign n6635 = ~n6372;
  assign n6507 = ~n6337;
  assign n6605 = ~n6356;
  assign n6607 = ~n5271;
  assign n6612 = ~n5213;
  assign n6611 = ~n6108;
  assign n6609 = ~n6399;
  assign n5729 = ~n6107;
  assign n5733 = ~n6407;
  assign n6460 = ~n5275;
  assign n6786 = ~n6344;
  assign n5553 = ~n4994;
  assign n6615 = ~n6367;
  assign n6459 = ~n6412;
  assign n5737 = ~n5221;
  assign n6677 = ~n6185;
  assign n6618 = ~n6370;
  assign n6617 = ~n6369;
  assign n5844 = ~n5319;
  assign n6788 = ~n6414;
  assign n5531 = ~n5297;
  assign n5461 = ~n6383;
  assign n6584 = ~n6310;
  assign n6619 = ~n6103;
  assign n4120 = ~n3898;
  assign n5751 = ~n5030;
  assign n6672 = ~n5293;
  assign n5499 = ~n6143;
  assign n5541 = ~n6157;
  assign n5525 = ~n5000;
  assign n5723 = ~n5211;
  assign n5785 = ~n6419;
  assign n6630 = ~n6374;
  assign n6629 = ~n6373;
  assign n6585 = ~n6417;
  assign n6636 = ~n5239;
  assign n5759 = ~n5245;
  assign n6631 = ~n6361;
  assign n5555 = ~n5106;
  assign n6473 = ~n6269;
  assign n5761 = ~n5247;
  assign n6625 = ~n6128;
  assign n6633 = ~n6387;
  assign n6787 = ~n6165;
  assign n6797 = ~n6376;
  assign n5767 = ~n6375;
  assign n5763 = ~n6117;
  assign n6683 = ~n6115;
  assign n6799 = ~n6060;
  assign n5813 = ~n5167;
  assign n5755 = ~n6403;
  assign n6614 = ~n6096;
  assign n6689 = ~n6079;
  assign n6639 = ~n6327;
  assign n5771 = ~n5146;
  assign n6642 = ~n6394;
  assign n6641 = ~n6393;
  assign n6613 = ~n5008;
  assign n6644 = ~n5279;
  assign n6643 = ~n6416;
  assign n6645 = ~n6073;
  assign n5769 = ~n6095;
  assign n6648 = ~n6392;
  assign n6647 = ~n6391;
  assign n5821 = ~n6431;
  assign n6550 = ~n6132;
  assign n5781 = ~n5006;
  assign n6807 = ~n6396;
  assign n6649 = ~n6390;
  assign n5669 = ~n5251;
  assign n6710 = ~n6061;
  assign n6512 = ~n6100;
  assign n6809 = ~n6398;
  assign n6511 = ~n6099;
  assign n5793 = ~n6397;
  assign n6651 = ~n6085;
  assign n5795 = ~n5229;
  assign n6697 = ~n6440;
  assign n5797 = ~n6439;
  assign n5643 = ~n5155;
  assign n6654 = ~n6438;
  assign n5791 = ~n5014;
  assign n6655 = ~n6433;
  assign n6653 = ~n6437;
  assign n5747 = ~n6413;
  assign n5801 = ~n5303;
  assign n6684 = ~n6116;
  assign n6657 = ~n6075;
  assign n6801 = ~n5012;
  assign n6662 = ~n6402;
  assign n6661 = ~n6401;
  assign n6659 = ~n6379;
  assign n6803 = ~n6339;
  assign n6592 = ~n6288;
  assign n5807 = ~n5078;
  assign n6591 = ~n6287;
  assign n5809 = ~n5267;
  assign n6663 = ~n6083;
  assign n6620 = ~n6104;
  assign n6665 = ~n6305;
  assign n5739 = ~n5283;
  assign n5679 = ~n6275;
  assign n6535 = ~n6321;
  assign n5777 = ~n4998;
  assign n5811 = ~n5287;
  assign n5339 = ~n6105;
  assign n6782 = ~n6405;
  assign n6602 = ~n6366;
  assign n5815 = ~n6429;
  assign n5757 = ~n5289;
  assign n5835 = ~n5243;
  assign n6634 = ~n6388;
  assign n6588 = ~n6124;
  assign n6622 = ~n6436;
  assign n6621 = ~n6435;
  assign n6667 = ~n6293;
  assign n5819 = ~n5026;
  assign n6740 = ~n6432;
  assign n6674 = ~n5032;
  assign n6673 = ~n6110;
  assign n6558 = ~n6262;
  assign n5823 = ~n6109;
  assign n6675 = ~n6331;
  assign n5827 = ~n4990;
  assign n5825 = ~n6145;
  assign n6785 = ~n6251;
  assign n6721 = ~n4988;
  assign n6680 = ~n6112;
  assign n5829 = ~n6081;
  assign n6679 = ~n6111;
  assign n6656 = ~n6434;
  assign n6820 = ~n6212;
  assign n5837 = ~n5054;
  assign n6784 = ~n6053;
  assign n6685 = ~n6088;
  assign n5839 = ~n5080;
  assign n5645 = ~n6087;
  assign n6688 = ~n6120;
  assign n5731 = ~n5235;
  assign n6668 = ~n7021;
  assign n7007 = n6048 & n7008;
  assign n6696 = ~n7006;
  assign n4459 = ~n4431;
  assign n6694 = ~n4979;
  assign n6690 = ~n6080;
  assign n4461 = ~n4435;
  assign n6692 = ~n4983;
  assign n4116 = ~n4349;
  assign n6698 = ~n4987;
  assign n4118 = ~n3906;
  assign n6474 = ~n7970;
  assign n6978 = ~n5018;
  assign n5343 = ~n7989;
  assign n5480 = ~n7990;
  assign n5359 = ~n7991;
  assign n6963 = ~n6207;
  assign n5327 = ~n7992;
  assign n4529 = ~n4946;
  assign n5336 = ~n7993;
  assign n6964 = ~n6395;
  assign n7001 = ~n5295;
  assign n6993 = ~n5241;
  assign n6987 = ~n5048;
  assign n5385 = ~n7994;
  assign n6955 = ~n6089;
  assign n4340 = ~n4006;
  assign n5392 = ~n7995;
  assign n5467 = ~n7996;
  assign n6953 = ~n7997;
  assign n3773 = n4963 ^ n4964;
  assign n4487 = n4965 ^ n3888;
  assign n3221 = n4966 ^ n4967;
  assign n2959 = n4968 ^ n3898;
  assign n3777 = n4969 ^ n4126;
  assign n2703 = n4970 ^ n3728;
  assign n2705 = n4971 ^ n4972;
  assign n2641 = n4973 ^ n4974;
  assign n2637 = n4975 ^ n3896;
  assign n4416 = n4976 ^ n4977;
  assign n4948 = n4978 ^ n4979;
  assign n2870 = n4980 ^ n4981;
  assign n2621 = n4982 ^ n4983;
  assign n4508 = n4984 ^ n4985;
  assign n3787 = n4986 ^ n4987;
  assign n4473 = n4988 ^ n4989;
  assign n4472 = n4990 ^ n4991;
  assign n4229 = n4992 ^ n4993;
  assign n4485 = n4994 ^ n4995;
  assign n3286 = n4996 ^ n4997;
  assign n4469 = n4998 ^ n4999;
  assign n3288 = n5000 ^ n5001;
  assign n2957 = n5002 ^ n5003;
  assign n4225 = n5004 ^ n5005;
  assign n3213 = n5006 ^ n5007;
  assign n4231 = n5008 ^ n5009;
  assign n3841 = n5010 ^ n5011;
  assign n3874 = n5012 ^ n5013;
  assign n4477 = n5014 ^ n5015;
  assign n4486 = n5016 ^ n5017;
  assign n3289 = n5018 ^ n5019;
  assign n4482 = n5020 ^ n5021;
  assign n4484 = n5022 ^ n5023;
  assign n3217 = n5024 ^ n5025;
  assign n3752 = n5026 ^ n5027;
  assign n3547 = n5028 ^ n5029;
  assign n4515 = n5030 ^ n5031;
  assign n4483 = n5032 ^ n5033;
  assign n4470 = n5034 ^ n5035;
  assign n3762 = n5036 ^ n5037;
  assign n3302 = n5038 ^ n5039;
  assign n3844 = n5040 ^ n5041;
  assign n3757 = n5042 ^ n5043;
  assign n4491 = n5044 ^ n5045;
  assign n4490 = n5046 ^ n5047;
  assign n4489 = n5048 ^ n5049;
  assign n4488 = n5050 ^ n5051;
  assign n4236 = n5052 ^ n5053;
  assign n3218 = n5054 ^ n5055;
  assign n3549 = n5056 ^ n5057;
  assign n4421 = n5058 ^ n5059;
  assign n4420 = n5060 ^ n5061;
  assign n4531 = n5062 ^ n5063;
  assign n4530 = n5064 ^ n5065;
  assign n3760 = n5066 ^ n5067;
  assign n3303 = n5068 ^ n5069;
  assign n3759 = n5070 ^ n5071;
  assign n4426 = n5072 ^ n5073;
  assign n4417 = n5074 ^ n5075;
  assign n4589 = n5076 ^ n5077;
  assign n3210 = n5078 ^ n5079;
  assign n4500 = n5080 ^ n5081;
  assign n4221 = n5082 ^ n5083;
  assign n4227 = n5084 ^ n5085;
  assign n4493 = n5086 ^ n5087;
  assign n3769 = n5088 ^ n5089;
  assign n3208 = n5090 ^ n5091;
  assign n4492 = n5092 ^ n5093;
  assign n3300 = n5094 ^ n5095;
  assign n3306 = n5096 ^ n5097;
  assign n3765 = n5098 ^ n5099;
  assign n4466 = n5100 ^ n5101;
  assign n4465 = n5102 ^ n5103;
  assign n2623 = n5104 ^ n5105;
  assign n3308 = n5106 ^ n5107;
  assign n4468 = n5108 ^ n5109;
  assign n3767 = n5110 ^ n5111;
  assign n4467 = n5112 ^ n5113;
  assign n3310 = n5114 ^ n5115;
  assign n3771 = n5116 ^ n5117;
  assign n4495 = n5118 ^ n5119;
  assign n4494 = n5120 ^ n5121;
  assign n3225 = n5122 ^ n5123;
  assign n4506 = n5124 ^ n5125;
  assign n4243 = n5126 ^ n5127;
  assign n4505 = n5128 ^ n5129;
  assign n4497 = n5130 ^ n5131;
  assign n4945 = n5132 ^ n5133;
  assign n4496 = n5134 ^ n5135;
  assign n4241 = n5136 ^ n5137;
  assign n4471 = n5138 ^ n5139;
  assign n4239 = n5140 ^ n5141;
  assign n3227 = n5142 ^ n5143;
  assign n3552 = n5144 ^ n5145;
  assign n3751 = n5146 ^ n5147;
  assign n4499 = n5148 ^ n5149;
  assign n4498 = n5150 ^ n5151;
  assign n4525 = n4941 ^ n5154;
  assign n3233 = n5155 ^ n5156;
  assign n3312 = n5157 ^ n5158;
  assign n4502 = n5159 ^ n5160;
  assign n4501 = n5161 ^ n5162;
  assign n3297 = n5163 ^ n5164;
  assign n3778 = n5165 ^ n5166;
  assign n4265 = n5167 ^ n5168;
  assign n4250 = n5169 ^ n5170;
  assign n3237 = n5171 ^ n5172;
  assign n3556 = n5173 ^ n5174;
  assign n3554 = n5175 ^ n5176;
  assign n4418 = n5177 ^ n5178;
  assign n4514 = n5179 ^ n5180;
  assign n4504 = n5181 ^ n5182;
  assign n3781 = n5183 ^ n5184;
  assign n4513 = n5185 ^ n5186;
  assign n4503 = n5187 ^ n5188;
  assign n4255 = n5189 ^ n5190;
  assign n3314 = n5191 ^ n5192;
  assign n3318 = n5193 ^ n5194;
  assign n2985 = n5195 ^ n5196;
  assign n4261 = n5197 ^ n5198;
  assign n3229 = n5199 ^ n5200;
  assign n4246 = n5201 ^ n5202;
  assign n4507 = n5203 ^ n5204;
  assign n4512 = n5205 ^ n5206;
  assign n3783 = n5207 ^ n5208;
  assign n3837 = n5209 ^ n5210;
  assign n4248 = n5211 ^ n5212;
  assign n3234 = n5213 ^ n5214;
  assign n4511 = n5215 ^ n5216;
  assign n3848 = n5217 ^ n5218;
  assign n4510 = n5219 ^ n5220;
  assign n3316 = n5221 ^ n5222;
  assign n3789 = n5223 ^ n5224;
  assign n4519 = n5225 ^ n5226;
  assign n3839 = n5227 ^ n5228;
  assign n4517 = n5229 ^ n5230;
  assign n4521 = n5231 ^ n5232;
  assign n3791 = n5233 ^ n5234;
  assign n4520 = n5235 ^ n5236;
  assign n4419 = n5237 ^ n5238;
  assign n4509 = n5239 ^ n5240;
  assign n2631 = n5241 ^ n5242;
  assign n3322 = n5243 ^ n5244;
  assign n4257 = n5245 ^ n5246;
  assign n3240 = n5247 ^ n5248;
  assign n3324 = n5249 ^ n5250;
  assign n3294 = n5251 ^ n5252;
  assign n2961 = n5253 ^ n5254;
  assign n4252 = n5255 ^ n5256;
  assign n4259 = n5257 ^ n5258;
  assign n4263 = n5259 ^ n5260;
  assign n3320 = n5261 ^ n5262;
  assign n4522 = n5263 ^ n5264;
  assign n3292 = n5265 ^ n5266;
  assign n3792 = n5267 ^ n5268;
  assign n4233 = n5269 ^ n5270;
  assign n4474 = n5271 ^ n5272;
  assign n3214 = n5273 ^ n5274;
  assign n3747 = n5275 ^ n5276;
  assign n4223 = n5277 ^ n5278;
  assign n4479 = n5279 ^ n5280;
  assign n4478 = n5281 ^ n5282;
  assign n3249 = n5283 ^ n5284;
  assign n4518 = n5285 ^ n5286;
  assign n2711 = n5287 ^ n5288;
  assign n3784 = n5289 ^ n5290;
  assign n3755 = n5291 ^ n5292;
  assign n2806 = n5293 ^ n5294;
  assign n2319 = n5295 ^ n5296;
  assign n4481 = n5297 ^ n5298;
  assign n4476 = n5299 ^ n5300;
  assign n4480 = n5301 ^ n5302;
  assign n3749 = n5303 ^ n5304;
  assign n4475 = n5305 ^ n5306;
  assign n5316 = n5141 & n5140;
  assign n5317 = n5256 & n5255;
  assign n4341 = ~n3296;
  assign n4942 = ~n4427;
  assign n4342 = ~n3904;
  assign n4943 = ~n4516;
  assign n4344 = ~n3243;
  assign n4944 = ~n4523;
  assign n4343 = ~n3326;
  assign n4112 = ~n5154;
  assign n5308 = ~n4981;
  assign n5309 = ~n5141;
  assign n4114 = ~n3918;
  assign n5312 = ~n4985;
  assign n5313 = ~n5256;
  assign n5845 = n6441 & n6442;
  assign n5846 = n6443 & n6444;
  assign n5847 = n6445 & n6446;
  assign n5848 = n6447 & n6448;
  assign n5849 = n6449 & n6450;
  assign n5850 = n6451 & n6452;
  assign n5851 = n6453 & n6454;
  assign n5852 = n6455 & n6456;
  assign n5853 = n6457 & n6458;
  assign n5854 = n6459 & n6460;
  assign n5855 = n6461 & n6462;
  assign n5856 = n6463 & n6464;
  assign n5857 = n6465 & n6466;
  assign n5858 = n6467 & n6468;
  assign n5859 = n6469 & n6470;
  assign n5860 = n6471 & n6472;
  assign n5861 = n6473 & n6474;
  assign n5862 = n6475 & n6476;
  assign n5863 = n6477 & n6478;
  assign n5864 = n6479 & n6480;
  assign n5865 = n6481 & n6482;
  assign n5866 = n6483 & n6484;
  assign n5867 = n6485 & n6486;
  assign n5868 = n6487 & n6488;
  assign n5869 = n6489 & n6490;
  assign n5870 = n6491 & n6492;
  assign n5871 = n6493 & n6494;
  assign n5872 = n6495 & n6496;
  assign n5873 = n6497 & n6498;
  assign n5874 = n6499 & n6500;
  assign n5875 = n6501 & n6502;
  assign n5876 = n6503 & n6504;
  assign n5877 = n6505 & n6506;
  assign n5878 = n6507 & n6508;
  assign n5879 = n6509 & n6510;
  assign n5880 = n6511 & n6512;
  assign n5881 = n6513 & n6514;
  assign n5882 = n6515 & n6516;
  assign n5883 = n6517 & n6518;
  assign n5884 = n6519 & n6520;
  assign n5885 = n6521 & n6522;
  assign n5886 = n6523 & n6524;
  assign n5887 = n6525 & n6526;
  assign n5888 = n6527 & n6528;
  assign n5889 = n6529 & n6530;
  assign n5890 = n6531 & n6532;
  assign n5891 = n6533 & n6534;
  assign n5892 = n6535 & n6536;
  assign n5893 = n6537 & n6538;
  assign n5894 = n6539 & n6540;
  assign n5895 = n6541 & n6542;
  assign n5896 = n6543 & n6544;
  assign n5897 = n6545 & n6546;
  assign n5898 = n6547 & n6548;
  assign n5899 = n6549 & n6550;
  assign n5900 = n6551 & n6552;
  assign n5901 = n6553 & n6554;
  assign n5902 = n6555 & n6556;
  assign n5903 = n6557 & n6558;
  assign n5904 = n6559 & n6560;
  assign n5905 = n6561 & n6562;
  assign n5906 = n6563 & n6564;
  assign n5907 = n6565 & n6566;
  assign n5908 = n6567 & n6568;
  assign n5909 = n6569 & n6570;
  assign n5910 = n6571 & n6572;
  assign n5911 = n6573 & n6574;
  assign n5912 = n6575 & n6576;
  assign n5913 = n6577 & n6578;
  assign n5914 = n6579 & n6580;
  assign n5915 = n6581 & n6582;
  assign n5916 = n6583 & n6584;
  assign n5917 = n6585 & n6586;
  assign n5918 = n6587 & n6588;
  assign n5919 = n6589 & n6590;
  assign n5920 = n6591 & n6592;
  assign n5921 = n6593 & n6594;
  assign n5922 = n6595 & n6596;
  assign n5923 = n6597 & n6598;
  assign n5924 = n6599 & n6600;
  assign n5925 = n6601 & n6602;
  assign n5926 = n6603 & n6604;
  assign n5927 = n6605 & n6606;
  assign n5928 = n6607 & n6608;
  assign n5929 = n6609 & n6610;
  assign n5930 = n6611 & n6612;
  assign n5931 = n6613 & n6614;
  assign n5932 = n6615 & n6616;
  assign n5933 = n6617 & n6618;
  assign n5934 = n6619 & n6620;
  assign n5935 = n6621 & n6622;
  assign n5936 = n6623 & n6624;
  assign n5937 = n6625 & n6626;
  assign n5938 = n6627 & n6628;
  assign n5939 = n6629 & n6630;
  assign n5940 = n6631 & n6632;
  assign n5941 = n6633 & n6634;
  assign n5942 = n6635 & n6636;
  assign n5943 = n6637 & n6638;
  assign n5944 = n6639 & n6640;
  assign n5945 = n6641 & n6642;
  assign n5946 = n6643 & n6644;
  assign n5947 = n6645 & n6646;
  assign n5948 = n6647 & n6648;
  assign n5949 = n6649 & n6650;
  assign n5950 = n6651 & n6652;
  assign n5951 = n6653 & n6654;
  assign n5952 = n6655 & n6656;
  assign n5953 = n6657 & n6658;
  assign n5954 = n6659 & n6660;
  assign n5955 = n6661 & n6662;
  assign n5956 = n6663 & n6664;
  assign n5957 = n6665 & n6666;
  assign n5958 = n6667 & n6668;
  assign n5959 = n6669 & n6670;
  assign n5960 = n6671 & n6672;
  assign n5961 = n6673 & n6674;
  assign n5962 = n6675 & n6676;
  assign n5963 = n6677 & n6678;
  assign n5964 = n6679 & n6680;
  assign n5965 = n6681 & n6682;
  assign n5966 = n6683 & n6684;
  assign n5967 = n6685 & n6686;
  assign n5968 = n6687 & n6688;
  assign n5969 = n6689 & n6690;
  assign n5970 = n6691 & n6692;
  assign n5971 = n6693 & n6694;
  assign n5972 = n6695 & n6696;
  assign n5973 = n6697 & n6698;
  assign n5974 = n6699 & n6700;
  assign n5975 = n4346 & n6701;
  assign n5976 = n4345 & n6702;
  assign n5977 = n4348 & n6703;
  assign n5978 = n3728 & n6704;
  assign n5979 = n4972 & n6705;
  assign n5980 = n6706 & n6707;
  assign n5981 = n4122 & n6708;
  assign n5982 = n6709 & n6710;
  assign n5983 = n4120 & n6711;
  assign n5984 = n6712 & n5082;
  assign n3933 = n6713 & n6093;
  assign n5985 = n6714 & n6198;
  assign n5986 = n6715 & n5018;
  assign n5987 = n6716 & n3888;
  assign n5988 = n6717 & n6089;
  assign n5989 = n6719 & n33;
  assign n5554 = ~n6720;
  assign n5990 = n6721 & n6082;
  assign n5568 = ~n6722;
  assign n5991 = n6723 & n6160;
  assign n5572 = ~n6724;
  assign n5576 = ~n6725;
  assign n5992 = n6726 & n3890;
  assign n5993 = n6727 & n6423;
  assign n5994 = n6728 & n6227;
  assign n5804 = ~n6729;
  assign n4032 = ~n6730;
  assign n5586 = ~n6731;
  assign n5995 = n6732 & n6242;
  assign n5996 = n6733 & n6260;
  assign n5997 = n6734 & n6207;
  assign n5596 = ~n6737;
  assign n5998 = n6738 & n5028;
  assign n5999 = n6739 & n5175;
  assign n6000 = n6740 & n5295;
  assign n5602 = ~n6741;
  assign n6001 = n6742 & n6304;
  assign n3966 = n6743 & n6219;
  assign n6002 = n6744 & n5068;
  assign n6003 = n6745 & n6308;
  assign n5614 = ~n6746;
  assign n6004 = n6747 & n6247;
  assign n6005 = n6748 & n4967;
  assign n5840 = ~n6749;
  assign n5706 = ~n6750;
  assign n6006 = n6751 & n6192;
  assign n5624 = ~n6752;
  assign n6007 = n6753 & n5249;
  assign n5548 = ~n6754;
  assign n6008 = n6755 & n6273;
  assign n6009 = n6756 & n6236;
  assign n5642 = ~n6757;
  assign n5646 = ~n6758;
  assign n6010 = n6759 & n6315;
  assign n5654 = ~n6760;
  assign n6011 = n6761 & n5173;
  assign n5650 = ~n6762;
  assign n5666 = ~n6763;
  assign n5660 = ~n6764;
  assign n5320 = n6766 & n6311;
  assign n5152 = n6767 & n6267;
  assign n6012 = n6768 & n4963;
  assign n6013 = n6769 & n6320;
  assign n6014 = n6770 & n6428;
  assign n6015 = n6771 & n6352;
  assign n5682 = ~n6772;
  assign n5734 = ~n6773;
  assign n6016 = n6774 & n6358;
  assign n5540 = ~n6775;
  assign n6017 = n6776 & n6282;
  assign n5700 = ~n6777;
  assign n5696 = ~n6778;
  assign n5708 = ~n6779;
  assign n5686 = ~n6780;
  assign n6018 = n6781 & n6092;
  assign n6019 = n6782 & n6406;
  assign n5720 = ~n6783;
  assign n6020 = n6784 & n6054;
  assign n6021 = n6785 & n6252;
  assign n3992 = n6786 & n6343;
  assign n6022 = n6787 & n6166;
  assign n6023 = n6788 & n5277;
  assign n5746 = ~n6790;
  assign n5748 = ~n6791;
  assign n5556 = ~n6792;
  assign n5752 = ~n6793;
  assign n6024 = n6794 & n6404;
  assign n6025 = n6795 & n6118;
  assign n5754 = ~n6796;
  assign n6026 = n6797 & n5241;
  assign n6027 = n6799 & n4974;
  assign n5524 = ~n6800;
  assign n6028 = n6801 & n6346;
  assign n5762 = ~n6802;
  assign n6029 = n6803 & n6340;
  assign n6030 = n6804 & n5048;
  assign n6031 = n6805 & n6149;
  assign n6032 = n6806 & n6221;
  assign n6033 = n6807 & n6395;
  assign n5780 = ~n6808;
  assign n6034 = n6809 & n5299;
  assign n5792 = ~n6810;
  assign n5786 = ~n6811;
  assign n6035 = n6812 & n5209;
  assign n6036 = n6813 & n6425;
  assign n5810 = ~n6814;
  assign n5726 = ~n6815;
  assign n6037 = n6817 & n5052;
  assign n5824 = ~n6818;
  assign n5828 = ~n6819;
  assign n5318 = n6820 & n6211;
  assign n6038 = n5841 & n6052;
  assign n6039 = n6821 & n6158;
  assign n6040 = n4126 & n6184;
  assign n6041 = n4347 & n6057;
  assign n6042 = n6821 & n6059;
  assign n6043 = n4972 & n6053;
  assign n6044 = n4124 & n6106;
  assign n6045 = n6706 & n6060;
  assign n6046 = n6709 & n33;
  assign n4443 = ~n6822;
  assign n3484 = ~n6823;
  assign n5838 = ~n6824;
  assign n5522 = ~n6825;
  assign n5670 = ~n6826;
  assign n5542 = ~n6827;
  assign n5526 = ~n6828;
  assign n5816 = ~n6829;
  assign n4453 = ~n6830;
  assign n5534 = ~n6831;
  assign n5538 = ~n6832;
  assign n5558 = ~n6833;
  assign n5546 = ~n6834;
  assign n5550 = ~n6835;
  assign n5346 = ~n6836;
  assign n5692 = ~n6837;
  assign n5562 = ~n6838;
  assign n5560 = ~n6839;
  assign n5698 = ~n6840;
  assign n5566 = ~n6841;
  assign n5722 = ~n6842;
  assign n5774 = ~n6843;
  assign n5570 = ~n6844;
  assign n4439 = ~n6845;
  assign n5574 = ~n6846;
  assign n4026 = ~n6847;
  assign n5578 = ~n6848;
  assign n5580 = ~n6849;
  assign n5582 = ~n6850;
  assign n5584 = ~n6851;
  assign n4036 = ~n6852;
  assign n5588 = ~n6853;
  assign n5590 = ~n6854;
  assign n5592 = ~n6855;
  assign n5594 = ~n6856;
  assign n5598 = ~n6857;
  assign n5600 = ~n6858;
  assign n5606 = ~n6859;
  assign n5604 = ~n6860;
  assign n5608 = ~n6861;
  assign n5552 = ~n6862;
  assign n5612 = ~n6863;
  assign n5528 = ~n6864;
  assign n5616 = ~n6865;
  assign n4447 = ~n6866;
  assign n4102 = ~n6867;
  assign n5618 = ~n6868;
  assign n4044 = ~n6869;
  assign n5620 = ~n6870;
  assign n5622 = ~n6871;
  assign n5626 = ~n6872;
  assign n5628 = ~n6873;
  assign n5630 = ~n6874;
  assign n5636 = ~n6875;
  assign n5634 = ~n6876;
  assign n5638 = ~n6877;
  assign n5640 = ~n6878;
  assign n5307 = ~n6879;
  assign n5648 = ~n6880;
  assign n5652 = ~n6881;
  assign n5632 = ~n6882;
  assign n5658 = ~n6883;
  assign n5662 = ~n6884;
  assign n5532 = ~n6885;
  assign n5738 = ~n6886;
  assign n5842 = ~n6887;
  assign n5674 = ~n6888;
  assign n5678 = ~n6889;
  assign n5676 = ~n6890;
  assign n5680 = ~n6891;
  assign n5672 = ~n6892;
  assign n5684 = ~n6893;
  assign n5808 = ~n6894;
  assign n5688 = ~n6895;
  assign n5690 = ~n6896;
  assign n5832 = ~n6897;
  assign n5694 = ~n6898;
  assign n5724 = ~n6899;
  assign n5702 = ~n6900;
  assign n5704 = ~n6901;
  assign n5710 = ~n6902;
  assign n5712 = ~n6903;
  assign n5714 = ~n6904;
  assign n5716 = ~n6905;
  assign n5564 = ~n6906;
  assign n5311 = ~n6907;
  assign n5830 = ~n6908;
  assign n5834 = ~n6909;
  assign n5728 = ~n6910;
  assign n5730 = ~n6911;
  assign n5732 = ~n6912;
  assign n5644 = ~n6913;
  assign n5736 = ~n6914;
  assign n5742 = ~n6915;
  assign n5740 = ~n6916;
  assign n5744 = ~n6917;
  assign n5750 = ~n6918;
  assign n5784 = ~n6919;
  assign n5756 = ~n6920;
  assign n5758 = ~n6921;
  assign n5760 = ~n6922;
  assign n4457 = ~n6923;
  assign n5770 = ~n6924;
  assign n5772 = ~n6925;
  assign n5768 = ~n6926;
  assign n5782 = ~n6927;
  assign n5776 = ~n6928;
  assign n5788 = ~n6929;
  assign n5794 = ~n6930;
  assign n5790 = ~n6931;
  assign n5796 = ~n6932;
  assign n5798 = ~n6933;
  assign n5544 = ~n6934;
  assign n5530 = ~n6935;
  assign n5800 = ~n6936;
  assign n5802 = ~n6937;
  assign n4455 = ~n6938;
  assign n5806 = ~n6939;
  assign n5664 = ~n6940;
  assign n5812 = ~n6941;
  assign n5814 = ~n6942;
  assign n5668 = ~n6943;
  assign n5718 = ~n6944;
  assign n5818 = ~n6945;
  assign n5822 = ~n6946;
  assign n5826 = ~n6947;
  assign n5778 = ~n6948;
  assign n5656 = ~n6949;
  assign n5836 = ~n6950;
  assign n5764 = ~n6951;
  assign n6718 = n6955 & n6090;
  assign n6735 = n6963 & n6208;
  assign n6736 = n6964 & n6396;
  assign n6765 = n6978 & n6114;
  assign n6789 = n6987 & n6140;
  assign n6798 = n6993 & n6376;
  assign n6816 = n7001 & n6432;
  assign n6952 = ~n7007;
  assign n6047 = n6953 & n7008;
  assign n2617 = n4420 ^ n4421;
  assign n3758 = n4426 ^ n4427;
  assign n2639 = n2319 ^ n2806;
  assign n3764 = n4465 ^ n4466;
  assign n3766 = n4467 ^ n4468;
  assign n3763 = n4469 ^ n4470;
  assign n3803 = n4174 ^ n4471;
  assign n3795 = n4472 ^ n4473;
  assign n3746 = n4223 ^ n4474;
  assign n3797 = n3554 ^ n4418;
  assign n3748 = n4475 ^ n4476;
  assign n3799 = n4477 ^ n3874;
  assign n3750 = n4478 ^ n4479;
  assign n2948 = n4480 ^ n4481;
  assign n3753 = n4482 ^ n4483;
  assign n3754 = n4484 ^ n4485;
  assign n2615 = n4486 ^ n4487;
  assign n2613 = n4488 ^ n4489;
  assign n3756 = n4490 ^ n4491;
  assign n3768 = n4492 ^ n4493;
  assign n3770 = n4494 ^ n4495;
  assign n3772 = n4496 ^ n4497;
  assign n3774 = n4498 ^ n4499;
  assign n3776 = n4221 ^ n4500;
  assign n3779 = n4501 ^ n4502;
  assign n3780 = n4503 ^ n4504;
  assign n3230 = n4505 ^ n4506;
  assign n2625 = n4507 ^ n4508;
  assign n3805 = n4509 ^ n4419;
  assign n2946 = n4510 ^ n4511;
  assign n3782 = n3837 ^ n4512;
  assign n3238 = n4513 ^ n4514;
  assign n3785 = n4515 ^ n4516;
  assign n3786 = n4517 ^ n4518;
  assign n3788 = n3839 ^ n4519;
  assign n3790 = n4520 ^ n4521;
  assign n3793 = n4522 ^ n4523;
  assign n3761 = n4530 ^ n4531;
  assign n3801 = n4589 ^ n4417;
  assign n4572 = n3759 & n4942;
  assign n4592 = n4515 & n4943;
  assign n4594 = n4522 & n4944;
  assign n4598 = n3777 & n4500;
  assign n4600 = n4482 & n4483;
  assign n4601 = n4945 & n4946;
  assign n4602 = n4491 & n3757;
  assign n4603 = n4420 & n4421;
  assign n4604 = n4466 & n3765;
  assign n4605 = n3767 & n4468;
  assign n4606 = n4495 & n3771;
  assign n4608 = n3787 & n4518;
  assign n4609 = n4501 & n4502;
  assign n4610 = n4513 & n4514;
  assign n4611 = n4480 & n4481;
  assign n4612 = n4508 & n4507;
  assign n4613 = n3755 & n4485;
  assign n4614 = n3791 & n4521;
  assign n4615 = n3747 & n4474;
  assign n4616 = n3751 & n4479;
  assign n4597 = ~n3773;
  assign n4599 = ~n4487;
  assign n4413 = ~n3221;
  assign n2977 = ~n2959;
  assign n4574 = ~n3777;
  assign n2979 = ~n2641;
  assign n2981 = ~n2637;
  assign n4269 = ~n4416;
  assign n4527 = ~n4948;
  assign n2905 = ~n2870;
  assign n2697 = ~n2621;
  assign n4552 = ~n4508;
  assign n4557 = ~n3787;
  assign n4562 = ~n4473;
  assign n4566 = ~n4472;
  assign n4289 = ~n4229;
  assign n4537 = ~n4485;
  assign n3635 = ~n3286;
  assign n4565 = ~n4469;
  assign n2971 = ~n2957;
  assign n4293 = ~n4225;
  assign n4377 = ~n3213;
  assign n3519 = ~n4231;
  assign n4267 = ~n3841;
  assign n4310 = ~n3874;
  assign n3394 = ~n4477;
  assign n4563 = ~n4486;
  assign n4532 = ~n4482;
  assign n4197 = ~n4484;
  assign n4271 = ~n3217;
  assign n4195 = ~n3752;
  assign n4591 = ~n4515;
  assign n4533 = ~n4483;
  assign n4564 = ~n4470;
  assign n3637 = ~n3302;
  assign n4316 = ~n3844;
  assign n4539 = ~n3757;
  assign n4538 = ~n4491;
  assign n4199 = ~n4490;
  assign n4568 = ~n4489;
  assign n4567 = ~n4488;
  assign n4384 = ~n4236;
  assign n3521 = ~n3218;
  assign n4541 = ~n4421;
  assign n4540 = ~n4420;
  assign n4570 = ~n4531;
  assign n4569 = ~n4530;
  assign n3813 = ~n3760;
  assign n3563 = ~n3303;
  assign n4571 = ~n3759;
  assign n4201 = ~n4426;
  assign n4273 = ~n4417;
  assign n3524 = ~n4589;
  assign n3517 = ~n3210;
  assign n4573 = ~n4500;
  assign n4275 = ~n4227;
  assign n4576 = ~n4493;
  assign n4575 = ~n3769;
  assign n3816 = ~n4492;
  assign n3641 = ~n3300;
  assign n3639 = ~n3306;
  assign n4543 = ~n3765;
  assign n4542 = ~n4466;
  assign n4203 = ~n4465;
  assign n2973 = ~n2623;
  assign n4545 = ~n4468;
  assign n4544 = ~n3767;
  assign n4205 = ~n4467;
  assign n4547 = ~n3771;
  assign n4546 = ~n4495;
  assign n4207 = ~n4494;
  assign n4392 = ~n3225;
  assign n4579 = ~n4506;
  assign n3527 = ~n4243;
  assign n4577 = ~n4505;
  assign n4578 = ~n4497;
  assign n4528 = ~n4945;
  assign n3821 = ~n4496;
  assign n4277 = ~n4241;
  assign n3494 = ~n4471;
  assign n4279 = ~n3227;
  assign n4560 = ~n3751;
  assign n4580 = ~n4499;
  assign n3823 = ~n4498;
  assign n4397 = ~n3233;
  assign n3643 = ~n3312;
  assign n4549 = ~n4502;
  assign n4548 = ~n4501;
  assign n3407 = ~n3297;
  assign n4209 = ~n3778;
  assign n3542 = ~n4265;
  assign n3531 = ~n4250;
  assign n4283 = ~n3237;
  assign n4281 = ~n4418;
  assign n4551 = ~n4514;
  assign n4583 = ~n4504;
  assign n4582 = ~n3781;
  assign n4550 = ~n4513;
  assign n3826 = ~n4503;
  assign n4400 = ~n4255;
  assign n3645 = ~n3314;
  assign n3647 = ~n3318;
  assign n3168 = ~n2985;
  assign n4285 = ~n4261;
  assign n4287 = ~n3229;
  assign n3534 = ~n4246;
  assign n4553 = ~n4507;
  assign n4585 = ~n4512;
  assign n4584 = ~n3783;
  assign n4291 = ~n4248;
  assign n3536 = ~n3234;
  assign n4587 = ~n4511;
  assign n3865 = ~n3848;
  assign n4586 = ~n4510;
  assign n3650 = ~n3316;
  assign n4590 = ~n3789;
  assign n4588 = ~n4519;
  assign n4215 = ~n4517;
  assign n4555 = ~n4521;
  assign n4554 = ~n3791;
  assign n4211 = ~n4520;
  assign n4295 = ~n4419;
  assign n3538 = ~n4509;
  assign n2804 = ~n2631;
  assign n3652 = ~n3322;
  assign n4297 = ~n4257;
  assign n3540 = ~n3240;
  assign n3654 = ~n3294;
  assign n2975 = ~n2961;
  assign n3656 = ~n4259;
  assign n4299 = ~n4263;
  assign n4593 = ~n4522;
  assign n4217 = ~n3792;
  assign n4409 = ~n4233;
  assign n4559 = ~n4474;
  assign n4558 = ~n3747;
  assign n4561 = ~n4479;
  assign n4219 = ~n4478;
  assign n4301 = ~n3249;
  assign n4556 = ~n4518;
  assign n2802 = ~n2711;
  assign n4213 = ~n3784;
  assign n4536 = ~n3755;
  assign n2701 = ~n2806;
  assign n4535 = ~n4481;
  assign n4596 = ~n4476;
  assign n4534 = ~n4480;
  assign n4595 = ~n3749;
  assign n3833 = ~n4475;
  assign n3775 = n5152 ^ n5153;
  assign n4949 = n5307 & n5308;
  assign n4950 = n5309 & n5310;
  assign n4951 = n5311 & n5312;
  assign n4952 = n5313 & n5314;
  assign n4060 = ~n5316;
  assign n4086 = ~n5317;
  assign n3900 = n5318 ^ n5319;
  assign n3924 = n5320 ^ n5321;
  assign n5322 = n5522 & n5523;
  assign n5323 = n5524 & n5525;
  assign n5324 = n5526 & n5527;
  assign n5325 = n5528 & n5529;
  assign n5328 = n5530 & n5531;
  assign n5329 = n5532 & n5533;
  assign n5330 = n5534 & n5535;
  assign n5332 = n5538 & n5539;
  assign n5333 = n5540 & n5541;
  assign n5334 = n5542 & n5543;
  assign n5337 = n5544 & n5545;
  assign n5340 = n5546 & n5547;
  assign n5341 = n5548 & n5549;
  assign n5344 = n5550 & n5551;
  assign n5349 = n5552 & n5553;
  assign n5350 = n5554 & n5555;
  assign n5351 = n5556 & n5557;
  assign n5352 = n5558 & n5559;
  assign n5353 = n5560 & n5561;
  assign n5354 = n5562 & n5563;
  assign n5355 = n5564 & n5565;
  assign n5356 = n5566 & n5567;
  assign n5357 = n5568 & n5569;
  assign n5360 = n5570 & n5571;
  assign n5363 = n5572 & n5573;
  assign n5364 = n5574 & n5575;
  assign n5365 = n5576 & n5577;
  assign n5368 = n5578 & n5579;
  assign n5369 = n5580 & n5581;
  assign n5370 = n5582 & n5583;
  assign n5371 = n5584 & n5585;
  assign n5372 = n5586 & n5587;
  assign n5373 = n5588 & n5589;
  assign n5374 = n5590 & n5591;
  assign n5375 = n5592 & n5593;
  assign n5376 = n5594 & n5595;
  assign n5377 = n5596 & n5597;
  assign n5378 = n5598 & n5599;
  assign n5379 = n5600 & n5601;
  assign n5380 = n5602 & n5603;
  assign n5381 = n5604 & n5605;
  assign n5382 = n5606 & n5607;
  assign n5383 = n5608 & n5609;
  assign n5387 = n5612 & n5613;
  assign n5388 = n5614 & n5615;
  assign n5389 = n5616 & n5617;
  assign n5390 = n5618 & n5619;
  assign n5393 = n5620 & n5621;
  assign n5394 = n5622 & n5623;
  assign n5395 = n5624 & n5625;
  assign n5396 = n5626 & n5627;
  assign n5397 = n5628 & n5629;
  assign n5398 = n5630 & n5631;
  assign n5399 = n5632 & n5633;
  assign n5400 = n5634 & n5635;
  assign n5401 = n5636 & n5637;
  assign n5402 = n5638 & n5639;
  assign n5403 = n5640 & n5641;
  assign n5404 = n5642 & n5643;
  assign n5405 = n5644 & n5645;
  assign n5406 = n5646 & n5647;
  assign n5407 = n5648 & n5649;
  assign n5408 = n5650 & n5651;
  assign n5409 = n5652 & n5653;
  assign n5410 = n5654 & n5655;
  assign n5411 = n5656 & n5657;
  assign n5412 = n5658 & n5659;
  assign n5413 = n5660 & n5661;
  assign n5414 = n5662 & n5663;
  assign n5415 = n5664 & n5665;
  assign n5416 = n5666 & n5667;
  assign n5417 = n5668 & n5669;
  assign n5418 = n5670 & n5671;
  assign n5419 = n5672 & n5673;
  assign n5420 = n5674 & n5675;
  assign n5421 = n5676 & n5677;
  assign n5422 = n5678 & n5679;
  assign n5423 = n5680 & n5681;
  assign n5424 = n5682 & n5683;
  assign n5425 = n5684 & n5685;
  assign n5426 = n5686 & n5687;
  assign n5427 = n5688 & n5689;
  assign n5430 = n5690 & n5691;
  assign n5431 = n5692 & n5693;
  assign n5432 = n5694 & n5695;
  assign n5433 = n5696 & n5697;
  assign n5434 = n5698 & n5699;
  assign n5435 = n5700 & n5701;
  assign n5436 = n5702 & n5703;
  assign n5437 = n5704 & n5705;
  assign n5438 = n5706 & n5707;
  assign n5439 = n5708 & n5709;
  assign n5440 = n5710 & n5711;
  assign n5441 = n5712 & n5713;
  assign n5442 = n5714 & n5715;
  assign n5443 = n5716 & n5717;
  assign n5444 = n5718 & n5719;
  assign n5445 = n5720 & n5721;
  assign n5446 = n5722 & n5723;
  assign n5447 = n5724 & n5725;
  assign n5448 = n5726 & n5727;
  assign n5449 = n5728 & n5729;
  assign n5450 = n5730 & n5731;
  assign n5451 = n5732 & n5733;
  assign n5452 = n5734 & n5735;
  assign n5453 = n5736 & n5737;
  assign n5454 = n5738 & n5739;
  assign n5455 = n5740 & n5741;
  assign n5456 = n5742 & n5743;
  assign n5459 = n5744 & n5745;
  assign n5462 = n5746 & n5747;
  assign n5463 = n5748 & n5749;
  assign n5464 = n5750 & n5751;
  assign n5465 = n5752 & n5753;
  assign n5468 = n5754 & n5755;
  assign n5469 = n5756 & n5757;
  assign n5470 = n5758 & n5759;
  assign n5471 = n5760 & n5761;
  assign n5472 = n5762 & n5763;
  assign n5473 = n5764 & n5765;
  assign n5475 = n5768 & n5769;
  assign n5476 = n5770 & n5771;
  assign n5477 = n5772 & n5773;
  assign n5478 = n5774 & n5775;
  assign n5481 = n5776 & n5777;
  assign n5482 = n5778 & n5779;
  assign n5483 = n5780 & n5781;
  assign n5484 = n5782 & n5783;
  assign n5485 = n5784 & n5785;
  assign n5486 = n5786 & n5787;
  assign n5487 = n5788 & n5789;
  assign n5488 = n5790 & n5791;
  assign n5489 = n5792 & n5793;
  assign n5490 = n5794 & n5795;
  assign n5491 = n5796 & n5797;
  assign n5492 = n5798 & n5799;
  assign n5493 = n5800 & n5801;
  assign n5494 = n5802 & n5803;
  assign n5495 = n5804 & n5805;
  assign n5496 = n5806 & n5807;
  assign n5497 = n5808 & n5809;
  assign n5500 = n5810 & n5811;
  assign n5501 = n5812 & n5813;
  assign n5502 = n5814 & n5815;
  assign n5503 = n5816 & n5817;
  assign n5504 = n5818 & n5819;
  assign n5506 = n5822 & n5823;
  assign n5507 = n5824 & n5825;
  assign n5508 = n5826 & n5827;
  assign n5509 = n5828 & n5829;
  assign n5510 = n5830 & n5831;
  assign n5511 = n5832 & n5833;
  assign n5512 = n5834 & n5835;
  assign n5513 = n5836 & n5837;
  assign n5514 = n5838 & n5839;
  assign n5515 = n5840 & n5841;
  assign n5516 = n5152 & n5842;
  assign n5517 = n5320 & n5843;
  assign n5519 = n5318 & n5844;
  assign n4423 = ~n5845;
  assign n4620 = ~n5846;
  assign n4626 = ~n5847;
  assign n4874 = ~n5848;
  assign n4628 = ~n5849;
  assign n5326 = ~n5850;
  assign n4630 = ~n5851;
  assign n4656 = ~n5852;
  assign n5335 = ~n5853;
  assign n4836 = ~n5854;
  assign n5342 = ~n5855;
  assign n4648 = ~n5856;
  assign n5347 = ~n5857;
  assign n4646 = ~n5858;
  assign n4634 = ~n5859;
  assign n4660 = ~n5860;
  assign n5361 = ~n5861;
  assign n4688 = ~n5862;
  assign n4654 = ~n5863;
  assign n4662 = ~n5864;
  assign n4666 = ~n5865;
  assign n5358 = ~n5866;
  assign n4668 = ~n5867;
  assign n4638 = ~n5868;
  assign n4674 = ~n5869;
  assign n4676 = ~n5870;
  assign n4678 = ~n5871;
  assign n4680 = ~n5872;
  assign n4690 = ~n5873;
  assign n4692 = ~n5874;
  assign n4696 = ~n5875;
  assign n4698 = ~n5876;
  assign n4700 = ~n5877;
  assign n4820 = ~n5878;
  assign n4702 = ~n5879;
  assign n4890 = ~n5880;
  assign n4704 = ~n5881;
  assign n4706 = ~n5882;
  assign n4712 = ~n5883;
  assign n4642 = ~n5884;
  assign n4714 = ~n5885;
  assign n4716 = ~n5886;
  assign n4720 = ~n5887;
  assign n4722 = ~n5888;
  assign n4724 = ~n5889;
  assign n4726 = ~n5890;
  assign n4730 = ~n5891;
  assign n4916 = ~n5892;
  assign n4732 = ~n5893;
  assign n4734 = ~n5894;
  assign n4736 = ~n5895;
  assign n4740 = ~n5896;
  assign n4742 = ~n5897;
  assign n4748 = ~n5898;
  assign n4640 = ~n5899;
  assign n4750 = ~n5900;
  assign n4756 = ~n5901;
  assign n4822 = ~n5902;
  assign n4758 = ~n5903;
  assign n4760 = ~n5904;
  assign n4766 = ~n5905;
  assign n4768 = ~n5906;
  assign n4772 = ~n5907;
  assign n4774 = ~n5908;
  assign n4776 = ~n5909;
  assign n4778 = ~n5910;
  assign n4784 = ~n5911;
  assign n4786 = ~n5912;
  assign n4788 = ~n5913;
  assign n4792 = ~n5914;
  assign n4796 = ~n5915;
  assign n4800 = ~n5916;
  assign n4860 = ~n5917;
  assign n4902 = ~n5918;
  assign n4804 = ~n5919;
  assign n4908 = ~n5920;
  assign n4806 = ~n5921;
  assign n4808 = ~n5922;
  assign n4810 = ~n5923;
  assign n4886 = ~n5924;
  assign n4814 = ~n5925;
  assign n4425 = ~n5926;
  assign n4824 = ~n5927;
  assign n4826 = ~n5928;
  assign n4828 = ~n5929;
  assign n4830 = ~n5930;
  assign n4876 = ~n5931;
  assign n4838 = ~n5932;
  assign n4840 = ~n5933;
  assign n4848 = ~n5934;
  assign n4922 = ~n5935;
  assign n4852 = ~n5936;
  assign n4854 = ~n5937;
  assign n5466 = ~n5938;
  assign n4858 = ~n5939;
  assign n4864 = ~n5940;
  assign n4868 = ~n5941;
  assign n4844 = ~n5942;
  assign n4920 = ~n5943;
  assign n4872 = ~n5944;
  assign n4880 = ~n5945;
  assign n4878 = ~n5946;
  assign n5479 = ~n5947;
  assign n4882 = ~n5948;
  assign n4888 = ~n5949;
  assign n4894 = ~n5950;
  assign n4900 = ~n5951;
  assign n4918 = ~n5952;
  assign n5384 = ~n5953;
  assign n4904 = ~n5954;
  assign n4906 = ~n5955;
  assign n4910 = ~n5956;
  assign n4914 = ~n5957;
  assign n5457 = ~n5958;
  assign n5391 = ~n5959;
  assign n4938 = ~n5960;
  assign n4926 = ~n5961;
  assign n4930 = ~n5962;
  assign n4932 = ~n5963;
  assign n4934 = ~n5964;
  assign n4936 = ~n5965;
  assign n4896 = ~n5966;
  assign n4940 = ~n5967;
  assign n4816 = ~n5968;
  assign n3674 = ~n5969;
  assign n4708 = ~n5970;
  assign n4644 = ~n5971;
  assign n4451 = ~n5972;
  assign n4850 = ~n5973;
  assign n3707 = ~n5974;
  assign n3423 = ~n5975;
  assign n3435 = ~n5976;
  assign n3445 = ~n5977;
  assign n5428 = ~n5978;
  assign n4790 = ~n5979;
  assign n4812 = ~n5980;
  assign n5460 = ~n5981;
  assign n3478 = ~n5982;
  assign n5498 = ~n5983;
  assign n4686 = ~n5984;
  assign n4337 = ~n3933;
  assign n4622 = ~n5985;
  assign n4632 = ~n5986;
  assign n4449 = ~n5987;
  assign n4618 = ~n5988;
  assign n3671 = ~n5989;
  assign n4664 = ~n5990;
  assign n4670 = ~n5991;
  assign n4445 = ~n5992;
  assign n4684 = ~n5993;
  assign n4682 = ~n5994;
  assign n4694 = ~n5995;
  assign n4754 = ~n5996;
  assign n3438 = ~n5997;
  assign n4672 = ~n5998;
  assign n4710 = ~n5999;
  assign n4924 = ~n6000;
  assign n4658 = ~n6001;
  assign n4338 = ~n3966;
  assign n4866 = ~n6002;
  assign n4764 = ~n6003;
  assign n4718 = ~n6004;
  assign n3443 = ~n6005;
  assign n4728 = ~n6006;
  assign n4738 = ~n6007;
  assign n4744 = ~n6008;
  assign n4746 = ~n6009;
  assign n4752 = ~n6010;
  assign n4762 = ~n6011;
  assign n5518 = ~n5320;
  assign n3453 = ~n6012;
  assign n4770 = ~n6013;
  assign n4782 = ~n6014;
  assign n4780 = ~n6015;
  assign n4794 = ~n6016;
  assign n4798 = ~n6017;
  assign n4636 = ~n6018;
  assign n4846 = ~n6019;
  assign n3462 = ~n6020;
  assign n4832 = ~n6021;
  assign n4339 = ~n3992;
  assign n4834 = ~n6022;
  assign n4842 = ~n6023;
  assign n4856 = ~n6024;
  assign n4862 = ~n6025;
  assign n4870 = ~n6026;
  assign n3472 = ~n6027;
  assign n4898 = ~n6028;
  assign n4818 = ~n6029;
  assign n4624 = ~n6030;
  assign n4884 = ~n6031;
  assign n4652 = ~n6032;
  assign n3476 = ~n6033;
  assign n4892 = ~n6034;
  assign n4802 = ~n6035;
  assign n4912 = ~n6036;
  assign n4928 = ~n6037;
  assign n5520 = ~n5318;
  assign n4066 = ~n6038;
  assign n4650 = ~n6039;
  assign n5366 = ~n6040;
  assign n3432 = ~n6041;
  assign n4046 = ~n6042;
  assign n4082 = ~n6043;
  assign n5338 = ~n6044;
  assign n4094 = ~n6045;
  assign n4052 = ~n6046;
  assign n12376 = n6047 ^ n6048;
  assign n5521 = ~n6718;
  assign n4038 = ~n6735;
  assign n4100 = ~n6736;
  assign n5536 = ~n6765;
  assign n5610 = ~n6789;
  assign n5766 = ~n6798;
  assign n5820 = ~n6816;
  assign n4357 = n6952 & n6953;
  assign n2029 = n3746 ^ n3747;
  assign n2850 = n3748 ^ n3749;
  assign n2996 = n3750 ^ n3751;
  assign n1952 = n3752 ^ n3753;
  assign n2999 = n3754 ^ n3755;
  assign n2168 = n3756 ^ n3757;
  assign n1672 = n3758 ^ n3759;
  assign n1716 = n3760 ^ n3761;
  assign n2821 = n3762 ^ n3763;
  assign n1923 = n3764 ^ n3765;
  assign n1842 = n3766 ^ n3767;
  assign n2362 = n3768 ^ n3769;
  assign n2741 = n3770 ^ n3771;
  assign n2138 = n3772 ^ n3773;
  assign n2852 = n3774 ^ n3775;
  assign n1425 = n3776 ^ n3777;
  assign n2176 = n3778 ^ n3779;
  assign n2180 = n3780 ^ n3781;
  assign n2824 = n3782 ^ n3783;
  assign n2857 = n3784 ^ n3785;
  assign n1966 = n3786 ^ n3787;
  assign n2438 = n3788 ^ n3789;
  assign n3003 = n3790 ^ n3791;
  assign n1754 = n3792 ^ n3793;
  assign n2942 = n2705 ^ n3168;
  assign n4360 = n4528 & n4529;
  assign n4361 = n4532 & n4533;
  assign n4362 = n4534 & n4535;
  assign n4363 = n4536 & n4537;
  assign n4364 = n4538 & n4539;
  assign n4365 = n4540 & n4541;
  assign n4366 = n4542 & n4543;
  assign n4367 = n4544 & n4545;
  assign n4368 = n4546 & n4547;
  assign n4369 = n4548 & n4549;
  assign n4370 = n4550 & n4551;
  assign n4371 = n4552 & n4553;
  assign n4372 = n4554 & n4555;
  assign n4373 = n4556 & n4557;
  assign n4374 = n4558 & n4559;
  assign n4375 = n4560 & n4561;
  assign n4376 = n4472 & n4562;
  assign n4378 = n4563 & n4487;
  assign n4379 = n4469 & n4564;
  assign n4380 = n4565 & n4470;
  assign n4381 = n4566 & n4473;
  assign n4382 = n4567 & n4489;
  assign n4383 = n4488 & n4568;
  assign n4385 = n4569 & n4531;
  assign n4386 = n4530 & n4570;
  assign n4387 = n4571 & n4427;
  assign n4200 = ~n4572;
  assign n4388 = n4573 & n4574;
  assign n4389 = n4575 & n4493;
  assign n4390 = n3769 & n4576;
  assign n4391 = n4577 & n4506;
  assign n4393 = n4578 & n3773;
  assign n4394 = n4505 & n4579;
  assign n4395 = n3775 & n4580;
  assign n4398 = n4582 & n4504;
  assign n4399 = n3781 & n4583;
  assign n4401 = n4584 & n4512;
  assign n4402 = n3783 & n4585;
  assign n4403 = n4586 & n4511;
  assign n4404 = n4510 & n4587;
  assign n4405 = n4588 & n3789;
  assign n4406 = n4519 & n4590;
  assign n4407 = n4591 & n4516;
  assign n4212 = ~n4592;
  assign n4408 = n4593 & n4523;
  assign n4216 = ~n4594;
  assign n4410 = n4595 & n4476;
  assign n4411 = n3749 & n4596;
  assign n4412 = n4497 & n4597;
  assign n4220 = ~n4598;
  assign n4414 = n4599 & n4486;
  assign n4194 = ~n4600;
  assign n3173 = ~n4601;
  assign n4198 = ~n4602;
  assign n2669 = ~n4603;
  assign n4202 = ~n4604;
  assign n4204 = ~n4605;
  assign n4206 = ~n4606;
  assign n4214 = ~n4608;
  assign n4208 = ~n4609;
  assign n3557 = ~n4610;
  assign n2969 = ~n4611;
  assign n2685 = ~n4612;
  assign n4196 = ~n4613;
  assign n4210 = ~n4614;
  assign n4222 = ~n4615;
  assign n4218 = ~n4616;
  assign n4581 = ~n3775;
  assign n4422 = ~n4949;
  assign n3449 = ~n4950;
  assign n4424 = ~n4951;
  assign n3468 = ~n4952;
  assign n4815 = ~n5322;
  assign n4635 = ~n5323;
  assign n4619 = ~n5324;
  assign n4625 = ~n5325;
  assign n4524 = n5326 & n5327;
  assign n4919 = ~n5328;
  assign n4627 = ~n5329;
  assign n4629 = ~n5330;
  assign n4633 = ~n5332;
  assign n4649 = ~n5333;
  assign n4637 = ~n5334;
  assign n4430 = n5335 & n5336;
  assign n4639 = ~n5337;
  assign n4953 = n5338 & n5339;
  assign n4643 = ~n5340;
  assign n4621 = ~n5341;
  assign n4947 = n5342 & n5343;
  assign n4645 = ~n5344;
  assign n4432 = n5347 & n5348;
  assign n4885 = ~n5349;
  assign n4651 = ~n5350;
  assign n4685 = ~n5351;
  assign n4641 = ~n5352;
  assign n4687 = ~n5353;
  assign n4653 = ~n5354;
  assign n4661 = ~n5355;
  assign n4659 = ~n5356;
  assign n4865 = ~n5357;
  assign n4434 = n5358 & n5359;
  assign n4665 = ~n5360;
  assign n4428 = n5361 & n5362;
  assign n4657 = ~n5363;
  assign n4667 = ~n5364;
  assign n4669 = ~n5365;
  assign n4955 = n5366 & n5367;
  assign n4675 = ~n5368;
  assign n4673 = ~n5369;
  assign n4677 = ~n5370;
  assign n4679 = ~n5371;
  assign n4681 = ~n5372;
  assign n4695 = ~n5373;
  assign n4691 = ~n5374;
  assign n4697 = ~n5375;
  assign n4699 = ~n5376;
  assign n4693 = ~n5377;
  assign n4701 = ~n5378;
  assign n4689 = ~n5379;
  assign n4683 = ~n5380;
  assign n4703 = ~n5381;
  assign n4707 = ~n5382;
  assign n4705 = ~n5383;
  assign n4004 = n5384 & n5385;
  assign n4711 = ~n5387;
  assign n4709 = ~n5388;
  assign n4713 = ~n5389;
  assign n4715 = ~n5390;
  assign n4436 = n5391 & n5392;
  assign n4719 = ~n5393;
  assign n4721 = ~n5394;
  assign n4727 = ~n5395;
  assign n4729 = ~n5396;
  assign n4725 = ~n5397;
  assign n4731 = ~n5398;
  assign n4733 = ~n5399;
  assign n4723 = ~n5400;
  assign n4739 = ~n5401;
  assign n4741 = ~n5402;
  assign n4735 = ~n5403;
  assign n4743 = ~n5404;
  assign n4939 = ~n5405;
  assign n4745 = ~n5406;
  assign n4749 = ~n5407;
  assign n4737 = ~n5408;
  assign n4747 = ~n5409;
  assign n4753 = ~n5410;
  assign n4755 = ~n5411;
  assign n4757 = ~n5412;
  assign n4751 = ~n5413;
  assign n4759 = ~n5414;
  assign n4909 = ~n5415;
  assign n4761 = ~n5416;
  assign n4917 = ~n5417;
  assign n4655 = ~n5418;
  assign n4767 = ~n5419;
  assign n4771 = ~n5420;
  assign n4773 = ~n5421;
  assign n4775 = ~n5422;
  assign n4777 = ~n5423;
  assign n4763 = ~n5424;
  assign n4783 = ~n5425;
  assign n4781 = ~n5426;
  assign n4785 = ~n5427;
  assign n4956 = n5428 & n5429;
  assign n4787 = ~n5430;
  assign n4791 = ~n5431;
  assign n4795 = ~n5432;
  assign n4793 = ~n5433;
  assign n4647 = ~n5434;
  assign n4797 = ~n5435;
  assign n4799 = ~n5436;
  assign n4789 = ~n5437;
  assign n4769 = ~n5438;
  assign n4801 = ~n5439;
  assign n4803 = ~n5440;
  assign n4805 = ~n5441;
  assign n4807 = ~n5442;
  assign n4809 = ~n5443;
  assign n4813 = ~n5444;
  assign n4817 = ~n5445;
  assign n4819 = ~n5446;
  assign n4823 = ~n5447;
  assign n4671 = ~n5448;
  assign n4829 = ~n5449;
  assign n4827 = ~n5450;
  assign n4825 = ~n5451;
  assign n4779 = ~n5452;
  assign n4837 = ~n5453;
  assign n4913 = ~n5454;
  assign n4835 = ~n5455;
  assign n4839 = ~n5456;
  assign n3169 = n5457 & n5458;
  assign n4843 = ~n5459;
  assign n4957 = n5460 & n5461;
  assign n4841 = ~n5462;
  assign n4831 = ~n5463;
  assign n4847 = ~n5464;
  assign n4845 = ~n5465;
  assign n3989 = n5466 & n5467;
  assign n4855 = ~n5468;
  assign n4857 = ~n5469;
  assign n4859 = ~n5470;
  assign n4863 = ~n5471;
  assign n4861 = ~n5472;
  assign n4867 = ~n5473;
  assign n4875 = ~n5475;
  assign n4871 = ~n5476;
  assign n4879 = ~n5477;
  assign n4877 = ~n5478;
  assign n4958 = n5479 & n5480;
  assign n4873 = ~n5481;
  assign n4881 = ~n5482;
  assign n4883 = ~n5483;
  assign n4853 = ~n5484;
  assign n4851 = ~n5485;
  assign n4833 = ~n5486;
  assign n4887 = ~n5487;
  assign n4889 = ~n5488;
  assign n4891 = ~n5489;
  assign n4893 = ~n5490;
  assign n4849 = ~n5491;
  assign n4895 = ~n5492;
  assign n4899 = ~n5493;
  assign n4905 = ~n5494;
  assign n4897 = ~n5495;
  assign n4903 = ~n5496;
  assign n4907 = ~n5497;
  assign n4959 = n5498 & n5499;
  assign n4911 = ~n5500;
  assign n4915 = ~n5501;
  assign n4937 = ~n5502;
  assign n4921 = ~n5503;
  assign n4901 = ~n5504;
  assign n4925 = ~n5506;
  assign n4927 = ~n5507;
  assign n4929 = ~n5508;
  assign n4663 = ~n5509;
  assign n4811 = ~n5510;
  assign n4933 = ~n5511;
  assign n4821 = ~n5512;
  assign n4935 = ~n5513;
  assign n4931 = ~n5514;
  assign n4717 = ~n5515;
  assign n4960 = n4451 & n5346;
  assign n4765 = ~n5516;
  assign n3459 = ~n5517;
  assign n4961 = n5518 & n5321;
  assign n3490 = ~n5519;
  assign n4962 = n5520 & n5319;
  assign n5315 = n5521 & n4977;
  assign n5331 = n5536 & n5537;
  assign n5386 = n5610 & n5611;
  assign n5474 = n5766 & n5767;
  assign n5505 = n5820 & n5821;
  assign n5345 = ~n4357;
  assign n3004 = ~n2850;
  assign n2836 = ~n2996;
  assign n1758 = ~n1952;
  assign n2838 = ~n2999;
  assign n2828 = ~n2168;
  assign n1750 = ~n1672;
  assign n1889 = ~n1716;
  assign n2830 = ~n2821;
  assign n1760 = ~n1923;
  assign n1972 = ~n1842;
  assign n2513 = ~n2362;
  assign n2840 = ~n2741;
  assign n2844 = ~n2138;
  assign n3005 = ~n2852;
  assign n2288 = ~n2176;
  assign n3006 = ~n2180;
  assign n2009 = ~n2824;
  assign n3007 = ~n2857;
  assign n1618 = ~n1966;
  assign n2509 = ~n2438;
  assign n2834 = ~n3003;
  assign n1950 = ~n1754;
  assign n3809 = n4194 & n4195;
  assign n3810 = n4196 & n4197;
  assign n3811 = n4198 & n4199;
  assign n3814 = n4200 & n4201;
  assign n3817 = n4202 & n4203;
  assign n3818 = n4204 & n4205;
  assign n3819 = n4206 & n4207;
  assign n3824 = n4208 & n4209;
  assign n3827 = n4210 & n4211;
  assign n3828 = n4212 & n4213;
  assign n3829 = n4214 & n4215;
  assign n3830 = n4216 & n4217;
  assign n3831 = n4218 & n4219;
  assign n3835 = n4220 & n4221;
  assign n3840 = n4222 & n4223;
  assign n3808 = ~n4360;
  assign n3251 = ~n4361;
  assign n2421 = ~n4362;
  assign n3253 = ~n4363;
  assign n3255 = ~n4364;
  assign n2099 = ~n4365;
  assign n3261 = ~n4366;
  assign n3263 = ~n4367;
  assign n3265 = ~n4368;
  assign n3267 = ~n4369;
  assign n3043 = ~n4370;
  assign n2115 = ~n4371;
  assign n3269 = ~n4372;
  assign n3273 = ~n4373;
  assign n3277 = ~n4374;
  assign n3279 = ~n4375;
  assign n3807 = ~n4376;
  assign n2095 = ~n4378;
  assign n3834 = ~n4379;
  assign n3175 = ~n4380;
  assign n3171 = ~n4381;
  assign n2097 = ~n4382;
  assign n2667 = ~n4383;
  assign n3177 = ~n4385;
  assign n3812 = ~n4386;
  assign n3257 = ~n4387;
  assign n3259 = ~n4388;
  assign n3179 = ~n4389;
  assign n3815 = ~n4390;
  assign n2952 = ~n4391;
  assign n3181 = ~n4393;
  assign n3405 = ~n4394;
  assign n3183 = ~n4395;
  assign n3185 = ~n4398;
  assign n3825 = ~n4399;
  assign n3187 = ~n4401;
  assign n3836 = ~n4402;
  assign n2414 = ~n4403;
  assign n2967 = ~n4404;
  assign n3189 = ~n4405;
  assign n3838 = ~n4406;
  assign n3271 = ~n4407;
  assign n3275 = ~n4408;
  assign n3191 = ~n4410;
  assign n3832 = ~n4411;
  assign n3820 = ~n4412;
  assign n2661 = ~n4414;
  assign n3794 = n4422 & n4423;
  assign n2656 = n4424 & n4425;
  assign n2725 = n4428 ^ n4429;
  assign n3842 = n4430 ^ n4431;
  assign n2875 = n4432 ^ n4433;
  assign n3846 = n4434 ^ n4435;
  assign n3850 = n4436 ^ n4437;
  assign n3207 = n4524 ^ n4525;
  assign n4396 = n4581 & n4499;
  assign n3985 = n4619 & n4620;
  assign n3958 = n4621 & n4622;
  assign n3934 = n4625 & n4626;
  assign n4230 = n4627 & n4628;
  assign n3942 = n4629 & n4630;
  assign n3941 = n4633 & n4634;
  assign n3986 = n4635 & n4636;
  assign n3903 = n4637 & n4638;
  assign n3944 = n4639 & n4640;
  assign n3943 = n4641 & n4642;
  assign n4415 = n4643 & n4644;
  assign n3333 = n4645 & n4646;
  assign n3957 = n4647 & n4648;
  assign n2888 = n4649 & n4650;
  assign n3962 = n4651 & n4652;
  assign n3365 = n4653 & n4654;
  assign n3347 = n4655 & n4656;
  assign n4237 = n4657 & n4658;
  assign n3961 = n4659 & n4660;
  assign n4234 = n4661 & n4662;
  assign n3905 = n4663 & n4664;
  assign n3945 = n4665 & n4666;
  assign n3845 = n4667 & n4668;
  assign n3335 = n4669 & n4670;
  assign n3927 = n4671 & n4672;
  assign n4235 = n4673 & n4674;
  assign n3950 = n4675 & n4676;
  assign n3949 = n4677 & n4678;
  assign n3337 = n4679 & n4680;
  assign n3349 = n4681 & n4682;
  assign n3919 = n4683 & n4684;
  assign n3889 = n4685 & n4686;
  assign n3937 = n4687 & n4688;
  assign n3913 = n4689 & n4690;
  assign n3907 = n4691 & n4692;
  assign n3964 = n4693 & n4694;
  assign n3345 = n4695 & n4696;
  assign n3960 = n4697 & n4698;
  assign n3959 = n4699 & n4700;
  assign n3909 = n4701 & n4702;
  assign n3963 = n4703 & n4704;
  assign n3891 = n4705 & n4706;
  assign n3800 = n4707 & n4708;
  assign n4226 = n4709 & n4710;
  assign n3341 = n4711 & n4712;
  assign n3965 = n4713 & n4714;
  assign n3351 = n4715 & n4716;
  assign n2647 = n4717 & n4718;
  assign n3972 = n4719 & n4720;
  assign n3343 = n4721 & n4722;
  assign n3911 = n4723 & n4724;
  assign n3971 = n4725 & n4726;
  assign n3954 = n4727 & n4728;
  assign n3953 = n4729 & n4730;
  assign n3955 = n4731 & n4732;
  assign n3956 = n4733 & n4734;
  assign n3353 = n4735 & n4736;
  assign n3921 = n4737 & n4738;
  assign n3968 = n4739 & n4740;
  assign n3967 = n4741 & n4742;
  assign n3976 = n4743 & n4744;
  assign n3970 = n4745 & n4746;
  assign n3975 = n4747 & n4748;
  assign n3969 = n4749 & n4750;
  assign n3327 = n4751 & n4752;
  assign n4238 = n4753 & n4754;
  assign n3355 = n4755 & n4756;
  assign n3974 = n4757 & n4758;
  assign n3973 = n4759 & n4760;
  assign n4242 = n4761 & n4762;
  assign n4335 = n4763 & n4764;
  assign n4240 = n4765 & n4766;
  assign n3367 = n4767 & n4768;
  assign n4254 = n4769 & n4770;
  assign n3978 = n4771 & n4772;
  assign n3915 = n4773 & n4774;
  assign n3977 = n4775 & n4776;
  assign n3357 = n4777 & n4778;
  assign n3893 = n4779 & n4780;
  assign n3982 = n4781 & n4782;
  assign n4244 = n4783 & n4784;
  assign n3981 = n4785 & n4786;
  assign n3361 = n4787 & n4788;
  assign n3796 = n4789 & n4790;
  assign n3917 = n4791 & n4792;
  assign n4249 = n4793 & n4794;
  assign n3359 = n4795 & n4796;
  assign n3980 = n4797 & n4798;
  assign n3979 = n4799 & n4800;
  assign n4253 = n4801 & n4802;
  assign n3923 = n4803 & n4804;
  assign n3984 = n4805 & n4806;
  assign n3983 = n4807 & n4808;
  assign n3993 = n4809 & n4810;
  assign n4260 = n4811 & n4812;
  assign n3994 = n4813 & n4814;
  assign n4228 = n4815 & n4816;
  assign n3363 = n4817 & n4818;
  assign n3988 = n4819 & n4820;
  assign n3895 = n4821 & n4822;
  assign n3987 = n4823 & n4824;
  assign n4002 = n4825 & n4826;
  assign n3371 = n4827 & n4828;
  assign n4245 = n4829 & n4830;
  assign n3901 = n4831 & n4832;
  assign n4336 = n4833 & n4834;
  assign n4001 = n4835 & n4836;
  assign n3991 = n4837 & n4838;
  assign n3369 = n4839 & n4840;
  assign n3377 = n4841 & n4842;
  assign n4247 = n4843 & n4844;
  assign n3948 = n4845 & n4846;
  assign n4251 = n4847 & n4848;
  assign n4262 = n4849 & n4850;
  assign n3375 = n4851 & n4852;
  assign n3897 = n4853 & n4854;
  assign n3947 = n4855 & n4856;
  assign n3990 = n4857 & n4858;
  assign n3996 = n4859 & n4860;
  assign n3940 = n4861 & n4862;
  assign n3995 = n4863 & n4864;
  assign n3946 = n4865 & n4866;
  assign n3373 = n4867 & n4868;
  assign n3999 = n4871 & n4872;
  assign n3939 = n4873 & n4874;
  assign n3929 = n4875 & n4876;
  assign n4000 = n4877 & n4878;
  assign n3564 = n4879 & n4880;
  assign n4256 = n4881 & n4882;
  assign n4008 = n4883 & n4884;
  assign n3938 = n4885 & n4886;
  assign n3925 = n4887 & n4888;
  assign n3383 = n4889 & n4890;
  assign n3931 = n4891 & n4892;
  assign n4258 = n4893 & n4894;
  assign n4010 = n4895 & n4896;
  assign n4007 = n4897 & n4898;
  assign n3385 = n4899 & n4900;
  assign n3936 = n4901 & n4902;
  assign n4009 = n4903 & n4904;
  assign n4003 = n4905 & n4906;
  assign n3379 = n4907 & n4908;
  assign n4232 = n4909 & n4910;
  assign n3998 = n4911 & n4912;
  assign n4005 = n4913 & n4914;
  assign n3381 = n4915 & n4916;
  assign n3997 = n4917 & n4918;
  assign n3952 = n4919 & n4920;
  assign n3951 = n4921 & n4922;
  assign n3935 = n4925 & n4926;
  assign n3887 = n4927 & n4928;
  assign n3387 = n4929 & n4930;
  assign n3339 = n4931 & n4932;
  assign n3329 = n4933 & n4934;
  assign n3331 = n4935 & n4936;
  assign n4264 = n4937 & n4938;
  assign n3899 = n4939 & n4940;
  assign n4462 = n4524 & n4941;
  assign n4463 = n4430 & n4431;
  assign n4464 = n4434 & n4435;
  assign n4607 = n4947 & n4948;
  assign n4440 = ~n4524;
  assign n4458 = ~n4430;
  assign n4448 = ~n4953;
  assign n4526 = ~n4947;
  assign n4442 = ~n4432;
  assign n4460 = ~n4434;
  assign n4438 = ~n4428;
  assign n4444 = ~n4955;
  assign n4106 = ~n4004;
  assign n4456 = ~n4436;
  assign n4446 = ~n4956;
  assign n2965 = ~n3169;
  assign n4452 = ~n4957;
  assign n4092 = ~n3989;
  assign n3617 = ~n4958;
  assign n4454 = ~n4959;
  assign n4358 = ~n4960;
  assign n4072 = ~n4961;
  assign n4110 = ~n4962;
  assign n4617 = ~n5315;
  assign n4631 = ~n5331;
  assign n4954 = n5345 & n5346;
  assign n4623 = ~n5386;
  assign n4869 = ~n5474;
  assign n4923 = ~n5505;
  assign n2232 = n3794 ^ n3795;
  assign n2162 = n3796 ^ n3797;
  assign n2170 = n3800 ^ n3801;
  assign n3250 = ~n3809;
  assign n3252 = ~n3810;
  assign n3254 = ~n3811;
  assign n3522 = n3812 & n3813;
  assign n3256 = ~n3814;
  assign n3525 = n3815 & n3816;
  assign n3260 = ~n3817;
  assign n3262 = ~n3818;
  assign n3264 = ~n3819;
  assign n3528 = n3820 & n3821;
  assign n3266 = ~n3824;
  assign n3532 = n3825 & n3826;
  assign n3268 = ~n3827;
  assign n3270 = ~n3828;
  assign n3272 = ~n3829;
  assign n3274 = ~n3830;
  assign n3278 = ~n3831;
  assign n3543 = n3832 & n3833;
  assign n3204 = n3808 & n3173;
  assign n3545 = n3834 & n3762;
  assign n3258 = ~n3835;
  assign n3559 = n3836 & n3837;
  assign n3560 = n3838 & n3839;
  assign n3276 = ~n3840;
  assign n3283 = n3841 ^ n3842;
  assign n2442 = n3845 ^ n3846;
  assign n3332 = n3887 ^ n3888;
  assign n3340 = n3889 ^ n3890;
  assign n3342 = n3891 ^ n3892;
  assign n3368 = n3893 ^ n3894;
  assign n3372 = n3895 ^ n3896;
  assign n3323 = n3897 ^ n3898;
  assign n2605 = n3899 ^ n3900;
  assign n2316 = n3901 ^ n3902;
  assign n3290 = n3903 ^ n3904;
  assign n3388 = n3905 ^ n3906;
  assign n3304 = n3907 ^ n3908;
  assign n2619 = n3909 ^ n3910;
  assign n3231 = n3911 ^ n3912;
  assign n2607 = n3913 ^ n3914;
  assign n3239 = n3915 ^ n3916;
  assign n3360 = n3917 ^ n3918;
  assign n3298 = n3919 ^ n3920;
  assign n3245 = n3921 ^ n3922;
  assign n2246 = n3923 ^ n3924;
  assign n3247 = n3925 ^ n3926;
  assign n2526 = n3927 ^ n3928;
  assign n2611 = n3929 ^ n3930;
  assign n2609 = n3931 ^ n3932;
  assign n3287 = n3933 ^ n3934;
  assign n3330 = n3935 ^ n3936;
  assign n3366 = n3937 ^ n3938;
  assign n3293 = n3939 ^ n3940;
  assign n3295 = n3941 ^ n3942;
  assign n3334 = n3943 ^ n3944;
  assign n3336 = n3945 ^ n3946;
  assign n3376 = n3947 ^ n3948;
  assign n3338 = n3949 ^ n3950;
  assign n3325 = n3951 ^ n3952;
  assign n3344 = n3953 ^ n3954;
  assign n3299 = n3955 ^ n3956;
  assign n3301 = n3957 ^ n3958;
  assign n3346 = n3959 ^ n3960;
  assign n3348 = n3961 ^ n3962;
  assign n3350 = n3963 ^ n3964;
  assign n3352 = n3965 ^ n3966;
  assign n3305 = n3967 ^ n3968;
  assign n3307 = n3969 ^ n3970;
  assign n3354 = n3971 ^ n3972;
  assign n3356 = n3973 ^ n3974;
  assign n3309 = n3975 ^ n3976;
  assign n3358 = n3977 ^ n3978;
  assign n3311 = n3979 ^ n3980;
  assign n3362 = n3981 ^ n3982;
  assign n3313 = n3983 ^ n3984;
  assign n3285 = n3985 ^ n3986;
  assign n3364 = n3987 ^ n3988;
  assign n3315 = n3989 ^ n3990;
  assign n3370 = n3991 ^ n3992;
  assign n3317 = n3993 ^ n3994;
  assign n3374 = n3995 ^ n3996;
  assign n3319 = n3997 ^ n3998;
  assign n3321 = n3999 ^ n4000;
  assign n3378 = n4001 ^ n4002;
  assign n3380 = n4003 ^ n4004;
  assign n3382 = n4005 ^ n4006;
  assign n3384 = n4007 ^ n4008;
  assign n3386 = n4009 ^ n4010;
  assign n3209 = n4226 ^ n4227;
  assign n3211 = n4228 ^ n4229;
  assign n3212 = n4230 ^ n4231;
  assign n3215 = n4232 ^ n4233;
  assign n3216 = n4234 ^ n3547;
  assign n3219 = n4235 ^ n4236;
  assign n3220 = n4237 ^ n3549;
  assign n3223 = n4238 ^ n4239;
  assign n3222 = n4240 ^ n4241;
  assign n3224 = n4242 ^ n4243;
  assign n3226 = n4244 ^ n3552;
  assign n3228 = n4245 ^ n4246;
  assign n3235 = n4247 ^ n4248;
  assign n3232 = n4249 ^ n4250;
  assign n2629 = n4251 ^ n4252;
  assign n3236 = n4253 ^ n3556;
  assign n3244 = n4254 ^ n4255;
  assign n3241 = n4256 ^ n4257;
  assign n3242 = n4258 ^ n4259;
  assign n2633 = n4260 ^ n4261;
  assign n3246 = n4262 ^ n4263;
  assign n3248 = n4264 ^ n4265;
  assign n3328 = n4335 ^ n4136;
  assign n3291 = n4336 ^ n4139;
  assign n3806 = ~n3794;
  assign n2679 = ~n2656;
  assign n4128 = n3934 & n4337;
  assign n4134 = n3965 & n4338;
  assign n4141 = n3991 & n4339;
  assign n4144 = n4005 & n4340;
  assign n4145 = n3942 & n4341;
  assign n4146 = n3903 & n4342;
  assign n4147 = n3952 & n4343;
  assign n4148 = n4258 & n4344;
  assign n4149 = n3891 & n4345;
  assign n4150 = n4336 & n4346;
  assign n4151 = n3327 & n4347;
  assign n4152 = n3367 & n4348;
  assign n4153 = n3985 & n3986;
  assign n4154 = n3339 & n3890;
  assign n4155 = n3997 & n3998;
  assign n4156 = n3943 & n3944;
  assign n4157 = n3365 & n3938;
  assign n4158 = n3347 & n3962;
  assign n4159 = n3957 & n3958;
  assign n4160 = n3945 & n3946;
  assign n4161 = n3949 & n3950;
  assign n4162 = n3960 & n3345;
  assign n4163 = n3964 & n3349;
  assign n4164 = n3383 & n4008;
  assign n4165 = n3967 & n3968;
  assign n4166 = n3971 & n3972;
  assign n4167 = n3953 & n3954;
  assign n4168 = n3887 & n3888;
  assign n4169 = n3956 & n3955;
  assign n4170 = n3385 & n4010;
  assign n4171 = n3969 & n3970;
  assign n4172 = n3975 & n3976;
  assign n4173 = n3974 & n3355;
  assign n4175 = n3977 & n3978;
  assign n4176 = n3981 & n3982;
  assign n4177 = n3917 & n3918;
  assign n4178 = n3979 & n3980;
  assign n4179 = n3983 & n3984;
  assign n4180 = n3994 & n3993;
  assign n4181 = n3988 & n3363;
  assign n4182 = n3895 & n3896;
  assign n4183 = n4001 & n4002;
  assign n4184 = n3375 & n3948;
  assign n4185 = n3995 & n3996;
  assign n4186 = n3564 & n4349;
  assign n4187 = n3897 & n3898;
  assign n4188 = n4000 & n3999;
  assign n4189 = n3939 & n3940;
  assign n4190 = n4003 & n4004;
  assign n4191 = n3990 & n3989;
  assign n4192 = n3387 & n3906;
  assign n4193 = n3935 & n3936;
  assign n2426 = ~n2725;
  assign n3015 = ~n2875;
  assign n3565 = n3617 ^ n4116;
  assign n3872 = ~n3850;
  assign n12377 = n4357 ^ n4358;
  assign n3513 = ~n3207;
  assign n2944 = n2965 ^ n2703;
  assign n4309 = n4230 & n4377;
  assign n4311 = n4235 & n4384;
  assign n4312 = n4242 & n4392;
  assign n3822 = ~n4396;
  assign n4313 = n4249 & n4397;
  assign n4314 = n4254 & n4400;
  assign n4315 = n4232 & n4409;
  assign n4317 = n4237 & n4413;
  assign n4318 = n4228 & n4229;
  assign n4320 = n4415 & n4416;
  assign n4321 = n4234 & n3217;
  assign n4322 = n3800 & n4417;
  assign n4323 = n4226 & n4227;
  assign n4324 = n4240 & n4241;
  assign n4325 = n4244 & n3227;
  assign n4326 = n4253 & n3237;
  assign n4327 = n3796 & n4418;
  assign n4328 = n4260 & n4261;
  assign n4329 = n4245 & n3229;
  assign n4330 = n4247 & n4248;
  assign n4332 = n4256 & n4257;
  assign n4333 = n4262 & n4263;
  assign n4334 = n4264 & n3249;
  assign n4350 = n4438 & n4439;
  assign n4039 = ~n3985;
  assign n4012 = ~n3958;
  assign n4127 = ~n3934;
  assign n4303 = ~n4230;
  assign n4351 = n4440 & n4441;
  assign n4129 = ~n3942;
  assign n3569 = ~n3941;
  assign n4040 = ~n3986;
  assign n4130 = ~n3903;
  assign n4014 = ~n3944;
  assign n4013 = ~n3943;
  assign n4268 = ~n4415;
  assign n3571 = ~n3333;
  assign n4352 = n4442 & n4443;
  assign n4011 = ~n3957;
  assign n2913 = ~n2888;
  assign n4020 = ~n3962;
  assign n4017 = ~n3365;
  assign n4019 = ~n3347;
  assign n4302 = ~n4237;
  assign n3615 = ~n3961;
  assign n4270 = ~n4234;
  assign n3631 = ~n3905;
  assign n4021 = ~n3945;
  assign n4024 = ~n3845;
  assign n3573 = ~n3335;
  assign n4051 = ~n3927;
  assign n2648 = n4444 & n4445;
  assign n4304 = ~n4235;
  assign n4028 = ~n3950;
  assign n4027 = ~n3949;
  assign n3575 = ~n3337;
  assign n4030 = ~n3349;
  assign n4025 = ~n3919;
  assign n3567 = ~n3889;
  assign n3609 = ~n3937;
  assign n4031 = ~n3913;
  assign n4035 = ~n3907;
  assign n4029 = ~n3964;
  assign n4034 = ~n3345;
  assign n4033 = ~n3960;
  assign n3802 = n4446 & n4447;
  assign n3577 = ~n3959;
  assign n4037 = ~n3909;
  assign n3579 = ~n3963;
  assign n4132 = ~n3891;
  assign n4272 = ~n3800;
  assign n4274 = ~n4226;
  assign n3581 = ~n3341;
  assign n4133 = ~n3965;
  assign n3583 = ~n3351;
  assign n3011 = ~n2647;
  assign n4042 = ~n3972;
  assign n3587 = ~n3343;
  assign n4043 = ~n3911;
  assign n4041 = ~n3971;
  assign n4054 = ~n3954;
  assign n4053 = ~n3953;
  assign n4058 = ~n3955;
  assign n4057 = ~n3956;
  assign n3585 = ~n3353;
  assign n4045 = ~n3921;
  assign n4048 = ~n3968;
  assign n4047 = ~n3967;
  assign n4050 = ~n3976;
  assign n4056 = ~n3970;
  assign n4049 = ~n3975;
  assign n4055 = ~n3969;
  assign n3798 = n4448 & n4449;
  assign n4135 = ~n3327;
  assign n4059 = ~n4238;
  assign n4062 = ~n3355;
  assign n4061 = ~n3974;
  assign n3589 = ~n3973;
  assign n4305 = ~n4242;
  assign n3591 = ~n4335;
  assign n4276 = ~n4240;
  assign n4137 = ~n3367;
  assign n4306 = ~n4254;
  assign n4064 = ~n3978;
  assign n4065 = ~n3915;
  assign n4063 = ~n3977;
  assign n3593 = ~n3357;
  assign n3595 = ~n3893;
  assign n4068 = ~n3982;
  assign n4278 = ~n4244;
  assign n4067 = ~n3981;
  assign n3597 = ~n3361;
  assign n4280 = ~n3796;
  assign n4113 = ~n3917;
  assign n4307 = ~n4249;
  assign n3599 = ~n3359;
  assign n4070 = ~n3980;
  assign n4069 = ~n3979;
  assign n4282 = ~n4253;
  assign n4071 = ~n3923;
  assign n4074 = ~n3984;
  assign n4073 = ~n3983;
  assign n4076 = ~n3993;
  assign n4284 = ~n4260;
  assign n4075 = ~n3994;
  assign n4288 = ~n4228;
  assign n4078 = ~n3363;
  assign n4077 = ~n3988;
  assign n4121 = ~n3895;
  assign n3601 = ~n3987;
  assign n4080 = ~n4002;
  assign n3603 = ~n3371;
  assign n4286 = ~n4245;
  assign n4081 = ~n3901;
  assign n4138 = ~n4336;
  assign n4079 = ~n4001;
  assign n4140 = ~n3991;
  assign n3605 = ~n3369;
  assign n3607 = ~n3377;
  assign n4290 = ~n4247;
  assign n3847 = n4452 & n4453;
  assign n4084 = ~n3948;
  assign n4085 = ~n4251;
  assign n4298 = ~n4262;
  assign n4083 = ~n3375;
  assign n4119 = ~n3897;
  assign n3611 = ~n3947;
  assign n4091 = ~n3990;
  assign n4090 = ~n3996;
  assign n4088 = ~n3940;
  assign n4089 = ~n3995;
  assign n4022 = ~n3946;
  assign n3613 = ~n3373;
  assign n4096 = ~n3999;
  assign n4087 = ~n3939;
  assign n4093 = ~n3929;
  assign n4095 = ~n4000;
  assign n4115 = ~n3564;
  assign n4296 = ~n4256;
  assign n4098 = ~n4008;
  assign n4018 = ~n3938;
  assign n4099 = ~n3925;
  assign n4097 = ~n3383;
  assign n4101 = ~n3931;
  assign n4142 = ~n4258;
  assign n4104 = ~n4010;
  assign n3619 = ~n4007;
  assign n4103 = ~n3385;
  assign n4108 = ~n3936;
  assign n3621 = ~n4009;
  assign n4105 = ~n4003;
  assign n3623 = ~n3379;
  assign n3843 = n4454 & n4455;
  assign n4308 = ~n4232;
  assign n4016 = ~n3998;
  assign n4143 = ~n4005;
  assign n3625 = ~n3381;
  assign n4354 = n4456 & n4457;
  assign n4015 = ~n3997;
  assign n4131 = ~n3952;
  assign n3627 = ~n3951;
  assign n4107 = ~n3935;
  assign n4123 = ~n3887;
  assign n4117 = ~n3387;
  assign n4125 = ~n3339;
  assign n3629 = ~n3329;
  assign n3633 = ~n3331;
  assign n4300 = ~n4264;
  assign n4109 = ~n3899;
  assign n4355 = n4458 & n4459;
  assign n4356 = n4460 & n4461;
  assign n4111 = ~n4462;
  assign n4266 = ~n4463;
  assign n4023 = ~n4464;
  assign n4359 = n4526 & n4527;
  assign n2765 = ~n4607;
  assign n3284 = n4617 & n4618;
  assign n2645 = n4623 & n4624;
  assign n4224 = n4631 & n4632;
  assign n3804 = n4869 & n4870;
  assign n3849 = n4923 & n4924;
  assign n4450 = ~n4954;
  assign n1817 = n3208 ^ n3209;
  assign n2997 = n3210 ^ n3211;
  assign n1674 = n3212 ^ n3213;
  assign n2995 = n3214 ^ n3215;
  assign n1670 = n3216 ^ n3217;
  assign n1921 = n3218 ^ n3219;
  assign n2826 = n3220 ^ n3221;
  assign n2321 = n3222 ^ n3223;
  assign n2477 = n3224 ^ n3225;
  assign n2406 = n3226 ^ n3227;
  assign n2178 = n3228 ^ n3229;
  assign n1752 = n3230 ^ n3231;
  assign n2156 = n3232 ^ n3233;
  assign n2367 = n3234 ^ n3235;
  assign n1676 = n3236 ^ n3237;
  assign n1848 = n3238 ^ n3239;
  assign n2479 = n3240 ^ n3241;
  assign n2184 = n3242 ^ n3243;
  assign n2739 = n3244 ^ n3245;
  assign n1963 = n3246 ^ n3247;
  assign n1660 = n3248 ^ n3249;
  assign n2185 = n3250 & n3251;
  assign n2445 = n3252 & n3253;
  assign n2892 = n3254 & n3255;
  assign n2556 = n3256 & n3257;
  assign n2820 = n3258 & n3259;
  assign n2255 = n3260 & n3261;
  assign n2032 = n3262 & n3263;
  assign n2449 = n3264 & n3265;
  assign n2055 = n3266 & n3267;
  assign n2295 = n3268 & n3269;
  assign n2822 = n3270 & n3271;
  assign n2561 = n3272 & n3273;
  assign n2193 = n3274 & n3275;
  assign n2880 = n3276 & n3277;
  assign n3002 = n3278 & n3279;
  assign n3195 = n3283 & n3284;
  assign n2871 = n3285 ^ n3286;
  assign n2370 = n3287 ^ n3288;
  assign n3018 = n3289 ^ n3290;
  assign n2889 = n3291 ^ n3292;
  assign n2763 = n3293 ^ n3294;
  assign n2530 = n2316 ^ n2711;
  assign n2440 = n3295 ^ n3296;
  assign n2532 = n3297 ^ n3298;
  assign n2172 = n3299 ^ n3300;
  assign n2031 = n3301 ^ n3302;
  assign n2534 = n3303 ^ n3304;
  assign n2877 = n3305 ^ n3306;
  assign n2540 = n3307 ^ n3308;
  assign n2182 = n3309 ^ n3310;
  assign n2887 = n3311 ^ n3312;
  assign n2546 = n3313 ^ n3314;
  assign n2248 = n3315 ^ n3316;
  assign n2879 = n3317 ^ n3318;
  assign n2528 = n3319 ^ n3320;
  assign n2158 = n3321 ^ n3322;
  assign n2873 = n3323 ^ n3324;
  assign n2230 = n3325 ^ n3326;
  assign n2524 = n3327 ^ n3328;
  assign n2234 = n3329 ^ n3330;
  assign n2164 = n3331 ^ n3332;
  assign n2998 = n3333 ^ n3334;
  assign n2885 = n3335 ^ n3336;
  assign n2883 = n3337 ^ n3338;
  assign n2240 = n3339 ^ n3340;
  assign n2238 = n3341 ^ n3342;
  assign n2538 = n3343 ^ n3344;
  assign n2536 = n3345 ^ n3346;
  assign n2376 = n3347 ^ n3348;
  assign n2242 = n3349 ^ n3350;
  assign n2876 = n3351 ^ n3352;
  assign n2244 = n3353 ^ n3354;
  assign n2174 = n3355 ^ n3356;
  assign n3000 = n3357 ^ n3358;
  assign n2542 = n3359 ^ n3360;
  assign n2548 = n3361 ^ n3362;
  assign n2544 = n3363 ^ n3364;
  assign n2874 = n3365 ^ n3366;
  assign n3008 = n3367 ^ n3368;
  assign n2550 = n3369 ^ n3370;
  assign n2878 = n3371 ^ n3372;
  assign n3001 = n3373 ^ n3374;
  assign n2522 = n3375 ^ n3376;
  assign n2881 = n3377 ^ n3378;
  assign n2552 = n3379 ^ n3380;
  assign n2891 = n3381 ^ n3382;
  assign n2236 = n3383 ^ n3384;
  assign n2761 = n3385 ^ n3386;
  assign n2516 = n3387 ^ n3388;
  assign n2286 = ~n2170;
  assign n3176 = ~n3522;
  assign n3178 = ~n3525;
  assign n3180 = ~n3528;
  assign n3184 = ~n3532;
  assign n3190 = ~n3543;
  assign n3174 = ~n3545;
  assign n3414 = n3239 & n3557;
  assign n3186 = ~n3559;
  assign n3188 = ~n3560;
  assign n3418 = n3304 & n3563;
  assign n3420 = n3298 & n3297;
  assign n3192 = ~n3283;
  assign n2954 = ~n2442;
  assign n2371 = n3564 ^ n3565;
  assign n2801 = ~n2605;
  assign n3419 = ~n3304;
  assign n2803 = ~n2619;
  assign n3404 = ~n3231;
  assign n2805 = ~n2607;
  assign n3406 = ~n3298;
  assign n3016 = ~n2526;
  assign n3014 = ~n2611;
  assign n2983 = ~n2609;
  assign n1768 = n3798 ^ n3799;
  assign n1954 = n3802 ^ n3803;
  assign n2823 = n3804 ^ n3805;
  assign n3514 = n3806 & n3807;
  assign n3529 = n3822 & n3823;
  assign n2872 = n3843 ^ n3844;
  assign n3282 = ~n3223;
  assign n2909 = ~n2629;
  assign n2627 = n3847 ^ n3848;
  assign n2635 = n3849 ^ n3850;
  assign n3667 = n4011 & n4012;
  assign n3668 = n4013 & n4014;
  assign n3669 = n4015 & n4016;
  assign n3672 = n4017 & n4018;
  assign n3675 = n4019 & n4020;
  assign n3676 = n4021 & n4022;
  assign n3677 = n4023 & n4024;
  assign n3678 = n4025 & n4026;
  assign n3679 = n4027 & n4028;
  assign n3680 = n4029 & n4030;
  assign n3681 = n4031 & n4032;
  assign n3682 = n4033 & n4034;
  assign n3683 = n4035 & n4036;
  assign n3684 = n4037 & n4038;
  assign n3685 = n4039 & n4040;
  assign n3686 = n4041 & n4042;
  assign n3687 = n4043 & n4044;
  assign n3688 = n4045 & n4046;
  assign n3689 = n4047 & n4048;
  assign n3690 = n4049 & n4050;
  assign n3691 = n4051 & n4052;
  assign n3692 = n4053 & n4054;
  assign n3693 = n4055 & n4056;
  assign n3694 = n4057 & n4058;
  assign n3695 = n4059 & n4060;
  assign n3696 = n4061 & n4062;
  assign n3697 = n4063 & n4064;
  assign n3698 = n4065 & n4066;
  assign n3699 = n4067 & n4068;
  assign n3700 = n4069 & n4070;
  assign n3701 = n4071 & n4072;
  assign n3702 = n4073 & n4074;
  assign n3703 = n4075 & n4076;
  assign n3704 = n4077 & n4078;
  assign n3705 = n4079 & n4080;
  assign n3708 = n4081 & n4082;
  assign n3709 = n4083 & n4084;
  assign n3710 = n4085 & n4086;
  assign n3711 = n4087 & n4088;
  assign n3712 = n4089 & n4090;
  assign n3713 = n4091 & n4092;
  assign n3714 = n4093 & n4094;
  assign n3715 = n4095 & n4096;
  assign n3716 = n4097 & n4098;
  assign n3717 = n4099 & n4100;
  assign n3718 = n4101 & n4102;
  assign n3719 = n4103 & n4104;
  assign n3720 = n4105 & n4106;
  assign n3721 = n4107 & n4108;
  assign n3722 = n4109 & n4110;
  assign n3723 = n4111 & n4112;
  assign n3724 = n4113 & n4114;
  assign n3725 = n4115 & n4116;
  assign n3726 = n4117 & n4118;
  assign n3729 = n4119 & n4120;
  assign n3730 = n4121 & n4122;
  assign n3731 = n4123 & n4124;
  assign n3732 = n4125 & n4126;
  assign n3733 = n4127 & n3933;
  assign n3658 = ~n4128;
  assign n3734 = n4129 & n3296;
  assign n3735 = n4130 & n3904;
  assign n3736 = n4131 & n3326;
  assign n3737 = n4132 & n3892;
  assign n3738 = n4133 & n3966;
  assign n3582 = ~n4134;
  assign n3739 = n4135 & n4136;
  assign n3740 = n4137 & n3894;
  assign n3741 = n4138 & n4139;
  assign n3742 = n4140 & n3992;
  assign n3604 = ~n4141;
  assign n3743 = n4142 & n3243;
  assign n3744 = n4143 & n4006;
  assign n3624 = ~n4144;
  assign n3568 = ~n4145;
  assign n3661 = ~n4146;
  assign n3626 = ~n4147;
  assign n3655 = ~n4148;
  assign n3580 = ~n4149;
  assign n3666 = ~n4150;
  assign n3590 = ~n4151;
  assign n3594 = ~n4152;
  assign n3634 = ~n4153;
  assign n3566 = ~n4154;
  assign n3660 = ~n4155;
  assign n3570 = ~n4156;
  assign n3608 = ~n4157;
  assign n3614 = ~n4158;
  assign n3636 = ~n4159;
  assign n3572 = ~n4160;
  assign n3574 = ~n4161;
  assign n3576 = ~n4162;
  assign n3578 = ~n4163;
  assign n3618 = ~n4164;
  assign n3638 = ~n4165;
  assign n3584 = ~n4166;
  assign n3586 = ~n4167;
  assign n3632 = ~n4168;
  assign n3640 = ~n4169;
  assign n3620 = ~n4170;
  assign n3662 = ~n4171;
  assign n3663 = ~n4172;
  assign n3588 = ~n4173;
  assign n3745 = n3802 & n4174;
  assign n3592 = ~n4175;
  assign n3596 = ~n4176;
  assign n3598 = ~n4177;
  assign n3642 = ~n4178;
  assign n3644 = ~n4179;
  assign n3646 = ~n4180;
  assign n3600 = ~n4181;
  assign n3602 = ~n4182;
  assign n3606 = ~n4183;
  assign n3610 = ~n4184;
  assign n3612 = ~n4185;
  assign n3616 = ~n4186;
  assign n3664 = ~n4187;
  assign n3651 = ~n4188;
  assign n3653 = ~n4189;
  assign n3622 = ~n4190;
  assign n3649 = ~n4191;
  assign n3630 = ~n4192;
  assign n3628 = ~n4193;
  assign n3206 = n4224 ^ n4225;
  assign n3851 = n4266 & n4267;
  assign n3852 = n4268 & n4269;
  assign n3853 = n4270 & n4271;
  assign n3854 = n4272 & n4273;
  assign n3855 = n4274 & n4275;
  assign n3856 = n4276 & n4277;
  assign n3857 = n4278 & n4279;
  assign n3858 = n4280 & n4281;
  assign n3859 = n4282 & n4283;
  assign n3860 = n4284 & n4285;
  assign n3861 = n4286 & n4287;
  assign n3862 = n4288 & n4289;
  assign n3863 = n4290 & n4291;
  assign n3868 = n4296 & n4297;
  assign n3869 = n4298 & n4299;
  assign n3870 = n4300 & n4301;
  assign n3875 = n4302 & n3221;
  assign n3876 = n4303 & n3213;
  assign n3877 = n4304 & n4236;
  assign n3878 = n4305 & n3225;
  assign n3879 = n4306 & n4255;
  assign n3880 = n4307 & n3233;
  assign n3882 = n4308 & n4233;
  assign n3518 = ~n4309;
  assign n3883 = n3798 & n4310;
  assign n3520 = ~n4311;
  assign n3526 = ~n4312;
  assign n3530 = ~n4313;
  assign n3558 = ~n4314;
  assign n3562 = ~n4315;
  assign n3884 = n3843 & n4316;
  assign n3548 = ~n4317;
  assign n3516 = ~n4318;
  assign n1985 = ~n4320;
  assign n3546 = ~n4321;
  assign n3523 = ~n4322;
  assign n3550 = ~n4323;
  assign n3281 = ~n4324;
  assign n3551 = ~n4325;
  assign n3885 = n3850 & n3849;
  assign n3555 = ~n4326;
  assign n3553 = ~n4327;
  assign n2681 = ~n4328;
  assign n3533 = ~n4329;
  assign n3535 = ~n4330;
  assign n3886 = n3847 & n3848;
  assign n3539 = ~n4332;
  assign n3561 = ~n4333;
  assign n3541 = ~n4334;
  assign n3706 = ~n4350;
  assign n3425 = ~n4351;
  assign n3670 = ~n4352;
  assign n2665 = ~n2648;
  assign n3727 = ~n3802;
  assign n3873 = ~n3798;
  assign n3864 = ~n3847;
  assign n3881 = ~n3843;
  assign n3673 = ~n4354;
  assign n3390 = ~n4355;
  assign n3429 = ~n4356;
  assign n2262 = ~n4359;
  assign n4319 = n4224 & n4225;
  assign n4331 = n3804 & n4419;
  assign n3193 = ~n3284;
  assign n2659 = ~n2645;
  assign n4292 = ~n4224;
  assign n4353 = n4450 & n4451;
  assign n4294 = ~n3804;
  assign n3871 = ~n3849;
  assign n1626 = n2820 ^ n2821;
  assign n1820 = n2822 ^ n2823;
  assign n2022 = n2295 ^ n2824;
  assign n2444 = n2870 ^ n2871;
  assign n2454 = n2872 ^ n2873;
  assign n2446 = n2874 ^ n2875;
  assign n2450 = n2876 ^ n2877;
  assign n2458 = n2878 ^ n2879;
  assign n2437 = n2880 ^ n2881;
  assign n2452 = n2888 ^ n2889;
  assign n1819 = n2995 ^ n2996;
  assign n1829 = n2997 ^ n2850;
  assign n1831 = n1670 ^ n1952;
  assign n1833 = n2998 ^ n2999;
  assign n1838 = n1674 ^ n1768;
  assign n2405 = n3000 ^ n2852;
  assign n1823 = n3001 ^ n2857;
  assign n1827 = n3002 ^ n3003;
  assign n2848 = n2997 & n3004;
  assign n2853 = n3000 & n3005;
  assign n2855 = n2546 & n3006;
  assign n2858 = n3001 & n3007;
  assign n2859 = n2998 & n2999;
  assign n2860 = n2556 & n2168;
  assign n2861 = n2820 & n2821;
  assign n2862 = n2321 & n2741;
  assign n2863 = n2995 & n2996;
  assign n2864 = n2477 & n2138;
  assign n2866 = n2544 & n2178;
  assign n2867 = n2156 & n3008;
  assign n2868 = n2822 & n2823;
  assign n2869 = n3002 & n3003;
  assign n2919 = n2238 & n3011;
  assign n2928 = n2236 & n3014;
  assign n2929 = n2445 & n3015;
  assign n2930 = n2185 & n3016;
  assign n2931 = n2871 & n2870;
  assign n2933 = n2889 & n2888;
  assign n2934 = n2172 & n2538;
  assign n2937 = n2248 & n2629;
  assign n2938 = n2879 & n2878;
  assign n2939 = n2158 & n2522;
  assign n2940 = n2880 & n2881;
  assign n1885 = ~n1817;
  assign n2849 = ~n2997;
  assign n2835 = ~n2995;
  assign n2085 = ~n1921;
  assign n2846 = ~n2826;
  assign n2839 = ~n2321;
  assign n2843 = ~n2477;
  assign n2842 = ~n2178;
  assign n1951 = ~n1752;
  assign n2847 = ~n2156;
  assign n2514 = ~n2367;
  assign n1973 = ~n1848;
  assign n2507 = ~n2479;
  assign n2757 = ~n2184;
  assign n2511 = ~n2739;
  assign n1533 = ~n1963;
  assign n2081 = ~n1660;
  assign n2917 = ~n2185;
  assign n2762 = n3174 & n3175;
  assign n2916 = ~n2445;
  assign n2336 = ~n2892;
  assign n2447 = n3176 & n3177;
  assign n2827 = ~n2556;
  assign n2829 = ~n2820;
  assign n2257 = n3178 & n3179;
  assign n2302 = ~n2255;
  assign n2268 = ~n2032;
  assign n2341 = ~n2449;
  assign n2187 = n3180 & n3181;
  assign n2306 = ~n2055;
  assign n2455 = n3184 & n3185;
  assign n1955 = n3186 & n3187;
  assign n3048 = n3188 & n3189;
  assign n2079 = ~n2295;
  assign n2831 = ~n2822;
  assign n2330 = ~n2561;
  assign n2282 = ~n2193;
  assign n2902 = ~n2880;
  assign n2833 = ~n3002;
  assign n2760 = n3190 & n3191;
  assign n3063 = n3192 & n3193;
  assign n1347 = ~n3195;
  assign n2904 = ~n2871;
  assign n2568 = ~n2370;
  assign n2897 = ~n3018;
  assign n2912 = ~n2889;
  assign n2772 = ~n2763;
  assign n2922 = ~n2440;
  assign n2906 = ~n2172;
  assign n2052 = ~n2031;
  assign n2923 = ~n2877;
  assign n2789 = ~n2540;
  assign n2790 = ~n2182;
  assign n2901 = ~n2887;
  assign n2854 = ~n2546;
  assign n2908 = ~n2248;
  assign n2914 = ~n2879;
  assign n2785 = ~n2528;
  assign n2910 = ~n2158;
  assign n2083 = ~n2230;
  assign n2794 = ~n2524;
  assign n2310 = ~n2234;
  assign n2585 = ~n2164;
  assign n2837 = ~n2998;
  assign n2355 = ~n2885;
  assign n2570 = ~n2883;
  assign n2314 = ~n2240;
  assign n2927 = ~n2238;
  assign n2907 = ~n2538;
  assign n2573 = ~n2536;
  assign n2571 = ~n2376;
  assign n2312 = ~n2242;
  assign n2924 = ~n2876;
  assign n2899 = ~n2244;
  assign n2575 = ~n2174;
  assign n2851 = ~n3000;
  assign n2577 = ~n2542;
  assign n2579 = ~n2548;
  assign n2841 = ~n2544;
  assign n2505 = ~n2874;
  assign n2520 = ~n3008;
  assign n2791 = ~n2550;
  assign n2915 = ~n2878;
  assign n2856 = ~n3001;
  assign n2911 = ~n2522;
  assign n2903 = ~n2881;
  assign n2582 = ~n2552;
  assign n2925 = ~n2891;
  assign n2926 = ~n2236;
  assign n2775 = ~n2761;
  assign n2359 = ~n2516;
  assign n2759 = n3206 ^ n3207;
  assign n3194 = n3281 & n3282;
  assign n3197 = n3404 & n3405;
  assign n3198 = n3406 & n3407;
  assign n3042 = ~n3414;
  assign n2671 = ~n3418;
  assign n3200 = n3419 & n3303;
  assign n2683 = ~n3420;
  assign n2699 = ~n2371;
  assign n1949 = ~n1768;
  assign n1766 = ~n1954;
  assign n2832 = ~n2823;
  assign n3170 = ~n3514;
  assign n3391 = n3516 & n3517;
  assign n3392 = n3518 & n3519;
  assign n3395 = n3520 & n3521;
  assign n3396 = n3523 & n3524;
  assign n3397 = n3526 & n3527;
  assign n3182 = ~n3529;
  assign n3398 = n3530 & n3531;
  assign n3399 = n3533 & n3534;
  assign n3400 = n3535 & n3536;
  assign n3402 = n3539 & n3540;
  assign n3403 = n3541 & n3542;
  assign n3408 = n3546 & n3547;
  assign n3409 = n3548 & n3549;
  assign n3410 = n3550 & n3208;
  assign n3411 = n3551 & n3552;
  assign n3412 = n3553 & n3554;
  assign n3413 = n3555 & n3556;
  assign n3415 = n3558 & n3245;
  assign n3416 = n3561 & n3247;
  assign n3417 = n3562 & n3214;
  assign n3421 = n3566 & n3567;
  assign n3426 = n3568 & n3569;
  assign n3427 = n3570 & n3571;
  assign n3430 = n3572 & n3573;
  assign n3433 = n3574 & n3575;
  assign n3436 = n3576 & n3577;
  assign n3439 = n3578 & n3579;
  assign n3440 = n3580 & n3581;
  assign n3441 = n3582 & n3583;
  assign n3446 = n3584 & n3585;
  assign n3447 = n3586 & n3587;
  assign n3450 = n3588 & n3589;
  assign n3451 = n3590 & n3591;
  assign n3454 = n3592 & n3593;
  assign n3455 = n3594 & n3595;
  assign n3456 = n3596 & n3597;
  assign n3457 = n3598 & n3599;
  assign n3460 = n3600 & n3601;
  assign n3463 = n3602 & n3603;
  assign n3464 = n3604 & n3605;
  assign n3465 = n3606 & n3607;
  assign n3466 = n3608 & n3609;
  assign n3469 = n3610 & n3611;
  assign n3470 = n3612 & n3613;
  assign n3473 = n3614 & n3615;
  assign n3474 = n3616 & n3617;
  assign n3479 = n3618 & n3619;
  assign n3480 = n3620 & n3621;
  assign n3481 = n3622 & n3623;
  assign n3482 = n3624 & n3625;
  assign n3485 = n3626 & n3627;
  assign n3486 = n3628 & n3629;
  assign n3487 = n3630 & n3631;
  assign n3488 = n3632 & n3633;
  assign n3491 = n3634 & n3635;
  assign n3492 = n3636 & n3637;
  assign n3495 = n3638 & n3639;
  assign n3496 = n3640 & n3641;
  assign n3497 = n3642 & n3643;
  assign n3498 = n3644 & n3645;
  assign n3499 = n3646 & n3647;
  assign n3500 = n3649 & n3650;
  assign n3501 = n3651 & n3652;
  assign n3502 = n3653 & n3654;
  assign n3503 = n3655 & n3656;
  assign n3504 = n3658 & n3288;
  assign n3505 = n3660 & n3320;
  assign n3506 = n3661 & n3289;
  assign n3507 = n3662 & n3308;
  assign n3508 = n3663 & n3310;
  assign n3509 = n3664 & n3324;
  assign n3510 = n3666 & n3292;
  assign n3067 = ~n3667;
  assign n3075 = ~n3668;
  assign n3077 = ~n3669;
  assign n2642 = n3670 & n3671;
  assign n3079 = ~n3672;
  assign n2890 = n3673 & n3674;
  assign n3081 = ~n3675;
  assign n3157 = ~n3676;
  assign n3428 = ~n3677;
  assign n3422 = ~n3678;
  assign n3085 = ~n3679;
  assign n3083 = ~n3680;
  assign n3431 = ~n3681;
  assign n3087 = ~n3682;
  assign n3434 = ~n3683;
  assign n3437 = ~n3684;
  assign n3065 = ~n3685;
  assign n3093 = ~n3686;
  assign n3444 = ~n3687;
  assign n3442 = ~n3688;
  assign n3095 = ~n3689;
  assign n3097 = ~n3690;
  assign n3483 = ~n3691;
  assign n3099 = ~n3692;
  assign n3101 = ~n3693;
  assign n3103 = ~n3694;
  assign n3448 = ~n3695;
  assign n3107 = ~n3696;
  assign n3111 = ~n3697;
  assign n3452 = ~n3698;
  assign n3113 = ~n3699;
  assign n3117 = ~n3700;
  assign n3458 = ~n3701;
  assign n3119 = ~n3702;
  assign n3121 = ~n3703;
  assign n3123 = ~n3704;
  assign n3127 = ~n3705;
  assign n3201 = n3706 & n3707;
  assign n3461 = ~n3708;
  assign n3135 = ~n3709;
  assign n3467 = ~n3710;
  assign n3137 = ~n3711;
  assign n3139 = ~n3712;
  assign n3141 = ~n3713;
  assign n3471 = ~n3714;
  assign n3143 = ~n3715;
  assign n3147 = ~n3716;
  assign n3475 = ~n3717;
  assign n3477 = ~n3718;
  assign n3149 = ~n3719;
  assign n3153 = ~n3720;
  assign n3161 = ~n3721;
  assign n3489 = ~n3722;
  assign n3424 = ~n3723;
  assign n3115 = ~n3724;
  assign n3145 = ~n3725;
  assign n3167 = ~n3726;
  assign n3511 = n3727 & n3728;
  assign n3133 = ~n3729;
  assign n3125 = ~n3730;
  assign n3165 = ~n3731;
  assign n3163 = ~n3732;
  assign n3069 = ~n3733;
  assign n3071 = ~n3734;
  assign n3073 = ~n3735;
  assign n3159 = ~n3736;
  assign n3089 = ~n3737;
  assign n3091 = ~n3738;
  assign n3105 = ~n3739;
  assign n3109 = ~n3740;
  assign n3129 = ~n3741;
  assign n3131 = ~n3742;
  assign n3151 = ~n3743;
  assign n3155 = ~n3744;
  assign n3493 = ~n3745;
  assign n3544 = n2262 & n2765;
  assign n3389 = ~n3851;
  assign n1632 = ~n3852;
  assign n3060 = ~n3853;
  assign n3027 = ~n3854;
  assign n3029 = ~n3855;
  assign n2895 = ~n3856;
  assign n3035 = ~n3857;
  assign n3037 = ~n3858;
  assign n3041 = ~n3859;
  assign n2111 = ~n3860;
  assign n3045 = ~n3861;
  assign n3062 = ~n3862;
  assign n3047 = ~n3863;
  assign n3648 = n3864 & n3865;
  assign n3052 = ~n3868;
  assign n3054 = ~n3869;
  assign n3058 = ~n3870;
  assign n3657 = n3871 & n3872;
  assign n3659 = n3873 & n3874;
  assign n3023 = ~n3875;
  assign n3021 = ~n3876;
  assign n3025 = ~n3877;
  assign n3031 = ~n3878;
  assign n3033 = ~n3879;
  assign n3039 = ~n3880;
  assign n3665 = n3881 & n3844;
  assign n3056 = ~n3882;
  assign n3393 = ~n3883;
  assign n3013 = ~n3884;
  assign n2695 = ~n3885;
  assign n2687 = ~n3886;
  assign n3866 = n4292 & n4293;
  assign n3867 = n4294 & n4295;
  assign n3512 = ~n4319;
  assign n3537 = ~n4331;
  assign n3205 = ~n4353;
  assign n990 = n2405 ^ n2406;
  assign n1441 = n2437 ^ n2438;
  assign n1401 = n2445 ^ n2446;
  assign n1789 = n2449 ^ n2450;
  assign n1852 = n1955 ^ n1676;
  assign n2471 = ~n2454;
  assign n2324 = n2760 ^ n2761;
  assign n2165 = n2762 ^ n2763;
  assign n2742 = n2827 & n2828;
  assign n2743 = n2829 & n2830;
  assign n2744 = n2831 & n2832;
  assign n2745 = n2833 & n2834;
  assign n2746 = n2835 & n2836;
  assign n2747 = n2837 & n2838;
  assign n2748 = n2839 & n2840;
  assign n2749 = n2841 & n2842;
  assign n2750 = n2843 & n2844;
  assign n2752 = n2847 & n2520;
  assign n1856 = ~n2848;
  assign n2753 = n2849 & n2850;
  assign n2754 = n2851 & n2852;
  assign n2737 = ~n2853;
  assign n2755 = n2854 & n2180;
  assign n2734 = ~n2855;
  assign n2756 = n2856 & n2857;
  assign n1971 = ~n2858;
  assign n1905 = ~n2859;
  assign n2728 = ~n2860;
  assign n1662 = ~n2861;
  assign n2731 = ~n2862;
  assign n1879 = ~n2863;
  assign n2025 = ~n2864;
  assign n2736 = ~n2866;
  assign n2027 = ~n2867;
  assign n1877 = ~n2868;
  assign n1911 = ~n2869;
  assign n2460 = n2890 ^ n2891;
  assign n2773 = n2902 & n2903;
  assign n2776 = n2904 & n2905;
  assign n2777 = n2906 & n2907;
  assign n2778 = n2908 & n2909;
  assign n2779 = n2910 & n2911;
  assign n2780 = n2912 & n2913;
  assign n2781 = n2914 & n2915;
  assign n2782 = n2916 & n2875;
  assign n2783 = n2917 & n2526;
  assign n2040 = ~n2919;
  assign n2787 = n2923 & n2876;
  assign n2788 = n2877 & n2924;
  assign n2792 = n2890 & n2925;
  assign n2793 = n2926 & n2611;
  assign n2795 = n2927 & n2647;
  assign n2501 = ~n2928;
  assign n2504 = ~n2929;
  assign n2485 = ~n2930;
  assign n2796 = n2760 & n2761;
  assign n2483 = ~n2931;
  assign n2797 = n2763 & n2762;
  assign n2481 = ~n2933;
  assign n2487 = ~n2934;
  assign n2493 = ~n2937;
  assign n2495 = ~n2938;
  assign n2499 = ~n2939;
  assign n2508 = ~n2940;
  assign n2921 = n3013 & n2873;
  assign n2771 = ~n2762;
  assign n2767 = ~n2447;
  assign n2300 = ~n2257;
  assign n2271 = ~n2187;
  assign n1843 = n3042 & n3043;
  assign n2491 = ~n2455;
  assign n1756 = ~n1955;
  assign n2469 = ~n3048;
  assign n2774 = ~n2760;
  assign n1097 = ~n3063;
  assign n2503 = ~n2759;
  assign n3019 = n3170 & n3171;
  assign n2740 = n3182 & n3183;
  assign n2894 = ~n3194;
  assign n2951 = ~n3197;
  assign n2109 = ~n3198;
  assign n2101 = ~n3200;
  assign n65 = n3201 ^ n3202;
  assign n12378 = n3204 ^ n3205;
  assign n3017 = n3389 & n3390;
  assign n3061 = ~n3391;
  assign n3020 = ~n3392;
  assign n3196 = n3393 & n3394;
  assign n3024 = ~n3395;
  assign n3026 = ~n3396;
  assign n3030 = ~n3397;
  assign n3038 = ~n3398;
  assign n3044 = ~n3399;
  assign n3046 = ~n3400;
  assign n3051 = ~n3402;
  assign n3057 = ~n3403;
  assign n3199 = n1632 & n1985;
  assign n3059 = ~n3408;
  assign n3022 = ~n3409;
  assign n3028 = ~n3410;
  assign n3034 = ~n3411;
  assign n3036 = ~n3412;
  assign n3040 = ~n3413;
  assign n3032 = ~n3415;
  assign n3053 = ~n3416;
  assign n3055 = ~n3417;
  assign n3162 = ~n3421;
  assign n2943 = n3422 & n3423;
  assign n2956 = n3424 & n3425;
  assign n3070 = ~n3426;
  assign n3074 = ~n3427;
  assign n2893 = n3428 & n3429;
  assign n3156 = ~n3430;
  assign n2958 = n3431 & n3432;
  assign n3084 = ~n3433;
  assign n2884 = n3434 & n3435;
  assign n3086 = ~n3436;
  assign n2882 = n3437 & n3438;
  assign n3082 = ~n3439;
  assign n3088 = ~n3440;
  assign n3090 = ~n3441;
  assign n2825 = n3442 & n3443;
  assign n2652 = n3444 & n3445;
  assign n3092 = ~n3446;
  assign n3098 = ~n3447;
  assign n2259 = n3448 & n3449;
  assign n3106 = ~n3450;
  assign n3104 = ~n3451;
  assign n2655 = n3452 & n3453;
  assign n3110 = ~n3454;
  assign n3108 = ~n3455;
  assign n3112 = ~n3456;
  assign n3114 = ~n3457;
  assign n2886 = n3458 & n3459;
  assign n3122 = ~n3460;
  assign n2941 = n3461 & n3462;
  assign n3124 = ~n3463;
  assign n3130 = ~n3464;
  assign n3126 = ~n3465;
  assign n3078 = ~n3466;
  assign n2945 = n3467 & n3468;
  assign n3134 = ~n3469;
  assign n3138 = ~n3470;
  assign n2061 = n3471 & n3472;
  assign n3080 = ~n3473;
  assign n3144 = ~n3474;
  assign n2960 = n3475 & n3476;
  assign n2059 = n3477 & n3478;
  assign n3146 = ~n3479;
  assign n3148 = ~n3480;
  assign n3152 = ~n3481;
  assign n3154 = ~n3482;
  assign n2251 = n3483 & n3484;
  assign n3158 = ~n3485;
  assign n3160 = ~n3486;
  assign n3166 = ~n3487;
  assign n3164 = ~n3488;
  assign n2947 = n3489 & n3490;
  assign n3064 = ~n3491;
  assign n3066 = ~n3492;
  assign n3203 = n3493 & n3494;
  assign n3094 = ~n3495;
  assign n3102 = ~n3496;
  assign n3116 = ~n3497;
  assign n3118 = ~n3498;
  assign n3120 = ~n3499;
  assign n3140 = ~n3500;
  assign n3142 = ~n3501;
  assign n3136 = ~n3502;
  assign n3150 = ~n3503;
  assign n3068 = ~n3504;
  assign n3076 = ~n3505;
  assign n3072 = ~n3506;
  assign n3100 = ~n3507;
  assign n3096 = ~n3508;
  assign n3132 = ~n3509;
  assign n3128 = ~n3510;
  assign n2663 = ~n2642;
  assign n3012 = ~n2890;
  assign n2963 = ~n3511;
  assign n3280 = n3512 & n3513;
  assign n3401 = n3537 & n3538;
  assign n2819 = ~n3544;
  assign n2119 = ~n3648;
  assign n2130 = ~n3657;
  assign n2950 = ~n3659;
  assign n2497 = ~n3665;
  assign n3515 = n3205 & n3808;
  assign n3010 = ~n3866;
  assign n3050 = ~n3867;
  assign n1273 = ~n990;
  assign n1592 = ~n1441;
  assign n1960 = ~n1789;
  assign n2353 = n2504 & n2505;
  assign n2357 = n2508 & n2509;
  assign n2155 = n2469 ^ n2520;
  assign n2472 = n2737 & n2406;
  assign n2320 = n2740 ^ n2741;
  assign n2144 = ~n2742;
  assign n1367 = ~n2743;
  assign n1512 = ~n2744;
  assign n1544 = ~n2745;
  assign n1496 = ~n2746;
  assign n1535 = ~n2747;
  assign n2148 = ~n2748;
  assign n2154 = ~n2749;
  assign n2465 = ~n2750;
  assign n2468 = ~n2752;
  assign n1500 = ~n2753;
  assign n2150 = ~n2754;
  assign n2152 = ~n2755;
  assign n1590 = ~n2756;
  assign n2580 = n2771 & n2772;
  assign n2220 = ~n2773;
  assign n2583 = n2774 & n2775;
  assign n2198 = ~n2776;
  assign n2204 = ~n2777;
  assign n2210 = ~n2778;
  assign n2217 = ~n2779;
  assign n2224 = ~n2780;
  assign n2212 = ~n2781;
  assign n2586 = n1097 & n1347;
  assign n2200 = ~n2782;
  assign n2202 = ~n2783;
  assign n2042 = ~n2787;
  assign n2340 = ~n2788;
  assign n2348 = ~n2792;
  assign n2222 = ~n2793;
  assign n2338 = ~n2795;
  assign n2351 = ~n2796;
  assign n2226 = ~n2797;
  assign n2436 = n2825 ^ n2826;
  assign n2441 = n2882 ^ n2883;
  assign n2448 = n2884 ^ n2885;
  assign n2456 = n2886 ^ n2887;
  assign n2439 = n2892 ^ n2893;
  assign n2475 = n2894 & n2895;
  assign n2496 = ~n2921;
  assign n2786 = n2893 & n2922;
  assign n2798 = n2884 & n2447;
  assign n1341 = n2941 ^ n2942;
  assign n1957 = n2943 ^ n2944;
  assign n2474 = n2945 ^ n2946;
  assign n2160 = n2947 ^ n2948;
  assign n1744 = n2951 & n2952;
  assign n1875 = ~n1843;
  assign n2369 = n2956 ^ n2957;
  assign n2374 = n2958 ^ n2959;
  assign n2372 = n2960 ^ n2961;
  assign n2865 = n2825 & n2826;
  assign n2920 = n3012 & n2891;
  assign n2932 = n3017 & n3018;
  assign n2935 = n2655 & n2244;
  assign n2936 = n2886 & n2887;
  assign n2196 = ~n3019;
  assign n2377 = n3020 & n3021;
  assign n2451 = n3022 & n3023;
  assign n2553 = n3024 & n3025;
  assign n2555 = n3026 & n3027;
  assign n2373 = n3028 & n3029;
  assign n2539 = n3030 & n3031;
  assign n2435 = n3032 & n3033;
  assign n2557 = n3034 & n3035;
  assign n2732 = ~n2740;
  assign n2249 = n3036 & n3037;
  assign n2559 = n3038 & n3039;
  assign n2476 = n3040 & n3041;
  assign n2545 = n3044 & n3045;
  assign n2543 = n3046 & n3047;
  assign n2057 = n3051 & n3052;
  assign n2141 = n3053 & n3054;
  assign n2521 = n3055 & n3056;
  assign n2459 = n3057 & n3058;
  assign n2525 = n3059 & n3060;
  assign n2323 = n3061 & n3062;
  assign n2955 = n2882 & n2442;
  assign n2604 = n3064 & n3065;
  assign n2453 = n3066 & n3067;
  assign n2443 = n3068 & n3069;
  assign n2253 = n3070 & n3071;
  assign n2758 = n3072 & n3073;
  assign n2644 = n3074 & n3075;
  assign n2523 = n3076 & n3077;
  assign n2643 = n3078 & n3079;
  assign n2614 = n3080 & n3081;
  assign n2649 = n3082 & n3083;
  assign n2612 = n3084 & n3085;
  assign n2616 = n3086 & n3087;
  assign n2533 = n3088 & n3089;
  assign n2620 = n3090 & n3091;
  assign n2646 = n3092 & n3093;
  assign n2537 = n3094 & n3095;
  assign n2653 = n3096 & n3097;
  assign n2618 = n3098 & n3099;
  assign n2799 = n3100 & n3101;
  assign n2535 = n3102 & n3103;
  assign n2606 = n3104 & n3105;
  assign n2622 = n3106 & n3107;
  assign n2560 = n3108 & n3109;
  assign n2558 = n3110 & n3111;
  assign n2654 = n3112 & n3113;
  assign n2651 = n3114 & n3115;
  assign n2650 = n3116 & n3117;
  assign n2541 = n3118 & n3119;
  assign n2189 = n3120 & n3121;
  assign n2657 = n3122 & n3123;
  assign n2547 = n3124 & n3125;
  assign n2632 = n3126 & n3127;
  assign n2531 = n3128 & n3129;
  assign n2624 = n3130 & n3131;
  assign n2738 = n3132 & n3133;
  assign n2626 = n3134 & n3135;
  assign n2527 = n3136 & n3137;
  assign n2628 = n3138 & n3139;
  assign n2549 = n3140 & n3141;
  assign n2457 = n3142 & n3143;
  assign n2630 = n3144 & n3145;
  assign n2640 = n3146 & n3147;
  assign n2636 = n3148 & n3149;
  assign n2478 = n3150 & n3151;
  assign n2562 = n3152 & n3153;
  assign n2551 = n3154 & n3155;
  assign n2554 = n3156 & n3157;
  assign n2634 = n3158 & n3159;
  assign n2608 = n3160 & n3161;
  assign n2529 = n3162 & n3163;
  assign n2610 = n3164 & n3165;
  assign n2638 = n3166 & n3167;
  assign n2986 = n2941 & n3168;
  assign n2987 = n2956 & n2957;
  assign n2988 = n2958 & n2959;
  assign n2989 = n2943 & n3169;
  assign n2990 = n2259 & n2623;
  assign n2991 = n2061 & n2641;
  assign n2992 = n2960 & n2961;
  assign n2993 = n2059 & n2637;
  assign n2994 = n2251 & n2609;
  assign n2896 = ~n3017;
  assign n2949 = ~n3196;
  assign n1979 = ~n3199;
  assign n2964 = ~n2943;
  assign n2970 = ~n2956;
  assign n2918 = ~n2893;
  assign n2976 = ~n2958;
  assign n2766 = ~n2884;
  assign n2953 = ~n2882;
  assign n2845 = ~n2825;
  assign n2673 = ~n2652;
  assign n2972 = ~n2259;
  assign n2898 = ~n2655;
  assign n2900 = ~n2886;
  assign n2984 = ~n2941;
  assign n2966 = ~n2945;
  assign n2978 = ~n2061;
  assign n2974 = ~n2960;
  assign n2980 = ~n2059;
  assign n2982 = ~n2251;
  assign n2968 = ~n2947;
  assign n2962 = ~n3203;
  assign n3009 = ~n3280;
  assign n3049 = ~n3401;
  assign n3172 = ~n3515;
  assign n1214 = n2155 ^ n2156;
  assign n1190 = n2320 ^ n2321;
  assign n1306 = n2323 ^ n2324;
  assign n2269 = n2340 & n2341;
  assign n2199 = ~n2353;
  assign n2219 = ~n2357;
  assign n2227 = n2369 ^ n2370;
  assign n1958 = n2371 ^ n2372;
  assign n2030 = n2373 ^ n2374;
  assign n1567 = n2435 ^ n2436;
  assign n1443 = n2439 ^ n2440;
  assign n1782 = n2441 ^ n2442;
  assign n1962 = n2443 ^ n2444;
  assign n1575 = n2447 ^ n2448;
  assign n1965 = n2451 ^ n2452;
  assign n1792 = n2453 ^ n2454;
  assign n1385 = n2455 ^ n2456;
  assign n1439 = n2457 ^ n2458;
  assign n1486 = n2459 ^ n2460;
  assign n2326 = n2468 & n2469;
  assign n2149 = ~n2472;
  assign n1850 = n2474 ^ n2367;
  assign n1624 = n2475 ^ n2362;
  assign n2137 = n2476 ^ n2477;
  assign n2142 = n2478 ^ n2479;
  assign n2139 = n2496 & n2497;
  assign n2364 = n2475 & n2513;
  assign n2365 = n2474 & n2514;
  assign n2368 = n2160 & n2516;
  assign n2157 = n2521 ^ n2522;
  assign n2159 = n2196 ^ n2359;
  assign n2161 = n2523 ^ n2524;
  assign n2186 = n2525 ^ n2526;
  assign n1656 = n2527 ^ n2528;
  assign n2166 = n2529 ^ n2530;
  assign n1977 = n2531 ^ n2532;
  assign n1404 = n2533 ^ n2534;
  assign n2169 = n2535 ^ n2536;
  assign n2171 = n2537 ^ n2538;
  assign n2188 = n2539 ^ n2540;
  assign n2175 = n2541 ^ n2542;
  assign n2177 = n2543 ^ n2544;
  assign n2179 = n2545 ^ n2546;
  assign n2190 = n2547 ^ n2548;
  assign n2192 = n2549 ^ n2550;
  assign n2194 = n2551 ^ n2552;
  assign n2163 = n2553 ^ n2554;
  assign n2167 = n2555 ^ n2556;
  assign n2173 = n2557 ^ n2558;
  assign n2181 = n2559 ^ n2560;
  assign n2183 = n2561 ^ n2562;
  assign n1860 = ~n2580;
  assign n2047 = ~n2583;
  assign n1381 = ~n2586;
  assign n2231 = n2604 ^ n2605;
  assign n2250 = n2606 ^ n2607;
  assign n2252 = n2608 ^ n2609;
  assign n2235 = n2610 ^ n2611;
  assign n1902 = n2612 ^ n2613;
  assign n1528 = n2614 ^ n2615;
  assign n1658 = n2616 ^ n2617;
  assign n2256 = n2618 ^ n2619;
  assign n2258 = n2620 ^ n2621;
  assign n2260 = n2622 ^ n2623;
  assign n2013 = n2624 ^ n2625;
  assign n2294 = n2626 ^ n2627;
  assign n2247 = n2628 ^ n2629;
  assign n2058 = n2630 ^ n2631;
  assign n1919 = n2632 ^ n2633;
  assign n1343 = n2634 ^ n2635;
  assign n2060 = n2636 ^ n2637;
  assign n2229 = n2638 ^ n2639;
  assign n2062 = n2640 ^ n2641;
  assign n2233 = n2642 ^ n2643;
  assign n2254 = n2644 ^ n2645;
  assign n2237 = n2646 ^ n2647;
  assign n2239 = n2648 ^ n2649;
  assign n2056 = n2650 ^ n2651;
  assign n2241 = n2652 ^ n2653;
  assign n2243 = n2654 ^ n2655;
  assign n2245 = n2656 ^ n2657;
  assign n2463 = n2731 & n2732;
  assign n2473 = n2453 & n2454;
  assign n2140 = n2738 ^ n2739;
  assign n2515 = n2562 & n2757;
  assign n2517 = n2758 & n2759;
  assign n2518 = n2478 & n2479;
  assign n2519 = n2738 & n2739;
  assign n2564 = n2766 & n2767;
  assign n2361 = ~n2475;
  assign n2592 = n2527 & n2785;
  assign n2335 = ~n2786;
  assign n2593 = n2539 & n2789;
  assign n2594 = n2560 & n2790;
  assign n2595 = n2549 & n2791;
  assign n2596 = n2523 & n2794;
  assign n2597 = n2554 & n2164;
  assign n2354 = ~n2798;
  assign n2598 = n2535 & n2536;
  assign n2599 = n2799 & n2376;
  assign n2600 = n2558 & n2174;
  assign n2601 = n2541 & n2542;
  assign n2602 = n2189 & n2548;
  assign n2603 = n2551 & n2552;
  assign n1358 = ~n1341;
  assign n1764 = ~n1957;
  assign n2366 = ~n2474;
  assign n2358 = ~n2160;
  assign n1638 = ~n1744;
  assign n2712 = n2604 & n2801;
  assign n2713 = n2529 & n2802;
  assign n2714 = n2618 & n2803;
  assign n2715 = n2630 & n2804;
  assign n2716 = n2606 & n2805;
  assign n2717 = n2253 & n2645;
  assign n2718 = n2643 & n2642;
  assign n2719 = n2649 & n2648;
  assign n2720 = n2620 & n2621;
  assign n2721 = n2653 & n2652;
  assign n2722 = n2650 & n2651;
  assign n2723 = n2657 & n2656;
  assign n2726 = n2638 & n2806;
  assign n2751 = n2845 & n2846;
  assign n2729 = ~n2865;
  assign n2768 = n2896 & n2897;
  assign n2769 = n2898 & n2899;
  assign n2770 = n2900 & n2901;
  assign n2784 = n2918 & n2440;
  assign n2045 = ~n2920;
  assign n947 = ~n2932;
  assign n2488 = ~n2935;
  assign n2490 = ~n2936;
  assign n2381 = ~n2377;
  assign n2378 = n2949 & n2950;
  assign n2480 = ~n2451;
  assign n2265 = ~n2553;
  assign n2727 = ~n2555;
  assign n2566 = ~n2373;
  assign n2588 = ~n2539;
  assign n2730 = ~n2435;
  assign n2275 = ~n2557;
  assign n2304 = ~n2249;
  assign n2273 = ~n2559;
  assign n2464 = ~n2476;
  assign n2733 = ~n2545;
  assign n2735 = ~n2543;
  assign n2308 = ~n2057;
  assign n2328 = ~n2141;
  assign n2498 = ~n2521;
  assign n2347 = ~n2459;
  assign n2484 = ~n2525;
  assign n2350 = ~n2323;
  assign n2800 = n2953 & n2954;
  assign n2569 = ~n2955;
  assign n2706 = ~n2604;
  assign n2470 = ~n2453;
  assign n2482 = ~n2443;
  assign n2658 = ~n2253;
  assign n2502 = ~n2758;
  assign n2297 = ~n2644;
  assign n2587 = ~n2523;
  assign n2662 = ~n2643;
  assign n2660 = ~n2614;
  assign n2664 = ~n2649;
  assign n2666 = ~n2612;
  assign n2668 = ~n2616;
  assign n2670 = ~n2533;
  assign n2724 = n2962 & n2963;
  assign n2696 = ~n2620;
  assign n2337 = ~n2646;
  assign n2486 = ~n2537;
  assign n2672 = ~n2653;
  assign n2707 = ~n2618;
  assign n2375 = ~n2799;
  assign n2572 = ~n2535;
  assign n2708 = ~n2606;
  assign n2674 = ~n2622;
  assign n2589 = ~n2560;
  assign n2574 = ~n2558;
  assign n2489 = ~n2654;
  assign n2676 = ~n2651;
  assign n2677 = ~n2650;
  assign n2576 = ~n2541;
  assign n2578 = ~n2189;
  assign n2678 = ~n2657;
  assign n2277 = ~n2547;
  assign n2680 = ~n2632;
  assign n2682 = ~n2531;
  assign n2684 = ~n2624;
  assign n2807 = n2964 & n2965;
  assign n2510 = ~n2738;
  assign n2686 = ~n2626;
  assign n2808 = n2966 & n2967;
  assign n2590 = ~n2527;
  assign n2492 = ~n2628;
  assign n2591 = ~n2549;
  assign n2494 = ~n2457;
  assign n2709 = ~n2630;
  assign n2689 = ~n2640;
  assign n2690 = ~n2636;
  assign n2506 = ~n2478;
  assign n2512 = ~n2562;
  assign n2581 = ~n2551;
  assign n2584 = ~n2554;
  assign n2694 = ~n2634;
  assign n2692 = ~n2608;
  assign n2710 = ~n2529;
  assign n2500 = ~n2610;
  assign n2700 = ~n2638;
  assign n2809 = n2968 & n2969;
  assign n2810 = n2970 & n2971;
  assign n2811 = n2972 & n2973;
  assign n2812 = n2974 & n2975;
  assign n2813 = n2976 & n2977;
  assign n2814 = n2978 & n2979;
  assign n2815 = n2980 & n2981;
  assign n2816 = n2982 & n2983;
  assign n2817 = n2984 & n2985;
  assign n2704 = ~n2986;
  assign n2567 = ~n2987;
  assign n2565 = ~n2988;
  assign n2702 = ~n2989;
  assign n2675 = ~n2990;
  assign n2688 = ~n2991;
  assign n2698 = ~n2992;
  assign n2691 = ~n2993;
  assign n2693 = ~n2994;
  assign n2228 = n3009 & n3010;
  assign n2191 = n3049 & n3050;
  assign n2818 = n3172 & n3173;
  assign n1247 = ~n1214;
  assign n1573 = n2030 ^ n2031;
  assign n1840 = n2055 ^ n2056;
  assign n1822 = n2057 ^ n2058;
  assign n1718 = n2059 ^ n2060;
  assign n1835 = n2061 ^ n2062;
  assign n1061 = ~n1190;
  assign n1379 = n2137 ^ n2138;
  assign n1337 = n2139 ^ n2140;
  assign n1289 = n2141 ^ n2142;
  assign n1576 = n2149 & n2150;
  assign n1400 = n2157 ^ n2158;
  assign n1711 = n2159 ^ n2160;
  assign n1790 = n2161 ^ n2162;
  assign n1693 = n2163 ^ n2164;
  assign n1571 = n2165 ^ n2166;
  assign n1783 = n2167 ^ n2168;
  assign n1785 = n2169 ^ n2170;
  assign n1787 = n2171 ^ n2172;
  assign n1383 = n2173 ^ n2174;
  assign n1191 = n2175 ^ n2176;
  assign n1691 = n2177 ^ n2178;
  assign n1262 = n2179 ^ n2180;
  assign n1287 = n2181 ^ n2182;
  assign n1216 = n2183 ^ n2184;
  assign n1307 = n2185 ^ n2186;
  assign n1596 = ~n1306;
  assign n1695 = n2187 ^ n2188;
  assign n1446 = n2189 ^ n2190;
  assign n1449 = n2191 ^ n2192;
  assign n1304 = n2193 ^ n2194;
  assign n1828 = n2199 & n2200;
  assign n1529 = n2219 & n2220;
  assign n2053 = n2227 & n2228;
  assign n2054 = n2030 & n2031;
  assign n1825 = n2229 ^ n2230;
  assign n1975 = n2231 ^ n2232;
  assign n1622 = n2233 ^ n2234;
  assign n1620 = n2235 ^ n2236;
  assign n1445 = n2237 ^ n2238;
  assign n1310 = n2239 ^ n2240;
  assign n1312 = n2241 ^ n2242;
  assign n1844 = n2243 ^ n2244;
  assign n1846 = n2245 ^ n2246;
  assign n1821 = n2247 ^ n2248;
  assign n1816 = n2249 ^ n2250;
  assign n1818 = n2251 ^ n2252;
  assign n1714 = n2253 ^ n2254;
  assign n1784 = n2255 ^ n2256;
  assign n1786 = n2257 ^ n2258;
  assign n1788 = n2259 ^ n2260;
  assign n1628 = n1638 ^ n1425;
  assign n2041 = ~n2269;
  assign n2089 = n1528 & n1921;
  assign n2090 = n2294 & n2295;
  assign n2091 = n1343 & n1660;
  assign n2092 = n2229 & n2230;
  assign n2048 = ~n2227;
  assign n1490 = ~n1958;
  assign n2051 = ~n2030;
  assign n1477 = ~n1567;
  assign n1564 = ~n1443;
  assign n1798 = ~n1782;
  assign n1794 = ~n1962;
  assign n1600 = ~n1575;
  assign n1804 = ~n1965;
  assign n1602 = ~n1385;
  assign n1609 = ~n1439;
  assign n2026 = ~n2326;
  assign n2263 = n2335 & n2336;
  assign n2266 = n2337 & n2338;
  assign n2213 = ~n2139;
  assign n2280 = n2347 & n2348;
  assign n2283 = n2350 & n2351;
  assign n2284 = n2354 & n2355;
  assign n2289 = n2358 & n2359;
  assign n2292 = n2361 & n2362;
  assign n1640 = ~n2364;
  assign n1510 = ~n2365;
  assign n2293 = n2366 & n2367;
  assign n2195 = ~n2368;
  assign n2225 = ~n2166;
  assign n1883 = ~n1977;
  assign n2033 = n2375 ^ n2376;
  assign n2028 = n2377 ^ n2378;
  assign n2011 = ~n1902;
  assign n2084 = ~n1528;
  assign n1668 = ~n1658;
  assign n2015 = ~n2013;
  assign n2023 = ~n2294;
  assign n1762 = ~n1919;
  assign n2080 = ~n1343;
  assign n2082 = ~n2229;
  assign n2147 = ~n2463;
  assign n2325 = n2464 & n2465;
  assign n2331 = n2470 & n2471;
  assign n1858 = ~n2473;
  assign n2332 = n2480 & n2481;
  assign n2333 = n2482 & n2483;
  assign n2334 = n2484 & n2485;
  assign n2339 = n2486 & n2487;
  assign n2342 = n2488 & n2489;
  assign n2343 = n2490 & n2491;
  assign n2344 = n2492 & n2493;
  assign n2345 = n2494 & n2495;
  assign n2346 = n2498 & n2499;
  assign n2349 = n2500 & n2501;
  assign n2352 = n2502 & n2503;
  assign n2356 = n2506 & n2507;
  assign n2360 = n2510 & n2511;
  assign n2363 = n2512 & n2184;
  assign n2329 = ~n2515;
  assign n606 = ~n2517;
  assign n2327 = ~n2518;
  assign n2214 = ~n2519;
  assign n2038 = ~n2564;
  assign n2379 = n2565 & n2566;
  assign n2382 = n2567 & n2568;
  assign n2383 = n2569 & n2570;
  assign n2384 = n2375 & n2571;
  assign n2385 = n2572 & n2573;
  assign n2386 = n2574 & n2575;
  assign n2387 = n2576 & n2577;
  assign n2388 = n2578 & n2579;
  assign n2389 = n2581 & n2582;
  assign n2390 = n2584 & n2585;
  assign n2391 = n2587 & n2524;
  assign n2392 = n2588 & n2540;
  assign n2393 = n2589 & n2182;
  assign n2394 = n2590 & n2528;
  assign n2395 = n2591 & n2550;
  assign n1664 = ~n2592;
  assign n2270 = ~n2593;
  assign n2272 = ~n2594;
  assign n2278 = ~n2595;
  assign n2291 = ~n2596;
  assign n2264 = ~n2597;
  assign n2396 = n2378 & n2377;
  assign n2285 = ~n2598;
  assign n2267 = ~n2599;
  assign n2274 = ~n2600;
  assign n2287 = ~n2601;
  assign n2276 = ~n2602;
  assign n2281 = ~n2603;
  assign n2397 = n2658 & n2659;
  assign n2398 = n2660 & n2661;
  assign n2399 = n2662 & n2663;
  assign n2400 = n2664 & n2665;
  assign n2401 = n2666 & n2667;
  assign n2402 = n2668 & n2669;
  assign n2403 = n2670 & n2671;
  assign n2404 = n2672 & n2673;
  assign n2407 = n2674 & n2675;
  assign n2408 = n2676 & n2677;
  assign n2409 = n2678 & n2679;
  assign n2410 = n2680 & n2681;
  assign n2411 = n2682 & n2683;
  assign n2412 = n2684 & n2685;
  assign n2415 = n2686 & n2687;
  assign n2416 = n2688 & n2689;
  assign n2417 = n2690 & n2691;
  assign n2418 = n2692 & n2693;
  assign n2419 = n2694 & n2695;
  assign n2422 = n2696 & n2697;
  assign n2423 = n2698 & n2699;
  assign n2424 = n2700 & n2701;
  assign n2427 = n2702 & n2703;
  assign n2428 = n2704 & n2705;
  assign n2429 = n2706 & n2605;
  assign n2430 = n2707 & n2619;
  assign n2431 = n2708 & n2607;
  assign n2432 = n2709 & n2631;
  assign n2433 = n2710 & n2711;
  assign n2290 = ~n2712;
  assign n2315 = ~n2713;
  assign n2301 = ~n2714;
  assign n2307 = ~n2715;
  assign n2303 = ~n2716;
  assign n2296 = ~n2717;
  assign n2309 = ~n2718;
  assign n2313 = ~n2719;
  assign n2299 = ~n2720;
  assign n2311 = ~n2721;
  assign n2305 = ~n2722;
  assign n2317 = ~n2723;
  assign n2434 = n2724 & n2725;
  assign n2318 = ~n2726;
  assign n2461 = n2727 & n2728;
  assign n2462 = n2729 & n2730;
  assign n2466 = n2733 & n2734;
  assign n2467 = n2735 & n2736;
  assign n2146 = ~n2751;
  assign n768 = ~n2768;
  assign n2206 = ~n2769;
  assign n2208 = ~n2770;
  assign n2036 = ~n2784;
  assign n2380 = ~n2378;
  assign n2069 = ~n2800;
  assign n2425 = ~n2724;
  assign n2117 = ~n2807;
  assign n2413 = ~n2808;
  assign n2420 = ~n2809;
  assign n2064 = ~n2810;
  assign n2105 = ~n2811;
  assign n2124 = ~n2812;
  assign n2066 = ~n2813;
  assign n2121 = ~n2814;
  assign n2126 = ~n2815;
  assign n2128 = ~n2816;
  assign n2113 = ~n2817;
  assign n12379 = n2818 ^ n2819;
  assign n2049 = ~n2228;
  assign n2279 = ~n2191;
  assign n2764 = ~n2818;
  assign n998 = n1782 ^ n1783;
  assign n1145 = n1784 ^ n1785;
  assign n1291 = n1786 ^ n1787;
  assign n1551 = n1788 ^ n1789;
  assign n1451 = n1816 ^ n1817;
  assign n1220 = n1818 ^ n1819;
  assign n1461 = n1820 ^ n1821;
  assign n1387 = n1822 ^ n1823;
  assign n1095 = n1828 ^ n1829;
  assign n1457 = n1843 ^ n1844;
  assign n1781 = n1289 & n1958;
  assign n1808 = n1788 & n1960;
  assign n1811 = n1216 & n1963;
  assign n1812 = n1783 & n1782;
  assign n1813 = n1787 & n1786;
  assign n1815 = n1304 & n1966;
  assign n1887 = n1822 & n1971;
  assign n1890 = n1445 & n1972;
  assign n1896 = n1816 & n1817;
  assign n1899 = n1844 & n1843;
  assign n1873 = ~n1840;
  assign n1732 = ~n1718;
  assign n1881 = ~n1835;
  assign n1016 = ~n1379;
  assign n942 = n2022 ^ n2023;
  assign n1245 = ~n1337;
  assign n1780 = ~n1289;
  assign n1409 = ~n1576;
  assign n1491 = n2026 & n2027;
  assign n1516 = ~n1400;
  assign n1594 = ~n1711;
  assign n925 = n2028 ^ n2029;
  assign n967 = ~n1790;
  assign n1703 = ~n1693;
  assign n1606 = ~n1571;
  assign n1797 = ~n1783;
  assign n1805 = ~n1785;
  assign n1799 = ~n1787;
  assign n1598 = ~n1383;
  assign n999 = ~n1191;
  assign n1796 = ~n1691;
  assign n1275 = ~n1262;
  assign n1301 = ~n1287;
  assign n1801 = ~n1216;
  assign n940 = n2032 ^ n2033;
  assign n1809 = ~n1695;
  assign n1604 = ~n1446;
  assign n1475 = ~n1449;
  assign n1802 = ~n1304;
  assign n1855 = ~n1828;
  assign n1531 = n2041 & n2042;
  assign n1644 = ~n1529;
  assign n2007 = n2048 & n2049;
  assign n2010 = n2051 & n2052;
  assign n471 = ~n2053;
  assign n1634 = ~n2054;
  assign n1871 = ~n1975;
  assign n1646 = ~n1622;
  assign n1740 = ~n1620;
  assign n1893 = ~n1445;
  assign n1333 = ~n1310;
  assign n1335 = ~n1312;
  assign n1874 = ~n1844;
  assign n1891 = ~n1846;
  assign n1876 = ~n1821;
  assign n1884 = ~n1816;
  assign n1878 = ~n1818;
  assign n1725 = ~n1714;
  assign n1806 = ~n1784;
  assign n1800 = ~n1786;
  assign n1807 = ~n1788;
  assign n2016 = n2023 & n2079;
  assign n2017 = n2080 & n2081;
  assign n2018 = n2082 & n2083;
  assign n2019 = n2084 & n2085;
  assign n1537 = ~n2089;
  assign n2008 = ~n2090;
  assign n1666 = ~n2091;
  assign n1546 = ~n2092;
  assign n1550 = n2147 & n2148;
  assign n2034 = n2195 & n2196;
  assign n2043 = n2213 & n2214;
  assign n2050 = n2225 & n2226;
  assign n2035 = ~n2263;
  assign n2067 = n2264 & n2265;
  assign n2039 = ~n2266;
  assign n2070 = n2267 & n2268;
  assign n2071 = n2270 & n2271;
  assign n2072 = n2272 & n2273;
  assign n2073 = n2274 & n2275;
  assign n2074 = n2276 & n2277;
  assign n2075 = n2278 & n2279;
  assign n2044 = ~n2280;
  assign n2076 = n2281 & n2282;
  assign n2046 = ~n2283;
  assign n2037 = ~n2284;
  assign n2077 = n2285 & n2286;
  assign n2078 = n2287 & n2288;
  assign n1869 = ~n2289;
  assign n2086 = n2290 & n2232;
  assign n2087 = n2291 & n2162;
  assign n1353 = ~n2292;
  assign n1864 = ~n2293;
  assign n2093 = n2296 & n2297;
  assign n2102 = n2299 & n2300;
  assign n2103 = n2301 & n2302;
  assign n2106 = n2303 & n2304;
  assign n2107 = n2305 & n2306;
  assign n2122 = n2307 & n2308;
  assign n2131 = n2309 & n2310;
  assign n2132 = n2311 & n2312;
  assign n2133 = n2313 & n2314;
  assign n2134 = n2315 & n2316;
  assign n2135 = n2317 & n2246;
  assign n2136 = n2318 & n2319;
  assign n2024 = ~n2325;
  assign n2215 = n2327 & n2328;
  assign n2218 = n2329 & n2330;
  assign n1494 = ~n2331;
  assign n2223 = ~n2332;
  assign n2197 = ~n2333;
  assign n2201 = ~n2334;
  assign n2203 = ~n2339;
  assign n2205 = ~n2342;
  assign n2207 = ~n2343;
  assign n2209 = ~n2344;
  assign n2211 = ~n2345;
  assign n2216 = ~n2346;
  assign n2221 = ~n2349;
  assign n523 = ~n2352;
  assign n1968 = ~n2356;
  assign n1862 = ~n2360;
  assign n854 = n768 & n947;
  assign n1970 = ~n2363;
  assign n2065 = ~n2379;
  assign n2298 = n2380 & n2381;
  assign n2063 = ~n2382;
  assign n2068 = ~n2383;
  assign n1989 = ~n2384;
  assign n1991 = ~n2385;
  assign n1997 = ~n2386;
  assign n1999 = ~n2387;
  assign n2001 = ~n2388;
  assign n2006 = ~n2389;
  assign n1983 = ~n2390;
  assign n1987 = ~n2391;
  assign n1993 = ~n2392;
  assign n1995 = ~n2393;
  assign n1373 = ~n2394;
  assign n2003 = ~n2395;
  assign n2088 = ~n2396;
  assign n1925 = ~n2397;
  assign n2094 = ~n2398;
  assign n1927 = ~n2399;
  assign n1929 = ~n2400;
  assign n2096 = ~n2401;
  assign n2098 = ~n2402;
  assign n2100 = ~n2403;
  assign n1933 = ~n2404;
  assign n2104 = ~n2407;
  assign n1939 = ~n2408;
  assign n1941 = ~n2409;
  assign n2110 = ~n2410;
  assign n2108 = ~n2411;
  assign n2114 = ~n2412;
  assign n2012 = n2413 & n2414;
  assign n2118 = ~n2415;
  assign n2120 = ~n2416;
  assign n2125 = ~n2417;
  assign n2127 = ~n2418;
  assign n2129 = ~n2419;
  assign n1824 = n2420 & n2421;
  assign n1931 = ~n2422;
  assign n2123 = ~n2423;
  assign n1947 = ~n2424;
  assign n2322 = n2425 & n2426;
  assign n2116 = ~n2427;
  assign n2112 = ~n2428;
  assign n1981 = ~n2429;
  assign n1935 = ~n2430;
  assign n1937 = ~n2431;
  assign n1943 = ~n2432;
  assign n1945 = ~n2433;
  assign n70 = ~n2434;
  assign n2143 = ~n2461;
  assign n2145 = ~n2462;
  assign n2151 = ~n2466;
  assign n2153 = ~n2467;
  assign n2563 = n2764 & n2765;
  assign n732 = n1550 ^ n1551;
  assign n1243 = ~n1220;
  assign n1471 = ~n1461;
  assign n1473 = ~n1387;
  assign n1183 = ~n1095;
  assign n1689 = n1780 & n1490;
  assign n1679 = ~n1781;
  assign n1698 = n1797 & n1798;
  assign n1699 = n1799 & n1800;
  assign n1700 = n1801 & n1533;
  assign n1701 = n1802 & n1618;
  assign n1706 = n1805 & n1784;
  assign n1707 = n1785 & n1806;
  assign n1708 = n1807 & n1789;
  assign n1560 = ~n1808;
  assign n1295 = ~n1811;
  assign n965 = ~n1812;
  assign n1241 = ~n1813;
  assign n1563 = ~n1815;
  assign n1569 = n1824 ^ n1825;
  assign n1719 = n1855 & n1856;
  assign n1727 = n1874 & n1875;
  assign n1728 = n1876 & n1877;
  assign n1729 = n1878 & n1879;
  assign n1734 = n1884 & n1885;
  assign n1589 = ~n1887;
  assign n1232 = ~n1890;
  assign n1741 = n1893 & n1842;
  assign n1224 = ~n1896;
  assign n1586 = ~n1899;
  assign n1588 = ~n1491;
  assign n944 = ~n925;
  assign n1636 = ~n1531;
  assign n437 = ~n2007;
  assign n1915 = n2008 & n2009;
  assign n1349 = ~n2010;
  assign n1690 = n2012 ^ n2013;
  assign n1642 = ~n2016;
  assign n1375 = ~n2017;
  assign n1914 = ~n2018;
  assign n1907 = ~n2019;
  assign n1561 = ~n1550;
  assign n1694 = n2024 & n2025;
  assign n1868 = ~n2034;
  assign n1713 = n2035 & n2036;
  assign n1692 = n2037 & n2038;
  assign n1715 = n2039 & n2040;
  assign n1861 = ~n2043;
  assign n2004 = n2044 & n2045;
  assign n1717 = n2046 & n2047;
  assign n1859 = ~n2050;
  assign n1961 = n2063 & n2064;
  assign n1791 = n2065 & n2066;
  assign n1982 = ~n2067;
  assign n1901 = n2068 & n2069;
  assign n1988 = ~n2070;
  assign n1992 = ~n2071;
  assign n1994 = ~n2072;
  assign n1996 = ~n2073;
  assign n2000 = ~n2074;
  assign n2002 = ~n2075;
  assign n2005 = ~n2076;
  assign n1990 = ~n2077;
  assign n1998 = ~n2078;
  assign n1980 = ~n2086;
  assign n1986 = ~n2087;
  assign n2020 = n2088 & n2029;
  assign n2021 = n2012 & n2013;
  assign n1924 = ~n2093;
  assign n1837 = n2094 & n2095;
  assign n1830 = n2096 & n2097;
  assign n1832 = n2098 & n2099;
  assign n1920 = n2100 & n2101;
  assign n1930 = ~n2102;
  assign n1934 = ~n2103;
  assign n1922 = n2104 & n2105;
  assign n1936 = ~n2106;
  assign n1938 = ~n2107;
  assign n1956 = n2108 & n2109;
  assign n1751 = n2110 & n2111;
  assign n1189 = n2112 & n2113;
  assign n1845 = n2114 & n2115;
  assign n1953 = n2116 & n2117;
  assign n1851 = n2118 & n2119;
  assign n1918 = n2120 & n2121;
  assign n1942 = ~n2122;
  assign n1565 = n2123 & n2124;
  assign n1854 = n2125 & n2126;
  assign n1826 = n2127 & n2128;
  assign n1753 = n2129 & n2130;
  assign n1926 = ~n2131;
  assign n1932 = ~n2132;
  assign n1928 = ~n2133;
  assign n1944 = ~n2134;
  assign n1940 = ~n2135;
  assign n1946 = ~n2136;
  assign n1487 = n2143 & n2144;
  assign n1964 = n2145 & n2146;
  assign n1578 = n2151 & n2152;
  assign n1458 = n2153 & n2154;
  assign n1974 = n2197 & n2198;
  assign n1629 = n2201 & n2202;
  assign n1836 = n2203 & n2204;
  assign n1841 = n2205 & n2206;
  assign n1839 = n2207 & n2208;
  assign n1849 = n2209 & n2210;
  assign n1847 = n2211 & n2212;
  assign n1967 = ~n2215;
  assign n1853 = n2216 & n2217;
  assign n1969 = ~n2218;
  assign n1834 = n2221 & n2222;
  assign n1976 = n2223 & n2224;
  assign n588 = n523 & n606;
  assign n1909 = ~n2298;
  assign n2014 = ~n2012;
  assign n1913 = ~n1824;
  assign n67 = ~n2322;
  assign n2261 = ~n2563;
  assign n1256 = ~n732;
  assign n1464 = n1560 & n1561;
  assign n1482 = n1565 & n1387;
  assign n1267 = n1589 & n1590;
  assign n1377 = ~n1689;
  assign n1048 = n1690 ^ n1691;
  assign n1293 = n1692 ^ n1693;
  assign n1147 = n1694 ^ n1695;
  assign n829 = ~n1698;
  assign n1074 = ~n1699;
  assign n1463 = ~n1700;
  assign n1395 = ~n1701;
  assign n956 = ~n1706;
  assign n1103 = ~n1707;
  assign n1389 = ~n1708;
  assign n1469 = ~n1569;
  assign n1402 = n1713 ^ n1714;
  assign n1403 = n1715 ^ n1716;
  assign n1399 = n1717 ^ n1718;
  assign n1499 = ~n1719;
  assign n1322 = ~n1727;
  assign n1511 = ~n1728;
  assign n1495 = ~n1729;
  assign n1498 = ~n1734;
  assign n1649 = n437 & n471;
  assign n1503 = ~n1741;
  assign n1492 = n1751 ^ n1752;
  assign n1485 = n1753 ^ n1754;
  assign n1141 = n1189 ^ n1790;
  assign n1167 = n1791 ^ n1792;
  assign n1709 = n1694 & n1809;
  assign n1712 = n1692 & n1693;
  assign n1218 = n1826 ^ n1827;
  assign n996 = n1830 ^ n1831;
  assign n1442 = n1832 ^ n1833;
  assign n1440 = n1834 ^ n1835;
  assign n1453 = n1836 ^ n1672;
  assign n1023 = n1837 ^ n1838;
  assign n1455 = n1839 ^ n1840;
  assign n1444 = n1841 ^ n1842;
  assign n1459 = n1845 ^ n1846;
  assign n1447 = n1847 ^ n1848;
  assign n1448 = n1849 ^ n1850;
  assign n1043 = n1851 ^ n1852;
  assign n1438 = n1853 ^ n1854;
  assign n1142 = n1859 & n1860;
  assign n1566 = n1861 & n1862;
  assign n1568 = n1868 & n1869;
  assign n1738 = n1715 & n1889;
  assign n1739 = n1845 & n1891;
  assign n1742 = n1717 & n1718;
  assign n1743 = n1713 & n1714;
  assign n1488 = n1901 ^ n1902;
  assign n1748 = n1913 & n1914;
  assign n1641 = ~n1915;
  assign n1530 = n1918 ^ n1919;
  assign n1527 = n1920 ^ n1921;
  assign n1532 = n1922 ^ n1923;
  assign n1621 = n1924 & n1925;
  assign n1630 = n1926 & n1927;
  assign n1570 = n1928 & n1929;
  assign n1452 = n1930 & n1931;
  assign n1625 = n1932 & n1933;
  assign n1657 = n1934 & n1935;
  assign n1572 = n1936 & n1937;
  assign n1577 = n1938 & n1939;
  assign n1579 = n1940 & n1941;
  assign n1460 = n1942 & n1943;
  assign n1655 = n1944 & n1945;
  assign n1659 = n1946 & n1947;
  assign n1771 = n1837 & n1949;
  assign n1772 = n1753 & n1950;
  assign n1773 = n1751 & n1951;
  assign n1774 = n1830 & n1952;
  assign n1775 = n1922 & n1923;
  assign n1776 = n1953 & n1954;
  assign n1777 = n1851 & n1955;
  assign n1778 = n1918 & n1919;
  assign n1779 = n1956 & n1957;
  assign n1810 = n1961 & n1962;
  assign n1814 = n1964 & n1965;
  assign n1705 = ~n1694;
  assign n1580 = n1967 & n1968;
  assign n1867 = n1969 & n1970;
  assign n1892 = n1847 & n1973;
  assign n1894 = n1834 & n1835;
  assign n1895 = n1974 & n1975;
  assign n1897 = n1976 & n1977;
  assign n1898 = n1839 & n1840;
  assign n1900 = n1854 & n1853;
  assign n1710 = n1980 & n1981;
  assign n1619 = n1982 & n1983;
  assign n1450 = n1986 & n1987;
  assign n1724 = ~n1713;
  assign n1702 = ~n1692;
  assign n1735 = ~n1715;
  assign n1574 = n1988 & n1989;
  assign n1344 = n1990 & n1991;
  assign n1088 = n1992 & n1993;
  assign n1627 = n1994 & n1995;
  assign n1623 = n1996 & n1997;
  assign n1454 = n1998 & n1999;
  assign n1456 = n2000 & n2001;
  assign n1222 = n2002 & n2003;
  assign n1562 = ~n2004;
  assign n1912 = n2005 & n2006;
  assign n1731 = ~n1717;
  assign n1917 = n1901 & n2011;
  assign n1793 = ~n1961;
  assign n1857 = ~n1791;
  assign n1916 = ~n1901;
  assign n1948 = n2014 & n2015;
  assign n1908 = ~n2020;
  assign n1795 = ~n2021;
  assign n1767 = ~n1837;
  assign n1757 = ~n1830;
  assign n1904 = ~n1832;
  assign n1906 = ~n1920;
  assign n1759 = ~n1922;
  assign n1763 = ~n1956;
  assign n1770 = ~n1751;
  assign n1112 = ~n1189;
  assign n1886 = ~n1845;
  assign n1765 = ~n1953;
  assign n1755 = ~n1851;
  assign n1761 = ~n1918;
  assign n1472 = ~n1565;
  assign n1865 = ~n1854;
  assign n1910 = ~n1826;
  assign n1769 = ~n1753;
  assign n1959 = n67 & n70;
  assign n1582 = ~n1487;
  assign n1803 = ~n1964;
  assign n1411 = ~n1578;
  assign n1507 = ~n1458;
  assign n1870 = ~n1974;
  assign n1407 = ~n1629;
  assign n1431 = ~n1836;
  assign n1502 = ~n1841;
  assign n1872 = ~n1839;
  assign n1863 = ~n1849;
  assign n1888 = ~n1847;
  assign n1866 = ~n1853;
  assign n1880 = ~n1834;
  assign n1882 = ~n1976;
  assign n1978 = n2261 & n2262;
  assign n837 = n1399 ^ n1400;
  assign n883 = n1401 ^ n1402;
  assign n857 = n1403 ^ n1404;
  assign n1398 = n1048 & n1222;
  assign n701 = n1438 ^ n1439;
  assign n1264 = n1440 ^ n1441;
  assign n1259 = n1442 ^ n1443;
  assign n914 = n1444 ^ n1445;
  assign n1125 = n1446 ^ n1447;
  assign n1266 = n1448 ^ n1449;
  assign n722 = n1450 ^ n1451;
  assign n911 = n1452 ^ n1453;
  assign n783 = n1454 ^ n1455;
  assign n871 = n1456 ^ n1457;
  assign n1261 = n1458 ^ n1459;
  assign n1268 = n1460 ^ n1461;
  assign n1388 = ~n1464;
  assign n1414 = n1472 & n1473;
  assign n1392 = ~n1482;
  assign n1169 = n1485 ^ n1486;
  assign n1260 = n1487 ^ n1488;
  assign n1286 = n1491 ^ n1492;
  assign n1217 = n1495 & n1496;
  assign n1219 = n1499 & n1500;
  assign n1421 = n1502 & n1503;
  assign n1265 = n1511 & n1512;
  assign n1391 = ~n1267;
  assign n853 = n1527 ^ n1528;
  assign n1213 = n1529 ^ n1530;
  assign n1290 = n1531 ^ n1532;
  assign n1467 = n1562 & n1563;
  assign n1478 = n1442 & n1564;
  assign n1480 = n1448 & n1449;
  assign n1481 = n1460 & n1461;
  assign n1483 = n1566 & n1567;
  assign n1484 = n1568 & n1569;
  assign n1437 = ~n1048;
  assign n1139 = n1570 ^ n1571;
  assign n1164 = n1572 ^ n1573;
  assign n1063 = n1574 ^ n1575;
  assign n1382 = n1576 ^ n1577;
  assign n1384 = n1578 ^ n1579;
  assign n1386 = n1580 ^ n1565;
  assign n1303 = n1562 ^ n1618;
  assign n1093 = n1619 ^ n1620;
  assign n1308 = n1621 ^ n1622;
  assign n1361 = n1623 ^ n1624;
  assign n1309 = n1625 ^ n1626;
  assign n1311 = n1627 ^ n1628;
  assign n1305 = n1629 ^ n1630;
  assign n1281 = n1641 & n1642;
  assign n473 = ~n1649;
  assign n1340 = n1655 ^ n1656;
  assign n1345 = n1657 ^ n1658;
  assign n1342 = n1659 ^ n1660;
  assign n1162 = ~n1167;
  assign n1607 = n1702 & n1703;
  assign n1611 = n1705 & n1695;
  assign n1152 = ~n1709;
  assign n1612 = n1710 & n1711;
  assign n1613 = n1630 & n1306;
  assign n1228 = ~n1712;
  assign n1614 = n1570 & n1571;
  assign n1615 = n1574 & n1575;
  assign n1616 = n1577 & n1383;
  assign n1617 = n1579 & n1385;
  assign n1239 = ~n1218;
  assign n1479 = ~n1442;
  assign n1041 = ~n1023;
  assign n1474 = ~n1448;
  assign n1099 = ~n1142;
  assign n1476 = ~n1566;
  assign n1468 = ~n1568;
  assign n1647 = n1724 & n1725;
  assign n1648 = n1731 & n1732;
  assign n1651 = n1735 & n1716;
  assign n1526 = ~n1738;
  assign n1506 = ~n1739;
  assign n1652 = n1619 & n1740;
  assign n1515 = ~n1742;
  assign n1653 = n1621 & n1622;
  assign n1525 = ~n1743;
  assign n1654 = n1627 & n1744;
  assign n1545 = ~n1748;
  assign n1677 = n1452 & n1750;
  assign n1678 = n1657 & n1658;
  assign n1645 = ~n1621;
  assign n1595 = ~n1630;
  assign n1605 = ~n1570;
  assign n1671 = ~n1452;
  assign n1661 = ~n1625;
  assign n1667 = ~n1657;
  assign n1633 = ~n1572;
  assign n1597 = ~n1577;
  assign n1601 = ~n1579;
  assign n1680 = n1755 & n1756;
  assign n1470 = ~n1460;
  assign n1663 = ~n1655;
  assign n1665 = ~n1659;
  assign n1681 = n1757 & n1758;
  assign n1682 = n1759 & n1760;
  assign n1683 = n1761 & n1762;
  assign n1684 = n1763 & n1764;
  assign n1685 = n1765 & n1766;
  assign n1686 = n1767 & n1768;
  assign n1687 = n1769 & n1754;
  assign n1688 = n1770 & n1752;
  assign n1673 = ~n1771;
  assign n1610 = ~n1772;
  assign n1587 = ~n1773;
  assign n1669 = ~n1774;
  assign n1635 = ~n1775;
  assign n79 = ~n1776;
  assign n1675 = ~n1777;
  assign n1643 = ~n1778;
  assign n84 = ~n1779;
  assign n1696 = n1793 & n1794;
  assign n1697 = n1795 & n1796;
  assign n1704 = n1803 & n1804;
  assign n427 = ~n1810;
  assign n98 = ~n1814;
  assign n1720 = n1857 & n1858;
  assign n1721 = n1863 & n1864;
  assign n1722 = n1865 & n1866;
  assign n1393 = ~n1580;
  assign n1489 = ~n1867;
  assign n1723 = n1870 & n1871;
  assign n1726 = n1872 & n1873;
  assign n1730 = n1880 & n1881;
  assign n1733 = n1882 & n1883;
  assign n1736 = n1886 & n1846;
  assign n1737 = n1888 & n1848;
  assign n1603 = ~n1892;
  assign n1591 = ~n1894;
  assign n421 = ~n1895;
  assign n91 = ~n1897;
  assign n1583 = ~n1898;
  assign n1608 = ~n1900;
  assign n1593 = ~n1710;
  assign n1650 = ~n1619;
  assign n1497 = ~n1450;
  assign n1745 = n1904 & n1905;
  assign n1746 = n1906 & n1907;
  assign n1263 = n1908 & n1909;
  assign n1599 = ~n1574;
  assign n1433 = ~n1344;
  assign n1072 = ~n1088;
  assign n1637 = ~n1627;
  assign n1639 = ~n1623;
  assign n1584 = ~n1454;
  assign n1585 = ~n1456;
  assign n1436 = ~n1222;
  assign n1747 = n1910 & n1911;
  assign n1462 = ~n1912;
  assign n1749 = n1916 & n1902;
  assign n1581 = ~n1917;
  assign n1466 = ~n1948;
  assign n72 = ~n1959;
  assign n12380 = n1978 ^ n1979;
  assign n1984 = ~n1978;
  assign n1051 = n1213 ^ n1214;
  assign n984 = n1217 ^ n1218;
  assign n982 = n1219 ^ n1220;
  assign n575 = n1259 ^ n1260;
  assign n1014 = n1261 ^ n1262;
  assign n736 = n1263 ^ n1264;
  assign n972 = n1265 ^ n1266;
  assign n969 = n1267 ^ n1268;
  assign n1025 = n1286 ^ n1287;
  assign n885 = n1290 ^ n1291;
  assign n1212 = n1286 & n1287;
  assign n1201 = n1303 ^ n1304;
  assign n790 = ~n837;
  assign n835 = n1305 ^ n1306;
  assign n781 = n1307 ^ n1308;
  assign n980 = ~n883;
  assign n988 = n1309 ^ n1310;
  assign n862 = ~n857;
  assign n1127 = n1311 ^ n1312;
  assign n1124 = n1281 ^ n1043;
  assign n1251 = n1213 & n1214;
  assign n1253 = n1217 & n1218;
  assign n1254 = n1219 & n1220;
  assign n1143 = n1340 ^ n1341;
  assign n1170 = n1342 ^ n1343;
  assign n797 = n1344 ^ n1345;
  assign n1258 = n1361 & n732;
  assign n1283 = n1264 & n1263;
  assign n1284 = n783 & n990;
  assign n1282 = n1261 & n1262;
  assign n1285 = n871 & n1379;
  assign n851 = n1382 ^ n1383;
  assign n800 = n1384 ^ n1385;
  assign n1193 = n1386 ^ n1387;
  assign n1128 = n1388 & n1389;
  assign n1299 = n1392 & n1393;
  assign n1271 = ~n1398;
  assign n642 = ~n701;
  assign n1278 = ~n1264;
  assign n919 = ~n914;
  assign n1280 = ~n1125;
  assign n670 = ~n722;
  assign n917 = ~n911;
  assign n1272 = ~n783;
  assign n1276 = ~n871;
  assign n1274 = ~n1261;
  assign n1134 = ~n1414;
  assign n1338 = n1309 & n1310;
  assign n1339 = n1311 & n1312;
  assign n1160 = ~n1169;
  assign n1300 = ~n1286;
  assign n1238 = ~n1217;
  assign n1242 = ~n1219;
  assign n1231 = ~n1421;
  assign n1297 = ~n1265;
  assign n1360 = n1340 & n1341;
  assign n864 = ~n853;
  assign n1246 = ~n1213;
  assign n1240 = ~n1290;
  assign n1396 = n1436 & n1437;
  assign n1405 = n1462 & n1463;
  assign n1394 = ~n1467;
  assign n1412 = n1468 & n1469;
  assign n1413 = n1470 & n1471;
  assign n1415 = n1474 & n1475;
  assign n1416 = n1476 & n1477;
  assign n1397 = ~n1478;
  assign n1418 = n1479 & n1443;
  assign n1057 = ~n1480;
  assign n1390 = ~n1481;
  assign n105 = ~n1483;
  assign n406 = ~n1484;
  assign n1083 = ~n1164;
  assign n1065 = n1072 ^ n940;
  assign n1288 = n1489 ^ n1490;
  assign n1420 = n1497 & n1498;
  assign n1422 = n1506 & n1507;
  assign n1423 = n1515 & n1516;
  assign n1427 = n1525 & n1401;
  assign n1428 = n1526 & n1404;
  assign n929 = ~n1361;
  assign n1332 = ~n1309;
  assign n1334 = ~n1311;
  assign n1215 = n1462 ^ n1533;
  assign n1378 = ~n1281;
  assign n1171 = n1545 & n1546;
  assign n1357 = ~n1340;
  assign n1501 = n1581 & n1582;
  assign n1504 = n1583 & n1584;
  assign n1505 = n1585 & n1586;
  assign n1508 = n1587 & n1588;
  assign n1513 = n1591 & n1592;
  assign n1514 = n1593 & n1594;
  assign n1517 = n1595 & n1596;
  assign n1518 = n1597 & n1598;
  assign n1519 = n1599 & n1600;
  assign n1520 = n1601 & n1602;
  assign n1521 = n1603 & n1604;
  assign n1522 = n1605 & n1606;
  assign n1069 = ~n1607;
  assign n1523 = n1608 & n1609;
  assign n1524 = n1610 & n1486;
  assign n936 = ~n1611;
  assign n415 = ~n1612;
  assign n1406 = ~n1613;
  assign n1101 = ~n1614;
  assign n1076 = ~n1615;
  assign n1408 = ~n1616;
  assign n1410 = ~n1617;
  assign n1538 = n1633 & n1634;
  assign n1539 = n1635 & n1636;
  assign n1540 = n1637 & n1638;
  assign n1541 = n1639 & n1640;
  assign n1542 = n1643 & n1644;
  assign n1547 = n1645 & n1646;
  assign n1226 = ~n1647;
  assign n1237 = ~n1648;
  assign n1548 = n1650 & n1620;
  assign n1230 = ~n1651;
  assign n1109 = ~n1652;
  assign n1426 = ~n1653;
  assign n1424 = ~n1654;
  assign n1549 = n1661 & n1662;
  assign n1552 = n1663 & n1664;
  assign n1553 = n1665 & n1666;
  assign n1554 = n1667 & n1668;
  assign n1555 = n1669 & n1670;
  assign n1556 = n1671 & n1672;
  assign n1557 = n1673 & n1674;
  assign n1558 = n1675 & n1676;
  assign n1430 = ~n1677;
  assign n1432 = ~n1678;
  assign n1559 = n1489 & n1679;
  assign n1371 = ~n1680;
  assign n1365 = ~n1681;
  assign n1351 = ~n1682;
  assign n1355 = ~n1683;
  assign n81 = ~n1684;
  assign n74 = ~n1685;
  assign n1363 = ~n1686;
  assign n1314 = ~n1687;
  assign n1324 = ~n1688;
  assign n424 = ~n1696;
  assign n1465 = ~n1697;
  assign n95 = ~n1704;
  assign n1493 = ~n1720;
  assign n1509 = ~n1721;
  assign n1329 = ~n1722;
  assign n417 = ~n1723;
  assign n1320 = ~n1726;
  assign n1331 = ~n1730;
  assign n88 = ~n1733;
  assign n1235 = ~n1736;
  assign n1327 = ~n1737;
  assign n1534 = ~n1745;
  assign n1536 = ~n1746;
  assign n1277 = ~n1263;
  assign n1543 = ~n1747;
  assign n1317 = ~n1749;
  assign n1903 = n1984 & n1985;
  assign n887 = n1124 ^ n1125;
  assign n813 = n1142 ^ n1143;
  assign n1091 = n1170 & n1171;
  assign n1121 = n851 & n1190;
  assign n1122 = n800 & n1191;
  assign n963 = ~n575;
  assign n897 = ~n972;
  assign n899 = ~n969;
  assign n1037 = ~n885;
  assign n859 = ~n1212;
  assign n1136 = ~n1201;
  assign n788 = ~n835;
  assign n746 = ~n781;
  assign n1105 = n1215 ^ n1216;
  assign n1064 = n1231 & n1232;
  assign n1178 = n1238 & n1239;
  assign n1179 = n1240 & n1241;
  assign n1180 = n1242 & n1243;
  assign n1182 = n1246 & n1247;
  assign n1156 = ~n1251;
  assign n992 = ~n1253;
  assign n1002 = ~n1254;
  assign n1158 = ~n1170;
  assign n806 = ~n797;
  assign n1188 = n929 & n1256;
  assign n823 = ~n1258;
  assign n1195 = n1272 & n1273;
  assign n1196 = n1274 & n1275;
  assign n1197 = n1276 & n1016;
  assign n1198 = n1277 & n1278;
  assign n1199 = n1280 & n1281;
  assign n841 = ~n1282;
  assign n753 = ~n1283;
  assign n974 = ~n1284;
  assign n1110 = ~n1285;
  assign n1119 = n1288 ^ n1289;
  assign n1115 = ~n851;
  assign n1116 = ~n800;
  assign n1114 = ~n1193;
  assign n889 = ~n1128;
  assign n1133 = ~n1299;
  assign n1209 = n1300 & n1301;
  assign n1248 = n1332 & n1333;
  assign n1249 = n1334 & n1335;
  assign n1004 = ~n1338;
  assign n1154 = ~n1339;
  assign n1257 = n1357 & n1358;
  assign n950 = ~n1360;
  assign n1279 = n1378 & n1125;
  assign n1298 = n1390 & n1391;
  assign n1104 = n1394 & n1395;
  assign n1031 = ~n1396;
  assign n1302 = n1397 & n1260;
  assign n1294 = ~n1405;
  assign n1315 = n1406 & n1407;
  assign n1318 = n1408 & n1409;
  assign n1325 = n1410 & n1411;
  assign n403 = ~n1412;
  assign n1132 = ~n1413;
  assign n1296 = ~n1415;
  assign n102 = ~n1416;
  assign n1130 = ~n1418;
  assign n1223 = ~n1420;
  assign n1234 = ~n1422;
  assign n1236 = ~n1423;
  assign n1356 = n1424 & n1425;
  assign n1359 = n1426 & n1307;
  assign n1225 = ~n1427;
  assign n1229 = ~n1428;
  assign n1368 = n1430 & n1431;
  assign n1369 = n1432 & n1433;
  assign n1157 = ~n1171;
  assign n1013 = n1465 & n1466;
  assign n1417 = n424 & n427;
  assign n1419 = n95 & n98;
  assign n1336 = n1493 & n1494;
  assign n1316 = ~n1501;
  assign n1319 = ~n1504;
  assign n1321 = ~n1505;
  assign n1323 = ~n1508;
  assign n1221 = n1509 & n1510;
  assign n1330 = ~n1513;
  assign n410 = ~n1514;
  assign n1203 = ~n1517;
  assign n1205 = ~n1518;
  assign n876 = ~n1519;
  assign n1207 = ~n1520;
  assign n1326 = ~n1521;
  assign n954 = ~n1522;
  assign n1328 = ~n1523;
  assign n418 = n417 & n421;
  assign n1313 = ~n1524;
  assign n1429 = n88 & n91;
  assign n1165 = n1534 & n1535;
  assign n1292 = n1536 & n1537;
  assign n1348 = ~n1538;
  assign n1350 = ~n1539;
  assign n1176 = ~n1540;
  assign n1352 = ~n1541;
  assign n1354 = ~n1542;
  assign n1089 = n1543 & n1544;
  assign n1173 = ~n1547;
  assign n902 = ~n1548;
  assign n1366 = ~n1549;
  assign n1372 = ~n1552;
  assign n1374 = ~n1553;
  assign n1187 = ~n1554;
  assign n1364 = ~n1555;
  assign n1185 = ~n1556;
  assign n1362 = ~n1557;
  assign n1370 = ~n1558;
  assign n1434 = n74 & n79;
  assign n1435 = n81 & n84;
  assign n1376 = ~n1559;
  assign n1631 = ~n1903;
  assign n932 = n1013 ^ n1014;
  assign n904 = ~n887;
  assign n764 = ~n813;
  assign n856 = n1064 ^ n1065;
  assign n1011 = n1064 & n1088;
  assign n399 = ~n1091;
  assign n1049 = n1104 & n1105;
  assign n1038 = n1115 & n1061;
  assign n1039 = n1116 & n999;
  assign n959 = ~n1121;
  assign n961 = ~n1122;
  assign n968 = n1133 & n1134;
  assign n1080 = n1157 & n1158;
  assign n1060 = ~n1105;
  assign n1071 = ~n1064;
  assign n802 = ~n1178;
  assign n1073 = ~n1179;
  assign n816 = ~n1180;
  assign n938 = ~n1182;
  assign n957 = ~n1188;
  assign n785 = ~n1195;
  assign n1029 = ~n1196;
  assign n894 = ~n1197;
  assign n600 = ~n1198;
  assign n1042 = ~n1199;
  assign n1035 = ~n1119;
  assign n1055 = ~n1209;
  assign n1053 = n1165 ^ n996;
  assign n1047 = n1221 ^ n1222;
  assign n1163 = n1223 & n1224;
  assign n926 = n1225 & n1226;
  assign n1062 = n1229 & n1230;
  assign n1177 = n1234 & n1235;
  assign n985 = n1236 & n1237;
  assign n818 = ~n1248;
  assign n934 = ~n1249;
  assign n1098 = ~n1257;
  assign n843 = ~n1279;
  assign n1022 = n1292 ^ n1293;
  assign n1118 = n1294 & n1295;
  assign n1208 = n1296 & n1297;
  assign n1131 = ~n1298;
  assign n1059 = ~n1104;
  assign n1210 = n403 & n406;
  assign n1129 = ~n1302;
  assign n1211 = n102 & n105;
  assign n1200 = n1313 & n1314;
  assign n1202 = ~n1315;
  assign n1052 = n1316 & n1317;
  assign n1204 = ~n1318;
  assign n1233 = n1319 & n1320;
  assign n1146 = n1321 & n1322;
  assign n1126 = n1323 & n1324;
  assign n1206 = ~n1325;
  assign n687 = n1326 & n1327;
  assign n886 = n1328 & n1329;
  assign n1050 = n1330 & n1331;
  assign n1250 = n410 & n415;
  assign n1252 = n1336 & n1337;
  assign n1166 = n1348 & n1349;
  assign n1144 = n1350 & n1351;
  assign n1120 = n1352 & n1353;
  assign n1024 = n1354 & n1355;
  assign n1175 = ~n1356;
  assign n1172 = ~n1359;
  assign n1092 = n1362 & n1363;
  assign n1094 = n1364 & n1365;
  assign n1138 = n1366 & n1367;
  assign n1184 = ~n1368;
  assign n1186 = ~n1369;
  assign n1269 = n1370 & n1371;
  assign n1140 = n1372 & n1373;
  assign n1168 = n1374 & n1375;
  assign n1192 = n1376 & n1377;
  assign n1028 = ~n1013;
  assign n429 = ~n1417;
  assign n100 = ~n1419;
  assign n1244 = ~n1336;
  assign n1270 = ~n1221;
  assign n93 = ~n1429;
  assign n1149 = ~n1165;
  assign n1227 = ~n1292;
  assign n1067 = ~n1089;
  assign n77 = ~n1434;
  assign n86 = ~n1435;
  assign n1380 = n1631 & n1632;
  assign n720 = n856 ^ n857;
  assign n612 = n886 ^ n887;
  assign n868 = n856 & n857;
  assign n873 = ~n932;
  assign n908 = n968 & n969;
  assign n910 = n886 & n887;
  assign n861 = ~n856;
  assign n939 = ~n1011;
  assign n718 = n1022 ^ n1023;
  assign n833 = n1024 ^ n1025;
  assign n975 = n1028 & n1029;
  assign n825 = ~n1038;
  assign n827 = ~n1039;
  assign n979 = n1042 & n1043;
  assign n906 = n1047 ^ n1048;
  assign n379 = ~n1049;
  assign n573 = n1050 ^ n1051;
  assign n792 = n1052 ^ n1053;
  assign n898 = ~n968;
  assign n994 = n1059 & n1060;
  assign n852 = n1062 ^ n1063;
  assign n1007 = n1071 & n1072;
  assign n769 = n1073 & n1074;
  assign n396 = ~n1080;
  assign n1012 = n985 & n1089;
  assign n924 = n1092 ^ n1093;
  assign n927 = n1094 ^ n1095;
  assign n1018 = n1098 & n1099;
  assign n1044 = n1118 & n1119;
  assign n1045 = n1022 & n1023;
  assign n1046 = n1120 & n885;
  assign n751 = n1126 ^ n1127;
  assign n884 = n1128 ^ n1120;
  assign n708 = n1129 & n1130;
  assign n971 = n1131 & n1132;
  assign n711 = n1138 ^ n1139;
  assign n810 = n1140 ^ n1141;
  assign n912 = n1144 ^ n1145;
  assign n913 = n1146 ^ n1147;
  assign n1085 = n1163 & n1164;
  assign n1086 = n1052 & n1165;
  assign n1087 = n1166 & n1167;
  assign n1090 = n1168 & n1169;
  assign n986 = n1067 ^ n942;
  assign n981 = n1172 & n1173;
  assign n1082 = ~n1163;
  assign n1006 = ~n926;
  assign n1075 = ~n1062;
  assign n987 = n1175 & n1176;
  assign n960 = ~n1177;
  assign n1066 = ~n985;
  assign n1107 = n1094 & n1183;
  assign n997 = n1184 & n1185;
  assign n663 = n1186 & n1187;
  assign n1117 = n1140 & n1189;
  assign n1123 = n1192 & n1193;
  assign n1137 = n1200 & n1201;
  assign n1040 = ~n1022;
  assign n1034 = ~n1118;
  assign n983 = n1202 & n1203;
  assign n1150 = n1204 & n1205;
  assign n989 = n1206 & n1207;
  assign n1056 = ~n1208;
  assign n408 = ~n1210;
  assign n107 = ~n1211;
  assign n1135 = ~n1200;
  assign n1148 = ~n1052;
  assign n1174 = n1227 & n1228;
  assign n958 = ~n1233;
  assign n1151 = ~n1146;
  assign n1153 = ~n1126;
  assign n696 = ~n687;
  assign n903 = ~n886;
  assign n1155 = ~n1050;
  assign n1181 = n1244 & n1245;
  assign n413 = ~n1250;
  assign n114 = ~n1252;
  assign n1161 = ~n1166;
  assign n1102 = ~n1144;
  assign n1036 = ~n1120;
  assign n1054 = ~n1024;
  assign n1108 = ~n1092;
  assign n1106 = ~n1094;
  assign n1100 = ~n1138;
  assign n1015 = ~n1269;
  assign n1111 = ~n1140;
  assign n1159 = ~n1168;
  assign n1194 = n1270 & n1271;
  assign n1113 = ~n1192;
  assign n12381 = n1380 ^ n1381;
  assign n1346 = ~n1380;
  assign n621 = n852 ^ n853;
  assign n807 = n861 & n862;
  assign n738 = ~n868;
  assign n709 = n792 ^ n883;
  assign n716 = n884 ^ n885;
  assign n847 = n898 & n899;
  assign n848 = n903 & n904;
  assign n357 = ~n908;
  assign n635 = ~n910;
  assign n770 = n911 ^ n912;
  assign n772 = n913 ^ n914;
  assign n869 = n852 & n853;
  assign n734 = n924 ^ n925;
  assign n780 = n926 ^ n927;
  assign n877 = n939 & n940;
  assign n880 = n396 & n399;
  assign n891 = n958 & n959;
  assign n892 = n960 & n961;
  assign n909 = n971 & n972;
  assign n778 = ~n833;
  assign n840 = ~n975;
  assign n842 = ~n979;
  assign n921 = n708 & n980;
  assign n922 = n912 & n911;
  assign n923 = n913 & n914;
  assign n845 = ~n906;
  assign n834 = n981 ^ n982;
  assign n836 = n983 ^ n984;
  assign n838 = n985 ^ n986;
  assign n552 = ~n573;
  assign n796 = n987 ^ n988;
  assign n782 = n989 ^ n990;
  assign n375 = ~n994;
  assign n946 = n924 & n925;
  assign n863 = ~n852;
  assign n798 = n997 ^ n998;
  assign n799 = n960 ^ n999;
  assign n757 = ~n1007;
  assign n740 = ~n769;
  assign n941 = ~n1012;
  assign n943 = ~n924;
  assign n870 = n1015 ^ n1016;
  assign n949 = ~n1018;
  assign n970 = n663 & n575;
  assign n976 = n1034 & n1035;
  assign n977 = n1036 & n1037;
  assign n978 = n1040 & n1041;
  assign n372 = ~n1044;
  assign n691 = ~n1045;
  assign n888 = ~n1046;
  assign n699 = ~n751;
  assign n920 = ~n708;
  assign n993 = n1054 & n1055;
  assign n907 = n1056 & n1057;
  assign n896 = ~n971;
  assign n850 = n958 ^ n1061;
  assign n655 = ~n711;
  assign n762 = ~n810;
  assign n916 = ~n912;
  assign n918 = ~n913;
  assign n1000 = n1066 & n1067;
  assign n1008 = n1075 & n1076;
  assign n1009 = n1082 & n1083;
  assign n126 = ~n1085;
  assign n995 = ~n1086;
  assign n119 = ~n1087;
  assign n393 = ~n1090;
  assign n1001 = ~n981;
  assign n1019 = n1100 & n1101;
  assign n1020 = n1102 & n1103;
  assign n1003 = ~n987;
  assign n1021 = n1106 & n1095;
  assign n1005 = ~n1107;
  assign n964 = ~n997;
  assign n1026 = n1108 & n1109;
  assign n962 = ~n663;
  assign n1027 = n1015 & n1110;
  assign n1032 = n1111 & n1112;
  assign n1033 = n1113 & n1114;
  assign n966 = ~n1117;
  assign n365 = ~n1123;
  assign n1058 = n1135 & n1136;
  assign n385 = ~n1137;
  assign n991 = ~n983;
  assign n1070 = n1148 & n1149;
  assign n928 = ~n1150;
  assign n1077 = n1151 & n1152;
  assign n1078 = n1153 & n1154;
  assign n973 = ~n989;
  assign n1079 = n1155 & n1156;
  assign n1081 = n1159 & n1160;
  assign n1084 = n1161 & n1162;
  assign n1068 = ~n1174;
  assign n109 = ~n1181;
  assign n1030 = ~n1194;
  assign n1255 = n1346 & n1347;
  assign n503 = n708 ^ n709;
  assign n647 = n769 ^ n770;
  assign n609 = n780 ^ n781;
  assign n713 = n782 ^ n783;
  assign n749 = n780 & n781;
  assign n668 = n797 ^ n798;
  assign n728 = n799 ^ n800;
  assign n626 = ~n807;
  assign n649 = n834 ^ n835;
  assign n651 = n836 ^ n837;
  assign n653 = n838 ^ n701;
  assign n658 = ~n716;
  assign n727 = n840 & n841;
  assign n581 = n842 & n843;
  assign n354 = ~n847;
  assign n542 = ~n848;
  assign n793 = n834 & n835;
  assign n794 = n836 & n837;
  assign n730 = n850 ^ n851;
  assign n808 = n863 & n864;
  assign n377 = n375 & n379;
  assign n811 = n798 & n797;
  assign n602 = ~n869;
  assign n688 = n870 ^ n871;
  assign n745 = ~n780;
  assign n756 = ~n877;
  assign n401 = ~n880;
  assign n839 = n888 & n889;
  assign n824 = ~n891;
  assign n826 = ~n892;
  assign n846 = n896 & n897;
  assign n849 = n906 & n907;
  assign n350 = ~n909;
  assign n860 = n916 & n917;
  assign n865 = n918 & n919;
  assign n867 = n920 & n883;
  assign n791 = ~n921;
  assign n631 = ~n922;
  assign n614 = ~n923;
  assign n787 = ~n834;
  assign n789 = ~n836;
  assign n595 = ~n838;
  assign n742 = ~n796;
  assign n731 = n928 ^ n929;
  assign n878 = n941 & n942;
  assign n879 = n943 & n944;
  assign n598 = ~n946;
  assign n805 = ~n798;
  assign n809 = n949 & n950;
  assign n890 = n928 & n957;
  assign n895 = n962 & n963;
  assign n900 = n964 & n965;
  assign n905 = n966 & n967;
  assign n679 = ~n970;
  assign n915 = n973 & n974;
  assign n368 = ~n976;
  assign n774 = ~n977;
  assign n586 = ~n978;
  assign n930 = n991 & n992;
  assign n858 = ~n993;
  assign n844 = ~n907;
  assign n945 = n995 & n996;
  assign n759 = ~n1000;
  assign n948 = n1001 & n1002;
  assign n951 = n1003 & n1004;
  assign n952 = n1005 & n1006;
  assign n875 = ~n1008;
  assign n123 = ~n1009;
  assign n953 = ~n1019;
  assign n955 = ~n1020;
  assign n820 = ~n1021;
  assign n901 = ~n1026;
  assign n893 = ~n1027;
  assign n931 = n1030 & n1031;
  assign n831 = ~n1032;
  assign n361 = ~n1033;
  assign n382 = ~n1058;
  assign n733 = n1068 & n1069;
  assign n804 = ~n1070;
  assign n935 = ~n1077;
  assign n933 = ~n1078;
  assign n937 = ~n1079;
  assign n389 = ~n1081;
  assign n116 = ~n1084;
  assign n1010 = n109 & n114;
  assign n1096 = ~n1255;
  assign n484 = ~n503;
  assign n582 = n687 ^ n688;
  assign n605 = ~n647;
  assign n685 = n727 & n728;
  assign n666 = n731 ^ n732;
  assign n660 = ~n713;
  assign n547 = n733 ^ n734;
  assign n700 = n745 & n746;
  assign n538 = ~n749;
  assign n702 = n688 & n687;
  assign n683 = ~n728;
  assign n620 = n756 & n757;
  assign n726 = n354 & n357;
  assign n682 = ~n727;
  assign n633 = ~n581;
  assign n743 = n787 & n788;
  assign n744 = n789 & n790;
  assign n747 = n791 & n792;
  assign n674 = ~n793;
  assign n676 = ~n794;
  assign n681 = ~n730;
  assign n760 = n805 & n806;
  assign n550 = ~n808;
  assign n765 = n809 & n810;
  assign n693 = ~n811;
  assign n695 = ~n688;
  assign n665 = n824 & n825;
  assign n712 = n826 & n827;
  assign n773 = ~n839;
  assign n786 = n844 & n845;
  assign n347 = ~n846;
  assign n370 = n368 & n372;
  assign n343 = ~n849;
  assign n750 = n858 & n859;
  assign n739 = ~n860;
  assign n776 = ~n865;
  assign n672 = ~n867;
  assign n717 = n875 & n876;
  assign n758 = ~n878;
  assign n755 = ~n879;
  assign n821 = n123 & n126;
  assign n761 = ~n809;
  assign n822 = ~n890;
  assign n771 = n893 & n894;
  assign n567 = ~n895;
  assign n828 = ~n900;
  assign n735 = n901 & n902;
  assign n363 = n361 & n365;
  assign n830 = ~n905;
  assign n784 = ~n915;
  assign n866 = n382 & n385;
  assign n801 = ~n930;
  assign n874 = n931 & n932;
  assign n795 = n933 & n934;
  assign n719 = n935 & n936;
  assign n832 = n937 & n938;
  assign n390 = n389 & n393;
  assign n803 = ~n945;
  assign n881 = n116 & n119;
  assign n815 = ~n948;
  assign n817 = ~n951;
  assign n819 = ~n952;
  assign n812 = n953 & n954;
  assign n667 = n955 & n956;
  assign n872 = ~n931;
  assign n754 = ~n733;
  assign n112 = ~n1010;
  assign n1017 = n1096 & n1097;
  assign n486 = n581 ^ n582;
  assign n559 = n620 ^ n621;
  assign n619 = n665 & n666;
  assign n557 = n667 ^ n668;
  assign n637 = n682 & n683;
  assign n329 = ~n685;
  assign n616 = ~n666;
  assign n515 = ~n547;
  assign n640 = n695 & n696;
  assign n628 = ~n700;
  assign n632 = ~n702;
  assign n601 = ~n620;
  assign n661 = n712 & n713;
  assign n493 = n717 ^ n718;
  assign n561 = n719 ^ n720;
  assign n359 = ~n726;
  assign n569 = n735 ^ n736;
  assign n694 = n739 & n740;
  assign n563 = ~n743;
  assign n565 = ~n744;
  assign n671 = ~n747;
  assign n703 = n750 & n751;
  assign n705 = n754 & n755;
  assign n611 = n758 & n759;
  assign n591 = ~n760;
  assign n706 = n761 & n762;
  assign n140 = ~n765;
  assign n495 = n771 ^ n772;
  assign n646 = n773 & n774;
  assign n615 = ~n665;
  assign n659 = ~n712;
  assign n725 = n347 & n350;
  assign n729 = n784 & n785;
  assign n340 = ~n786;
  assign n748 = n795 & n796;
  assign n652 = n801 & n802;
  assign n608 = n803 & n804;
  assign n698 = ~n750;
  assign n766 = n812 & n813;
  assign n650 = n815 & n816;
  assign n710 = n817 & n818;
  assign n648 = n819 & n820;
  assign n690 = ~n717;
  assign n128 = ~n821;
  assign n715 = n822 & n823;
  assign n662 = n828 & n829;
  assign n721 = n830 & n831;
  assign n779 = n832 & n833;
  assign n775 = ~n771;
  assign n752 = ~n735;
  assign n387 = ~n866;
  assign n814 = n872 & n873;
  assign n336 = ~n874;
  assign n741 = ~n795;
  assign n737 = ~n719;
  assign n777 = ~n832;
  assign n121 = ~n881;
  assign n763 = ~n812;
  assign n692 = ~n667;
  assign n855 = ~n1017;
  assign n475 = ~n486;
  assign n529 = ~n559;
  assign n576 = n601 & n602;
  assign n555 = n608 ^ n609;
  assign n461 = n611 ^ n612;
  assign n583 = n615 & n616;
  assign n309 = ~n619;
  assign n526 = ~n557;
  assign n592 = n632 & n633;
  assign n326 = ~n637;
  assign n540 = ~n640;
  assign n607 = n646 & n647;
  assign n491 = n648 ^ n649;
  assign n505 = n650 ^ n651;
  assign n507 = n652 ^ n653;
  assign n618 = n659 & n660;
  assign n322 = ~n661;
  assign n574 = n662 ^ n663;
  assign n466 = ~n493;
  assign n531 = ~n561;
  assign n554 = n671 & n672;
  assign n544 = ~n569;
  assign n638 = n690 & n691;
  assign n639 = n692 & n693;
  assign n630 = ~n694;
  assign n643 = n698 & n699;
  assign n644 = n652 & n701;
  assign n168 = ~n703;
  assign n597 = ~n705;
  assign n634 = ~n611;
  assign n137 = ~n706;
  assign n656 = n710 & n711;
  assign n664 = n715 & n716;
  assign n464 = ~n495;
  assign n677 = n721 & n722;
  assign n604 = ~n646;
  assign n352 = ~n725;
  assign n684 = n340 & n343;
  assign n686 = n729 & n730;
  assign n680 = ~n729;
  assign n689 = n737 & n738;
  assign n697 = n741 & n742;
  assign n163 = ~n748;
  assign n641 = ~n652;
  assign n704 = n752 & n753;
  assign n627 = ~n608;
  assign n707 = n763 & n764;
  assign n147 = ~n766;
  assign n675 = ~n650;
  assign n654 = ~n710;
  assign n673 = ~n648;
  assign n657 = ~n715;
  assign n723 = n775 & n776;
  assign n724 = n777 & n778;
  assign n678 = ~n662;
  assign n669 = ~n721;
  assign n175 = ~n779;
  assign n333 = ~n814;
  assign n12382 = n854 ^ n855;
  assign n882 = n855 & n947;
  assign n524 = n554 & n555;
  assign n545 = n326 & n329;
  assign n518 = n574 ^ n575;
  assign n549 = ~n576;
  assign n521 = ~n555;
  assign n454 = ~n461;
  assign n305 = ~n583;
  assign n539 = ~n592;
  assign n568 = n597 & n598;
  assign n577 = n604 & n605;
  assign n578 = n137 & n140;
  assign n294 = ~n607;
  assign n477 = ~n491;
  assign n480 = ~n505;
  assign n482 = ~n507;
  assign n319 = ~n618;
  assign n520 = ~n554;
  assign n587 = n627 & n628;
  assign n556 = n630 & n631;
  assign n593 = n634 & n635;
  assign n585 = ~n638;
  assign n590 = ~n639;
  assign n603 = n641 & n642;
  assign n165 = ~n643;
  assign n594 = ~n644;
  assign n610 = n654 & n655;
  assign n156 = ~n656;
  assign n617 = n657 & n658;
  assign n302 = ~n664;
  assign n622 = n669 & n670;
  assign n623 = n673 & n674;
  assign n624 = n675 & n676;
  assign n133 = ~n677;
  assign n629 = n678 & n679;
  assign n636 = n680 & n681;
  assign n345 = ~n684;
  assign n316 = ~n686;
  assign n625 = ~n689;
  assign n158 = ~n697;
  assign n645 = n333 & n336;
  assign n599 = ~n704;
  assign n144 = ~n707;
  assign n613 = ~n723;
  assign n172 = ~n724;
  assign n767 = ~n882;
  assign n500 = n520 & n521;
  assign n266 = ~n524;
  assign n307 = n305 & n309;
  assign n494 = n539 & n540;
  assign n331 = ~n545;
  assign n492 = n549 & n550;
  assign n497 = ~n518;
  assign n532 = n319 & n322;
  assign n533 = n556 & n557;
  assign n548 = n568 & n569;
  assign n543 = ~n568;
  assign n291 = ~n577;
  assign n142 = ~n578;
  assign n546 = n585 & n586;
  assign n537 = ~n587;
  assign n517 = n590 & n591;
  assign n525 = ~n556;
  assign n541 = ~n593;
  assign n570 = n594 & n595;
  assign n571 = n165 & n168;
  assign n572 = n599 & n600;
  assign n512 = ~n603;
  assign n579 = n144 & n147;
  assign n151 = ~n610;
  assign n560 = n613 & n614;
  assign n298 = ~n617;
  assign n584 = n172 & n175;
  assign n130 = ~n622;
  assign n562 = ~n623;
  assign n564 = ~n624;
  assign n558 = n625 & n626;
  assign n566 = ~n629;
  assign n312 = ~n636;
  assign n596 = n158 & n163;
  assign n338 = ~n645;
  assign n714 = n767 & n768;
  assign n467 = n492 & n493;
  assign n468 = n494 & n495;
  assign n263 = ~n500;
  assign n463 = ~n494;
  assign n499 = n517 & n518;
  assign n465 = ~n492;
  assign n501 = n291 & n294;
  assign n508 = n525 & n526;
  assign n324 = ~n532;
  assign n287 = ~n533;
  assign n490 = n537 & n538;
  assign n485 = n541 & n542;
  assign n513 = n543 & n544;
  assign n516 = n546 & n547;
  assign n189 = ~n548;
  assign n527 = n151 & n156;
  assign n300 = n298 & n302;
  assign n534 = n558 & n559;
  assign n535 = n560 & n561;
  assign n536 = n130 & n133;
  assign n504 = n562 & n563;
  assign n506 = n564 & n565;
  assign n502 = n566 & n567;
  assign n314 = n312 & n316;
  assign n514 = ~n546;
  assign n496 = ~n517;
  assign n511 = ~n570;
  assign n170 = ~n571;
  assign n553 = n572 & n573;
  assign n551 = ~n572;
  assign n149 = ~n579;
  assign n530 = ~n560;
  assign n177 = ~n584;
  assign n528 = ~n558;
  assign n161 = ~n596;
  assign n589 = ~n714;
  assign n447 = n463 & n464;
  assign n448 = n465 & n466;
  assign n203 = ~n467;
  assign n224 = ~n468;
  assign n452 = n263 & n266;
  assign n459 = n485 & n486;
  assign n462 = n490 & n491;
  assign n469 = n496 & n497;
  assign n280 = ~n499;
  assign n296 = ~n501;
  assign n487 = n502 & n503;
  assign n488 = n504 & n505;
  assign n489 = n506 & n507;
  assign n284 = ~n508;
  assign n460 = n511 & n512;
  assign n476 = ~n490;
  assign n474 = ~n485;
  assign n186 = ~n513;
  assign n498 = n514 & n515;
  assign n196 = ~n516;
  assign n154 = ~n527;
  assign n509 = n528 & n529;
  assign n510 = n530 & n531;
  assign n210 = ~n534;
  assign n217 = ~n535;
  assign n135 = ~n536;
  assign n479 = ~n504;
  assign n481 = ~n506;
  assign n483 = ~n502;
  assign n519 = n551 & n552;
  assign n182 = ~n553;
  assign n12383 = n588 ^ n589;
  assign n580 = n589 & n606;
  assign n221 = ~n447;
  assign n200 = ~n448;
  assign n268 = ~n452;
  assign n443 = n284 & n287;
  assign n231 = ~n459;
  assign n446 = n460 & n461;
  assign n261 = ~n462;
  assign n449 = n186 & n189;
  assign n277 = ~n469;
  assign n455 = n474 & n475;
  assign n456 = n476 & n477;
  assign n478 = n479 & n480;
  assign n457 = n481 & n482;
  assign n458 = n483 & n484;
  assign n273 = ~n487;
  assign n254 = ~n488;
  assign n247 = ~n489;
  assign n453 = ~n460;
  assign n193 = ~n498;
  assign n207 = ~n509;
  assign n214 = ~n510;
  assign n179 = ~n519;
  assign n522 = ~n580;
  assign n431 = n200 & n203;
  assign n432 = n221 & n224;
  assign n435 = n277 & n280;
  assign n289 = ~n443;
  assign n238 = ~n446;
  assign n191 = ~n449;
  assign n441 = n193 & n196;
  assign n442 = n453 & n454;
  assign n228 = ~n455;
  assign n256 = ~n456;
  assign n242 = ~n457;
  assign n270 = ~n458;
  assign n444 = n207 & n210;
  assign n445 = n214 & n217;
  assign n450 = n179 & n182;
  assign n249 = ~n478;
  assign n472 = n522 & n523;
  assign n205 = ~n431;
  assign n226 = ~n432;
  assign n282 = ~n435;
  assign n433 = n228 & n231;
  assign n434 = n256 & n261;
  assign n198 = ~n441;
  assign n438 = n242 & n247;
  assign n439 = n249 & n254;
  assign n440 = n270 & n273;
  assign n235 = ~n442;
  assign n212 = ~n444;
  assign n219 = ~n445;
  assign n184 = ~n450;
  assign n12384 = n472 ^ n473;
  assign n470 = ~n472;
  assign n233 = ~n433;
  assign n430 = n235 & n238;
  assign n259 = ~n434;
  assign n245 = ~n438;
  assign n252 = ~n439;
  assign n275 = ~n440;
  assign n451 = n470 & n471;
  assign n240 = ~n430;
  assign n436 = ~n451;
  assign n428 = n436 & n437;
  assign n12385 = n428 ^ n429;
  assign n426 = ~n428;
  assign n425 = n426 & n427;
  assign n423 = ~n425;
  assign n422 = n423 & n424;
  assign n419 = ~n422;
  assign n12386 = n418 ^ n419;
  assign n420 = n419 & n421;
  assign n416 = ~n420;
  assign n412 = n416 & n417;
  assign n12387 = n412 ^ n413;
  assign n414 = ~n412;
  assign n411 = n414 & n415;
  assign n409 = ~n411;
  assign n407 = n409 & n410;
  assign n12388 = n407 ^ n408;
  assign n405 = ~n407;
  assign n404 = n405 & n406;
  assign n402 = ~n404;
  assign n400 = n402 & n403;
  assign n12389 = n400 ^ n401;
  assign n398 = ~n400;
  assign n397 = n398 & n399;
  assign n395 = ~n397;
  assign n394 = n395 & n396;
  assign n391 = ~n394;
  assign n12390 = n390 ^ n391;
  assign n392 = n391 & n393;
  assign n388 = ~n392;
  assign n386 = n388 & n389;
  assign n12391 = n386 ^ n387;
  assign n384 = ~n386;
  assign n383 = n384 & n385;
  assign n381 = ~n383;
  assign n380 = n381 & n382;
  assign n378 = ~n380;
  assign n12392 = n377 ^ n378;
  assign n376 = n378 & n379;
  assign n374 = ~n376;
  assign n373 = n374 & n375;
  assign n371 = ~n373;
  assign n12393 = n370 ^ n371;
  assign n369 = n371 & n372;
  assign n367 = ~n369;
  assign n366 = n367 & n368;
  assign n364 = ~n366;
  assign n12394 = n363 ^ n364;
  assign n362 = n364 & n365;
  assign n360 = ~n362;
  assign n358 = n360 & n361;
  assign n12395 = n358 ^ n359;
  assign n356 = ~n358;
  assign n355 = n356 & n357;
  assign n353 = ~n355;
  assign n351 = n353 & n354;
  assign n12396 = n351 ^ n352;
  assign n349 = ~n351;
  assign n348 = n349 & n350;
  assign n346 = ~n348;
  assign n344 = n346 & n347;
  assign n12397 = n344 ^ n345;
  assign n342 = ~n344;
  assign n341 = n342 & n343;
  assign n339 = ~n341;
  assign n337 = n339 & n340;
  assign n12398 = n337 ^ n338;
  assign n335 = ~n337;
  assign n334 = n335 & n336;
  assign n332 = ~n334;
  assign n330 = n332 & n333;
  assign n12399 = n330 ^ n331;
  assign n328 = ~n330;
  assign n327 = n328 & n329;
  assign n325 = ~n327;
  assign n323 = n325 & n326;
  assign n12400 = n323 ^ n324;
  assign n321 = ~n323;
  assign n320 = n321 & n322;
  assign n318 = ~n320;
  assign n317 = n318 & n319;
  assign n315 = ~n317;
  assign n12401 = n314 ^ n315;
  assign n313 = n315 & n316;
  assign n311 = ~n313;
  assign n310 = n311 & n312;
  assign n308 = ~n310;
  assign n12402 = n307 ^ n308;
  assign n306 = n308 & n309;
  assign n304 = ~n306;
  assign n303 = n304 & n305;
  assign n301 = ~n303;
  assign n12403 = n300 ^ n301;
  assign n299 = n301 & n302;
  assign n297 = ~n299;
  assign n295 = n297 & n298;
  assign n12404 = n295 ^ n296;
  assign n293 = ~n295;
  assign n292 = n293 & n294;
  assign n290 = ~n292;
  assign n288 = n290 & n291;
  assign n12405 = n288 ^ n289;
  assign n286 = ~n288;
  assign n285 = n286 & n287;
  assign n283 = ~n285;
  assign n281 = n283 & n284;
  assign n12406 = n281 ^ n282;
  assign n279 = ~n281;
  assign n278 = n279 & n280;
  assign n276 = ~n278;
  assign n274 = n276 & n277;
  assign n12407 = n274 ^ n275;
  assign n272 = ~n274;
  assign n271 = n272 & n273;
  assign n269 = ~n271;
  assign n267 = n269 & n270;
  assign n12408 = n267 ^ n268;
  assign n265 = ~n267;
  assign n264 = n265 & n266;
  assign n262 = ~n264;
  assign n258 = n262 & n263;
  assign n12409 = n258 ^ n259;
  assign n260 = ~n258;
  assign n257 = n260 & n261;
  assign n255 = ~n257;
  assign n251 = n255 & n256;
  assign n12410 = n251 ^ n252;
  assign n253 = ~n251;
  assign n250 = n253 & n254;
  assign n248 = ~n250;
  assign n244 = n248 & n249;
  assign n12411 = n244 ^ n245;
  assign n246 = ~n244;
  assign n243 = n246 & n247;
  assign n241 = ~n243;
  assign n239 = n241 & n242;
  assign n12412 = n239 ^ n240;
  assign n237 = ~n239;
  assign n236 = n237 & n238;
  assign n234 = ~n236;
  assign n232 = n234 & n235;
  assign n12413 = n232 ^ n233;
  assign n230 = ~n232;
  assign n229 = n230 & n231;
  assign n227 = ~n229;
  assign n225 = n227 & n228;
  assign n12414 = n225 ^ n226;
  assign n223 = ~n225;
  assign n222 = n223 & n224;
  assign n220 = ~n222;
  assign n218 = n220 & n221;
  assign n12415 = n218 ^ n219;
  assign n216 = ~n218;
  assign n215 = n216 & n217;
  assign n213 = ~n215;
  assign n211 = n213 & n214;
  assign n12416 = n211 ^ n212;
  assign n209 = ~n211;
  assign n208 = n209 & n210;
  assign n206 = ~n208;
  assign n204 = n206 & n207;
  assign n12417 = n204 ^ n205;
  assign n202 = ~n204;
  assign n201 = n202 & n203;
  assign n199 = ~n201;
  assign n197 = n199 & n200;
  assign n12418 = n197 ^ n198;
  assign n195 = ~n197;
  assign n194 = n195 & n196;
  assign n192 = ~n194;
  assign n190 = n192 & n193;
  assign n12419 = n190 ^ n191;
  assign n188 = ~n190;
  assign n187 = n188 & n189;
  assign n185 = ~n187;
  assign n183 = n185 & n186;
  assign n12420 = n183 ^ n184;
  assign n181 = ~n183;
  assign n180 = n181 & n182;
  assign n178 = ~n180;
  assign n176 = n178 & n179;
  assign n12421 = n176 ^ n177;
  assign n174 = ~n176;
  assign n173 = n174 & n175;
  assign n171 = ~n173;
  assign n169 = n171 & n172;
  assign n12422 = n169 ^ n170;
  assign n167 = ~n169;
  assign n166 = n167 & n168;
  assign n164 = ~n166;
  assign n160 = n164 & n165;
  assign n12423 = n160 ^ n161;
  assign n162 = ~n160;
  assign n159 = n162 & n163;
  assign n157 = ~n159;
  assign n153 = n157 & n158;
  assign n12424 = n153 ^ n154;
  assign n155 = ~n153;
  assign n152 = n155 & n156;
  assign n150 = ~n152;
  assign n148 = n150 & n151;
  assign n12425 = n148 ^ n149;
  assign n146 = ~n148;
  assign n145 = n146 & n147;
  assign n143 = ~n145;
  assign n141 = n143 & n144;
  assign n12426 = n141 ^ n142;
  assign n139 = ~n141;
  assign n138 = n139 & n140;
  assign n136 = ~n138;
  assign n134 = n136 & n137;
  assign n12427 = n134 ^ n135;
  assign n132 = ~n134;
  assign n131 = n132 & n133;
  assign n129 = ~n131;
  assign n127 = n129 & n130;
  assign n12428 = n127 ^ n128;
  assign n125 = ~n127;
  assign n124 = n125 & n126;
  assign n122 = ~n124;
  assign n120 = n122 & n123;
  assign n12429 = n120 ^ n121;
  assign n118 = ~n120;
  assign n117 = n118 & n119;
  assign n115 = ~n117;
  assign n111 = n115 & n116;
  assign n12430 = n111 ^ n112;
  assign n113 = ~n111;
  assign n110 = n113 & n114;
  assign n108 = ~n110;
  assign n106 = n108 & n109;
  assign n12431 = n106 ^ n107;
  assign n104 = ~n106;
  assign n103 = n104 & n105;
  assign n101 = ~n103;
  assign n99 = n101 & n102;
  assign n12432 = n99 ^ n100;
  assign n97 = ~n99;
  assign n96 = n97 & n98;
  assign n94 = ~n96;
  assign n92 = n94 & n95;
  assign n12433 = n92 ^ n93;
  assign n90 = ~n92;
  assign n89 = n90 & n91;
  assign n87 = ~n89;
  assign n85 = n87 & n88;
  assign n12434 = n85 ^ n86;
  assign n83 = ~n85;
  assign n82 = n83 & n84;
  assign n80 = ~n82;
  assign n76 = n80 & n81;
  assign n12435 = n76 ^ n77;
  assign n78 = ~n76;
  assign n75 = n78 & n79;
  assign n73 = ~n75;
  assign n71 = n73 & n74;
  assign n12436 = n71 ^ n72;
  assign n69 = ~n71;
  assign n68 = n69 & n70;
  assign n66 = ~n68;
  assign n64 = n66 & n67;
  assign n12437 = n64 ^ n65;
endmodule
