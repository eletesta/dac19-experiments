module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141;
  wire n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987;
  assign n148 = ~x8 & ~x10;
  assign n149 = ~x14 & ~x21;
  assign n150 = n148 & n149;
  assign n151 = ~x13 & n150;
  assign n152 = ~x4 & ~x9;
  assign n153 = ~x12 & n152;
  assign n154 = ~x7 & n153;
  assign n155 = n151 & n154;
  assign n156 = ~x6 & ~x7;
  assign n157 = x12 & x13;
  assign n158 = n156 & ~n157;
  assign n159 = ~x12 & ~x13;
  assign n160 = n159 ^ x9;
  assign n161 = n158 & ~n160;
  assign n162 = ~x9 & n159;
  assign n163 = x7 ^ x6;
  assign n164 = n162 & n163;
  assign n165 = ~n161 & ~n164;
  assign n166 = n155 & n165;
  assign n167 = ~x5 & ~x22;
  assign n168 = ~x11 & n167;
  assign n169 = ~x18 & ~x19;
  assign n170 = ~x16 & n169;
  assign n171 = n168 & n170;
  assign n172 = n166 & n171;
  assign n173 = ~x17 & n172;
  assign n174 = x54 & ~n173;
  assign n175 = ~x0 & ~n174;
  assign n176 = ~x13 & n149;
  assign n177 = ~x7 & n176;
  assign n178 = x13 & ~n149;
  assign n179 = x14 & x21;
  assign n180 = n148 & ~n179;
  assign n181 = ~n178 & n180;
  assign n182 = ~n177 & n181;
  assign n183 = x10 ^ x8;
  assign n184 = n176 & n183;
  assign n185 = ~n182 & ~n184;
  assign n186 = x7 & ~n151;
  assign n187 = ~n185 & ~n186;
  assign n188 = ~x6 & n170;
  assign n189 = n153 & n188;
  assign n190 = n187 & n189;
  assign n191 = ~x17 & x54;
  assign n192 = n168 & n191;
  assign n193 = n190 & n192;
  assign n194 = ~x9 & ~x11;
  assign n195 = n194 ^ n167;
  assign n196 = x54 & ~x56;
  assign n197 = n195 & n196;
  assign n198 = ~n193 & ~n197;
  assign n199 = ~n175 & n198;
  assign n200 = ~x3 & ~x129;
  assign n201 = ~n199 & n200;
  assign n202 = ~n172 & n191;
  assign n203 = ~x1 & n200;
  assign n204 = ~n202 & n203;
  assign n205 = ~x5 & n165;
  assign n206 = n191 & n200;
  assign n207 = n170 & n206;
  assign n208 = ~x11 & ~x22;
  assign n209 = ~x4 & n208;
  assign n210 = n150 & n209;
  assign n211 = n207 & n210;
  assign n212 = ~n205 & n211;
  assign n213 = x5 & ~n166;
  assign n214 = n212 & ~n213;
  assign n215 = ~n204 & ~n214;
  assign n216 = ~x42 & ~x44;
  assign n217 = ~x40 & n216;
  assign n218 = ~x38 & ~x50;
  assign n219 = n217 & n218;
  assign n220 = ~x41 & ~x46;
  assign n221 = ~x47 & ~x48;
  assign n222 = n220 & n221;
  assign n223 = ~x43 & n222;
  assign n224 = n219 & n223;
  assign n225 = ~x24 & ~x49;
  assign n226 = ~x45 & n225;
  assign n227 = n224 & n226;
  assign n228 = x82 & ~n227;
  assign n229 = x122 & x127;
  assign n230 = ~x82 & n229;
  assign n231 = ~n228 & ~n230;
  assign n232 = ~x15 & ~x20;
  assign n233 = x82 & ~n232;
  assign n234 = n231 & ~n233;
  assign n235 = x2 & ~n234;
  assign n236 = ~x2 & n232;
  assign n237 = n226 & n236;
  assign n238 = n223 & n237;
  assign n239 = x82 & ~n238;
  assign n240 = x82 & ~n218;
  assign n241 = ~n239 & ~n240;
  assign n242 = x82 & ~n217;
  assign n243 = n241 & ~n242;
  assign n244 = ~n229 & n243;
  assign n245 = ~x65 & n244;
  assign n246 = ~n235 & ~n245;
  assign n247 = ~x129 & ~n246;
  assign n248 = ~x61 & ~x118;
  assign n249 = ~x129 & n248;
  assign n250 = ~n173 & n249;
  assign n251 = ~x123 & ~x129;
  assign n252 = x0 & ~x113;
  assign n253 = n251 & n252;
  assign n254 = ~n250 & ~n253;
  assign n255 = n168 & n206;
  assign n256 = n190 & n255;
  assign n257 = x10 & n256;
  assign n258 = ~x54 & n200;
  assign n259 = x4 & n258;
  assign n260 = ~n257 & ~n259;
  assign n261 = ~x16 & n255;
  assign n262 = n166 & n261;
  assign n263 = ~x29 & ~x59;
  assign n264 = n169 & n263;
  assign n265 = n262 & n264;
  assign n266 = ~x25 & x28;
  assign n267 = n265 & n266;
  assign n268 = x5 & n258;
  assign n269 = ~n267 & ~n268;
  assign n270 = x25 & ~x28;
  assign n271 = n265 & n270;
  assign n272 = x6 & n258;
  assign n273 = ~n271 & ~n272;
  assign n274 = x8 & n256;
  assign n275 = x7 & n258;
  assign n276 = ~n274 & ~n275;
  assign n277 = x21 & n256;
  assign n278 = x8 & n258;
  assign n279 = ~n277 & ~n278;
  assign n280 = ~x5 & n207;
  assign n281 = n166 & n280;
  assign n282 = x11 & ~x22;
  assign n283 = n281 & n282;
  assign n284 = x9 & n258;
  assign n285 = ~n283 & ~n284;
  assign n286 = x14 & n256;
  assign n287 = x10 & n258;
  assign n288 = ~n286 & ~n287;
  assign n289 = ~x11 & x22;
  assign n290 = n281 & n289;
  assign n291 = x11 & n258;
  assign n292 = ~n290 & ~n291;
  assign n293 = x18 & ~x19;
  assign n294 = n262 & n293;
  assign n295 = x12 & n258;
  assign n296 = ~n294 & ~n295;
  assign n297 = x29 & x54;
  assign n298 = ~x59 & n297;
  assign n299 = ~x25 & ~x28;
  assign n300 = n298 & n299;
  assign n301 = n200 & n300;
  assign n302 = n173 & n301;
  assign n303 = x13 & n258;
  assign n304 = ~n302 & ~n303;
  assign n305 = x13 & n256;
  assign n306 = x14 & n258;
  assign n307 = ~n305 & ~n306;
  assign n308 = x15 & ~n231;
  assign n309 = ~x15 & n227;
  assign n310 = x82 & n309;
  assign n311 = ~x82 & ~n229;
  assign n312 = ~x70 & n311;
  assign n313 = ~n310 & ~n312;
  assign n314 = ~n308 & n313;
  assign n315 = ~x70 & ~n229;
  assign n316 = n236 & ~n315;
  assign n317 = ~x129 & ~n316;
  assign n318 = ~n314 & n317;
  assign n319 = x6 & n214;
  assign n320 = x16 & n258;
  assign n321 = ~n319 & ~n320;
  assign n322 = ~x29 & x59;
  assign n323 = n299 & n322;
  assign n324 = n206 & n323;
  assign n325 = n172 & n324;
  assign n326 = x17 & n258;
  assign n327 = ~n325 & ~n326;
  assign n328 = x16 & n169;
  assign n329 = n255 & n328;
  assign n330 = n166 & n329;
  assign n331 = x18 & n258;
  assign n332 = ~n330 & ~n331;
  assign n333 = x54 & n200;
  assign n334 = x17 & n333;
  assign n335 = n172 & n334;
  assign n336 = x19 & n258;
  assign n337 = ~n335 & ~n336;
  assign n338 = n309 ^ x20;
  assign n339 = x82 & ~n338;
  assign n340 = x20 & ~n311;
  assign n341 = ~x71 & ~n229;
  assign n342 = x2 & x82;
  assign n343 = ~n341 & ~n342;
  assign n344 = ~n340 & n343;
  assign n345 = ~x129 & ~n344;
  assign n346 = ~n339 & n345;
  assign n347 = ~x18 & x19;
  assign n348 = n262 & n347;
  assign n349 = x21 & n258;
  assign n350 = ~n348 & ~n349;
  assign n351 = n166 & n212;
  assign n352 = x22 & n258;
  assign n353 = ~n351 & ~n352;
  assign n354 = ~x23 & x55;
  assign n355 = x61 & ~x129;
  assign n356 = ~n354 & n355;
  assign n357 = x63 & n244;
  assign n358 = x82 & n224;
  assign n359 = ~x45 & n358;
  assign n360 = x82 & ~n359;
  assign n361 = x82 & ~n237;
  assign n362 = n229 & ~n361;
  assign n363 = ~x24 & ~n362;
  assign n364 = ~n360 & n363;
  assign n365 = x24 & ~n359;
  assign n366 = ~n364 & ~n365;
  assign n367 = ~x129 & ~n366;
  assign n368 = ~n357 & n367;
  assign n369 = x53 & x58;
  assign n370 = ~x85 & ~n369;
  assign n371 = ~x53 & ~x58;
  assign n372 = ~n370 & ~n371;
  assign n373 = ~x85 & n371;
  assign n374 = ~x26 & ~x27;
  assign n375 = ~n373 & n374;
  assign n376 = ~n372 & n375;
  assign n377 = x26 & x27;
  assign n378 = n373 & ~n377;
  assign n379 = ~n374 & n378;
  assign n380 = ~n376 & ~n379;
  assign n381 = ~x116 & ~n380;
  assign n382 = ~x95 & ~x100;
  assign n383 = ~x97 & n382;
  assign n384 = ~x110 & ~n383;
  assign n385 = n373 & n374;
  assign n386 = n384 & n385;
  assign n387 = ~x39 & ~x52;
  assign n388 = ~x51 & n387;
  assign n389 = x26 & x116;
  assign n390 = n388 & n389;
  assign n391 = n378 & ~n390;
  assign n392 = ~n386 & n391;
  assign n393 = ~n381 & ~n392;
  assign n394 = x27 & x116;
  assign n395 = ~n388 & n394;
  assign n396 = n200 & ~n395;
  assign n397 = x116 & ~n374;
  assign n398 = ~x25 & ~n397;
  assign n399 = n396 & ~n398;
  assign n400 = ~n393 & n399;
  assign n401 = ~x96 & ~x110;
  assign n402 = n401 ^ x116;
  assign n403 = ~x85 & n402;
  assign n404 = n403 ^ x116;
  assign n405 = x100 & n404;
  assign n406 = n200 & n374;
  assign n407 = n371 & n406;
  assign n408 = n405 & n407;
  assign n409 = ~n400 & ~n408;
  assign n410 = x116 & n388;
  assign n411 = n373 & ~n410;
  assign n412 = x26 & ~x27;
  assign n413 = n200 & n412;
  assign n414 = n411 & n413;
  assign n415 = ~n408 & ~n414;
  assign n416 = ~x26 & x27;
  assign n417 = n411 & n416;
  assign n418 = x85 & x116;
  assign n419 = ~x95 & ~n418;
  assign n420 = n371 & n374;
  assign n421 = ~n419 & n420;
  assign n422 = ~x100 & n421;
  assign n423 = n404 & n422;
  assign n424 = ~n417 & ~n423;
  assign n425 = n200 & ~n424;
  assign n426 = x28 & n381;
  assign n427 = ~x26 & x28;
  assign n428 = ~n384 & n427;
  assign n429 = ~n390 & ~n428;
  assign n430 = ~x27 & n373;
  assign n431 = ~n429 & n430;
  assign n432 = ~n426 & ~n431;
  assign n433 = ~n381 & n425;
  assign n434 = n432 & ~n433;
  assign n435 = n200 & ~n434;
  assign n436 = ~n384 & n385;
  assign n437 = ~n381 & ~n436;
  assign n438 = x29 & ~n437;
  assign n439 = n382 & n401;
  assign n440 = ~x58 & ~n439;
  assign n441 = x58 & ~x116;
  assign n442 = x97 & ~n441;
  assign n443 = ~n440 & n442;
  assign n444 = ~x53 & ~n443;
  assign n445 = x53 & x116;
  assign n446 = n370 & ~n445;
  assign n447 = n406 & n446;
  assign n448 = ~n444 & n447;
  assign n449 = ~n381 & n448;
  assign n450 = ~n438 & ~n449;
  assign n451 = n200 & ~n450;
  assign n452 = x60 ^ x30;
  assign n453 = x109 & n452;
  assign n454 = n453 ^ x30;
  assign n455 = ~x106 & ~n454;
  assign n456 = ~x88 & x106;
  assign n457 = ~x129 & ~n456;
  assign n458 = ~n455 & n457;
  assign n459 = x31 ^ x30;
  assign n460 = ~x109 & n459;
  assign n461 = n460 ^ x30;
  assign n462 = ~x106 & ~n461;
  assign n463 = ~x89 & x106;
  assign n464 = ~x129 & ~n463;
  assign n465 = ~n462 & n464;
  assign n466 = x32 ^ x31;
  assign n467 = ~x109 & n466;
  assign n468 = n467 ^ x31;
  assign n469 = ~x106 & ~n468;
  assign n470 = ~x99 & x106;
  assign n471 = ~x129 & ~n470;
  assign n472 = ~n469 & n471;
  assign n473 = x33 ^ x32;
  assign n474 = ~x109 & n473;
  assign n475 = n474 ^ x32;
  assign n476 = ~x106 & ~n475;
  assign n477 = ~x90 & x106;
  assign n478 = ~x129 & ~n477;
  assign n479 = ~n476 & n478;
  assign n480 = x34 ^ x33;
  assign n481 = ~x109 & n480;
  assign n482 = n481 ^ x33;
  assign n483 = ~x106 & ~n482;
  assign n484 = ~x91 & x106;
  assign n485 = ~x129 & ~n484;
  assign n486 = ~n483 & n485;
  assign n487 = x35 ^ x34;
  assign n488 = ~x109 & n487;
  assign n489 = n488 ^ x34;
  assign n490 = ~x106 & ~n489;
  assign n491 = ~x92 & x106;
  assign n492 = ~x129 & ~n491;
  assign n493 = ~n490 & n492;
  assign n494 = x36 ^ x35;
  assign n495 = ~x109 & n494;
  assign n496 = n495 ^ x35;
  assign n497 = ~x106 & ~n496;
  assign n498 = ~x98 & x106;
  assign n499 = ~x129 & ~n498;
  assign n500 = ~n497 & n499;
  assign n501 = x37 ^ x36;
  assign n502 = ~x109 & n501;
  assign n503 = n502 ^ x36;
  assign n504 = ~x106 & ~n503;
  assign n505 = ~x93 & x106;
  assign n506 = ~x129 & ~n505;
  assign n507 = ~n504 & n506;
  assign n508 = x74 ^ x38;
  assign n509 = ~n229 & ~n508;
  assign n510 = n509 ^ x38;
  assign n511 = n241 & ~n510;
  assign n512 = n217 ^ x38;
  assign n513 = x82 & ~n512;
  assign n514 = ~x129 & ~n513;
  assign n515 = ~n511 & n514;
  assign n516 = ~x51 & x109;
  assign n517 = ~x52 & n516;
  assign n518 = n517 ^ x39;
  assign n519 = ~x106 & ~n518;
  assign n520 = ~x129 & ~n519;
  assign n521 = ~x73 & ~n229;
  assign n522 = n241 & ~n521;
  assign n523 = ~n242 & ~n522;
  assign n524 = x82 & ~n216;
  assign n525 = ~n230 & ~n524;
  assign n526 = x40 & ~n525;
  assign n527 = ~n523 & ~n526;
  assign n528 = ~x129 & ~n527;
  assign n529 = ~x46 & n219;
  assign n530 = n529 ^ x41;
  assign n531 = x82 & ~n530;
  assign n532 = ~x129 & ~n531;
  assign n533 = x76 ^ x41;
  assign n534 = ~n229 & ~n533;
  assign n535 = n534 ^ x41;
  assign n536 = ~n239 & ~n535;
  assign n537 = n532 & ~n536;
  assign n538 = n216 & ~n243;
  assign n539 = x44 & x82;
  assign n540 = ~n230 & ~n539;
  assign n541 = x42 & ~n540;
  assign n542 = ~x72 & ~n229;
  assign n543 = ~n524 & n542;
  assign n544 = ~n541 & ~n543;
  assign n545 = ~n538 & n544;
  assign n546 = ~x129 & ~n545;
  assign n547 = n219 & n220;
  assign n548 = n547 ^ x43;
  assign n549 = x82 & ~n548;
  assign n550 = ~x129 & ~n549;
  assign n551 = x77 ^ x43;
  assign n552 = ~n229 & ~n551;
  assign n553 = n552 ^ x43;
  assign n554 = ~n239 & ~n553;
  assign n555 = n550 & ~n554;
  assign n556 = x67 ^ x44;
  assign n557 = ~n229 & ~n556;
  assign n558 = n557 ^ x44;
  assign n559 = n243 & ~n558;
  assign n560 = ~x129 & ~n539;
  assign n561 = ~n559 & n560;
  assign n562 = ~x68 & ~n229;
  assign n563 = ~n361 & ~n562;
  assign n564 = ~n360 & ~n563;
  assign n565 = x45 & ~n311;
  assign n566 = ~n358 & n565;
  assign n567 = ~n564 & ~n566;
  assign n568 = ~x129 & ~n567;
  assign n569 = x75 ^ x46;
  assign n570 = ~n229 & ~n569;
  assign n571 = n570 ^ x46;
  assign n572 = n243 & ~n571;
  assign n573 = n219 ^ x46;
  assign n574 = x82 & ~n573;
  assign n575 = ~x129 & ~n574;
  assign n576 = ~n572 & n575;
  assign n577 = ~x43 & n547;
  assign n578 = n577 ^ x47;
  assign n579 = x82 & ~n578;
  assign n580 = x64 ^ x47;
  assign n581 = ~n229 & ~n580;
  assign n582 = n581 ^ x47;
  assign n583 = ~n239 & ~n582;
  assign n584 = ~x129 & ~n583;
  assign n585 = ~n579 & n584;
  assign n586 = ~x47 & n577;
  assign n587 = n586 ^ x48;
  assign n588 = x82 & ~n587;
  assign n589 = x48 & ~n311;
  assign n590 = ~x62 & ~n229;
  assign n591 = ~n589 & ~n590;
  assign n592 = ~n361 & n591;
  assign n593 = ~x129 & ~n592;
  assign n594 = ~n588 & n593;
  assign n595 = ~x24 & n359;
  assign n596 = x49 & ~n311;
  assign n597 = ~n595 & n596;
  assign n598 = x82 & ~n236;
  assign n599 = ~x69 & ~n229;
  assign n600 = ~n598 & ~n599;
  assign n601 = ~n228 & ~n600;
  assign n602 = ~n597 & ~n601;
  assign n603 = ~x129 & ~n602;
  assign n604 = ~x66 & ~n229;
  assign n605 = n238 & ~n604;
  assign n606 = ~n230 & ~n240;
  assign n607 = ~n242 & n606;
  assign n608 = ~n605 & n607;
  assign n609 = ~x50 & ~n608;
  assign n610 = ~x38 & n217;
  assign n611 = n240 & n610;
  assign n612 = x66 & n311;
  assign n613 = ~x129 & ~n612;
  assign n614 = ~n611 & n613;
  assign n615 = ~n609 & n614;
  assign n616 = x109 ^ x51;
  assign n617 = ~x106 & ~n616;
  assign n618 = ~x129 & ~n617;
  assign n619 = n516 ^ x52;
  assign n620 = ~x106 & ~n619;
  assign n621 = ~x129 & ~n620;
  assign n622 = ~x129 & ~n244;
  assign n623 = x114 & ~x122;
  assign n624 = n251 & n623;
  assign n625 = ~n376 & ~n378;
  assign n626 = n200 & ~n625;
  assign n627 = ~n389 & ~n441;
  assign n628 = ~x94 & ~n627;
  assign n629 = ~x37 & ~x58;
  assign n630 = ~n389 & n629;
  assign n631 = ~n628 & ~n630;
  assign n632 = n626 & n631;
  assign n633 = x58 & x116;
  assign n634 = x60 ^ x57;
  assign n635 = n633 & n634;
  assign n636 = n635 ^ x57;
  assign n637 = n626 & n636;
  assign n638 = n388 & n397;
  assign n639 = ~n441 & ~n638;
  assign n640 = n626 & ~n639;
  assign n641 = x59 & ~n437;
  assign n642 = x96 & n386;
  assign n643 = ~n641 & ~n642;
  assign n644 = n200 & ~n643;
  assign n645 = ~x117 & ~x122;
  assign n646 = x123 ^ x60;
  assign n647 = n645 & n646;
  assign n648 = n647 ^ x60;
  assign n649 = ~x114 & ~x122;
  assign n650 = x123 & ~x129;
  assign n651 = n649 & n650;
  assign n652 = x132 & x133;
  assign n653 = x131 & n652;
  assign n654 = ~x138 & n653;
  assign n655 = x136 & ~x137;
  assign n656 = n654 & n655;
  assign n657 = ~x62 & ~n656;
  assign n658 = ~x129 & ~n657;
  assign n659 = x140 & n656;
  assign n660 = n658 & ~n659;
  assign n661 = ~x63 & ~n656;
  assign n662 = ~x129 & ~n661;
  assign n663 = x142 & n656;
  assign n664 = n662 & ~n663;
  assign n665 = ~x64 & ~n656;
  assign n666 = ~x129 & ~n665;
  assign n667 = x139 & n656;
  assign n668 = n666 & ~n667;
  assign n669 = ~x65 & ~n656;
  assign n670 = ~x129 & ~n669;
  assign n671 = x146 & n656;
  assign n672 = n670 & ~n671;
  assign n673 = ~x136 & ~x137;
  assign n674 = n654 & n673;
  assign n675 = ~x66 & ~n674;
  assign n676 = ~x129 & ~n675;
  assign n677 = x143 & n674;
  assign n678 = n676 & ~n677;
  assign n679 = ~x67 & ~n674;
  assign n680 = ~x129 & ~n679;
  assign n681 = x139 & n674;
  assign n682 = n680 & ~n681;
  assign n683 = ~x68 & ~n656;
  assign n684 = ~x129 & ~n683;
  assign n685 = x141 & n656;
  assign n686 = n684 & ~n685;
  assign n687 = ~x69 & ~n656;
  assign n688 = ~x129 & ~n687;
  assign n689 = x143 & n656;
  assign n690 = n688 & ~n689;
  assign n691 = ~x70 & ~n656;
  assign n692 = ~x129 & ~n691;
  assign n693 = x144 & n656;
  assign n694 = n692 & ~n693;
  assign n695 = ~x71 & ~n656;
  assign n696 = ~x129 & ~n695;
  assign n697 = x145 & n656;
  assign n698 = n696 & ~n697;
  assign n699 = ~x72 & ~n674;
  assign n700 = ~x129 & ~n699;
  assign n701 = x140 & n674;
  assign n702 = n700 & ~n701;
  assign n703 = ~x73 & ~n674;
  assign n704 = ~x129 & ~n703;
  assign n705 = x141 & n674;
  assign n706 = n704 & ~n705;
  assign n707 = ~x74 & ~n674;
  assign n708 = ~x129 & ~n707;
  assign n709 = x142 & n674;
  assign n710 = n708 & ~n709;
  assign n711 = ~x75 & ~n674;
  assign n712 = ~x129 & ~n711;
  assign n713 = x144 & n674;
  assign n714 = n712 & ~n713;
  assign n715 = ~x76 & ~n674;
  assign n716 = ~x129 & ~n715;
  assign n717 = x145 & n674;
  assign n718 = n716 & ~n717;
  assign n719 = ~x77 & ~n674;
  assign n720 = ~x129 & ~n719;
  assign n721 = x146 & n674;
  assign n722 = n720 & ~n721;
  assign n723 = ~x136 & x137;
  assign n724 = n654 & n723;
  assign n725 = ~x142 & n724;
  assign n726 = ~x129 & ~n725;
  assign n727 = ~x78 & ~n724;
  assign n728 = n726 & ~n727;
  assign n729 = ~x143 & n724;
  assign n730 = ~x129 & ~n729;
  assign n731 = ~x79 & ~n724;
  assign n732 = n730 & ~n731;
  assign n733 = ~x144 & n724;
  assign n734 = ~x129 & ~n733;
  assign n735 = ~x80 & ~n724;
  assign n736 = n734 & ~n735;
  assign n737 = ~x145 & n724;
  assign n738 = ~x129 & ~n737;
  assign n739 = ~x81 & ~n724;
  assign n740 = n738 & ~n739;
  assign n741 = ~x146 & n724;
  assign n742 = ~x129 & ~n741;
  assign n743 = ~x82 & ~n724;
  assign n744 = n742 & ~n743;
  assign n745 = x62 ^ x31;
  assign n746 = ~x137 & ~n745;
  assign n747 = n746 ^ x31;
  assign n748 = ~x138 & n747;
  assign n749 = ~x137 & x138;
  assign n750 = x89 & n749;
  assign n751 = x136 & ~n750;
  assign n752 = ~n748 & n751;
  assign n753 = x87 & ~x138;
  assign n754 = n723 & ~n753;
  assign n755 = ~x115 & x138;
  assign n756 = n754 & ~n755;
  assign n757 = x119 & x138;
  assign n758 = n673 & ~n757;
  assign n759 = ~x72 & ~x138;
  assign n760 = n758 & ~n759;
  assign n761 = ~n756 & ~n760;
  assign n762 = ~n752 & n761;
  assign n763 = ~x141 & n724;
  assign n764 = ~x129 & ~n763;
  assign n765 = ~x84 & ~n724;
  assign n766 = n764 & ~n765;
  assign n767 = x96 & n384;
  assign n768 = ~x85 & ~n767;
  assign n769 = n407 & ~n418;
  assign n770 = ~n768 & n769;
  assign n771 = ~x139 & n724;
  assign n772 = ~x129 & ~n771;
  assign n773 = ~x86 & ~n724;
  assign n774 = n772 & ~n773;
  assign n775 = ~x140 & n724;
  assign n776 = ~x129 & ~n775;
  assign n777 = ~x87 & ~n724;
  assign n778 = n776 & ~n777;
  assign n779 = x136 & x137;
  assign n780 = n654 & n779;
  assign n781 = ~x139 & n780;
  assign n782 = ~x129 & ~n781;
  assign n783 = ~x88 & ~n780;
  assign n784 = n782 & ~n783;
  assign n785 = ~x140 & n780;
  assign n786 = ~x129 & ~n785;
  assign n787 = ~x89 & ~n780;
  assign n788 = n786 & ~n787;
  assign n789 = ~x142 & n780;
  assign n790 = ~x129 & ~n789;
  assign n791 = ~x90 & ~n780;
  assign n792 = n790 & ~n791;
  assign n793 = ~x143 & n780;
  assign n794 = ~x129 & ~n793;
  assign n795 = ~x91 & ~n780;
  assign n796 = n794 & ~n795;
  assign n797 = ~x144 & n780;
  assign n798 = ~x129 & ~n797;
  assign n799 = ~x92 & ~n780;
  assign n800 = n798 & ~n799;
  assign n801 = ~x146 & n780;
  assign n802 = ~x129 & ~n801;
  assign n803 = ~x93 & ~n780;
  assign n804 = n802 & ~n803;
  assign n805 = x82 & x138;
  assign n806 = n673 & n805;
  assign n807 = n653 & n806;
  assign n808 = ~x142 & n807;
  assign n809 = ~x129 & ~n808;
  assign n810 = ~x94 & ~n807;
  assign n811 = n809 & ~n810;
  assign n812 = ~x3 & ~x110;
  assign n813 = n812 ^ n806;
  assign n814 = ~n653 & ~n813;
  assign n815 = n814 ^ n806;
  assign n816 = x95 & ~n815;
  assign n817 = x143 & n807;
  assign n818 = ~n816 & ~n817;
  assign n819 = ~x129 & ~n818;
  assign n820 = x96 & ~n815;
  assign n821 = x146 & n807;
  assign n822 = ~n820 & ~n821;
  assign n823 = ~x129 & ~n822;
  assign n824 = x97 & ~n815;
  assign n825 = x145 & n807;
  assign n826 = ~n824 & ~n825;
  assign n827 = ~x129 & ~n826;
  assign n828 = ~x145 & n780;
  assign n829 = ~x129 & ~n828;
  assign n830 = ~x98 & ~n780;
  assign n831 = n829 & ~n830;
  assign n832 = ~x141 & n780;
  assign n833 = ~x129 & ~n832;
  assign n834 = ~x99 & ~n780;
  assign n835 = n833 & ~n834;
  assign n836 = x100 & ~n815;
  assign n837 = x144 & n807;
  assign n838 = ~n836 & ~n837;
  assign n839 = ~x129 & ~n838;
  assign n840 = x37 & n779;
  assign n841 = x82 & n723;
  assign n842 = ~n840 & ~n841;
  assign n843 = ~x65 & n655;
  assign n844 = ~x138 & ~n843;
  assign n845 = n842 & n844;
  assign n846 = x93 & n655;
  assign n847 = x138 & ~n846;
  assign n848 = x96 & n723;
  assign n849 = n847 & ~n848;
  assign n850 = ~n845 & ~n849;
  assign n851 = x77 & ~x138;
  assign n852 = n673 & ~n851;
  assign n853 = ~x124 & x138;
  assign n854 = n852 & ~n853;
  assign n855 = ~n850 & ~n854;
  assign n856 = x34 & n779;
  assign n857 = ~x138 & ~n856;
  assign n858 = x79 & n723;
  assign n859 = n857 & ~n858;
  assign n860 = ~x69 & n655;
  assign n861 = ~x66 & n673;
  assign n862 = ~n860 & ~n861;
  assign n863 = n859 & n862;
  assign n864 = x95 & n723;
  assign n865 = x138 & ~n864;
  assign n866 = x91 & n655;
  assign n867 = n865 & ~n866;
  assign n868 = ~n863 & ~n867;
  assign n869 = x33 & n779;
  assign n870 = ~x63 & n655;
  assign n871 = ~n869 & ~n870;
  assign n872 = ~x74 & n673;
  assign n873 = n871 & ~n872;
  assign n874 = x78 & n723;
  assign n875 = ~x138 & ~n874;
  assign n876 = n873 & n875;
  assign n877 = x94 & n723;
  assign n878 = x138 & ~n877;
  assign n879 = x90 & n655;
  assign n880 = n878 & ~n879;
  assign n881 = ~n876 & ~n880;
  assign n882 = ~x73 & n673;
  assign n883 = ~x138 & ~n882;
  assign n884 = ~x68 & n655;
  assign n885 = n883 & ~n884;
  assign n886 = x32 & n779;
  assign n887 = x84 & n723;
  assign n888 = ~n886 & ~n887;
  assign n889 = n885 & n888;
  assign n890 = ~x112 & n723;
  assign n891 = x138 & ~n890;
  assign n892 = x99 & n655;
  assign n893 = n891 & ~n892;
  assign n894 = ~n889 & ~n893;
  assign n900 = x75 & n673;
  assign n901 = ~x80 & n723;
  assign n902 = ~n900 & ~n901;
  assign n903 = x70 & n655;
  assign n904 = ~x35 & n779;
  assign n905 = ~n903 & ~n904;
  assign n906 = n902 & n905;
  assign n895 = x125 & n673;
  assign n896 = x100 & n723;
  assign n897 = ~n895 & ~n896;
  assign n898 = x92 & n655;
  assign n899 = n897 & ~n898;
  assign n907 = n906 ^ n899;
  assign n908 = x138 & ~n907;
  assign n909 = n908 ^ n906;
  assign n910 = ~n386 & ~n418;
  assign n911 = n200 & ~n910;
  assign n912 = x71 ^ x36;
  assign n913 = ~x137 & ~n912;
  assign n914 = n913 ^ x36;
  assign n915 = ~x138 & n914;
  assign n916 = x98 & n749;
  assign n917 = ~n915 & ~n916;
  assign n918 = x136 & ~n917;
  assign n919 = x76 & ~x138;
  assign n920 = n673 & ~n919;
  assign n921 = ~x23 & x138;
  assign n922 = n920 & ~n921;
  assign n923 = ~x97 & x138;
  assign n924 = n723 & ~n923;
  assign n925 = ~x81 & ~x138;
  assign n926 = n924 & ~n925;
  assign n927 = ~n922 & ~n926;
  assign n928 = ~n918 & n927;
  assign n929 = x64 ^ x30;
  assign n930 = ~x137 & ~n929;
  assign n931 = n930 ^ x30;
  assign n932 = ~x138 & n931;
  assign n933 = x88 & n749;
  assign n934 = x136 & ~n933;
  assign n935 = ~n932 & n934;
  assign n936 = x120 & x138;
  assign n937 = n673 & ~n936;
  assign n938 = ~x67 & ~x138;
  assign n939 = n937 & ~n938;
  assign n940 = x111 & x138;
  assign n941 = n723 & ~n940;
  assign n942 = x86 & ~x138;
  assign n943 = n941 & ~n942;
  assign n944 = ~n939 & ~n943;
  assign n945 = ~n935 & n944;
  assign n946 = ~n388 & n416;
  assign n947 = ~n412 & ~n946;
  assign n948 = x116 & n200;
  assign n949 = ~n947 & n948;
  assign n950 = ~x53 & x97;
  assign n951 = x58 ^ x53;
  assign n952 = ~n950 & n951;
  assign n953 = n948 & n952;
  assign n954 = ~x129 & n653;
  assign n955 = ~x111 & ~n806;
  assign n956 = n954 & ~n955;
  assign n957 = ~x139 & n806;
  assign n958 = n956 & ~n957;
  assign n959 = x112 & ~n806;
  assign n960 = n954 & ~n959;
  assign n961 = ~x141 & n806;
  assign n962 = n960 & ~n961;
  assign n963 = ~n208 & n333;
  assign n964 = ~x113 & n258;
  assign n965 = ~n963 & ~n964;
  assign n966 = x115 & ~n806;
  assign n967 = n954 & ~n966;
  assign n968 = ~x140 & n806;
  assign n969 = n967 & ~n968;
  assign n970 = ~n154 & n333;
  assign n971 = x122 & ~x129;
  assign n972 = ~x54 & x118;
  assign n973 = ~n300 & ~n972;
  assign n974 = ~x129 & ~n973;
  assign n975 = ~x129 & ~n382;
  assign n976 = ~x120 & n812;
  assign n977 = ~x111 & ~x129;
  assign n978 = ~n976 & n977;
  assign n979 = x81 & x120;
  assign n980 = ~x129 & n979;
  assign n981 = ~x129 & ~x134;
  assign n982 = ~x129 & ~x135;
  assign n983 = x57 & ~x129;
  assign n984 = ~x96 & x125;
  assign n985 = ~x3 & ~n984;
  assign n986 = ~x129 & ~n985;
  assign n987 = ~x126 & n652;
  assign y0 = x108;
  assign y1 = x83;
  assign y2 = x104;
  assign y3 = x103;
  assign y4 = x102;
  assign y5 = x105;
  assign y6 = x107;
  assign y7 = x101;
  assign y8 = x126;
  assign y9 = x121;
  assign y10 = x1;
  assign y11 = x0;
  assign y12 = ~1'b0;
  assign y13 = x130;
  assign y14 = x128;
  assign y15 = ~n201;
  assign y16 = n215;
  assign y17 = n247;
  assign y18 = ~n254;
  assign y19 = ~n260;
  assign y20 = ~n269;
  assign y21 = ~n273;
  assign y22 = ~n276;
  assign y23 = ~n279;
  assign y24 = ~n285;
  assign y25 = ~n288;
  assign y26 = ~n292;
  assign y27 = ~n296;
  assign y28 = ~n304;
  assign y29 = ~n307;
  assign y30 = n318;
  assign y31 = ~n321;
  assign y32 = ~n327;
  assign y33 = ~n332;
  assign y34 = ~n337;
  assign y35 = n346;
  assign y36 = ~n350;
  assign y37 = ~n353;
  assign y38 = n356;
  assign y39 = n368;
  assign y40 = ~n409;
  assign y41 = ~n415;
  assign y42 = n425;
  assign y43 = n435;
  assign y44 = n451;
  assign y45 = n458;
  assign y46 = n465;
  assign y47 = n472;
  assign y48 = n479;
  assign y49 = n486;
  assign y50 = n493;
  assign y51 = n500;
  assign y52 = n507;
  assign y53 = n515;
  assign y54 = n520;
  assign y55 = n528;
  assign y56 = n537;
  assign y57 = n546;
  assign y58 = n555;
  assign y59 = n561;
  assign y60 = n568;
  assign y61 = n576;
  assign y62 = n585;
  assign y63 = n594;
  assign y64 = n603;
  assign y65 = n615;
  assign y66 = n618;
  assign y67 = n621;
  assign y68 = n448;
  assign y69 = ~n622;
  assign y70 = n624;
  assign y71 = n632;
  assign y72 = n637;
  assign y73 = n640;
  assign y74 = n644;
  assign y75 = n648;
  assign y76 = n651;
  assign y77 = ~n660;
  assign y78 = ~n664;
  assign y79 = ~n668;
  assign y80 = ~n672;
  assign y81 = ~n678;
  assign y82 = ~n682;
  assign y83 = ~n686;
  assign y84 = ~n690;
  assign y85 = ~n694;
  assign y86 = ~n698;
  assign y87 = ~n702;
  assign y88 = ~n706;
  assign y89 = ~n710;
  assign y90 = ~n714;
  assign y91 = ~n718;
  assign y92 = ~n722;
  assign y93 = n728;
  assign y94 = n732;
  assign y95 = n736;
  assign y96 = n740;
  assign y97 = n744;
  assign y98 = n762;
  assign y99 = n766;
  assign y100 = n770;
  assign y101 = n774;
  assign y102 = n778;
  assign y103 = n784;
  assign y104 = n788;
  assign y105 = n792;
  assign y106 = n796;
  assign y107 = n800;
  assign y108 = n804;
  assign y109 = n811;
  assign y110 = n819;
  assign y111 = n823;
  assign y112 = n827;
  assign y113 = n831;
  assign y114 = n835;
  assign y115 = n839;
  assign y116 = ~n855;
  assign y117 = n868;
  assign y118 = n881;
  assign y119 = n894;
  assign y120 = n909;
  assign y121 = n911;
  assign y122 = ~n928;
  assign y123 = n945;
  assign y124 = n949;
  assign y125 = n953;
  assign y126 = n958;
  assign y127 = n962;
  assign y128 = ~n965;
  assign y129 = ~n251;
  assign y130 = n969;
  assign y131 = n970;
  assign y132 = ~n971;
  assign y133 = n974;
  assign y134 = n975;
  assign y135 = n978;
  assign y136 = n980;
  assign y137 = ~n981;
  assign y138 = ~n982;
  assign y139 = n983;
  assign y140 = n986;
  assign y141 = n987;
endmodule
