module top(n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n363);
  input n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63;
  output n363;
  wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362;
  assign n341 = ~n59;
  assign n359 = ~n17;
  assign n349 = ~n28;
  assign n321 = ~n16;
  assign n360 = ~n49;
  assign n355 = ~n51;
  assign n362 = ~n14;
  assign n330 = ~n23;
  assign n358 = ~n1;
  assign n356 = ~n25;
  assign n226 = ~n46;
  assign n346 = ~n29;
  assign n261 = ~n40;
  assign n347 = ~n31;
  assign n342 = ~n34;
  assign n343 = ~n11;
  assign n333 = ~n30;
  assign n326 = ~n63;
  assign n334 = ~n2;
  assign n241 = ~n42;
  assign n246 = ~n58;
  assign n202 = ~n36;
  assign n323 = ~n15;
  assign n322 = ~n33;
  assign n357 = ~n7;
  assign n354 = ~n9;
  assign n340 = ~n12;
  assign n328 = ~n22;
  assign n345 = ~n55;
  assign n324 = ~n13;
  assign n238 = ~n52;
  assign n250 = ~n48;
  assign n167 = ~n44;
  assign n350 = ~n10;
  assign n337 = ~n5;
  assign n253 = ~n54;
  assign n352 = ~n43;
  assign n351 = ~n19;
  assign n200 = ~n37;
  assign n325 = ~n18;
  assign n248 = ~n38;
  assign n222 = ~n62;
  assign n339 = ~n61;
  assign n204 = ~n57;
  assign n224 = ~n60;
  assign n353 = ~n6;
  assign n338 = ~n21;
  assign n344 = ~n20;
  assign n198 = ~n56;
  assign n206 = ~n45;
  assign n336 = ~n26;
  assign n332 = ~n3;
  assign n361 = ~n27;
  assign n335 = ~n47;
  assign n243 = ~n50;
  assign n348 = ~n41;
  assign n275 = ~n0;
  assign n329 = ~n35;
  assign n331 = ~n53;
  assign n327 = ~n39;
  assign n280 = n321 & n48;
  assign n281 = n322 & n1;
  assign n283 = n323 & n47;
  assign n285 = n324 & n45;
  assign n307 = n325 & n50;
  assign n316 = n326 & n31;
  assign n308 = n327 & n7;
  assign n282 = n328 & n54;
  assign n314 = n329 & n3;
  assign n320 = n330 & n55;
  assign n284 = n331 & n21;
  assign n319 = n332 & n35;
  assign n287 = n333 & n62;
  assign n318 = n334 & n34;
  assign n288 = n335 & n15;
  assign n289 = n336 & n58;
  assign n290 = n337 & n37;
  assign n291 = n338 & n53;
  assign n292 = n339 & n29;
  assign n293 = n340 & n44;
  assign n294 = n341 & n27;
  assign n295 = n342 & n2;
  assign n296 = n343 & n43;
  assign n297 = n344 & n52;
  assign n313 = n345 & n23;
  assign n298 = n346 & n61;
  assign n302 = n347 & n63;
  assign n230 = n348 & n9;
  assign n299 = n349 & n60;
  assign n300 = n350 & n42;
  assign n301 = n351 & n51;
  assign n303 = n352 & n11;
  assign n312 = n353 & n38;
  assign n304 = n354 & n41;
  assign n305 = n355 & n19;
  assign n306 = n356 & n57;
  assign n309 = n357 & n39;
  assign n310 = n358 & n33;
  assign n311 = n359 & n49;
  assign n315 = n360 & n17;
  assign n317 = n361 & n59;
  assign n286 = n362 & n46;
  assign n78 = ~n280;
  assign n274 = ~n281;
  assign n277 = ~n282;
  assign n278 = ~n283;
  assign n188 = ~n284;
  assign n239 = ~n285;
  assign n279 = ~n286;
  assign n269 = ~n287;
  assign n139 = ~n288;
  assign n255 = ~n289;
  assign n251 = ~n290;
  assign n256 = ~n291;
  assign n186 = ~n292;
  assign n86 = ~n293;
  assign n141 = ~n294;
  assign n271 = ~n295;
  assign n258 = ~n296;
  assign n257 = ~n297;
  assign n262 = ~n298;
  assign n263 = ~n299;
  assign n259 = ~n300;
  assign n264 = ~n301;
  assign n268 = ~n302;
  assign n157 = ~n303;
  assign n260 = ~n304;
  assign n128 = ~n305;
  assign n244 = ~n306;
  assign n265 = ~n307;
  assign n180 = ~n308;
  assign n266 = ~n309;
  assign n272 = ~n310;
  assign n74 = ~n311;
  assign n267 = ~n312;
  assign n184 = ~n313;
  assign n270 = ~n314;
  assign n182 = ~n315;
  assign n130 = ~n316;
  assign n254 = ~n317;
  assign n273 = ~n318;
  assign n132 = ~n319;
  assign n276 = ~n320;
  assign n235 = n254 & n255;
  assign n227 = n256 & n257;
  assign n229 = n258 & n259;
  assign n231 = n260 & n261;
  assign n228 = n262 & n263;
  assign n76 = n264 & n265;
  assign n233 = n266 & n267;
  assign n148 = n268 & n269;
  assign n146 = n270 & n271;
  assign n191 = n272 & n273;
  assign n234 = n274 & n275;
  assign n150 = n276 & n277;
  assign n236 = n278 & n279;
  assign n237 = n256 & n20;
  assign n240 = n258 & n10;
  assign n242 = n264 & n18;
  assign n232 = n260 & n8;
  assign n247 = n266 & n6;
  assign n249 = n74 & n16;
  assign n221 = n268 & n30;
  assign n223 = n262 & n28;
  assign n252 = n276 & n22;
  assign n245 = n254 & n26;
  assign n225 = n278 & n14;
  assign n208 = n221 & n222;
  assign n209 = n223 & n224;
  assign n210 = n225 & n226;
  assign n72 = n150 & n227;
  assign n113 = n148 & n228;
  assign n211 = n229 & n230;
  assign n207 = n229 & n231;
  assign n212 = n229 & n232;
  assign n199 = n233 & n5;
  assign n213 = n234 & n32;
  assign n203 = n235 & n25;
  assign n205 = n236 & n13;
  assign n214 = n237 & n238;
  assign n84 = n236 & n239;
  assign n215 = n240 & n241;
  assign n216 = n242 & n243;
  assign n197 = n235 & n244;
  assign n217 = n245 & n246;
  assign n218 = n247 & n248;
  assign n219 = n249 & n250;
  assign n201 = n233 & n251;
  assign n220 = n252 & n253;
  assign n168 = n197 & n198;
  assign n189 = n199 & n200;
  assign n169 = n201 & n202;
  assign n192 = n203 & n204;
  assign n193 = n205 & n206;
  assign n166 = n84 & n12;
  assign n194 = n207 & n8;
  assign n195 = n197 & n24;
  assign n196 = n201 & n4;
  assign n119 = ~n208;
  assign n185 = ~n209;
  assign n165 = ~n210;
  assign n175 = ~n211;
  assign n177 = ~n207;
  assign n178 = ~n212;
  assign n190 = ~n213;
  assign n187 = ~n214;
  assign n176 = ~n215;
  assign n116 = ~n216;
  assign n159 = ~n217;
  assign n179 = ~n218;
  assign n181 = ~n219;
  assign n183 = ~n220;
  assign n153 = n166 & n167;
  assign n154 = n168 & n24;
  assign n155 = n169 & n4;
  assign n143 = n175 & n176;
  assign n170 = n177 & n178;
  assign n102 = n179 & n180;
  assign n171 = n181 & n182;
  assign n99 = n183 & n184;
  assign n172 = n185 & n186;
  assign n173 = n187 & n188;
  assign n160 = ~n168;
  assign n107 = ~n189;
  assign n162 = ~n169;
  assign n174 = n190 & n191;
  assign n158 = ~n192;
  assign n164 = ~n193;
  assign n156 = ~n194;
  assign n161 = ~n195;
  assign n163 = ~n196;
  assign n138 = ~n153;
  assign n140 = ~n154;
  assign n111 = ~n155;
  assign n142 = n156 & n157;
  assign n124 = n158 & n159;
  assign n151 = n160 & n161;
  assign n152 = n162 & n163;
  assign n126 = n164 & n165;
  assign n96 = ~n170;
  assign n144 = ~n171;
  assign n147 = ~n172;
  assign n149 = ~n173;
  assign n145 = ~n174;
  assign n125 = n138 & n139;
  assign n123 = n140 & n141;
  assign n91 = n142 & n143;
  assign n134 = n144 & n76;
  assign n135 = n145 & n146;
  assign n136 = n147 & n148;
  assign n137 = n149 & n150;
  assign n133 = ~n151;
  assign n131 = ~n152;
  assign n122 = n123 & n124;
  assign n81 = n125 & n126;
  assign n120 = n131 & n132;
  assign n70 = n133 & n113;
  assign n127 = ~n134;
  assign n121 = ~n135;
  assign n129 = ~n136;
  assign n104 = ~n137;
  assign n117 = n120 & n121;
  assign n112 = ~n122;
  assign n115 = n127 & n128;
  assign n118 = n129 & n130;
  assign n109 = n112 & n113;
  assign n114 = n115 & n116;
  assign n110 = ~n117;
  assign n67 = n118 & n119;
  assign n88 = ~n109;
  assign n106 = n110 & n111;
  assign n108 = ~n114;
  assign n101 = n106 & n107;
  assign n105 = n108 & n72;
  assign n100 = n101 & n102;
  assign n103 = ~n105;
  assign n95 = ~n100;
  assign n98 = n103 & n104;
  assign n94 = n95 & n96;
  assign n97 = n98 & n99;
  assign n90 = ~n94;
  assign n93 = ~n97;
  assign n89 = n90 & n91;
  assign n92 = n93 & n70;
  assign n85 = ~n89;
  assign n87 = ~n92;
  assign n83 = n85 & n86;
  assign n65 = n87 & n88;
  assign n82 = n83 & n84;
  assign n80 = ~n82;
  assign n79 = n80 & n81;
  assign n77 = ~n79;
  assign n75 = n77 & n78;
  assign n73 = n75 & n76;
  assign n71 = n73 & n74;
  assign n69 = n71 & n72;
  assign n68 = n69 & n70;
  assign n66 = ~n68;
  assign n64 = n66 & n67;
  assign n363 = n64 & n65;
endmodule
