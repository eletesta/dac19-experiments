module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127;
  wire n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759;
  assign n496 = x64 ^ x62;
  assign n497 = ~x129 & n496;
  assign n498 = n497 ^ x62;
  assign n493 = x63 ^ x61;
  assign n494 = ~x129 & n493;
  assign n495 = n494 ^ x61;
  assign n499 = n498 ^ n495;
  assign n500 = x128 & n499;
  assign n501 = n500 ^ n498;
  assign n487 = x56 ^ x54;
  assign n488 = ~x129 & n487;
  assign n489 = n488 ^ x54;
  assign n484 = x55 ^ x53;
  assign n485 = ~x129 & n484;
  assign n486 = n485 ^ x53;
  assign n490 = n489 ^ n486;
  assign n491 = x128 & n490;
  assign n492 = n491 ^ n489;
  assign n502 = n501 ^ n492;
  assign n503 = x131 & n502;
  assign n504 = n503 ^ n501;
  assign n475 = x60 ^ x58;
  assign n476 = ~x129 & n475;
  assign n477 = n476 ^ x58;
  assign n472 = x59 ^ x57;
  assign n473 = ~x129 & n472;
  assign n474 = n473 ^ x57;
  assign n478 = n477 ^ n474;
  assign n479 = x128 & n478;
  assign n480 = n479 ^ n477;
  assign n466 = x52 ^ x50;
  assign n467 = ~x129 & n466;
  assign n468 = n467 ^ x50;
  assign n463 = x51 ^ x49;
  assign n464 = ~x129 & n463;
  assign n465 = n464 ^ x49;
  assign n469 = n468 ^ n465;
  assign n470 = x128 & n469;
  assign n471 = n470 ^ n468;
  assign n481 = n480 ^ n471;
  assign n482 = x131 & n481;
  assign n483 = n482 ^ n480;
  assign n505 = n504 ^ n483;
  assign n506 = x130 & n505;
  assign n507 = n506 ^ n504;
  assign n451 = x32 ^ x30;
  assign n452 = ~x129 & n451;
  assign n453 = n452 ^ x30;
  assign n448 = x31 ^ x29;
  assign n449 = ~x129 & n448;
  assign n450 = n449 ^ x29;
  assign n454 = n453 ^ n450;
  assign n455 = x128 & n454;
  assign n456 = n455 ^ n453;
  assign n442 = x24 ^ x22;
  assign n443 = ~x129 & n442;
  assign n444 = n443 ^ x22;
  assign n439 = x23 ^ x21;
  assign n440 = ~x129 & n439;
  assign n441 = n440 ^ x21;
  assign n445 = n444 ^ n441;
  assign n446 = x128 & n445;
  assign n447 = n446 ^ n444;
  assign n457 = n456 ^ n447;
  assign n458 = x131 & n457;
  assign n459 = n458 ^ n456;
  assign n430 = x28 ^ x26;
  assign n431 = ~x129 & n430;
  assign n432 = n431 ^ x26;
  assign n427 = x27 ^ x25;
  assign n428 = ~x129 & n427;
  assign n429 = n428 ^ x25;
  assign n433 = n432 ^ n429;
  assign n434 = x128 & n433;
  assign n435 = n434 ^ n432;
  assign n421 = x20 ^ x18;
  assign n422 = ~x129 & n421;
  assign n423 = n422 ^ x18;
  assign n418 = x19 ^ x17;
  assign n419 = ~x129 & n418;
  assign n420 = n419 ^ x17;
  assign n424 = n423 ^ n420;
  assign n425 = x128 & n424;
  assign n426 = n425 ^ n423;
  assign n436 = n435 ^ n426;
  assign n437 = x131 & n436;
  assign n438 = n437 ^ n435;
  assign n460 = n459 ^ n438;
  assign n461 = x130 & n460;
  assign n462 = n461 ^ n459;
  assign n508 = n507 ^ n462;
  assign n509 = x133 & n508;
  assign n510 = n509 ^ n507;
  assign n403 = x48 ^ x46;
  assign n404 = ~x129 & n403;
  assign n405 = n404 ^ x46;
  assign n400 = x47 ^ x45;
  assign n401 = ~x129 & n400;
  assign n402 = n401 ^ x45;
  assign n406 = n405 ^ n402;
  assign n407 = x128 & n406;
  assign n408 = n407 ^ n405;
  assign n394 = x40 ^ x38;
  assign n395 = ~x129 & n394;
  assign n396 = n395 ^ x38;
  assign n391 = x39 ^ x37;
  assign n392 = ~x129 & n391;
  assign n393 = n392 ^ x37;
  assign n397 = n396 ^ n393;
  assign n398 = x128 & n397;
  assign n399 = n398 ^ n396;
  assign n409 = n408 ^ n399;
  assign n410 = x131 & n409;
  assign n411 = n410 ^ n408;
  assign n382 = x44 ^ x42;
  assign n383 = ~x129 & n382;
  assign n384 = n383 ^ x42;
  assign n379 = x43 ^ x41;
  assign n380 = ~x129 & n379;
  assign n381 = n380 ^ x41;
  assign n385 = n384 ^ n381;
  assign n386 = x128 & n385;
  assign n387 = n386 ^ n384;
  assign n373 = x36 ^ x34;
  assign n374 = ~x129 & n373;
  assign n375 = n374 ^ x34;
  assign n370 = x35 ^ x33;
  assign n371 = ~x129 & n370;
  assign n372 = n371 ^ x33;
  assign n376 = n375 ^ n372;
  assign n377 = x128 & n376;
  assign n378 = n377 ^ n375;
  assign n388 = n387 ^ n378;
  assign n389 = x131 & n388;
  assign n390 = n389 ^ n387;
  assign n412 = n411 ^ n390;
  assign n413 = x130 & n412;
  assign n414 = n413 ^ n411;
  assign n358 = x16 ^ x14;
  assign n359 = ~x129 & n358;
  assign n360 = n359 ^ x14;
  assign n355 = x15 ^ x13;
  assign n356 = ~x129 & n355;
  assign n357 = n356 ^ x13;
  assign n361 = n360 ^ n357;
  assign n362 = x128 & n361;
  assign n363 = n362 ^ n360;
  assign n349 = x8 ^ x6;
  assign n350 = ~x129 & n349;
  assign n351 = n350 ^ x6;
  assign n346 = x7 ^ x5;
  assign n347 = ~x129 & n346;
  assign n348 = n347 ^ x5;
  assign n352 = n351 ^ n348;
  assign n353 = x128 & n352;
  assign n354 = n353 ^ n351;
  assign n364 = n363 ^ n354;
  assign n365 = x131 & n364;
  assign n366 = n365 ^ n363;
  assign n337 = x12 ^ x10;
  assign n338 = ~x129 & n337;
  assign n339 = n338 ^ x10;
  assign n334 = x11 ^ x9;
  assign n335 = ~x129 & n334;
  assign n336 = n335 ^ x9;
  assign n340 = n339 ^ n336;
  assign n341 = x128 & n340;
  assign n342 = n341 ^ n339;
  assign n328 = x4 ^ x2;
  assign n329 = ~x129 & n328;
  assign n330 = n329 ^ x2;
  assign n325 = x3 ^ x1;
  assign n326 = ~x129 & n325;
  assign n327 = n326 ^ x1;
  assign n331 = n330 ^ n327;
  assign n332 = x128 & n331;
  assign n333 = n332 ^ n330;
  assign n343 = n342 ^ n333;
  assign n344 = x131 & n343;
  assign n345 = n344 ^ n342;
  assign n367 = n366 ^ n345;
  assign n368 = x130 & n367;
  assign n369 = n368 ^ n366;
  assign n415 = n414 ^ n369;
  assign n416 = x133 & n415;
  assign n417 = n416 ^ n414;
  assign n511 = n510 ^ n417;
  assign n512 = x132 & n511;
  assign n513 = n512 ^ n510;
  assign n307 = x126 ^ x0;
  assign n308 = x129 & n307;
  assign n309 = n308 ^ x0;
  assign n304 = x127 ^ x125;
  assign n305 = ~x129 & n304;
  assign n306 = n305 ^ x125;
  assign n310 = n309 ^ n306;
  assign n311 = x128 & n310;
  assign n312 = n311 ^ n309;
  assign n298 = x120 ^ x118;
  assign n299 = ~x129 & n298;
  assign n300 = n299 ^ x118;
  assign n295 = x119 ^ x117;
  assign n296 = ~x129 & n295;
  assign n297 = n296 ^ x117;
  assign n301 = n300 ^ n297;
  assign n302 = x128 & n301;
  assign n303 = n302 ^ n300;
  assign n313 = n312 ^ n303;
  assign n314 = x131 & n313;
  assign n315 = n314 ^ n312;
  assign n286 = x124 ^ x122;
  assign n287 = ~x129 & n286;
  assign n288 = n287 ^ x122;
  assign n283 = x123 ^ x121;
  assign n284 = ~x129 & n283;
  assign n285 = n284 ^ x121;
  assign n289 = n288 ^ n285;
  assign n290 = x128 & n289;
  assign n291 = n290 ^ n288;
  assign n277 = x116 ^ x114;
  assign n278 = ~x129 & n277;
  assign n279 = n278 ^ x114;
  assign n274 = x115 ^ x113;
  assign n275 = ~x129 & n274;
  assign n276 = n275 ^ x113;
  assign n280 = n279 ^ n276;
  assign n281 = x128 & n280;
  assign n282 = n281 ^ n279;
  assign n292 = n291 ^ n282;
  assign n293 = x131 & n292;
  assign n294 = n293 ^ n291;
  assign n316 = n315 ^ n294;
  assign n317 = x130 & n316;
  assign n318 = n317 ^ n315;
  assign n262 = x96 ^ x94;
  assign n263 = ~x129 & n262;
  assign n264 = n263 ^ x94;
  assign n259 = x95 ^ x93;
  assign n260 = ~x129 & n259;
  assign n261 = n260 ^ x93;
  assign n265 = n264 ^ n261;
  assign n266 = x128 & n265;
  assign n267 = n266 ^ n264;
  assign n253 = x88 ^ x86;
  assign n254 = ~x129 & n253;
  assign n255 = n254 ^ x86;
  assign n250 = x87 ^ x85;
  assign n251 = ~x129 & n250;
  assign n252 = n251 ^ x85;
  assign n256 = n255 ^ n252;
  assign n257 = x128 & n256;
  assign n258 = n257 ^ n255;
  assign n268 = n267 ^ n258;
  assign n269 = x131 & n268;
  assign n270 = n269 ^ n267;
  assign n241 = x92 ^ x90;
  assign n242 = ~x129 & n241;
  assign n243 = n242 ^ x90;
  assign n238 = x91 ^ x89;
  assign n239 = ~x129 & n238;
  assign n240 = n239 ^ x89;
  assign n244 = n243 ^ n240;
  assign n245 = x128 & n244;
  assign n246 = n245 ^ n243;
  assign n232 = x84 ^ x82;
  assign n233 = ~x129 & n232;
  assign n234 = n233 ^ x82;
  assign n229 = x83 ^ x81;
  assign n230 = ~x129 & n229;
  assign n231 = n230 ^ x81;
  assign n235 = n234 ^ n231;
  assign n236 = x128 & n235;
  assign n237 = n236 ^ n234;
  assign n247 = n246 ^ n237;
  assign n248 = x131 & n247;
  assign n249 = n248 ^ n246;
  assign n271 = n270 ^ n249;
  assign n272 = x130 & n271;
  assign n273 = n272 ^ n270;
  assign n319 = n318 ^ n273;
  assign n320 = x133 & n319;
  assign n321 = n320 ^ n318;
  assign n214 = x112 ^ x110;
  assign n215 = ~x129 & n214;
  assign n216 = n215 ^ x110;
  assign n211 = x111 ^ x109;
  assign n212 = ~x129 & n211;
  assign n213 = n212 ^ x109;
  assign n217 = n216 ^ n213;
  assign n218 = x128 & n217;
  assign n219 = n218 ^ n216;
  assign n205 = x104 ^ x102;
  assign n206 = ~x129 & n205;
  assign n207 = n206 ^ x102;
  assign n202 = x103 ^ x101;
  assign n203 = ~x129 & n202;
  assign n204 = n203 ^ x101;
  assign n208 = n207 ^ n204;
  assign n209 = x128 & n208;
  assign n210 = n209 ^ n207;
  assign n220 = n219 ^ n210;
  assign n221 = x131 & n220;
  assign n222 = n221 ^ n219;
  assign n193 = x108 ^ x106;
  assign n194 = ~x129 & n193;
  assign n195 = n194 ^ x106;
  assign n190 = x107 ^ x105;
  assign n191 = ~x129 & n190;
  assign n192 = n191 ^ x105;
  assign n196 = n195 ^ n192;
  assign n197 = x128 & n196;
  assign n198 = n197 ^ n195;
  assign n184 = x100 ^ x98;
  assign n185 = ~x129 & n184;
  assign n186 = n185 ^ x98;
  assign n181 = x99 ^ x97;
  assign n182 = ~x129 & n181;
  assign n183 = n182 ^ x97;
  assign n187 = n186 ^ n183;
  assign n188 = x128 & n187;
  assign n189 = n188 ^ n186;
  assign n199 = n198 ^ n189;
  assign n200 = x131 & n199;
  assign n201 = n200 ^ n198;
  assign n223 = n222 ^ n201;
  assign n224 = x130 & n223;
  assign n225 = n224 ^ n222;
  assign n169 = x80 ^ x78;
  assign n170 = ~x129 & n169;
  assign n171 = n170 ^ x78;
  assign n166 = x79 ^ x77;
  assign n167 = ~x129 & n166;
  assign n168 = n167 ^ x77;
  assign n172 = n171 ^ n168;
  assign n173 = x128 & n172;
  assign n174 = n173 ^ n171;
  assign n160 = x72 ^ x70;
  assign n161 = ~x129 & n160;
  assign n162 = n161 ^ x70;
  assign n157 = x71 ^ x69;
  assign n158 = ~x129 & n157;
  assign n159 = n158 ^ x69;
  assign n163 = n162 ^ n159;
  assign n164 = x128 & n163;
  assign n165 = n164 ^ n162;
  assign n175 = n174 ^ n165;
  assign n176 = x131 & n175;
  assign n177 = n176 ^ n174;
  assign n148 = x76 ^ x74;
  assign n149 = ~x129 & n148;
  assign n150 = n149 ^ x74;
  assign n145 = x75 ^ x73;
  assign n146 = ~x129 & n145;
  assign n147 = n146 ^ x73;
  assign n151 = n150 ^ n147;
  assign n152 = x128 & n151;
  assign n153 = n152 ^ n150;
  assign n139 = x68 ^ x66;
  assign n140 = ~x129 & n139;
  assign n141 = n140 ^ x66;
  assign n136 = x67 ^ x65;
  assign n137 = ~x129 & n136;
  assign n138 = n137 ^ x65;
  assign n142 = n141 ^ n138;
  assign n143 = x128 & n142;
  assign n144 = n143 ^ n141;
  assign n154 = n153 ^ n144;
  assign n155 = x131 & n154;
  assign n156 = n155 ^ n153;
  assign n178 = n177 ^ n156;
  assign n179 = x130 & n178;
  assign n180 = n179 ^ n177;
  assign n226 = n225 ^ n180;
  assign n227 = x133 & n226;
  assign n228 = n227 ^ n225;
  assign n322 = n321 ^ n228;
  assign n323 = x132 & n322;
  assign n324 = n323 ^ n321;
  assign n514 = n513 ^ n324;
  assign n515 = ~x134 & n514;
  assign n516 = n515 ^ n513;
  assign n781 = x65 ^ x63;
  assign n782 = ~x129 & n781;
  assign n783 = n782 ^ x63;
  assign n784 = n783 ^ n498;
  assign n785 = ~x128 & n784;
  assign n786 = n785 ^ n498;
  assign n775 = x57 ^ x55;
  assign n776 = ~x129 & n775;
  assign n777 = n776 ^ x55;
  assign n778 = n777 ^ n489;
  assign n779 = ~x128 & n778;
  assign n780 = n779 ^ n489;
  assign n787 = n786 ^ n780;
  assign n788 = x131 & n787;
  assign n789 = n788 ^ n786;
  assign n766 = x61 ^ x59;
  assign n767 = ~x129 & n766;
  assign n768 = n767 ^ x59;
  assign n769 = n768 ^ n477;
  assign n770 = ~x128 & n769;
  assign n771 = n770 ^ n477;
  assign n760 = x53 ^ x51;
  assign n761 = ~x129 & n760;
  assign n762 = n761 ^ x51;
  assign n763 = n762 ^ n468;
  assign n764 = ~x128 & n763;
  assign n765 = n764 ^ n468;
  assign n772 = n771 ^ n765;
  assign n773 = x131 & n772;
  assign n774 = n773 ^ n771;
  assign n790 = n789 ^ n774;
  assign n791 = x130 & n790;
  assign n792 = n791 ^ n789;
  assign n748 = x33 ^ x31;
  assign n749 = ~x129 & n748;
  assign n750 = n749 ^ x31;
  assign n751 = n750 ^ n453;
  assign n752 = ~x128 & n751;
  assign n753 = n752 ^ n453;
  assign n742 = x25 ^ x23;
  assign n743 = ~x129 & n742;
  assign n744 = n743 ^ x23;
  assign n745 = n744 ^ n444;
  assign n746 = ~x128 & n745;
  assign n747 = n746 ^ n444;
  assign n754 = n753 ^ n747;
  assign n755 = x131 & n754;
  assign n756 = n755 ^ n753;
  assign n733 = x29 ^ x27;
  assign n734 = ~x129 & n733;
  assign n735 = n734 ^ x27;
  assign n736 = n735 ^ n432;
  assign n737 = ~x128 & n736;
  assign n738 = n737 ^ n432;
  assign n727 = x21 ^ x19;
  assign n728 = ~x129 & n727;
  assign n729 = n728 ^ x19;
  assign n730 = n729 ^ n423;
  assign n731 = ~x128 & n730;
  assign n732 = n731 ^ n423;
  assign n739 = n738 ^ n732;
  assign n740 = x131 & n739;
  assign n741 = n740 ^ n738;
  assign n757 = n756 ^ n741;
  assign n758 = x130 & n757;
  assign n759 = n758 ^ n756;
  assign n793 = n792 ^ n759;
  assign n794 = x133 & n793;
  assign n795 = n794 ^ n792;
  assign n712 = x49 ^ x47;
  assign n713 = ~x129 & n712;
  assign n714 = n713 ^ x47;
  assign n715 = n714 ^ n405;
  assign n716 = ~x128 & n715;
  assign n717 = n716 ^ n405;
  assign n706 = x41 ^ x39;
  assign n707 = ~x129 & n706;
  assign n708 = n707 ^ x39;
  assign n709 = n708 ^ n396;
  assign n710 = ~x128 & n709;
  assign n711 = n710 ^ n396;
  assign n718 = n717 ^ n711;
  assign n719 = x131 & n718;
  assign n720 = n719 ^ n717;
  assign n697 = x45 ^ x43;
  assign n698 = ~x129 & n697;
  assign n699 = n698 ^ x43;
  assign n700 = n699 ^ n384;
  assign n701 = ~x128 & n700;
  assign n702 = n701 ^ n384;
  assign n691 = x37 ^ x35;
  assign n692 = ~x129 & n691;
  assign n693 = n692 ^ x35;
  assign n694 = n693 ^ n375;
  assign n695 = ~x128 & n694;
  assign n696 = n695 ^ n375;
  assign n703 = n702 ^ n696;
  assign n704 = x131 & n703;
  assign n705 = n704 ^ n702;
  assign n721 = n720 ^ n705;
  assign n722 = x130 & n721;
  assign n723 = n722 ^ n720;
  assign n679 = x17 ^ x15;
  assign n680 = ~x129 & n679;
  assign n681 = n680 ^ x15;
  assign n682 = n681 ^ n360;
  assign n683 = ~x128 & n682;
  assign n684 = n683 ^ n360;
  assign n673 = x9 ^ x7;
  assign n674 = ~x129 & n673;
  assign n675 = n674 ^ x7;
  assign n676 = n675 ^ n351;
  assign n677 = ~x128 & n676;
  assign n678 = n677 ^ n351;
  assign n685 = n684 ^ n678;
  assign n686 = x131 & n685;
  assign n687 = n686 ^ n684;
  assign n664 = x13 ^ x11;
  assign n665 = ~x129 & n664;
  assign n666 = n665 ^ x11;
  assign n667 = n666 ^ n339;
  assign n668 = ~x128 & n667;
  assign n669 = n668 ^ n339;
  assign n658 = x5 ^ x3;
  assign n659 = ~x129 & n658;
  assign n660 = n659 ^ x3;
  assign n661 = n660 ^ n330;
  assign n662 = ~x128 & n661;
  assign n663 = n662 ^ n330;
  assign n670 = n669 ^ n663;
  assign n671 = x131 & n670;
  assign n672 = n671 ^ n669;
  assign n688 = n687 ^ n672;
  assign n689 = x130 & n688;
  assign n690 = n689 ^ n687;
  assign n724 = n723 ^ n690;
  assign n725 = x133 & n724;
  assign n726 = n725 ^ n723;
  assign n796 = n795 ^ n726;
  assign n797 = x132 & n796;
  assign n798 = n797 ^ n795;
  assign n640 = x127 ^ x1;
  assign n641 = x129 & n640;
  assign n642 = n641 ^ x1;
  assign n643 = n642 ^ n309;
  assign n644 = ~x128 & n643;
  assign n645 = n644 ^ n309;
  assign n634 = x121 ^ x119;
  assign n635 = ~x129 & n634;
  assign n636 = n635 ^ x119;
  assign n637 = n636 ^ n300;
  assign n638 = ~x128 & n637;
  assign n639 = n638 ^ n300;
  assign n646 = n645 ^ n639;
  assign n647 = x131 & n646;
  assign n648 = n647 ^ n645;
  assign n625 = x125 ^ x123;
  assign n626 = ~x129 & n625;
  assign n627 = n626 ^ x123;
  assign n628 = n627 ^ n288;
  assign n629 = ~x128 & n628;
  assign n630 = n629 ^ n288;
  assign n619 = x117 ^ x115;
  assign n620 = ~x129 & n619;
  assign n621 = n620 ^ x115;
  assign n622 = n621 ^ n279;
  assign n623 = ~x128 & n622;
  assign n624 = n623 ^ n279;
  assign n631 = n630 ^ n624;
  assign n632 = x131 & n631;
  assign n633 = n632 ^ n630;
  assign n649 = n648 ^ n633;
  assign n650 = x130 & n649;
  assign n651 = n650 ^ n648;
  assign n607 = x97 ^ x95;
  assign n608 = ~x129 & n607;
  assign n609 = n608 ^ x95;
  assign n610 = n609 ^ n264;
  assign n611 = ~x128 & n610;
  assign n612 = n611 ^ n264;
  assign n601 = x89 ^ x87;
  assign n602 = ~x129 & n601;
  assign n603 = n602 ^ x87;
  assign n604 = n603 ^ n255;
  assign n605 = ~x128 & n604;
  assign n606 = n605 ^ n255;
  assign n613 = n612 ^ n606;
  assign n614 = x131 & n613;
  assign n615 = n614 ^ n612;
  assign n592 = x93 ^ x91;
  assign n593 = ~x129 & n592;
  assign n594 = n593 ^ x91;
  assign n595 = n594 ^ n243;
  assign n596 = ~x128 & n595;
  assign n597 = n596 ^ n243;
  assign n586 = x85 ^ x83;
  assign n587 = ~x129 & n586;
  assign n588 = n587 ^ x83;
  assign n589 = n588 ^ n234;
  assign n590 = ~x128 & n589;
  assign n591 = n590 ^ n234;
  assign n598 = n597 ^ n591;
  assign n599 = x131 & n598;
  assign n600 = n599 ^ n597;
  assign n616 = n615 ^ n600;
  assign n617 = x130 & n616;
  assign n618 = n617 ^ n615;
  assign n652 = n651 ^ n618;
  assign n653 = x133 & n652;
  assign n654 = n653 ^ n651;
  assign n571 = x113 ^ x111;
  assign n572 = ~x129 & n571;
  assign n573 = n572 ^ x111;
  assign n574 = n573 ^ n216;
  assign n575 = ~x128 & n574;
  assign n576 = n575 ^ n216;
  assign n565 = x105 ^ x103;
  assign n566 = ~x129 & n565;
  assign n567 = n566 ^ x103;
  assign n568 = n567 ^ n207;
  assign n569 = ~x128 & n568;
  assign n570 = n569 ^ n207;
  assign n577 = n576 ^ n570;
  assign n578 = x131 & n577;
  assign n579 = n578 ^ n576;
  assign n556 = x109 ^ x107;
  assign n557 = ~x129 & n556;
  assign n558 = n557 ^ x107;
  assign n559 = n558 ^ n195;
  assign n560 = ~x128 & n559;
  assign n561 = n560 ^ n195;
  assign n550 = x101 ^ x99;
  assign n551 = ~x129 & n550;
  assign n552 = n551 ^ x99;
  assign n553 = n552 ^ n186;
  assign n554 = ~x128 & n553;
  assign n555 = n554 ^ n186;
  assign n562 = n561 ^ n555;
  assign n563 = x131 & n562;
  assign n564 = n563 ^ n561;
  assign n580 = n579 ^ n564;
  assign n581 = x130 & n580;
  assign n582 = n581 ^ n579;
  assign n538 = x81 ^ x79;
  assign n539 = ~x129 & n538;
  assign n540 = n539 ^ x79;
  assign n541 = n540 ^ n171;
  assign n542 = ~x128 & n541;
  assign n543 = n542 ^ n171;
  assign n532 = x73 ^ x71;
  assign n533 = ~x129 & n532;
  assign n534 = n533 ^ x71;
  assign n535 = n534 ^ n162;
  assign n536 = ~x128 & n535;
  assign n537 = n536 ^ n162;
  assign n544 = n543 ^ n537;
  assign n545 = x131 & n544;
  assign n546 = n545 ^ n543;
  assign n523 = x77 ^ x75;
  assign n524 = ~x129 & n523;
  assign n525 = n524 ^ x75;
  assign n526 = n525 ^ n150;
  assign n527 = ~x128 & n526;
  assign n528 = n527 ^ n150;
  assign n517 = x69 ^ x67;
  assign n518 = ~x129 & n517;
  assign n519 = n518 ^ x67;
  assign n520 = n519 ^ n141;
  assign n521 = ~x128 & n520;
  assign n522 = n521 ^ n141;
  assign n529 = n528 ^ n522;
  assign n530 = x131 & n529;
  assign n531 = n530 ^ n528;
  assign n547 = n546 ^ n531;
  assign n548 = x130 & n547;
  assign n549 = n548 ^ n546;
  assign n583 = n582 ^ n549;
  assign n584 = x133 & n583;
  assign n585 = n584 ^ n582;
  assign n655 = n654 ^ n585;
  assign n656 = x132 & n655;
  assign n657 = n656 ^ n654;
  assign n799 = n798 ^ n657;
  assign n800 = ~x134 & n799;
  assign n801 = n800 ^ n798;
  assign n1066 = x66 ^ x64;
  assign n1067 = ~x129 & n1066;
  assign n1068 = n1067 ^ x64;
  assign n1069 = n1068 ^ n783;
  assign n1070 = ~x128 & n1069;
  assign n1071 = n1070 ^ n783;
  assign n1060 = x58 ^ x56;
  assign n1061 = ~x129 & n1060;
  assign n1062 = n1061 ^ x56;
  assign n1063 = n1062 ^ n777;
  assign n1064 = ~x128 & n1063;
  assign n1065 = n1064 ^ n777;
  assign n1072 = n1071 ^ n1065;
  assign n1073 = x131 & n1072;
  assign n1074 = n1073 ^ n1071;
  assign n1051 = x62 ^ x60;
  assign n1052 = ~x129 & n1051;
  assign n1053 = n1052 ^ x60;
  assign n1054 = n1053 ^ n768;
  assign n1055 = ~x128 & n1054;
  assign n1056 = n1055 ^ n768;
  assign n1045 = x54 ^ x52;
  assign n1046 = ~x129 & n1045;
  assign n1047 = n1046 ^ x52;
  assign n1048 = n1047 ^ n762;
  assign n1049 = ~x128 & n1048;
  assign n1050 = n1049 ^ n762;
  assign n1057 = n1056 ^ n1050;
  assign n1058 = x131 & n1057;
  assign n1059 = n1058 ^ n1056;
  assign n1075 = n1074 ^ n1059;
  assign n1076 = x130 & n1075;
  assign n1077 = n1076 ^ n1074;
  assign n1033 = x34 ^ x32;
  assign n1034 = ~x129 & n1033;
  assign n1035 = n1034 ^ x32;
  assign n1036 = n1035 ^ n750;
  assign n1037 = ~x128 & n1036;
  assign n1038 = n1037 ^ n750;
  assign n1027 = x26 ^ x24;
  assign n1028 = ~x129 & n1027;
  assign n1029 = n1028 ^ x24;
  assign n1030 = n1029 ^ n744;
  assign n1031 = ~x128 & n1030;
  assign n1032 = n1031 ^ n744;
  assign n1039 = n1038 ^ n1032;
  assign n1040 = x131 & n1039;
  assign n1041 = n1040 ^ n1038;
  assign n1018 = x30 ^ x28;
  assign n1019 = ~x129 & n1018;
  assign n1020 = n1019 ^ x28;
  assign n1021 = n1020 ^ n735;
  assign n1022 = ~x128 & n1021;
  assign n1023 = n1022 ^ n735;
  assign n1012 = x22 ^ x20;
  assign n1013 = ~x129 & n1012;
  assign n1014 = n1013 ^ x20;
  assign n1015 = n1014 ^ n729;
  assign n1016 = ~x128 & n1015;
  assign n1017 = n1016 ^ n729;
  assign n1024 = n1023 ^ n1017;
  assign n1025 = x131 & n1024;
  assign n1026 = n1025 ^ n1023;
  assign n1042 = n1041 ^ n1026;
  assign n1043 = x130 & n1042;
  assign n1044 = n1043 ^ n1041;
  assign n1078 = n1077 ^ n1044;
  assign n1079 = x133 & n1078;
  assign n1080 = n1079 ^ n1077;
  assign n997 = x50 ^ x48;
  assign n998 = ~x129 & n997;
  assign n999 = n998 ^ x48;
  assign n1000 = n999 ^ n714;
  assign n1001 = ~x128 & n1000;
  assign n1002 = n1001 ^ n714;
  assign n991 = x42 ^ x40;
  assign n992 = ~x129 & n991;
  assign n993 = n992 ^ x40;
  assign n994 = n993 ^ n708;
  assign n995 = ~x128 & n994;
  assign n996 = n995 ^ n708;
  assign n1003 = n1002 ^ n996;
  assign n1004 = x131 & n1003;
  assign n1005 = n1004 ^ n1002;
  assign n982 = x46 ^ x44;
  assign n983 = ~x129 & n982;
  assign n984 = n983 ^ x44;
  assign n985 = n984 ^ n699;
  assign n986 = ~x128 & n985;
  assign n987 = n986 ^ n699;
  assign n976 = x38 ^ x36;
  assign n977 = ~x129 & n976;
  assign n978 = n977 ^ x36;
  assign n979 = n978 ^ n693;
  assign n980 = ~x128 & n979;
  assign n981 = n980 ^ n693;
  assign n988 = n987 ^ n981;
  assign n989 = x131 & n988;
  assign n990 = n989 ^ n987;
  assign n1006 = n1005 ^ n990;
  assign n1007 = x130 & n1006;
  assign n1008 = n1007 ^ n1005;
  assign n964 = x18 ^ x16;
  assign n965 = ~x129 & n964;
  assign n966 = n965 ^ x16;
  assign n967 = n966 ^ n681;
  assign n968 = ~x128 & n967;
  assign n969 = n968 ^ n681;
  assign n958 = x10 ^ x8;
  assign n959 = ~x129 & n958;
  assign n960 = n959 ^ x8;
  assign n961 = n960 ^ n675;
  assign n962 = ~x128 & n961;
  assign n963 = n962 ^ n675;
  assign n970 = n969 ^ n963;
  assign n971 = x131 & n970;
  assign n972 = n971 ^ n969;
  assign n949 = x14 ^ x12;
  assign n950 = ~x129 & n949;
  assign n951 = n950 ^ x12;
  assign n952 = n951 ^ n666;
  assign n953 = ~x128 & n952;
  assign n954 = n953 ^ n666;
  assign n943 = x6 ^ x4;
  assign n944 = ~x129 & n943;
  assign n945 = n944 ^ x4;
  assign n946 = n945 ^ n660;
  assign n947 = ~x128 & n946;
  assign n948 = n947 ^ n660;
  assign n955 = n954 ^ n948;
  assign n956 = x131 & n955;
  assign n957 = n956 ^ n954;
  assign n973 = n972 ^ n957;
  assign n974 = x130 & n973;
  assign n975 = n974 ^ n972;
  assign n1009 = n1008 ^ n975;
  assign n1010 = x133 & n1009;
  assign n1011 = n1010 ^ n1008;
  assign n1081 = n1080 ^ n1011;
  assign n1082 = x132 & n1081;
  assign n1083 = n1082 ^ n1080;
  assign n925 = x2 ^ x0;
  assign n926 = ~x129 & n925;
  assign n927 = n926 ^ x0;
  assign n928 = n927 ^ n642;
  assign n929 = ~x128 & n928;
  assign n930 = n929 ^ n642;
  assign n919 = x122 ^ x120;
  assign n920 = ~x129 & n919;
  assign n921 = n920 ^ x120;
  assign n922 = n921 ^ n636;
  assign n923 = ~x128 & n922;
  assign n924 = n923 ^ n636;
  assign n931 = n930 ^ n924;
  assign n932 = x131 & n931;
  assign n933 = n932 ^ n930;
  assign n910 = x126 ^ x124;
  assign n911 = ~x129 & n910;
  assign n912 = n911 ^ x124;
  assign n913 = n912 ^ n627;
  assign n914 = ~x128 & n913;
  assign n915 = n914 ^ n627;
  assign n904 = x118 ^ x116;
  assign n905 = ~x129 & n904;
  assign n906 = n905 ^ x116;
  assign n907 = n906 ^ n621;
  assign n908 = ~x128 & n907;
  assign n909 = n908 ^ n621;
  assign n916 = n915 ^ n909;
  assign n917 = x131 & n916;
  assign n918 = n917 ^ n915;
  assign n934 = n933 ^ n918;
  assign n935 = x130 & n934;
  assign n936 = n935 ^ n933;
  assign n892 = x98 ^ x96;
  assign n893 = ~x129 & n892;
  assign n894 = n893 ^ x96;
  assign n895 = n894 ^ n609;
  assign n896 = ~x128 & n895;
  assign n897 = n896 ^ n609;
  assign n886 = x90 ^ x88;
  assign n887 = ~x129 & n886;
  assign n888 = n887 ^ x88;
  assign n889 = n888 ^ n603;
  assign n890 = ~x128 & n889;
  assign n891 = n890 ^ n603;
  assign n898 = n897 ^ n891;
  assign n899 = x131 & n898;
  assign n900 = n899 ^ n897;
  assign n877 = x94 ^ x92;
  assign n878 = ~x129 & n877;
  assign n879 = n878 ^ x92;
  assign n880 = n879 ^ n594;
  assign n881 = ~x128 & n880;
  assign n882 = n881 ^ n594;
  assign n871 = x86 ^ x84;
  assign n872 = ~x129 & n871;
  assign n873 = n872 ^ x84;
  assign n874 = n873 ^ n588;
  assign n875 = ~x128 & n874;
  assign n876 = n875 ^ n588;
  assign n883 = n882 ^ n876;
  assign n884 = x131 & n883;
  assign n885 = n884 ^ n882;
  assign n901 = n900 ^ n885;
  assign n902 = x130 & n901;
  assign n903 = n902 ^ n900;
  assign n937 = n936 ^ n903;
  assign n938 = x133 & n937;
  assign n939 = n938 ^ n936;
  assign n856 = x114 ^ x112;
  assign n857 = ~x129 & n856;
  assign n858 = n857 ^ x112;
  assign n859 = n858 ^ n573;
  assign n860 = ~x128 & n859;
  assign n861 = n860 ^ n573;
  assign n850 = x106 ^ x104;
  assign n851 = ~x129 & n850;
  assign n852 = n851 ^ x104;
  assign n853 = n852 ^ n567;
  assign n854 = ~x128 & n853;
  assign n855 = n854 ^ n567;
  assign n862 = n861 ^ n855;
  assign n863 = x131 & n862;
  assign n864 = n863 ^ n861;
  assign n841 = x110 ^ x108;
  assign n842 = ~x129 & n841;
  assign n843 = n842 ^ x108;
  assign n844 = n843 ^ n558;
  assign n845 = ~x128 & n844;
  assign n846 = n845 ^ n558;
  assign n835 = x102 ^ x100;
  assign n836 = ~x129 & n835;
  assign n837 = n836 ^ x100;
  assign n838 = n837 ^ n552;
  assign n839 = ~x128 & n838;
  assign n840 = n839 ^ n552;
  assign n847 = n846 ^ n840;
  assign n848 = x131 & n847;
  assign n849 = n848 ^ n846;
  assign n865 = n864 ^ n849;
  assign n866 = x130 & n865;
  assign n867 = n866 ^ n864;
  assign n823 = x82 ^ x80;
  assign n824 = ~x129 & n823;
  assign n825 = n824 ^ x80;
  assign n826 = n825 ^ n540;
  assign n827 = ~x128 & n826;
  assign n828 = n827 ^ n540;
  assign n817 = x74 ^ x72;
  assign n818 = ~x129 & n817;
  assign n819 = n818 ^ x72;
  assign n820 = n819 ^ n534;
  assign n821 = ~x128 & n820;
  assign n822 = n821 ^ n534;
  assign n829 = n828 ^ n822;
  assign n830 = x131 & n829;
  assign n831 = n830 ^ n828;
  assign n808 = x78 ^ x76;
  assign n809 = ~x129 & n808;
  assign n810 = n809 ^ x76;
  assign n811 = n810 ^ n525;
  assign n812 = ~x128 & n811;
  assign n813 = n812 ^ n525;
  assign n802 = x70 ^ x68;
  assign n803 = ~x129 & n802;
  assign n804 = n803 ^ x68;
  assign n805 = n804 ^ n519;
  assign n806 = ~x128 & n805;
  assign n807 = n806 ^ n519;
  assign n814 = n813 ^ n807;
  assign n815 = x131 & n814;
  assign n816 = n815 ^ n813;
  assign n832 = n831 ^ n816;
  assign n833 = x130 & n832;
  assign n834 = n833 ^ n831;
  assign n868 = n867 ^ n834;
  assign n869 = x133 & n868;
  assign n870 = n869 ^ n867;
  assign n940 = n939 ^ n870;
  assign n941 = x132 & n940;
  assign n942 = n941 ^ n939;
  assign n1084 = n1083 ^ n942;
  assign n1085 = ~x134 & n1084;
  assign n1086 = n1085 ^ n1083;
  assign n1258 = n1068 ^ n138;
  assign n1259 = x128 & n1258;
  assign n1260 = n1259 ^ n138;
  assign n1255 = n1062 ^ n474;
  assign n1256 = x128 & n1255;
  assign n1257 = n1256 ^ n474;
  assign n1261 = n1260 ^ n1257;
  assign n1262 = x131 & n1261;
  assign n1263 = n1262 ^ n1260;
  assign n1249 = n1053 ^ n495;
  assign n1250 = x128 & n1249;
  assign n1251 = n1250 ^ n495;
  assign n1246 = n1047 ^ n486;
  assign n1247 = x128 & n1246;
  assign n1248 = n1247 ^ n486;
  assign n1252 = n1251 ^ n1248;
  assign n1253 = x131 & n1252;
  assign n1254 = n1253 ^ n1251;
  assign n1264 = n1263 ^ n1254;
  assign n1265 = x130 & n1264;
  assign n1266 = n1265 ^ n1263;
  assign n1237 = n1035 ^ n372;
  assign n1238 = x128 & n1237;
  assign n1239 = n1238 ^ n372;
  assign n1234 = n1029 ^ n429;
  assign n1235 = x128 & n1234;
  assign n1236 = n1235 ^ n429;
  assign n1240 = n1239 ^ n1236;
  assign n1241 = x131 & n1240;
  assign n1242 = n1241 ^ n1239;
  assign n1228 = n1020 ^ n450;
  assign n1229 = x128 & n1228;
  assign n1230 = n1229 ^ n450;
  assign n1225 = n1014 ^ n441;
  assign n1226 = x128 & n1225;
  assign n1227 = n1226 ^ n441;
  assign n1231 = n1230 ^ n1227;
  assign n1232 = x131 & n1231;
  assign n1233 = n1232 ^ n1230;
  assign n1243 = n1242 ^ n1233;
  assign n1244 = x130 & n1243;
  assign n1245 = n1244 ^ n1242;
  assign n1267 = n1266 ^ n1245;
  assign n1268 = x133 & n1267;
  assign n1269 = n1268 ^ n1266;
  assign n1213 = n999 ^ n465;
  assign n1214 = x128 & n1213;
  assign n1215 = n1214 ^ n465;
  assign n1210 = n993 ^ n381;
  assign n1211 = x128 & n1210;
  assign n1212 = n1211 ^ n381;
  assign n1216 = n1215 ^ n1212;
  assign n1217 = x131 & n1216;
  assign n1218 = n1217 ^ n1215;
  assign n1204 = n984 ^ n402;
  assign n1205 = x128 & n1204;
  assign n1206 = n1205 ^ n402;
  assign n1201 = n978 ^ n393;
  assign n1202 = x128 & n1201;
  assign n1203 = n1202 ^ n393;
  assign n1207 = n1206 ^ n1203;
  assign n1208 = x131 & n1207;
  assign n1209 = n1208 ^ n1206;
  assign n1219 = n1218 ^ n1209;
  assign n1220 = x130 & n1219;
  assign n1221 = n1220 ^ n1218;
  assign n1192 = n966 ^ n420;
  assign n1193 = x128 & n1192;
  assign n1194 = n1193 ^ n420;
  assign n1189 = n960 ^ n336;
  assign n1190 = x128 & n1189;
  assign n1191 = n1190 ^ n336;
  assign n1195 = n1194 ^ n1191;
  assign n1196 = x131 & n1195;
  assign n1197 = n1196 ^ n1194;
  assign n1183 = n951 ^ n357;
  assign n1184 = x128 & n1183;
  assign n1185 = n1184 ^ n357;
  assign n1180 = n945 ^ n348;
  assign n1181 = x128 & n1180;
  assign n1182 = n1181 ^ n348;
  assign n1186 = n1185 ^ n1182;
  assign n1187 = x131 & n1186;
  assign n1188 = n1187 ^ n1185;
  assign n1198 = n1197 ^ n1188;
  assign n1199 = x130 & n1198;
  assign n1200 = n1199 ^ n1197;
  assign n1222 = n1221 ^ n1200;
  assign n1223 = x133 & n1222;
  assign n1224 = n1223 ^ n1221;
  assign n1270 = n1269 ^ n1224;
  assign n1271 = x132 & n1270;
  assign n1272 = n1271 ^ n1269;
  assign n1165 = n927 ^ n327;
  assign n1166 = x128 & n1165;
  assign n1167 = n1166 ^ n327;
  assign n1162 = n921 ^ n285;
  assign n1163 = x128 & n1162;
  assign n1164 = n1163 ^ n285;
  assign n1168 = n1167 ^ n1164;
  assign n1169 = x131 & n1168;
  assign n1170 = n1169 ^ n1167;
  assign n1156 = n912 ^ n306;
  assign n1157 = x128 & n1156;
  assign n1158 = n1157 ^ n306;
  assign n1153 = n906 ^ n297;
  assign n1154 = x128 & n1153;
  assign n1155 = n1154 ^ n297;
  assign n1159 = n1158 ^ n1155;
  assign n1160 = x131 & n1159;
  assign n1161 = n1160 ^ n1158;
  assign n1171 = n1170 ^ n1161;
  assign n1172 = x130 & n1171;
  assign n1173 = n1172 ^ n1170;
  assign n1144 = n894 ^ n183;
  assign n1145 = x128 & n1144;
  assign n1146 = n1145 ^ n183;
  assign n1141 = n888 ^ n240;
  assign n1142 = x128 & n1141;
  assign n1143 = n1142 ^ n240;
  assign n1147 = n1146 ^ n1143;
  assign n1148 = x131 & n1147;
  assign n1149 = n1148 ^ n1146;
  assign n1135 = n879 ^ n261;
  assign n1136 = x128 & n1135;
  assign n1137 = n1136 ^ n261;
  assign n1132 = n873 ^ n252;
  assign n1133 = x128 & n1132;
  assign n1134 = n1133 ^ n252;
  assign n1138 = n1137 ^ n1134;
  assign n1139 = x131 & n1138;
  assign n1140 = n1139 ^ n1137;
  assign n1150 = n1149 ^ n1140;
  assign n1151 = x130 & n1150;
  assign n1152 = n1151 ^ n1149;
  assign n1174 = n1173 ^ n1152;
  assign n1175 = x133 & n1174;
  assign n1176 = n1175 ^ n1173;
  assign n1120 = n858 ^ n276;
  assign n1121 = x128 & n1120;
  assign n1122 = n1121 ^ n276;
  assign n1117 = n852 ^ n192;
  assign n1118 = x128 & n1117;
  assign n1119 = n1118 ^ n192;
  assign n1123 = n1122 ^ n1119;
  assign n1124 = x131 & n1123;
  assign n1125 = n1124 ^ n1122;
  assign n1111 = n843 ^ n213;
  assign n1112 = x128 & n1111;
  assign n1113 = n1112 ^ n213;
  assign n1108 = n837 ^ n204;
  assign n1109 = x128 & n1108;
  assign n1110 = n1109 ^ n204;
  assign n1114 = n1113 ^ n1110;
  assign n1115 = x131 & n1114;
  assign n1116 = n1115 ^ n1113;
  assign n1126 = n1125 ^ n1116;
  assign n1127 = x130 & n1126;
  assign n1128 = n1127 ^ n1125;
  assign n1099 = n825 ^ n231;
  assign n1100 = x128 & n1099;
  assign n1101 = n1100 ^ n231;
  assign n1096 = n819 ^ n147;
  assign n1097 = x128 & n1096;
  assign n1098 = n1097 ^ n147;
  assign n1102 = n1101 ^ n1098;
  assign n1103 = x131 & n1102;
  assign n1104 = n1103 ^ n1101;
  assign n1090 = n810 ^ n168;
  assign n1091 = x128 & n1090;
  assign n1092 = n1091 ^ n168;
  assign n1087 = n804 ^ n159;
  assign n1088 = x128 & n1087;
  assign n1089 = n1088 ^ n159;
  assign n1093 = n1092 ^ n1089;
  assign n1094 = x131 & n1093;
  assign n1095 = n1094 ^ n1092;
  assign n1105 = n1104 ^ n1095;
  assign n1106 = x130 & n1105;
  assign n1107 = n1106 ^ n1104;
  assign n1129 = n1128 ^ n1107;
  assign n1130 = x133 & n1129;
  assign n1131 = n1130 ^ n1128;
  assign n1177 = n1176 ^ n1131;
  assign n1178 = x132 & n1177;
  assign n1179 = n1178 ^ n1176;
  assign n1273 = n1272 ^ n1179;
  assign n1274 = ~x134 & n1273;
  assign n1275 = n1274 ^ n1272;
  assign n1330 = n480 ^ n144;
  assign n1331 = ~x131 & n1330;
  assign n1332 = n1331 ^ n480;
  assign n1333 = n1332 ^ n504;
  assign n1334 = ~x130 & n1333;
  assign n1335 = n1334 ^ n504;
  assign n1324 = n435 ^ n378;
  assign n1325 = ~x131 & n1324;
  assign n1326 = n1325 ^ n435;
  assign n1327 = n1326 ^ n459;
  assign n1328 = ~x130 & n1327;
  assign n1329 = n1328 ^ n459;
  assign n1336 = n1335 ^ n1329;
  assign n1337 = x133 & n1336;
  assign n1338 = n1337 ^ n1335;
  assign n1315 = n471 ^ n387;
  assign n1316 = x131 & n1315;
  assign n1317 = n1316 ^ n471;
  assign n1318 = n1317 ^ n411;
  assign n1319 = ~x130 & n1318;
  assign n1320 = n1319 ^ n411;
  assign n1309 = n426 ^ n342;
  assign n1310 = x131 & n1309;
  assign n1311 = n1310 ^ n426;
  assign n1312 = n1311 ^ n366;
  assign n1313 = ~x130 & n1312;
  assign n1314 = n1313 ^ n366;
  assign n1321 = n1320 ^ n1314;
  assign n1322 = x133 & n1321;
  assign n1323 = n1322 ^ n1320;
  assign n1339 = n1338 ^ n1323;
  assign n1340 = x132 & n1339;
  assign n1341 = n1340 ^ n1338;
  assign n1297 = n333 ^ n291;
  assign n1298 = x131 & n1297;
  assign n1299 = n1298 ^ n333;
  assign n1300 = n1299 ^ n315;
  assign n1301 = ~x130 & n1300;
  assign n1302 = n1301 ^ n315;
  assign n1291 = n246 ^ n189;
  assign n1292 = ~x131 & n1291;
  assign n1293 = n1292 ^ n246;
  assign n1294 = n1293 ^ n270;
  assign n1295 = ~x130 & n1294;
  assign n1296 = n1295 ^ n270;
  assign n1303 = n1302 ^ n1296;
  assign n1304 = x133 & n1303;
  assign n1305 = n1304 ^ n1302;
  assign n1282 = n282 ^ n198;
  assign n1283 = x131 & n1282;
  assign n1284 = n1283 ^ n282;
  assign n1285 = n1284 ^ n222;
  assign n1286 = ~x130 & n1285;
  assign n1287 = n1286 ^ n222;
  assign n1276 = n237 ^ n153;
  assign n1277 = x131 & n1276;
  assign n1278 = n1277 ^ n237;
  assign n1279 = n1278 ^ n177;
  assign n1280 = ~x130 & n1279;
  assign n1281 = n1280 ^ n177;
  assign n1288 = n1287 ^ n1281;
  assign n1289 = x133 & n1288;
  assign n1290 = n1289 ^ n1287;
  assign n1306 = n1305 ^ n1290;
  assign n1307 = x132 & n1306;
  assign n1308 = n1307 ^ n1305;
  assign n1342 = n1341 ^ n1308;
  assign n1343 = ~x134 & n1342;
  assign n1344 = n1343 ^ n1341;
  assign n1399 = n771 ^ n522;
  assign n1400 = ~x131 & n1399;
  assign n1401 = n1400 ^ n771;
  assign n1402 = n1401 ^ n789;
  assign n1403 = ~x130 & n1402;
  assign n1404 = n1403 ^ n789;
  assign n1393 = n738 ^ n696;
  assign n1394 = ~x131 & n1393;
  assign n1395 = n1394 ^ n738;
  assign n1396 = n1395 ^ n756;
  assign n1397 = ~x130 & n1396;
  assign n1398 = n1397 ^ n756;
  assign n1405 = n1404 ^ n1398;
  assign n1406 = x133 & n1405;
  assign n1407 = n1406 ^ n1404;
  assign n1384 = n765 ^ n702;
  assign n1385 = x131 & n1384;
  assign n1386 = n1385 ^ n765;
  assign n1387 = n1386 ^ n720;
  assign n1388 = ~x130 & n1387;
  assign n1389 = n1388 ^ n720;
  assign n1378 = n732 ^ n669;
  assign n1379 = x131 & n1378;
  assign n1380 = n1379 ^ n732;
  assign n1381 = n1380 ^ n687;
  assign n1382 = ~x130 & n1381;
  assign n1383 = n1382 ^ n687;
  assign n1390 = n1389 ^ n1383;
  assign n1391 = x133 & n1390;
  assign n1392 = n1391 ^ n1389;
  assign n1408 = n1407 ^ n1392;
  assign n1409 = x132 & n1408;
  assign n1410 = n1409 ^ n1407;
  assign n1366 = n663 ^ n630;
  assign n1367 = x131 & n1366;
  assign n1368 = n1367 ^ n663;
  assign n1369 = n1368 ^ n648;
  assign n1370 = ~x130 & n1369;
  assign n1371 = n1370 ^ n648;
  assign n1360 = n597 ^ n555;
  assign n1361 = ~x131 & n1360;
  assign n1362 = n1361 ^ n597;
  assign n1363 = n1362 ^ n615;
  assign n1364 = ~x130 & n1363;
  assign n1365 = n1364 ^ n615;
  assign n1372 = n1371 ^ n1365;
  assign n1373 = x133 & n1372;
  assign n1374 = n1373 ^ n1371;
  assign n1351 = n624 ^ n561;
  assign n1352 = x131 & n1351;
  assign n1353 = n1352 ^ n624;
  assign n1354 = n1353 ^ n579;
  assign n1355 = ~x130 & n1354;
  assign n1356 = n1355 ^ n579;
  assign n1345 = n591 ^ n528;
  assign n1346 = x131 & n1345;
  assign n1347 = n1346 ^ n591;
  assign n1348 = n1347 ^ n546;
  assign n1349 = ~x130 & n1348;
  assign n1350 = n1349 ^ n546;
  assign n1357 = n1356 ^ n1350;
  assign n1358 = x133 & n1357;
  assign n1359 = n1358 ^ n1356;
  assign n1375 = n1374 ^ n1359;
  assign n1376 = x132 & n1375;
  assign n1377 = n1376 ^ n1374;
  assign n1411 = n1410 ^ n1377;
  assign n1412 = ~x134 & n1411;
  assign n1413 = n1412 ^ n1410;
  assign n1468 = n1056 ^ n807;
  assign n1469 = ~x131 & n1468;
  assign n1470 = n1469 ^ n1056;
  assign n1471 = n1470 ^ n1074;
  assign n1472 = ~x130 & n1471;
  assign n1473 = n1472 ^ n1074;
  assign n1462 = n1023 ^ n981;
  assign n1463 = ~x131 & n1462;
  assign n1464 = n1463 ^ n1023;
  assign n1465 = n1464 ^ n1041;
  assign n1466 = ~x130 & n1465;
  assign n1467 = n1466 ^ n1041;
  assign n1474 = n1473 ^ n1467;
  assign n1475 = x133 & n1474;
  assign n1476 = n1475 ^ n1473;
  assign n1453 = n1050 ^ n987;
  assign n1454 = x131 & n1453;
  assign n1455 = n1454 ^ n1050;
  assign n1456 = n1455 ^ n1005;
  assign n1457 = ~x130 & n1456;
  assign n1458 = n1457 ^ n1005;
  assign n1447 = n1017 ^ n954;
  assign n1448 = x131 & n1447;
  assign n1449 = n1448 ^ n1017;
  assign n1450 = n1449 ^ n972;
  assign n1451 = ~x130 & n1450;
  assign n1452 = n1451 ^ n972;
  assign n1459 = n1458 ^ n1452;
  assign n1460 = x133 & n1459;
  assign n1461 = n1460 ^ n1458;
  assign n1477 = n1476 ^ n1461;
  assign n1478 = x132 & n1477;
  assign n1479 = n1478 ^ n1476;
  assign n1435 = n948 ^ n915;
  assign n1436 = x131 & n1435;
  assign n1437 = n1436 ^ n948;
  assign n1438 = n1437 ^ n933;
  assign n1439 = ~x130 & n1438;
  assign n1440 = n1439 ^ n933;
  assign n1429 = n882 ^ n840;
  assign n1430 = ~x131 & n1429;
  assign n1431 = n1430 ^ n882;
  assign n1432 = n1431 ^ n900;
  assign n1433 = ~x130 & n1432;
  assign n1434 = n1433 ^ n900;
  assign n1441 = n1440 ^ n1434;
  assign n1442 = x133 & n1441;
  assign n1443 = n1442 ^ n1440;
  assign n1420 = n909 ^ n846;
  assign n1421 = x131 & n1420;
  assign n1422 = n1421 ^ n909;
  assign n1423 = n1422 ^ n864;
  assign n1424 = ~x130 & n1423;
  assign n1425 = n1424 ^ n864;
  assign n1414 = n876 ^ n813;
  assign n1415 = x131 & n1414;
  assign n1416 = n1415 ^ n876;
  assign n1417 = n1416 ^ n831;
  assign n1418 = ~x130 & n1417;
  assign n1419 = n1418 ^ n831;
  assign n1426 = n1425 ^ n1419;
  assign n1427 = x133 & n1426;
  assign n1428 = n1427 ^ n1425;
  assign n1444 = n1443 ^ n1428;
  assign n1445 = x132 & n1444;
  assign n1446 = n1445 ^ n1443;
  assign n1480 = n1479 ^ n1446;
  assign n1481 = ~x134 & n1480;
  assign n1482 = n1481 ^ n1479;
  assign n1537 = n1251 ^ n1089;
  assign n1538 = ~x131 & n1537;
  assign n1539 = n1538 ^ n1251;
  assign n1540 = n1539 ^ n1263;
  assign n1541 = ~x130 & n1540;
  assign n1542 = n1541 ^ n1263;
  assign n1531 = n1230 ^ n1203;
  assign n1532 = ~x131 & n1531;
  assign n1533 = n1532 ^ n1230;
  assign n1534 = n1533 ^ n1242;
  assign n1535 = ~x130 & n1534;
  assign n1536 = n1535 ^ n1242;
  assign n1543 = n1542 ^ n1536;
  assign n1544 = x133 & n1543;
  assign n1545 = n1544 ^ n1542;
  assign n1522 = n1248 ^ n1206;
  assign n1523 = x131 & n1522;
  assign n1524 = n1523 ^ n1248;
  assign n1525 = n1524 ^ n1218;
  assign n1526 = ~x130 & n1525;
  assign n1527 = n1526 ^ n1218;
  assign n1516 = n1227 ^ n1185;
  assign n1517 = x131 & n1516;
  assign n1518 = n1517 ^ n1227;
  assign n1519 = n1518 ^ n1197;
  assign n1520 = ~x130 & n1519;
  assign n1521 = n1520 ^ n1197;
  assign n1528 = n1527 ^ n1521;
  assign n1529 = x133 & n1528;
  assign n1530 = n1529 ^ n1527;
  assign n1546 = n1545 ^ n1530;
  assign n1547 = x132 & n1546;
  assign n1548 = n1547 ^ n1545;
  assign n1504 = n1182 ^ n1158;
  assign n1505 = x131 & n1504;
  assign n1506 = n1505 ^ n1182;
  assign n1507 = n1506 ^ n1170;
  assign n1508 = ~x130 & n1507;
  assign n1509 = n1508 ^ n1170;
  assign n1498 = n1137 ^ n1110;
  assign n1499 = ~x131 & n1498;
  assign n1500 = n1499 ^ n1137;
  assign n1501 = n1500 ^ n1149;
  assign n1502 = ~x130 & n1501;
  assign n1503 = n1502 ^ n1149;
  assign n1510 = n1509 ^ n1503;
  assign n1511 = x133 & n1510;
  assign n1512 = n1511 ^ n1509;
  assign n1489 = n1155 ^ n1113;
  assign n1490 = x131 & n1489;
  assign n1491 = n1490 ^ n1155;
  assign n1492 = n1491 ^ n1125;
  assign n1493 = ~x130 & n1492;
  assign n1494 = n1493 ^ n1125;
  assign n1483 = n1134 ^ n1092;
  assign n1484 = x131 & n1483;
  assign n1485 = n1484 ^ n1134;
  assign n1486 = n1485 ^ n1104;
  assign n1487 = ~x130 & n1486;
  assign n1488 = n1487 ^ n1104;
  assign n1495 = n1494 ^ n1488;
  assign n1496 = x133 & n1495;
  assign n1497 = n1496 ^ n1494;
  assign n1513 = n1512 ^ n1497;
  assign n1514 = x132 & n1513;
  assign n1515 = n1514 ^ n1512;
  assign n1549 = n1548 ^ n1515;
  assign n1550 = ~x134 & n1549;
  assign n1551 = n1550 ^ n1548;
  assign n1606 = n501 ^ n165;
  assign n1607 = ~x131 & n1606;
  assign n1608 = n1607 ^ n501;
  assign n1609 = n1608 ^ n1332;
  assign n1610 = ~x130 & n1609;
  assign n1611 = n1610 ^ n1332;
  assign n1600 = n456 ^ n399;
  assign n1601 = ~x131 & n1600;
  assign n1602 = n1601 ^ n456;
  assign n1603 = n1602 ^ n1326;
  assign n1604 = ~x130 & n1603;
  assign n1605 = n1604 ^ n1326;
  assign n1612 = n1611 ^ n1605;
  assign n1613 = x133 & n1612;
  assign n1614 = n1613 ^ n1611;
  assign n1591 = n492 ^ n408;
  assign n1592 = x131 & n1591;
  assign n1593 = n1592 ^ n492;
  assign n1594 = n1593 ^ n1317;
  assign n1595 = ~x130 & n1594;
  assign n1596 = n1595 ^ n1317;
  assign n1585 = n447 ^ n363;
  assign n1586 = x131 & n1585;
  assign n1587 = n1586 ^ n447;
  assign n1588 = n1587 ^ n1311;
  assign n1589 = ~x130 & n1588;
  assign n1590 = n1589 ^ n1311;
  assign n1597 = n1596 ^ n1590;
  assign n1598 = x133 & n1597;
  assign n1599 = n1598 ^ n1596;
  assign n1615 = n1614 ^ n1599;
  assign n1616 = x132 & n1615;
  assign n1617 = n1616 ^ n1614;
  assign n1573 = n354 ^ n312;
  assign n1574 = x131 & n1573;
  assign n1575 = n1574 ^ n354;
  assign n1576 = n1575 ^ n1299;
  assign n1577 = ~x130 & n1576;
  assign n1578 = n1577 ^ n1299;
  assign n1567 = n267 ^ n210;
  assign n1568 = ~x131 & n1567;
  assign n1569 = n1568 ^ n267;
  assign n1570 = n1569 ^ n1293;
  assign n1571 = ~x130 & n1570;
  assign n1572 = n1571 ^ n1293;
  assign n1579 = n1578 ^ n1572;
  assign n1580 = x133 & n1579;
  assign n1581 = n1580 ^ n1578;
  assign n1558 = n303 ^ n219;
  assign n1559 = x131 & n1558;
  assign n1560 = n1559 ^ n303;
  assign n1561 = n1560 ^ n1284;
  assign n1562 = ~x130 & n1561;
  assign n1563 = n1562 ^ n1284;
  assign n1552 = n258 ^ n174;
  assign n1553 = x131 & n1552;
  assign n1554 = n1553 ^ n258;
  assign n1555 = n1554 ^ n1278;
  assign n1556 = ~x130 & n1555;
  assign n1557 = n1556 ^ n1278;
  assign n1564 = n1563 ^ n1557;
  assign n1565 = x133 & n1564;
  assign n1566 = n1565 ^ n1563;
  assign n1582 = n1581 ^ n1566;
  assign n1583 = x132 & n1582;
  assign n1584 = n1583 ^ n1581;
  assign n1618 = n1617 ^ n1584;
  assign n1619 = ~x134 & n1618;
  assign n1620 = n1619 ^ n1617;
  assign n1675 = n786 ^ n537;
  assign n1676 = ~x131 & n1675;
  assign n1677 = n1676 ^ n786;
  assign n1678 = n1677 ^ n1401;
  assign n1679 = ~x130 & n1678;
  assign n1680 = n1679 ^ n1401;
  assign n1669 = n753 ^ n711;
  assign n1670 = ~x131 & n1669;
  assign n1671 = n1670 ^ n753;
  assign n1672 = n1671 ^ n1395;
  assign n1673 = ~x130 & n1672;
  assign n1674 = n1673 ^ n1395;
  assign n1681 = n1680 ^ n1674;
  assign n1682 = x133 & n1681;
  assign n1683 = n1682 ^ n1680;
  assign n1660 = n780 ^ n717;
  assign n1661 = x131 & n1660;
  assign n1662 = n1661 ^ n780;
  assign n1663 = n1662 ^ n1386;
  assign n1664 = ~x130 & n1663;
  assign n1665 = n1664 ^ n1386;
  assign n1654 = n747 ^ n684;
  assign n1655 = x131 & n1654;
  assign n1656 = n1655 ^ n747;
  assign n1657 = n1656 ^ n1380;
  assign n1658 = ~x130 & n1657;
  assign n1659 = n1658 ^ n1380;
  assign n1666 = n1665 ^ n1659;
  assign n1667 = x133 & n1666;
  assign n1668 = n1667 ^ n1665;
  assign n1684 = n1683 ^ n1668;
  assign n1685 = x132 & n1684;
  assign n1686 = n1685 ^ n1683;
  assign n1642 = n678 ^ n645;
  assign n1643 = x131 & n1642;
  assign n1644 = n1643 ^ n678;
  assign n1645 = n1644 ^ n1368;
  assign n1646 = ~x130 & n1645;
  assign n1647 = n1646 ^ n1368;
  assign n1636 = n612 ^ n570;
  assign n1637 = ~x131 & n1636;
  assign n1638 = n1637 ^ n612;
  assign n1639 = n1638 ^ n1362;
  assign n1640 = ~x130 & n1639;
  assign n1641 = n1640 ^ n1362;
  assign n1648 = n1647 ^ n1641;
  assign n1649 = x133 & n1648;
  assign n1650 = n1649 ^ n1647;
  assign n1627 = n639 ^ n576;
  assign n1628 = x131 & n1627;
  assign n1629 = n1628 ^ n639;
  assign n1630 = n1629 ^ n1353;
  assign n1631 = ~x130 & n1630;
  assign n1632 = n1631 ^ n1353;
  assign n1621 = n606 ^ n543;
  assign n1622 = x131 & n1621;
  assign n1623 = n1622 ^ n606;
  assign n1624 = n1623 ^ n1347;
  assign n1625 = ~x130 & n1624;
  assign n1626 = n1625 ^ n1347;
  assign n1633 = n1632 ^ n1626;
  assign n1634 = x133 & n1633;
  assign n1635 = n1634 ^ n1632;
  assign n1651 = n1650 ^ n1635;
  assign n1652 = x132 & n1651;
  assign n1653 = n1652 ^ n1650;
  assign n1687 = n1686 ^ n1653;
  assign n1688 = ~x134 & n1687;
  assign n1689 = n1688 ^ n1686;
  assign n1744 = n1071 ^ n822;
  assign n1745 = ~x131 & n1744;
  assign n1746 = n1745 ^ n1071;
  assign n1747 = n1746 ^ n1470;
  assign n1748 = ~x130 & n1747;
  assign n1749 = n1748 ^ n1470;
  assign n1738 = n1038 ^ n996;
  assign n1739 = ~x131 & n1738;
  assign n1740 = n1739 ^ n1038;
  assign n1741 = n1740 ^ n1464;
  assign n1742 = ~x130 & n1741;
  assign n1743 = n1742 ^ n1464;
  assign n1750 = n1749 ^ n1743;
  assign n1751 = x133 & n1750;
  assign n1752 = n1751 ^ n1749;
  assign n1729 = n1065 ^ n1002;
  assign n1730 = x131 & n1729;
  assign n1731 = n1730 ^ n1065;
  assign n1732 = n1731 ^ n1455;
  assign n1733 = ~x130 & n1732;
  assign n1734 = n1733 ^ n1455;
  assign n1723 = n1032 ^ n969;
  assign n1724 = x131 & n1723;
  assign n1725 = n1724 ^ n1032;
  assign n1726 = n1725 ^ n1449;
  assign n1727 = ~x130 & n1726;
  assign n1728 = n1727 ^ n1449;
  assign n1735 = n1734 ^ n1728;
  assign n1736 = x133 & n1735;
  assign n1737 = n1736 ^ n1734;
  assign n1753 = n1752 ^ n1737;
  assign n1754 = x132 & n1753;
  assign n1755 = n1754 ^ n1752;
  assign n1711 = n963 ^ n930;
  assign n1712 = x131 & n1711;
  assign n1713 = n1712 ^ n963;
  assign n1714 = n1713 ^ n1437;
  assign n1715 = ~x130 & n1714;
  assign n1716 = n1715 ^ n1437;
  assign n1705 = n897 ^ n855;
  assign n1706 = ~x131 & n1705;
  assign n1707 = n1706 ^ n897;
  assign n1708 = n1707 ^ n1431;
  assign n1709 = ~x130 & n1708;
  assign n1710 = n1709 ^ n1431;
  assign n1717 = n1716 ^ n1710;
  assign n1718 = x133 & n1717;
  assign n1719 = n1718 ^ n1716;
  assign n1696 = n924 ^ n861;
  assign n1697 = x131 & n1696;
  assign n1698 = n1697 ^ n924;
  assign n1699 = n1698 ^ n1422;
  assign n1700 = ~x130 & n1699;
  assign n1701 = n1700 ^ n1422;
  assign n1690 = n891 ^ n828;
  assign n1691 = x131 & n1690;
  assign n1692 = n1691 ^ n891;
  assign n1693 = n1692 ^ n1416;
  assign n1694 = ~x130 & n1693;
  assign n1695 = n1694 ^ n1416;
  assign n1702 = n1701 ^ n1695;
  assign n1703 = x133 & n1702;
  assign n1704 = n1703 ^ n1701;
  assign n1720 = n1719 ^ n1704;
  assign n1721 = x132 & n1720;
  assign n1722 = n1721 ^ n1719;
  assign n1756 = n1755 ^ n1722;
  assign n1757 = ~x134 & n1756;
  assign n1758 = n1757 ^ n1755;
  assign n1813 = n1260 ^ n1098;
  assign n1814 = ~x131 & n1813;
  assign n1815 = n1814 ^ n1260;
  assign n1816 = n1815 ^ n1539;
  assign n1817 = ~x130 & n1816;
  assign n1818 = n1817 ^ n1539;
  assign n1807 = n1239 ^ n1212;
  assign n1808 = ~x131 & n1807;
  assign n1809 = n1808 ^ n1239;
  assign n1810 = n1809 ^ n1533;
  assign n1811 = ~x130 & n1810;
  assign n1812 = n1811 ^ n1533;
  assign n1819 = n1818 ^ n1812;
  assign n1820 = x133 & n1819;
  assign n1821 = n1820 ^ n1818;
  assign n1798 = n1257 ^ n1215;
  assign n1799 = x131 & n1798;
  assign n1800 = n1799 ^ n1257;
  assign n1801 = n1800 ^ n1524;
  assign n1802 = ~x130 & n1801;
  assign n1803 = n1802 ^ n1524;
  assign n1792 = n1236 ^ n1194;
  assign n1793 = x131 & n1792;
  assign n1794 = n1793 ^ n1236;
  assign n1795 = n1794 ^ n1518;
  assign n1796 = ~x130 & n1795;
  assign n1797 = n1796 ^ n1518;
  assign n1804 = n1803 ^ n1797;
  assign n1805 = x133 & n1804;
  assign n1806 = n1805 ^ n1803;
  assign n1822 = n1821 ^ n1806;
  assign n1823 = x132 & n1822;
  assign n1824 = n1823 ^ n1821;
  assign n1780 = n1191 ^ n1167;
  assign n1781 = x131 & n1780;
  assign n1782 = n1781 ^ n1191;
  assign n1783 = n1782 ^ n1506;
  assign n1784 = ~x130 & n1783;
  assign n1785 = n1784 ^ n1506;
  assign n1774 = n1146 ^ n1119;
  assign n1775 = ~x131 & n1774;
  assign n1776 = n1775 ^ n1146;
  assign n1777 = n1776 ^ n1500;
  assign n1778 = ~x130 & n1777;
  assign n1779 = n1778 ^ n1500;
  assign n1786 = n1785 ^ n1779;
  assign n1787 = x133 & n1786;
  assign n1788 = n1787 ^ n1785;
  assign n1765 = n1164 ^ n1122;
  assign n1766 = x131 & n1765;
  assign n1767 = n1766 ^ n1164;
  assign n1768 = n1767 ^ n1491;
  assign n1769 = ~x130 & n1768;
  assign n1770 = n1769 ^ n1491;
  assign n1759 = n1143 ^ n1101;
  assign n1760 = x131 & n1759;
  assign n1761 = n1760 ^ n1143;
  assign n1762 = n1761 ^ n1485;
  assign n1763 = ~x130 & n1762;
  assign n1764 = n1763 ^ n1485;
  assign n1771 = n1770 ^ n1764;
  assign n1772 = x133 & n1771;
  assign n1773 = n1772 ^ n1770;
  assign n1789 = n1788 ^ n1773;
  assign n1790 = x132 & n1789;
  assign n1791 = n1790 ^ n1788;
  assign n1825 = n1824 ^ n1791;
  assign n1826 = ~x134 & n1825;
  assign n1827 = n1826 ^ n1824;
  assign n1861 = n1608 ^ n156;
  assign n1862 = x130 & n1861;
  assign n1863 = n1862 ^ n156;
  assign n1858 = n1602 ^ n390;
  assign n1859 = x130 & n1858;
  assign n1860 = n1859 ^ n390;
  assign n1864 = n1863 ^ n1860;
  assign n1865 = x133 & n1864;
  assign n1866 = n1865 ^ n1863;
  assign n1852 = n1593 ^ n483;
  assign n1853 = x130 & n1852;
  assign n1854 = n1853 ^ n483;
  assign n1849 = n1587 ^ n438;
  assign n1850 = x130 & n1849;
  assign n1851 = n1850 ^ n438;
  assign n1855 = n1854 ^ n1851;
  assign n1856 = x133 & n1855;
  assign n1857 = n1856 ^ n1854;
  assign n1867 = n1866 ^ n1857;
  assign n1868 = x132 & n1867;
  assign n1869 = n1868 ^ n1866;
  assign n1840 = n1575 ^ n345;
  assign n1841 = x130 & n1840;
  assign n1842 = n1841 ^ n345;
  assign n1837 = n1569 ^ n201;
  assign n1838 = x130 & n1837;
  assign n1839 = n1838 ^ n201;
  assign n1843 = n1842 ^ n1839;
  assign n1844 = x133 & n1843;
  assign n1845 = n1844 ^ n1842;
  assign n1831 = n1560 ^ n294;
  assign n1832 = x130 & n1831;
  assign n1833 = n1832 ^ n294;
  assign n1828 = n1554 ^ n249;
  assign n1829 = x130 & n1828;
  assign n1830 = n1829 ^ n249;
  assign n1834 = n1833 ^ n1830;
  assign n1835 = x133 & n1834;
  assign n1836 = n1835 ^ n1833;
  assign n1846 = n1845 ^ n1836;
  assign n1847 = x132 & n1846;
  assign n1848 = n1847 ^ n1845;
  assign n1870 = n1869 ^ n1848;
  assign n1871 = ~x134 & n1870;
  assign n1872 = n1871 ^ n1869;
  assign n1906 = n1677 ^ n531;
  assign n1907 = x130 & n1906;
  assign n1908 = n1907 ^ n531;
  assign n1903 = n1671 ^ n705;
  assign n1904 = x130 & n1903;
  assign n1905 = n1904 ^ n705;
  assign n1909 = n1908 ^ n1905;
  assign n1910 = x133 & n1909;
  assign n1911 = n1910 ^ n1908;
  assign n1897 = n1662 ^ n774;
  assign n1898 = x130 & n1897;
  assign n1899 = n1898 ^ n774;
  assign n1894 = n1656 ^ n741;
  assign n1895 = x130 & n1894;
  assign n1896 = n1895 ^ n741;
  assign n1900 = n1899 ^ n1896;
  assign n1901 = x133 & n1900;
  assign n1902 = n1901 ^ n1899;
  assign n1912 = n1911 ^ n1902;
  assign n1913 = x132 & n1912;
  assign n1914 = n1913 ^ n1911;
  assign n1885 = n1644 ^ n672;
  assign n1886 = x130 & n1885;
  assign n1887 = n1886 ^ n672;
  assign n1882 = n1638 ^ n564;
  assign n1883 = x130 & n1882;
  assign n1884 = n1883 ^ n564;
  assign n1888 = n1887 ^ n1884;
  assign n1889 = x133 & n1888;
  assign n1890 = n1889 ^ n1887;
  assign n1876 = n1629 ^ n633;
  assign n1877 = x130 & n1876;
  assign n1878 = n1877 ^ n633;
  assign n1873 = n1623 ^ n600;
  assign n1874 = x130 & n1873;
  assign n1875 = n1874 ^ n600;
  assign n1879 = n1878 ^ n1875;
  assign n1880 = x133 & n1879;
  assign n1881 = n1880 ^ n1878;
  assign n1891 = n1890 ^ n1881;
  assign n1892 = x132 & n1891;
  assign n1893 = n1892 ^ n1890;
  assign n1915 = n1914 ^ n1893;
  assign n1916 = ~x134 & n1915;
  assign n1917 = n1916 ^ n1914;
  assign n1951 = n1746 ^ n816;
  assign n1952 = x130 & n1951;
  assign n1953 = n1952 ^ n816;
  assign n1948 = n1740 ^ n990;
  assign n1949 = x130 & n1948;
  assign n1950 = n1949 ^ n990;
  assign n1954 = n1953 ^ n1950;
  assign n1955 = x133 & n1954;
  assign n1956 = n1955 ^ n1953;
  assign n1942 = n1731 ^ n1059;
  assign n1943 = x130 & n1942;
  assign n1944 = n1943 ^ n1059;
  assign n1939 = n1725 ^ n1026;
  assign n1940 = x130 & n1939;
  assign n1941 = n1940 ^ n1026;
  assign n1945 = n1944 ^ n1941;
  assign n1946 = x133 & n1945;
  assign n1947 = n1946 ^ n1944;
  assign n1957 = n1956 ^ n1947;
  assign n1958 = x132 & n1957;
  assign n1959 = n1958 ^ n1956;
  assign n1930 = n1713 ^ n957;
  assign n1931 = x130 & n1930;
  assign n1932 = n1931 ^ n957;
  assign n1927 = n1707 ^ n849;
  assign n1928 = x130 & n1927;
  assign n1929 = n1928 ^ n849;
  assign n1933 = n1932 ^ n1929;
  assign n1934 = x133 & n1933;
  assign n1935 = n1934 ^ n1932;
  assign n1921 = n1698 ^ n918;
  assign n1922 = x130 & n1921;
  assign n1923 = n1922 ^ n918;
  assign n1918 = n1692 ^ n885;
  assign n1919 = x130 & n1918;
  assign n1920 = n1919 ^ n885;
  assign n1924 = n1923 ^ n1920;
  assign n1925 = x133 & n1924;
  assign n1926 = n1925 ^ n1923;
  assign n1936 = n1935 ^ n1926;
  assign n1937 = x132 & n1936;
  assign n1938 = n1937 ^ n1935;
  assign n1960 = n1959 ^ n1938;
  assign n1961 = ~x134 & n1960;
  assign n1962 = n1961 ^ n1959;
  assign n1996 = n1815 ^ n1095;
  assign n1997 = x130 & n1996;
  assign n1998 = n1997 ^ n1095;
  assign n1993 = n1809 ^ n1209;
  assign n1994 = x130 & n1993;
  assign n1995 = n1994 ^ n1209;
  assign n1999 = n1998 ^ n1995;
  assign n2000 = x133 & n1999;
  assign n2001 = n2000 ^ n1998;
  assign n1987 = n1800 ^ n1254;
  assign n1988 = x130 & n1987;
  assign n1989 = n1988 ^ n1254;
  assign n1984 = n1794 ^ n1233;
  assign n1985 = x130 & n1984;
  assign n1986 = n1985 ^ n1233;
  assign n1990 = n1989 ^ n1986;
  assign n1991 = x133 & n1990;
  assign n1992 = n1991 ^ n1989;
  assign n2002 = n2001 ^ n1992;
  assign n2003 = x132 & n2002;
  assign n2004 = n2003 ^ n2001;
  assign n1975 = n1782 ^ n1188;
  assign n1976 = x130 & n1975;
  assign n1977 = n1976 ^ n1188;
  assign n1972 = n1776 ^ n1116;
  assign n1973 = x130 & n1972;
  assign n1974 = n1973 ^ n1116;
  assign n1978 = n1977 ^ n1974;
  assign n1979 = x133 & n1978;
  assign n1980 = n1979 ^ n1977;
  assign n1966 = n1767 ^ n1161;
  assign n1967 = x130 & n1966;
  assign n1968 = n1967 ^ n1161;
  assign n1963 = n1761 ^ n1140;
  assign n1964 = x130 & n1963;
  assign n1965 = n1964 ^ n1140;
  assign n1969 = n1968 ^ n1965;
  assign n1970 = x133 & n1969;
  assign n1971 = n1970 ^ n1968;
  assign n1981 = n1980 ^ n1971;
  assign n1982 = x132 & n1981;
  assign n1983 = n1982 ^ n1980;
  assign n2005 = n2004 ^ n1983;
  assign n2006 = ~x134 & n2005;
  assign n2007 = n2006 ^ n2004;
  assign n2014 = n414 ^ n180;
  assign n2015 = ~x133 & n2014;
  assign n2016 = n2015 ^ n414;
  assign n2017 = n2016 ^ n510;
  assign n2018 = ~x132 & n2017;
  assign n2019 = n2018 ^ n510;
  assign n2008 = n369 ^ n225;
  assign n2009 = x133 & n2008;
  assign n2010 = n2009 ^ n369;
  assign n2011 = n2010 ^ n321;
  assign n2012 = ~x132 & n2011;
  assign n2013 = n2012 ^ n321;
  assign n2020 = n2019 ^ n2013;
  assign n2021 = ~x134 & n2020;
  assign n2022 = n2021 ^ n2019;
  assign n2029 = n723 ^ n549;
  assign n2030 = ~x133 & n2029;
  assign n2031 = n2030 ^ n723;
  assign n2032 = n2031 ^ n795;
  assign n2033 = ~x132 & n2032;
  assign n2034 = n2033 ^ n795;
  assign n2023 = n690 ^ n582;
  assign n2024 = x133 & n2023;
  assign n2025 = n2024 ^ n690;
  assign n2026 = n2025 ^ n654;
  assign n2027 = ~x132 & n2026;
  assign n2028 = n2027 ^ n654;
  assign n2035 = n2034 ^ n2028;
  assign n2036 = ~x134 & n2035;
  assign n2037 = n2036 ^ n2034;
  assign n2044 = n1008 ^ n834;
  assign n2045 = ~x133 & n2044;
  assign n2046 = n2045 ^ n1008;
  assign n2047 = n2046 ^ n1080;
  assign n2048 = ~x132 & n2047;
  assign n2049 = n2048 ^ n1080;
  assign n2038 = n975 ^ n867;
  assign n2039 = x133 & n2038;
  assign n2040 = n2039 ^ n975;
  assign n2041 = n2040 ^ n939;
  assign n2042 = ~x132 & n2041;
  assign n2043 = n2042 ^ n939;
  assign n2050 = n2049 ^ n2043;
  assign n2051 = ~x134 & n2050;
  assign n2052 = n2051 ^ n2049;
  assign n2059 = n1221 ^ n1107;
  assign n2060 = ~x133 & n2059;
  assign n2061 = n2060 ^ n1221;
  assign n2062 = n2061 ^ n1269;
  assign n2063 = ~x132 & n2062;
  assign n2064 = n2063 ^ n1269;
  assign n2053 = n1200 ^ n1128;
  assign n2054 = x133 & n2053;
  assign n2055 = n2054 ^ n1200;
  assign n2056 = n2055 ^ n1176;
  assign n2057 = ~x132 & n2056;
  assign n2058 = n2057 ^ n1176;
  assign n2065 = n2064 ^ n2058;
  assign n2066 = ~x134 & n2065;
  assign n2067 = n2066 ^ n2064;
  assign n2074 = n1320 ^ n1281;
  assign n2075 = ~x133 & n2074;
  assign n2076 = n2075 ^ n1320;
  assign n2077 = n2076 ^ n1338;
  assign n2078 = ~x132 & n2077;
  assign n2079 = n2078 ^ n1338;
  assign n2068 = n1314 ^ n1287;
  assign n2069 = x133 & n2068;
  assign n2070 = n2069 ^ n1314;
  assign n2071 = n2070 ^ n1305;
  assign n2072 = ~x132 & n2071;
  assign n2073 = n2072 ^ n1305;
  assign n2080 = n2079 ^ n2073;
  assign n2081 = ~x134 & n2080;
  assign n2082 = n2081 ^ n2079;
  assign n2089 = n1389 ^ n1350;
  assign n2090 = ~x133 & n2089;
  assign n2091 = n2090 ^ n1389;
  assign n2092 = n2091 ^ n1407;
  assign n2093 = ~x132 & n2092;
  assign n2094 = n2093 ^ n1407;
  assign n2083 = n1383 ^ n1356;
  assign n2084 = x133 & n2083;
  assign n2085 = n2084 ^ n1383;
  assign n2086 = n2085 ^ n1374;
  assign n2087 = ~x132 & n2086;
  assign n2088 = n2087 ^ n1374;
  assign n2095 = n2094 ^ n2088;
  assign n2096 = ~x134 & n2095;
  assign n2097 = n2096 ^ n2094;
  assign n2104 = n1458 ^ n1419;
  assign n2105 = ~x133 & n2104;
  assign n2106 = n2105 ^ n1458;
  assign n2107 = n2106 ^ n1476;
  assign n2108 = ~x132 & n2107;
  assign n2109 = n2108 ^ n1476;
  assign n2098 = n1452 ^ n1425;
  assign n2099 = x133 & n2098;
  assign n2100 = n2099 ^ n1452;
  assign n2101 = n2100 ^ n1443;
  assign n2102 = ~x132 & n2101;
  assign n2103 = n2102 ^ n1443;
  assign n2110 = n2109 ^ n2103;
  assign n2111 = ~x134 & n2110;
  assign n2112 = n2111 ^ n2109;
  assign n2119 = n1527 ^ n1488;
  assign n2120 = ~x133 & n2119;
  assign n2121 = n2120 ^ n1527;
  assign n2122 = n2121 ^ n1545;
  assign n2123 = ~x132 & n2122;
  assign n2124 = n2123 ^ n1545;
  assign n2113 = n1521 ^ n1494;
  assign n2114 = x133 & n2113;
  assign n2115 = n2114 ^ n1521;
  assign n2116 = n2115 ^ n1512;
  assign n2117 = ~x132 & n2116;
  assign n2118 = n2117 ^ n1512;
  assign n2125 = n2124 ^ n2118;
  assign n2126 = ~x134 & n2125;
  assign n2127 = n2126 ^ n2124;
  assign n2134 = n1596 ^ n1557;
  assign n2135 = ~x133 & n2134;
  assign n2136 = n2135 ^ n1596;
  assign n2137 = n2136 ^ n1614;
  assign n2138 = ~x132 & n2137;
  assign n2139 = n2138 ^ n1614;
  assign n2128 = n1590 ^ n1563;
  assign n2129 = x133 & n2128;
  assign n2130 = n2129 ^ n1590;
  assign n2131 = n2130 ^ n1581;
  assign n2132 = ~x132 & n2131;
  assign n2133 = n2132 ^ n1581;
  assign n2140 = n2139 ^ n2133;
  assign n2141 = ~x134 & n2140;
  assign n2142 = n2141 ^ n2139;
  assign n2149 = n1665 ^ n1626;
  assign n2150 = ~x133 & n2149;
  assign n2151 = n2150 ^ n1665;
  assign n2152 = n2151 ^ n1683;
  assign n2153 = ~x132 & n2152;
  assign n2154 = n2153 ^ n1683;
  assign n2143 = n1659 ^ n1632;
  assign n2144 = x133 & n2143;
  assign n2145 = n2144 ^ n1659;
  assign n2146 = n2145 ^ n1650;
  assign n2147 = ~x132 & n2146;
  assign n2148 = n2147 ^ n1650;
  assign n2155 = n2154 ^ n2148;
  assign n2156 = ~x134 & n2155;
  assign n2157 = n2156 ^ n2154;
  assign n2164 = n1734 ^ n1695;
  assign n2165 = ~x133 & n2164;
  assign n2166 = n2165 ^ n1734;
  assign n2167 = n2166 ^ n1752;
  assign n2168 = ~x132 & n2167;
  assign n2169 = n2168 ^ n1752;
  assign n2158 = n1728 ^ n1701;
  assign n2159 = x133 & n2158;
  assign n2160 = n2159 ^ n1728;
  assign n2161 = n2160 ^ n1719;
  assign n2162 = ~x132 & n2161;
  assign n2163 = n2162 ^ n1719;
  assign n2170 = n2169 ^ n2163;
  assign n2171 = ~x134 & n2170;
  assign n2172 = n2171 ^ n2169;
  assign n2179 = n1803 ^ n1764;
  assign n2180 = ~x133 & n2179;
  assign n2181 = n2180 ^ n1803;
  assign n2182 = n2181 ^ n1821;
  assign n2183 = ~x132 & n2182;
  assign n2184 = n2183 ^ n1821;
  assign n2173 = n1797 ^ n1770;
  assign n2174 = x133 & n2173;
  assign n2175 = n2174 ^ n1797;
  assign n2176 = n2175 ^ n1788;
  assign n2177 = ~x132 & n2176;
  assign n2178 = n2177 ^ n1788;
  assign n2185 = n2184 ^ n2178;
  assign n2186 = ~x134 & n2185;
  assign n2187 = n2186 ^ n2184;
  assign n2194 = n1854 ^ n1830;
  assign n2195 = ~x133 & n2194;
  assign n2196 = n2195 ^ n1854;
  assign n2197 = n2196 ^ n1866;
  assign n2198 = ~x132 & n2197;
  assign n2199 = n2198 ^ n1866;
  assign n2188 = n1851 ^ n1833;
  assign n2189 = x133 & n2188;
  assign n2190 = n2189 ^ n1851;
  assign n2191 = n2190 ^ n1845;
  assign n2192 = ~x132 & n2191;
  assign n2193 = n2192 ^ n1845;
  assign n2200 = n2199 ^ n2193;
  assign n2201 = ~x134 & n2200;
  assign n2202 = n2201 ^ n2199;
  assign n2209 = n1899 ^ n1875;
  assign n2210 = ~x133 & n2209;
  assign n2211 = n2210 ^ n1899;
  assign n2212 = n2211 ^ n1911;
  assign n2213 = ~x132 & n2212;
  assign n2214 = n2213 ^ n1911;
  assign n2203 = n1896 ^ n1878;
  assign n2204 = x133 & n2203;
  assign n2205 = n2204 ^ n1896;
  assign n2206 = n2205 ^ n1890;
  assign n2207 = ~x132 & n2206;
  assign n2208 = n2207 ^ n1890;
  assign n2215 = n2214 ^ n2208;
  assign n2216 = ~x134 & n2215;
  assign n2217 = n2216 ^ n2214;
  assign n2224 = n1944 ^ n1920;
  assign n2225 = ~x133 & n2224;
  assign n2226 = n2225 ^ n1944;
  assign n2227 = n2226 ^ n1956;
  assign n2228 = ~x132 & n2227;
  assign n2229 = n2228 ^ n1956;
  assign n2218 = n1941 ^ n1923;
  assign n2219 = x133 & n2218;
  assign n2220 = n2219 ^ n1941;
  assign n2221 = n2220 ^ n1935;
  assign n2222 = ~x132 & n2221;
  assign n2223 = n2222 ^ n1935;
  assign n2230 = n2229 ^ n2223;
  assign n2231 = ~x134 & n2230;
  assign n2232 = n2231 ^ n2229;
  assign n2239 = n1989 ^ n1965;
  assign n2240 = ~x133 & n2239;
  assign n2241 = n2240 ^ n1989;
  assign n2242 = n2241 ^ n2001;
  assign n2243 = ~x132 & n2242;
  assign n2244 = n2243 ^ n2001;
  assign n2233 = n1986 ^ n1968;
  assign n2234 = x133 & n2233;
  assign n2235 = n2234 ^ n1986;
  assign n2236 = n2235 ^ n1980;
  assign n2237 = ~x132 & n2236;
  assign n2238 = n2237 ^ n1980;
  assign n2245 = n2244 ^ n2238;
  assign n2246 = ~x134 & n2245;
  assign n2247 = n2246 ^ n2244;
  assign n2254 = n507 ^ n273;
  assign n2255 = ~x133 & n2254;
  assign n2256 = n2255 ^ n507;
  assign n2257 = n2256 ^ n2016;
  assign n2258 = ~x132 & n2257;
  assign n2259 = n2258 ^ n2016;
  assign n2248 = n462 ^ n318;
  assign n2249 = x133 & n2248;
  assign n2250 = n2249 ^ n462;
  assign n2251 = n2250 ^ n2010;
  assign n2252 = ~x132 & n2251;
  assign n2253 = n2252 ^ n2010;
  assign n2260 = n2259 ^ n2253;
  assign n2261 = ~x134 & n2260;
  assign n2262 = n2261 ^ n2259;
  assign n2269 = n792 ^ n618;
  assign n2270 = ~x133 & n2269;
  assign n2271 = n2270 ^ n792;
  assign n2272 = n2271 ^ n2031;
  assign n2273 = ~x132 & n2272;
  assign n2274 = n2273 ^ n2031;
  assign n2263 = n759 ^ n651;
  assign n2264 = x133 & n2263;
  assign n2265 = n2264 ^ n759;
  assign n2266 = n2265 ^ n2025;
  assign n2267 = ~x132 & n2266;
  assign n2268 = n2267 ^ n2025;
  assign n2275 = n2274 ^ n2268;
  assign n2276 = ~x134 & n2275;
  assign n2277 = n2276 ^ n2274;
  assign n2284 = n1077 ^ n903;
  assign n2285 = ~x133 & n2284;
  assign n2286 = n2285 ^ n1077;
  assign n2287 = n2286 ^ n2046;
  assign n2288 = ~x132 & n2287;
  assign n2289 = n2288 ^ n2046;
  assign n2278 = n1044 ^ n936;
  assign n2279 = x133 & n2278;
  assign n2280 = n2279 ^ n1044;
  assign n2281 = n2280 ^ n2040;
  assign n2282 = ~x132 & n2281;
  assign n2283 = n2282 ^ n2040;
  assign n2290 = n2289 ^ n2283;
  assign n2291 = ~x134 & n2290;
  assign n2292 = n2291 ^ n2289;
  assign n2299 = n1266 ^ n1152;
  assign n2300 = ~x133 & n2299;
  assign n2301 = n2300 ^ n1266;
  assign n2302 = n2301 ^ n2061;
  assign n2303 = ~x132 & n2302;
  assign n2304 = n2303 ^ n2061;
  assign n2293 = n1245 ^ n1173;
  assign n2294 = x133 & n2293;
  assign n2295 = n2294 ^ n1245;
  assign n2296 = n2295 ^ n2055;
  assign n2297 = ~x132 & n2296;
  assign n2298 = n2297 ^ n2055;
  assign n2305 = n2304 ^ n2298;
  assign n2306 = ~x134 & n2305;
  assign n2307 = n2306 ^ n2304;
  assign n2314 = n1335 ^ n1296;
  assign n2315 = ~x133 & n2314;
  assign n2316 = n2315 ^ n1335;
  assign n2317 = n2316 ^ n2076;
  assign n2318 = ~x132 & n2317;
  assign n2319 = n2318 ^ n2076;
  assign n2308 = n1329 ^ n1302;
  assign n2309 = x133 & n2308;
  assign n2310 = n2309 ^ n1329;
  assign n2311 = n2310 ^ n2070;
  assign n2312 = ~x132 & n2311;
  assign n2313 = n2312 ^ n2070;
  assign n2320 = n2319 ^ n2313;
  assign n2321 = ~x134 & n2320;
  assign n2322 = n2321 ^ n2319;
  assign n2329 = n1404 ^ n1365;
  assign n2330 = ~x133 & n2329;
  assign n2331 = n2330 ^ n1404;
  assign n2332 = n2331 ^ n2091;
  assign n2333 = ~x132 & n2332;
  assign n2334 = n2333 ^ n2091;
  assign n2323 = n1398 ^ n1371;
  assign n2324 = x133 & n2323;
  assign n2325 = n2324 ^ n1398;
  assign n2326 = n2325 ^ n2085;
  assign n2327 = ~x132 & n2326;
  assign n2328 = n2327 ^ n2085;
  assign n2335 = n2334 ^ n2328;
  assign n2336 = ~x134 & n2335;
  assign n2337 = n2336 ^ n2334;
  assign n2344 = n1473 ^ n1434;
  assign n2345 = ~x133 & n2344;
  assign n2346 = n2345 ^ n1473;
  assign n2347 = n2346 ^ n2106;
  assign n2348 = ~x132 & n2347;
  assign n2349 = n2348 ^ n2106;
  assign n2338 = n1467 ^ n1440;
  assign n2339 = x133 & n2338;
  assign n2340 = n2339 ^ n1467;
  assign n2341 = n2340 ^ n2100;
  assign n2342 = ~x132 & n2341;
  assign n2343 = n2342 ^ n2100;
  assign n2350 = n2349 ^ n2343;
  assign n2351 = ~x134 & n2350;
  assign n2352 = n2351 ^ n2349;
  assign n2359 = n1542 ^ n1503;
  assign n2360 = ~x133 & n2359;
  assign n2361 = n2360 ^ n1542;
  assign n2362 = n2361 ^ n2121;
  assign n2363 = ~x132 & n2362;
  assign n2364 = n2363 ^ n2121;
  assign n2353 = n1536 ^ n1509;
  assign n2354 = x133 & n2353;
  assign n2355 = n2354 ^ n1536;
  assign n2356 = n2355 ^ n2115;
  assign n2357 = ~x132 & n2356;
  assign n2358 = n2357 ^ n2115;
  assign n2365 = n2364 ^ n2358;
  assign n2366 = ~x134 & n2365;
  assign n2367 = n2366 ^ n2364;
  assign n2374 = n1611 ^ n1572;
  assign n2375 = ~x133 & n2374;
  assign n2376 = n2375 ^ n1611;
  assign n2377 = n2376 ^ n2136;
  assign n2378 = ~x132 & n2377;
  assign n2379 = n2378 ^ n2136;
  assign n2368 = n1605 ^ n1578;
  assign n2369 = x133 & n2368;
  assign n2370 = n2369 ^ n1605;
  assign n2371 = n2370 ^ n2130;
  assign n2372 = ~x132 & n2371;
  assign n2373 = n2372 ^ n2130;
  assign n2380 = n2379 ^ n2373;
  assign n2381 = ~x134 & n2380;
  assign n2382 = n2381 ^ n2379;
  assign n2389 = n1680 ^ n1641;
  assign n2390 = ~x133 & n2389;
  assign n2391 = n2390 ^ n1680;
  assign n2392 = n2391 ^ n2151;
  assign n2393 = ~x132 & n2392;
  assign n2394 = n2393 ^ n2151;
  assign n2383 = n1674 ^ n1647;
  assign n2384 = x133 & n2383;
  assign n2385 = n2384 ^ n1674;
  assign n2386 = n2385 ^ n2145;
  assign n2387 = ~x132 & n2386;
  assign n2388 = n2387 ^ n2145;
  assign n2395 = n2394 ^ n2388;
  assign n2396 = ~x134 & n2395;
  assign n2397 = n2396 ^ n2394;
  assign n2404 = n1749 ^ n1710;
  assign n2405 = ~x133 & n2404;
  assign n2406 = n2405 ^ n1749;
  assign n2407 = n2406 ^ n2166;
  assign n2408 = ~x132 & n2407;
  assign n2409 = n2408 ^ n2166;
  assign n2398 = n1743 ^ n1716;
  assign n2399 = x133 & n2398;
  assign n2400 = n2399 ^ n1743;
  assign n2401 = n2400 ^ n2160;
  assign n2402 = ~x132 & n2401;
  assign n2403 = n2402 ^ n2160;
  assign n2410 = n2409 ^ n2403;
  assign n2411 = ~x134 & n2410;
  assign n2412 = n2411 ^ n2409;
  assign n2419 = n1818 ^ n1779;
  assign n2420 = ~x133 & n2419;
  assign n2421 = n2420 ^ n1818;
  assign n2422 = n2421 ^ n2181;
  assign n2423 = ~x132 & n2422;
  assign n2424 = n2423 ^ n2181;
  assign n2413 = n1812 ^ n1785;
  assign n2414 = x133 & n2413;
  assign n2415 = n2414 ^ n1812;
  assign n2416 = n2415 ^ n2175;
  assign n2417 = ~x132 & n2416;
  assign n2418 = n2417 ^ n2175;
  assign n2425 = n2424 ^ n2418;
  assign n2426 = ~x134 & n2425;
  assign n2427 = n2426 ^ n2424;
  assign n2434 = n1863 ^ n1839;
  assign n2435 = ~x133 & n2434;
  assign n2436 = n2435 ^ n1863;
  assign n2437 = n2436 ^ n2196;
  assign n2438 = ~x132 & n2437;
  assign n2439 = n2438 ^ n2196;
  assign n2428 = n1860 ^ n1842;
  assign n2429 = x133 & n2428;
  assign n2430 = n2429 ^ n1860;
  assign n2431 = n2430 ^ n2190;
  assign n2432 = ~x132 & n2431;
  assign n2433 = n2432 ^ n2190;
  assign n2440 = n2439 ^ n2433;
  assign n2441 = ~x134 & n2440;
  assign n2442 = n2441 ^ n2439;
  assign n2449 = n1908 ^ n1884;
  assign n2450 = ~x133 & n2449;
  assign n2451 = n2450 ^ n1908;
  assign n2452 = n2451 ^ n2211;
  assign n2453 = ~x132 & n2452;
  assign n2454 = n2453 ^ n2211;
  assign n2443 = n1905 ^ n1887;
  assign n2444 = x133 & n2443;
  assign n2445 = n2444 ^ n1905;
  assign n2446 = n2445 ^ n2205;
  assign n2447 = ~x132 & n2446;
  assign n2448 = n2447 ^ n2205;
  assign n2455 = n2454 ^ n2448;
  assign n2456 = ~x134 & n2455;
  assign n2457 = n2456 ^ n2454;
  assign n2464 = n1953 ^ n1929;
  assign n2465 = ~x133 & n2464;
  assign n2466 = n2465 ^ n1953;
  assign n2467 = n2466 ^ n2226;
  assign n2468 = ~x132 & n2467;
  assign n2469 = n2468 ^ n2226;
  assign n2458 = n1950 ^ n1932;
  assign n2459 = x133 & n2458;
  assign n2460 = n2459 ^ n1950;
  assign n2461 = n2460 ^ n2220;
  assign n2462 = ~x132 & n2461;
  assign n2463 = n2462 ^ n2220;
  assign n2470 = n2469 ^ n2463;
  assign n2471 = ~x134 & n2470;
  assign n2472 = n2471 ^ n2469;
  assign n2479 = n1998 ^ n1974;
  assign n2480 = ~x133 & n2479;
  assign n2481 = n2480 ^ n1998;
  assign n2482 = n2481 ^ n2241;
  assign n2483 = ~x132 & n2482;
  assign n2484 = n2483 ^ n2241;
  assign n2473 = n1995 ^ n1977;
  assign n2474 = x133 & n2473;
  assign n2475 = n2474 ^ n1995;
  assign n2476 = n2475 ^ n2235;
  assign n2477 = ~x132 & n2476;
  assign n2478 = n2477 ^ n2235;
  assign n2485 = n2484 ^ n2478;
  assign n2486 = ~x134 & n2485;
  assign n2487 = n2486 ^ n2484;
  assign n2491 = n2256 ^ n228;
  assign n2492 = x132 & n2491;
  assign n2493 = n2492 ^ n228;
  assign n2488 = n2250 ^ n417;
  assign n2489 = x132 & n2488;
  assign n2490 = n2489 ^ n417;
  assign n2494 = n2493 ^ n2490;
  assign n2495 = ~x134 & n2494;
  assign n2496 = n2495 ^ n2493;
  assign n2500 = n2271 ^ n585;
  assign n2501 = x132 & n2500;
  assign n2502 = n2501 ^ n585;
  assign n2497 = n2265 ^ n726;
  assign n2498 = x132 & n2497;
  assign n2499 = n2498 ^ n726;
  assign n2503 = n2502 ^ n2499;
  assign n2504 = ~x134 & n2503;
  assign n2505 = n2504 ^ n2502;
  assign n2509 = n2286 ^ n870;
  assign n2510 = x132 & n2509;
  assign n2511 = n2510 ^ n870;
  assign n2506 = n2280 ^ n1011;
  assign n2507 = x132 & n2506;
  assign n2508 = n2507 ^ n1011;
  assign n2512 = n2511 ^ n2508;
  assign n2513 = ~x134 & n2512;
  assign n2514 = n2513 ^ n2511;
  assign n2518 = n2301 ^ n1131;
  assign n2519 = x132 & n2518;
  assign n2520 = n2519 ^ n1131;
  assign n2515 = n2295 ^ n1224;
  assign n2516 = x132 & n2515;
  assign n2517 = n2516 ^ n1224;
  assign n2521 = n2520 ^ n2517;
  assign n2522 = ~x134 & n2521;
  assign n2523 = n2522 ^ n2520;
  assign n2527 = n2316 ^ n1290;
  assign n2528 = x132 & n2527;
  assign n2529 = n2528 ^ n1290;
  assign n2524 = n2310 ^ n1323;
  assign n2525 = x132 & n2524;
  assign n2526 = n2525 ^ n1323;
  assign n2530 = n2529 ^ n2526;
  assign n2531 = ~x134 & n2530;
  assign n2532 = n2531 ^ n2529;
  assign n2536 = n2331 ^ n1359;
  assign n2537 = x132 & n2536;
  assign n2538 = n2537 ^ n1359;
  assign n2533 = n2325 ^ n1392;
  assign n2534 = x132 & n2533;
  assign n2535 = n2534 ^ n1392;
  assign n2539 = n2538 ^ n2535;
  assign n2540 = ~x134 & n2539;
  assign n2541 = n2540 ^ n2538;
  assign n2545 = n2346 ^ n1428;
  assign n2546 = x132 & n2545;
  assign n2547 = n2546 ^ n1428;
  assign n2542 = n2340 ^ n1461;
  assign n2543 = x132 & n2542;
  assign n2544 = n2543 ^ n1461;
  assign n2548 = n2547 ^ n2544;
  assign n2549 = ~x134 & n2548;
  assign n2550 = n2549 ^ n2547;
  assign n2554 = n2361 ^ n1497;
  assign n2555 = x132 & n2554;
  assign n2556 = n2555 ^ n1497;
  assign n2551 = n2355 ^ n1530;
  assign n2552 = x132 & n2551;
  assign n2553 = n2552 ^ n1530;
  assign n2557 = n2556 ^ n2553;
  assign n2558 = ~x134 & n2557;
  assign n2559 = n2558 ^ n2556;
  assign n2563 = n2376 ^ n1566;
  assign n2564 = x132 & n2563;
  assign n2565 = n2564 ^ n1566;
  assign n2560 = n2370 ^ n1599;
  assign n2561 = x132 & n2560;
  assign n2562 = n2561 ^ n1599;
  assign n2566 = n2565 ^ n2562;
  assign n2567 = ~x134 & n2566;
  assign n2568 = n2567 ^ n2565;
  assign n2572 = n2391 ^ n1635;
  assign n2573 = x132 & n2572;
  assign n2574 = n2573 ^ n1635;
  assign n2569 = n2385 ^ n1668;
  assign n2570 = x132 & n2569;
  assign n2571 = n2570 ^ n1668;
  assign n2575 = n2574 ^ n2571;
  assign n2576 = ~x134 & n2575;
  assign n2577 = n2576 ^ n2574;
  assign n2581 = n2406 ^ n1704;
  assign n2582 = x132 & n2581;
  assign n2583 = n2582 ^ n1704;
  assign n2578 = n2400 ^ n1737;
  assign n2579 = x132 & n2578;
  assign n2580 = n2579 ^ n1737;
  assign n2584 = n2583 ^ n2580;
  assign n2585 = ~x134 & n2584;
  assign n2586 = n2585 ^ n2583;
  assign n2590 = n2421 ^ n1773;
  assign n2591 = x132 & n2590;
  assign n2592 = n2591 ^ n1773;
  assign n2587 = n2415 ^ n1806;
  assign n2588 = x132 & n2587;
  assign n2589 = n2588 ^ n1806;
  assign n2593 = n2592 ^ n2589;
  assign n2594 = ~x134 & n2593;
  assign n2595 = n2594 ^ n2592;
  assign n2599 = n2436 ^ n1836;
  assign n2600 = x132 & n2599;
  assign n2601 = n2600 ^ n1836;
  assign n2596 = n2430 ^ n1857;
  assign n2597 = x132 & n2596;
  assign n2598 = n2597 ^ n1857;
  assign n2602 = n2601 ^ n2598;
  assign n2603 = ~x134 & n2602;
  assign n2604 = n2603 ^ n2601;
  assign n2608 = n2451 ^ n1881;
  assign n2609 = x132 & n2608;
  assign n2610 = n2609 ^ n1881;
  assign n2605 = n2445 ^ n1902;
  assign n2606 = x132 & n2605;
  assign n2607 = n2606 ^ n1902;
  assign n2611 = n2610 ^ n2607;
  assign n2612 = ~x134 & n2611;
  assign n2613 = n2612 ^ n2610;
  assign n2617 = n2466 ^ n1926;
  assign n2618 = x132 & n2617;
  assign n2619 = n2618 ^ n1926;
  assign n2614 = n2460 ^ n1947;
  assign n2615 = x132 & n2614;
  assign n2616 = n2615 ^ n1947;
  assign n2620 = n2619 ^ n2616;
  assign n2621 = ~x134 & n2620;
  assign n2622 = n2621 ^ n2619;
  assign n2626 = n2481 ^ n1971;
  assign n2627 = x132 & n2626;
  assign n2628 = n2627 ^ n1971;
  assign n2623 = n2475 ^ n1992;
  assign n2624 = x132 & n2623;
  assign n2625 = n2624 ^ n1992;
  assign n2629 = n2628 ^ n2625;
  assign n2630 = ~x134 & n2629;
  assign n2631 = n2630 ^ n2628;
  assign n2632 = x134 & n514;
  assign n2633 = n2632 ^ n513;
  assign n2634 = x134 & n799;
  assign n2635 = n2634 ^ n798;
  assign n2636 = x134 & n1084;
  assign n2637 = n2636 ^ n1083;
  assign n2638 = x134 & n1273;
  assign n2639 = n2638 ^ n1272;
  assign n2640 = x134 & n1342;
  assign n2641 = n2640 ^ n1341;
  assign n2642 = x134 & n1411;
  assign n2643 = n2642 ^ n1410;
  assign n2644 = x134 & n1480;
  assign n2645 = n2644 ^ n1479;
  assign n2646 = x134 & n1549;
  assign n2647 = n2646 ^ n1548;
  assign n2648 = x134 & n1618;
  assign n2649 = n2648 ^ n1617;
  assign n2650 = x134 & n1687;
  assign n2651 = n2650 ^ n1686;
  assign n2652 = x134 & n1756;
  assign n2653 = n2652 ^ n1755;
  assign n2654 = x134 & n1825;
  assign n2655 = n2654 ^ n1824;
  assign n2656 = x134 & n1870;
  assign n2657 = n2656 ^ n1869;
  assign n2658 = x134 & n1915;
  assign n2659 = n2658 ^ n1914;
  assign n2660 = x134 & n1960;
  assign n2661 = n2660 ^ n1959;
  assign n2662 = x134 & n2005;
  assign n2663 = n2662 ^ n2004;
  assign n2664 = x134 & n2020;
  assign n2665 = n2664 ^ n2019;
  assign n2666 = x134 & n2035;
  assign n2667 = n2666 ^ n2034;
  assign n2668 = x134 & n2050;
  assign n2669 = n2668 ^ n2049;
  assign n2670 = x134 & n2065;
  assign n2671 = n2670 ^ n2064;
  assign n2672 = x134 & n2080;
  assign n2673 = n2672 ^ n2079;
  assign n2674 = x134 & n2095;
  assign n2675 = n2674 ^ n2094;
  assign n2676 = x134 & n2110;
  assign n2677 = n2676 ^ n2109;
  assign n2678 = x134 & n2125;
  assign n2679 = n2678 ^ n2124;
  assign n2680 = x134 & n2140;
  assign n2681 = n2680 ^ n2139;
  assign n2682 = x134 & n2155;
  assign n2683 = n2682 ^ n2154;
  assign n2684 = x134 & n2170;
  assign n2685 = n2684 ^ n2169;
  assign n2686 = x134 & n2185;
  assign n2687 = n2686 ^ n2184;
  assign n2688 = x134 & n2200;
  assign n2689 = n2688 ^ n2199;
  assign n2690 = x134 & n2215;
  assign n2691 = n2690 ^ n2214;
  assign n2692 = x134 & n2230;
  assign n2693 = n2692 ^ n2229;
  assign n2694 = x134 & n2245;
  assign n2695 = n2694 ^ n2244;
  assign n2696 = x134 & n2260;
  assign n2697 = n2696 ^ n2259;
  assign n2698 = x134 & n2275;
  assign n2699 = n2698 ^ n2274;
  assign n2700 = x134 & n2290;
  assign n2701 = n2700 ^ n2289;
  assign n2702 = x134 & n2305;
  assign n2703 = n2702 ^ n2304;
  assign n2704 = x134 & n2320;
  assign n2705 = n2704 ^ n2319;
  assign n2706 = x134 & n2335;
  assign n2707 = n2706 ^ n2334;
  assign n2708 = x134 & n2350;
  assign n2709 = n2708 ^ n2349;
  assign n2710 = x134 & n2365;
  assign n2711 = n2710 ^ n2364;
  assign n2712 = x134 & n2380;
  assign n2713 = n2712 ^ n2379;
  assign n2714 = x134 & n2395;
  assign n2715 = n2714 ^ n2394;
  assign n2716 = x134 & n2410;
  assign n2717 = n2716 ^ n2409;
  assign n2718 = x134 & n2425;
  assign n2719 = n2718 ^ n2424;
  assign n2720 = x134 & n2440;
  assign n2721 = n2720 ^ n2439;
  assign n2722 = x134 & n2455;
  assign n2723 = n2722 ^ n2454;
  assign n2724 = x134 & n2470;
  assign n2725 = n2724 ^ n2469;
  assign n2726 = x134 & n2485;
  assign n2727 = n2726 ^ n2484;
  assign n2728 = x134 & n2494;
  assign n2729 = n2728 ^ n2493;
  assign n2730 = x134 & n2503;
  assign n2731 = n2730 ^ n2502;
  assign n2732 = x134 & n2512;
  assign n2733 = n2732 ^ n2511;
  assign n2734 = x134 & n2521;
  assign n2735 = n2734 ^ n2520;
  assign n2736 = x134 & n2530;
  assign n2737 = n2736 ^ n2529;
  assign n2738 = x134 & n2539;
  assign n2739 = n2738 ^ n2538;
  assign n2740 = x134 & n2548;
  assign n2741 = n2740 ^ n2547;
  assign n2742 = x134 & n2557;
  assign n2743 = n2742 ^ n2556;
  assign n2744 = x134 & n2566;
  assign n2745 = n2744 ^ n2565;
  assign n2746 = x134 & n2575;
  assign n2747 = n2746 ^ n2574;
  assign n2748 = x134 & n2584;
  assign n2749 = n2748 ^ n2583;
  assign n2750 = x134 & n2593;
  assign n2751 = n2750 ^ n2592;
  assign n2752 = x134 & n2602;
  assign n2753 = n2752 ^ n2601;
  assign n2754 = x134 & n2611;
  assign n2755 = n2754 ^ n2610;
  assign n2756 = x134 & n2620;
  assign n2757 = n2756 ^ n2619;
  assign n2758 = x134 & n2629;
  assign n2759 = n2758 ^ n2628;
  assign y0 = n516;
  assign y1 = n801;
  assign y2 = n1086;
  assign y3 = n1275;
  assign y4 = n1344;
  assign y5 = n1413;
  assign y6 = n1482;
  assign y7 = n1551;
  assign y8 = n1620;
  assign y9 = n1689;
  assign y10 = n1758;
  assign y11 = n1827;
  assign y12 = n1872;
  assign y13 = n1917;
  assign y14 = n1962;
  assign y15 = n2007;
  assign y16 = n2022;
  assign y17 = n2037;
  assign y18 = n2052;
  assign y19 = n2067;
  assign y20 = n2082;
  assign y21 = n2097;
  assign y22 = n2112;
  assign y23 = n2127;
  assign y24 = n2142;
  assign y25 = n2157;
  assign y26 = n2172;
  assign y27 = n2187;
  assign y28 = n2202;
  assign y29 = n2217;
  assign y30 = n2232;
  assign y31 = n2247;
  assign y32 = n2262;
  assign y33 = n2277;
  assign y34 = n2292;
  assign y35 = n2307;
  assign y36 = n2322;
  assign y37 = n2337;
  assign y38 = n2352;
  assign y39 = n2367;
  assign y40 = n2382;
  assign y41 = n2397;
  assign y42 = n2412;
  assign y43 = n2427;
  assign y44 = n2442;
  assign y45 = n2457;
  assign y46 = n2472;
  assign y47 = n2487;
  assign y48 = n2496;
  assign y49 = n2505;
  assign y50 = n2514;
  assign y51 = n2523;
  assign y52 = n2532;
  assign y53 = n2541;
  assign y54 = n2550;
  assign y55 = n2559;
  assign y56 = n2568;
  assign y57 = n2577;
  assign y58 = n2586;
  assign y59 = n2595;
  assign y60 = n2604;
  assign y61 = n2613;
  assign y62 = n2622;
  assign y63 = n2631;
  assign y64 = n2633;
  assign y65 = n2635;
  assign y66 = n2637;
  assign y67 = n2639;
  assign y68 = n2641;
  assign y69 = n2643;
  assign y70 = n2645;
  assign y71 = n2647;
  assign y72 = n2649;
  assign y73 = n2651;
  assign y74 = n2653;
  assign y75 = n2655;
  assign y76 = n2657;
  assign y77 = n2659;
  assign y78 = n2661;
  assign y79 = n2663;
  assign y80 = n2665;
  assign y81 = n2667;
  assign y82 = n2669;
  assign y83 = n2671;
  assign y84 = n2673;
  assign y85 = n2675;
  assign y86 = n2677;
  assign y87 = n2679;
  assign y88 = n2681;
  assign y89 = n2683;
  assign y90 = n2685;
  assign y91 = n2687;
  assign y92 = n2689;
  assign y93 = n2691;
  assign y94 = n2693;
  assign y95 = n2695;
  assign y96 = n2697;
  assign y97 = n2699;
  assign y98 = n2701;
  assign y99 = n2703;
  assign y100 = n2705;
  assign y101 = n2707;
  assign y102 = n2709;
  assign y103 = n2711;
  assign y104 = n2713;
  assign y105 = n2715;
  assign y106 = n2717;
  assign y107 = n2719;
  assign y108 = n2721;
  assign y109 = n2723;
  assign y110 = n2725;
  assign y111 = n2727;
  assign y112 = n2729;
  assign y113 = n2731;
  assign y114 = n2733;
  assign y115 = n2735;
  assign y116 = n2737;
  assign y117 = n2739;
  assign y118 = n2741;
  assign y119 = n2743;
  assign y120 = n2745;
  assign y121 = n2747;
  assign y122 = n2749;
  assign y123 = n2751;
  assign y124 = n2753;
  assign y125 = n2755;
  assign y126 = n2757;
  assign y127 = n2759;
endmodule
