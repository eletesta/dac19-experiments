module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10;
  wire n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564;
  assign n11 = ~x5 & ~x6;
  assign n20 = ~x0 & x7;
  assign n21 = ~x2 & ~x8;
  assign n22 = x2 & x8;
  assign n23 = ~x9 & n22;
  assign n24 = ~n21 & ~n23;
  assign n25 = n20 & ~n24;
  assign n26 = x0 & x9;
  assign n27 = ~x2 & x8;
  assign n28 = n26 & n27;
  assign n29 = ~n25 & ~n28;
  assign n30 = ~x3 & ~n29;
  assign n31 = x8 & x9;
  assign n32 = x2 & ~x3;
  assign n33 = n31 & n32;
  assign n34 = ~x8 & ~x9;
  assign n35 = ~x2 & x3;
  assign n36 = n34 & n35;
  assign n37 = ~n33 & ~n36;
  assign n38 = ~x0 & ~n37;
  assign n39 = x3 & ~x9;
  assign n40 = x2 & ~n39;
  assign n41 = x0 & ~n35;
  assign n42 = ~n34 & n41;
  assign n43 = ~n40 & n42;
  assign n44 = ~n38 & ~n43;
  assign n45 = ~x7 & ~n44;
  assign n46 = ~n30 & ~n45;
  assign n47 = ~x1 & ~n46;
  assign n12 = ~x7 & ~x8;
  assign n13 = ~x2 & ~x3;
  assign n14 = ~x7 & ~x9;
  assign n15 = n13 & ~n14;
  assign n16 = ~x8 & x9;
  assign n17 = n16 ^ x0;
  assign n18 = n15 & n17;
  assign n19 = ~n12 & ~n18;
  assign n48 = n47 ^ n19;
  assign n49 = n11 & ~n48;
  assign n50 = ~x1 & ~x8;
  assign n51 = ~x3 & ~n50;
  assign n52 = ~x1 & x2;
  assign n53 = x8 & ~n52;
  assign n54 = x0 & ~n53;
  assign n55 = ~n51 & n54;
  assign n56 = ~x3 & ~n22;
  assign n57 = ~x8 & ~n52;
  assign n58 = ~n56 & ~n57;
  assign n59 = ~x1 & x8;
  assign n60 = ~x0 & ~n59;
  assign n61 = ~n58 & n60;
  assign n62 = ~x5 & ~x9;
  assign n63 = ~n61 & n62;
  assign n64 = ~n55 & n63;
  assign n65 = ~x5 & x8;
  assign n66 = x0 & x1;
  assign n67 = x8 & n66;
  assign n68 = ~x1 & ~x2;
  assign n69 = ~x5 & n68;
  assign n70 = x5 & ~x8;
  assign n71 = ~n13 & ~n70;
  assign n72 = ~n69 & n71;
  assign n73 = ~n67 & ~n72;
  assign n74 = ~n65 & ~n73;
  assign n75 = ~x5 & ~n35;
  assign n76 = ~x0 & ~x1;
  assign n77 = ~n70 & n76;
  assign n78 = ~n75 & n77;
  assign n79 = n31 & ~n32;
  assign n80 = x5 & x9;
  assign n81 = ~n26 & ~n80;
  assign n82 = ~n79 & n81;
  assign n83 = ~n78 & ~n82;
  assign n84 = ~n74 & n83;
  assign n85 = n13 & n76;
  assign n86 = x5 & n34;
  assign n87 = ~n85 & n86;
  assign n88 = x6 & ~x7;
  assign n89 = ~n87 & n88;
  assign n90 = ~n84 & n89;
  assign n91 = ~n64 & n90;
  assign n92 = x0 & ~x1;
  assign n93 = ~x1 & x9;
  assign n94 = n93 ^ x2;
  assign n95 = n92 & n94;
  assign n96 = n56 & ~n95;
  assign n97 = x0 & ~x2;
  assign n98 = ~x9 & n97;
  assign n99 = x2 & n16;
  assign n100 = ~n98 & ~n99;
  assign n101 = x1 & ~n100;
  assign n102 = x3 & ~n27;
  assign n103 = ~n101 & n102;
  assign n104 = ~n96 & ~n103;
  assign n105 = x9 ^ x0;
  assign n106 = x1 & ~n105;
  assign n107 = x8 & ~n106;
  assign n108 = x5 & ~x6;
  assign n109 = ~x7 & n108;
  assign n110 = ~n107 & n109;
  assign n111 = ~n104 & n110;
  assign n112 = ~n91 & ~n111;
  assign n113 = ~n49 & n112;
  assign n114 = ~x4 & ~n34;
  assign n115 = n85 & n114;
  assign n116 = x4 & ~n85;
  assign n117 = x6 ^ x5;
  assign n118 = x4 & n34;
  assign n119 = ~n117 & n118;
  assign n120 = ~n116 & ~n119;
  assign n121 = ~n115 & n120;
  assign n122 = ~n113 & n121;
  assign n138 = n22 & n92;
  assign n139 = n21 & n76;
  assign n140 = n14 & ~n139;
  assign n141 = ~n138 & n140;
  assign n123 = ~x3 & ~x9;
  assign n124 = ~x0 & x8;
  assign n125 = x1 & ~x2;
  assign n126 = n124 & n125;
  assign n127 = ~x7 & x8;
  assign n128 = ~n21 & ~n127;
  assign n129 = n92 & ~n128;
  assign n130 = ~n126 & ~n129;
  assign n131 = n123 & ~n130;
  assign n132 = ~n76 & ~n97;
  assign n133 = ~x3 & ~n68;
  assign n134 = n31 ^ x7;
  assign n135 = n133 & n134;
  assign n136 = ~n132 & n135;
  assign n137 = ~n131 & ~n136;
  assign n142 = n141 ^ n137;
  assign n143 = n11 & ~n142;
  assign n144 = ~x1 & ~x5;
  assign n145 = x9 ^ x3;
  assign n146 = x8 & n145;
  assign n147 = x0 & ~n34;
  assign n148 = ~x3 & ~n147;
  assign n149 = ~n146 & ~n148;
  assign n150 = n144 & ~n149;
  assign n151 = x1 & ~n145;
  assign n152 = ~x9 & ~n65;
  assign n153 = n151 & ~n152;
  assign n154 = x2 & ~n80;
  assign n155 = ~n153 & n154;
  assign n156 = ~n150 & n155;
  assign n157 = n13 & n66;
  assign n158 = ~x2 & ~n62;
  assign n159 = ~n157 & ~n158;
  assign n160 = x1 & ~n124;
  assign n161 = n80 & n160;
  assign n162 = ~n159 & ~n161;
  assign n163 = ~x3 & ~n76;
  assign n164 = n16 & n66;
  assign n165 = n163 & ~n164;
  assign n166 = n16 & n92;
  assign n167 = x3 & ~n80;
  assign n168 = ~n166 & n167;
  assign n169 = ~n165 & ~n168;
  assign n170 = n162 & ~n169;
  assign n171 = n88 & ~n170;
  assign n172 = ~n156 & n171;
  assign n173 = ~x3 & n138;
  assign n174 = x2 & x3;
  assign n175 = n16 & n174;
  assign n176 = ~n123 & ~n175;
  assign n177 = x1 & ~n176;
  assign n178 = ~n173 & ~n177;
  assign n179 = ~n31 & ~n93;
  assign n180 = x9 & ~n13;
  assign n181 = n179 & ~n180;
  assign n182 = ~x0 & n181;
  assign n183 = x1 & ~n27;
  assign n184 = ~x9 & ~n32;
  assign n185 = ~n183 & n184;
  assign n186 = ~n182 & ~n185;
  assign n187 = n178 & n186;
  assign n188 = n109 & ~n187;
  assign n189 = ~n172 & ~n188;
  assign n190 = ~n143 & n189;
  assign n191 = ~x0 & ~x6;
  assign n192 = ~x9 & ~n191;
  assign n193 = ~x3 & n68;
  assign n194 = ~n192 & n193;
  assign n195 = x4 & ~n194;
  assign n196 = ~n115 & ~n195;
  assign n197 = ~n190 & n196;
  assign n198 = ~x5 & x6;
  assign n199 = ~x6 & x9;
  assign n200 = ~n198 & ~n199;
  assign n201 = n59 & ~n200;
  assign n202 = ~n23 & n65;
  assign n203 = ~n124 & ~n202;
  assign n204 = ~n201 & n203;
  assign n205 = x2 & ~x5;
  assign n206 = ~x2 & ~x6;
  assign n207 = ~n205 & ~n206;
  assign n208 = ~x1 & n207;
  assign n209 = x1 & ~x9;
  assign n210 = n205 & n209;
  assign n211 = x5 & x6;
  assign n212 = ~x0 & ~n211;
  assign n213 = ~n158 & n212;
  assign n214 = ~n210 & n213;
  assign n215 = ~n208 & n214;
  assign n216 = ~n204 & ~n215;
  assign n217 = x1 & x6;
  assign n218 = ~x0 & n217;
  assign n219 = n205 & n218;
  assign n220 = n26 & ~n217;
  assign n221 = ~n219 & ~n220;
  assign n222 = x5 & n209;
  assign n223 = ~n207 & ~n222;
  assign n224 = x0 & ~n223;
  assign n225 = ~x0 & ~x9;
  assign n226 = ~n207 & n225;
  assign n227 = ~x8 & ~n226;
  assign n228 = ~n224 & n227;
  assign n229 = n221 & n228;
  assign n230 = ~n216 & ~n229;
  assign n231 = x3 & ~x4;
  assign n232 = ~n230 & n231;
  assign n233 = ~x2 & n76;
  assign n234 = ~x8 & n198;
  assign n235 = n233 & ~n234;
  assign n236 = n235 ^ x4;
  assign n237 = ~x3 & ~n236;
  assign n238 = ~n232 & ~n237;
  assign n272 = x1 & x9;
  assign n273 = x6 ^ x2;
  assign n274 = x8 ^ x6;
  assign n275 = n273 & n274;
  assign n276 = n275 ^ x2;
  assign n277 = n272 & ~n276;
  assign n278 = ~x0 & ~n277;
  assign n279 = ~x3 & x9;
  assign n280 = x0 & ~n21;
  assign n281 = n279 & ~n280;
  assign n266 = x1 & ~x6;
  assign n282 = x8 & ~x9;
  assign n283 = n266 & ~n282;
  assign n249 = x2 & ~x6;
  assign n284 = ~x3 & ~n249;
  assign n285 = ~n283 & n284;
  assign n286 = ~n281 & ~n285;
  assign n287 = ~n278 & ~n286;
  assign n288 = ~x7 & ~n287;
  assign n239 = n125 & n147;
  assign n240 = ~x6 & x8;
  assign n241 = ~x1 & ~n240;
  assign n242 = n98 & n241;
  assign n243 = ~x0 & x2;
  assign n244 = n31 & n243;
  assign n245 = ~n242 & ~n244;
  assign n246 = ~n239 & n245;
  assign n247 = ~x8 & ~n191;
  assign n248 = ~n206 & ~n247;
  assign n250 = x0 & ~n249;
  assign n251 = n209 & ~n250;
  assign n252 = ~n248 & n251;
  assign n253 = ~x9 & ~n22;
  assign n254 = ~x6 & ~n31;
  assign n255 = n76 & ~n254;
  assign n256 = ~n253 & n255;
  assign n257 = ~n252 & ~n256;
  assign n258 = n246 & n257;
  assign n259 = ~x5 & ~x7;
  assign n260 = x0 & n209;
  assign n261 = n11 & ~n16;
  assign n262 = ~n260 & n261;
  assign n263 = ~n259 & ~n262;
  assign n264 = ~x3 & ~n20;
  assign n265 = ~n123 & ~n264;
  assign n267 = ~x0 & n14;
  assign n268 = n266 & n267;
  assign n269 = ~n265 & ~n268;
  assign n270 = ~n263 & n269;
  assign n271 = ~n258 & n270;
  assign n289 = n288 ^ n271;
  assign n290 = ~n238 & n289;
  assign n291 = ~x0 & x5;
  assign n292 = ~n240 & n291;
  assign n293 = ~x5 & ~n282;
  assign n294 = x0 & ~n199;
  assign n295 = n293 & n294;
  assign n296 = ~n292 & ~n295;
  assign n297 = x1 & ~n296;
  assign n298 = x0 & x5;
  assign n299 = x1 & ~n298;
  assign n300 = ~x6 & n31;
  assign n301 = ~n299 & n300;
  assign n302 = n92 & ~n108;
  assign n303 = ~n293 & n302;
  assign n304 = ~n301 & ~n303;
  assign n305 = ~n297 & n304;
  assign n306 = ~n94 & ~n211;
  assign n307 = x3 & ~n306;
  assign n308 = ~n305 & n307;
  assign n309 = x2 & ~n34;
  assign n310 = x9 ^ x8;
  assign n311 = ~x2 & ~n310;
  assign n312 = x1 & ~n311;
  assign n313 = ~n309 & n312;
  assign n314 = ~x6 & n68;
  assign n315 = n34 & n314;
  assign n316 = ~n217 & ~n315;
  assign n317 = ~n313 & n316;
  assign n318 = n298 & ~n317;
  assign n319 = ~n93 & ~n124;
  assign n320 = x6 & ~n209;
  assign n321 = ~n319 & n320;
  assign n322 = ~x5 & ~n321;
  assign n323 = n31 & n76;
  assign n324 = ~x6 & ~n323;
  assign n325 = ~n249 & ~n324;
  assign n326 = n322 & n325;
  assign n327 = n22 & n272;
  assign n328 = ~x6 & ~n327;
  assign n329 = ~n217 & n291;
  assign n330 = x2 & n198;
  assign n331 = ~n329 & ~n330;
  assign n332 = ~n328 & ~n331;
  assign n333 = ~n124 & n210;
  assign n334 = ~x3 & ~n333;
  assign n335 = ~n332 & n334;
  assign n336 = ~n326 & n335;
  assign n337 = ~n318 & n336;
  assign n338 = ~n117 & n193;
  assign n339 = n338 ^ x4;
  assign n340 = ~x7 & ~n339;
  assign n341 = ~n337 & n340;
  assign n342 = ~n308 & n341;
  assign n343 = ~x7 & n211;
  assign n344 = n193 ^ x4;
  assign n345 = n233 & ~n344;
  assign n346 = x2 & ~x4;
  assign n347 = ~n76 & n346;
  assign n348 = ~n345 & ~n347;
  assign n349 = n343 & ~n348;
  assign n350 = n231 & ~n233;
  assign n351 = x4 & n85;
  assign n352 = ~n350 & ~n351;
  assign n353 = n343 & ~n352;
  assign n354 = ~x3 & ~x4;
  assign n378 = ~x7 & ~n327;
  assign n379 = x5 & ~n378;
  assign n380 = ~x2 & n259;
  assign n381 = n199 & n380;
  assign n382 = ~n379 & ~n381;
  assign n383 = ~n34 & n380;
  assign n384 = x6 & ~n383;
  assign n385 = x0 & ~n384;
  assign n386 = n382 & n385;
  assign n387 = ~x7 & ~n34;
  assign n388 = x2 & ~n387;
  assign n389 = n14 & n65;
  assign n367 = x7 & ~x8;
  assign n390 = x1 & ~n367;
  assign n391 = ~n389 & n390;
  assign n392 = ~n388 & n391;
  assign n393 = ~x2 & ~n14;
  assign n394 = ~n86 & ~n393;
  assign n395 = x7 & n31;
  assign n396 = ~x1 & ~n395;
  assign n397 = n394 & n396;
  assign n398 = ~n392 & ~n397;
  assign n399 = n386 & ~n398;
  assign n355 = n62 & ~n217;
  assign n356 = n127 & ~n355;
  assign n357 = x2 & ~n356;
  assign n358 = x5 & ~n266;
  assign n359 = ~n272 & ~n358;
  assign n360 = ~x7 & ~n359;
  assign n361 = ~x5 & ~n31;
  assign n362 = ~x1 & ~x6;
  assign n363 = ~n127 & n362;
  assign n364 = n361 & n363;
  assign n365 = ~n360 & ~n364;
  assign n366 = n357 & n365;
  assign n368 = ~x1 & n11;
  assign n369 = ~n367 & n368;
  assign n370 = ~n11 & ~n12;
  assign n371 = ~x9 & ~n370;
  assign n372 = ~n369 & n371;
  assign n373 = n12 & n217;
  assign n374 = ~x2 & ~n343;
  assign n375 = ~n373 & n374;
  assign n376 = ~n372 & n375;
  assign n377 = ~n366 & ~n376;
  assign n400 = n399 ^ n377;
  assign n401 = n354 & n400;
  assign n402 = ~n66 & n70;
  assign n403 = ~n125 & n402;
  assign n404 = ~n98 & n403;
  assign n405 = n93 & n243;
  assign n406 = x5 & x8;
  assign n407 = ~n209 & n406;
  assign n408 = ~n405 & n407;
  assign n409 = ~x4 & ~n408;
  assign n410 = ~n404 & n409;
  assign n411 = ~n211 & ~n410;
  assign n412 = ~n22 & ~n199;
  assign n413 = x0 & ~n412;
  assign n414 = ~x1 & ~n16;
  assign n415 = ~x2 & x6;
  assign n416 = n225 ^ n124;
  assign n417 = n415 & n416;
  assign n418 = n417 ^ n225;
  assign n419 = n414 & ~n418;
  assign n420 = ~n413 & n419;
  assign n421 = ~x0 & n31;
  assign n422 = ~n276 & n421;
  assign n423 = ~x2 & ~n124;
  assign n424 = n192 & n423;
  assign n425 = x1 & ~n424;
  assign n426 = ~n422 & n425;
  assign n427 = ~n420 & ~n426;
  assign n428 = ~x5 & n427;
  assign n429 = ~n411 & ~n428;
  assign n430 = ~n351 & ~n429;
  assign n431 = ~x7 & ~n354;
  assign n432 = ~n430 & n431;
  assign n433 = ~n401 & ~n432;
  assign n434 = ~n51 & ~n59;
  assign n435 = ~n179 & n434;
  assign n436 = x8 & n106;
  assign n437 = ~x3 & ~n436;
  assign n438 = ~n76 & ~n421;
  assign n439 = ~n437 & n438;
  assign n440 = ~n435 & n439;
  assign n441 = ~x2 & ~n440;
  assign n442 = n22 & n145;
  assign n443 = x0 & ~x8;
  assign n444 = ~n279 & n443;
  assign n445 = ~n35 & n444;
  assign n446 = ~n442 & ~n445;
  assign n447 = x1 & ~n446;
  assign n448 = n310 & n362;
  assign n449 = ~x0 & n13;
  assign n450 = n449 ^ x3;
  assign n451 = n448 & ~n450;
  assign n452 = n108 & ~n451;
  assign n453 = ~n447 & n452;
  assign n454 = ~n441 & n453;
  assign n471 = n34 & n163;
  assign n472 = ~n59 & n179;
  assign n473 = ~n471 & n472;
  assign n474 = ~n93 & n147;
  assign n475 = ~n473 & ~n474;
  assign n476 = ~x2 & ~n475;
  assign n477 = ~x0 & x3;
  assign n478 = ~n310 & n477;
  assign n479 = ~n309 & ~n478;
  assign n480 = ~x1 & ~n479;
  assign n481 = ~n33 & ~n480;
  assign n482 = ~n476 & n481;
  assign n483 = ~x4 & ~n482;
  assign n455 = x1 & ~n39;
  assign n456 = ~n243 & ~n279;
  assign n457 = n455 & ~n456;
  assign n458 = x3 & ~n93;
  assign n459 = n97 & ~n458;
  assign n460 = ~n457 & ~n459;
  assign n461 = x8 & ~n460;
  assign n462 = n32 & n272;
  assign n463 = ~n56 & ~n225;
  assign n464 = x3 & ~n21;
  assign n465 = ~x1 & ~n464;
  assign n466 = ~n463 & n465;
  assign n467 = ~n462 & ~n466;
  assign n468 = ~n461 & n467;
  assign n469 = ~x4 & ~n468;
  assign n470 = ~x6 & ~n469;
  assign n484 = n483 ^ n470;
  assign n485 = ~x5 & n484;
  assign n486 = ~n454 & ~n485;
  assign n487 = x7 & ~n451;
  assign n488 = n14 & n27;
  assign n489 = ~n367 & ~n488;
  assign n490 = x0 & n362;
  assign n491 = ~n489 & n490;
  assign n492 = ~n487 & ~n491;
  assign n493 = ~n116 & n492;
  assign n494 = ~n486 & n493;
  assign n495 = n259 & n351;
  assign n496 = ~n11 & ~n254;
  assign n497 = ~n26 & ~n222;
  assign n498 = n92 & ~n282;
  assign n499 = n319 & ~n498;
  assign n500 = n497 & n499;
  assign n501 = ~x2 & ~n500;
  assign n502 = ~x1 & ~n253;
  assign n503 = ~n361 & n502;
  assign n504 = n334 & ~n503;
  assign n505 = ~n501 & n504;
  assign n506 = ~n496 & n505;
  assign n507 = ~n76 & n472;
  assign n508 = n35 & n108;
  assign n509 = ~n323 & n508;
  assign n510 = ~n507 & n509;
  assign n511 = ~n233 & ~n362;
  assign n512 = ~x9 & ~n247;
  assign n513 = ~n511 & n512;
  assign n514 = x9 & n273;
  assign n515 = ~n160 & n514;
  assign n516 = ~n59 & n206;
  assign n517 = x3 & ~x5;
  assign n518 = ~n516 & n517;
  assign n519 = ~n515 & n518;
  assign n520 = ~n513 & n519;
  assign n521 = ~n510 & ~n520;
  assign n522 = ~n506 & n521;
  assign n523 = n11 & ~n31;
  assign n524 = ~x2 & ~n209;
  assign n525 = n76 & n309;
  assign n526 = ~n524 & ~n525;
  assign n527 = n523 & ~n526;
  assign n528 = x7 & ~n527;
  assign n529 = ~x4 & ~n528;
  assign n530 = ~n522 & n529;
  assign n531 = ~n495 & ~n530;
  assign n532 = ~n322 & ~n324;
  assign n533 = ~x1 & ~n34;
  assign n534 = n438 & ~n533;
  assign n535 = n11 & n534;
  assign n536 = ~n532 & ~n535;
  assign n537 = x5 ^ x2;
  assign n538 = n537 ^ x6;
  assign n539 = n211 & ~n538;
  assign n540 = n539 ^ n538;
  assign n541 = ~n536 & n540;
  assign n542 = x3 & ~x7;
  assign n543 = ~n541 & n542;
  assign n544 = n249 & n472;
  assign n545 = ~n11 & ~n68;
  assign n546 = ~n544 & n545;
  assign n547 = ~x9 & ~n124;
  assign n548 = n125 & ~n547;
  assign n549 = ~x2 & n92;
  assign n550 = ~x7 & ~n549;
  assign n551 = ~n548 & n550;
  assign n552 = ~n525 & ~n551;
  assign n553 = n22 & n93;
  assign n554 = ~x3 & ~n553;
  assign n555 = ~n338 & n554;
  assign n556 = ~n552 & n555;
  assign n557 = ~n546 & n556;
  assign n558 = ~n543 & ~n557;
  assign n559 = ~n344 & ~n558;
  assign n560 = n174 & n534;
  assign n561 = ~x4 & ~n560;
  assign n562 = ~x7 & n11;
  assign n563 = ~n116 & n562;
  assign n564 = ~n561 & n563;
  assign y0 = n122;
  assign y1 = n197;
  assign y2 = n290;
  assign y3 = n342;
  assign y4 = n349;
  assign y5 = n353;
  assign y6 = n433;
  assign y7 = ~n494;
  assign y8 = n531;
  assign y9 = n559;
  assign y10 = n564;
endmodule
