// Benchmark "top" written by ABC on Mon Nov 19 13:33:21 2018

module top ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127,
    po0, po1, po2, po3, po4, po5, po6, po7  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n448, n449, n450,
    n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
    n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
    n475, n476, n477, n479, n480, n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n495, n496, n499, n500, n501, n502, n503,
    n504;
  assign n138 = pi001 & ~pi002;
  assign n139 = ~n138 & ~pi003;
  assign n140 = ~n139 & ~pi004;
  assign n141 = ~n140 & ~pi005;
  assign n142 = ~n141 & ~pi006;
  assign n143 = ~n142 & ~pi007;
  assign n144 = ~n143 & ~pi008;
  assign n145 = ~n144 & ~pi009;
  assign n146 = ~n145 & ~pi010;
  assign n147 = ~n146 & ~pi011;
  assign n148 = ~n147 & ~pi012;
  assign n149 = ~n148 & ~pi013;
  assign n150 = ~n149 & ~pi014;
  assign n151 = ~n150 & ~pi015;
  assign n152 = ~n151 & ~pi016;
  assign n153 = ~n152 & ~pi017;
  assign n154 = ~n153 & ~pi018;
  assign n155 = ~n154 & ~pi019;
  assign n156 = ~n155 & ~pi020;
  assign n157 = ~n156 & ~pi021;
  assign n158 = ~n157 & ~pi022;
  assign n159 = ~n158 & ~pi023;
  assign n160 = ~n159 & ~pi024;
  assign n161 = ~n160 & ~pi025;
  assign n162 = ~n161 & ~pi026;
  assign n163 = ~n162 & ~pi027;
  assign n164 = ~n163 & ~pi028;
  assign n165 = ~n164 & ~pi029;
  assign n166 = ~n165 & ~pi030;
  assign n167 = ~n166 & ~pi031;
  assign n168 = ~n167 & ~pi032;
  assign n169 = ~n168 & ~pi033;
  assign n170 = ~n169 & ~pi034;
  assign n171 = ~n170 & ~pi035;
  assign n172 = ~n171 & ~pi036;
  assign n173 = ~n172 & ~pi037;
  assign n174 = ~n173 & ~pi038;
  assign n175 = ~n174 & ~pi039;
  assign n176 = ~n175 & ~pi040;
  assign n177 = ~n176 & ~pi041;
  assign n178 = ~n177 & ~pi042;
  assign n179 = ~n178 & ~pi043;
  assign n180 = ~n179 & ~pi044;
  assign n181 = ~n180 & ~pi045;
  assign n182 = ~n181 & ~pi046;
  assign n183 = ~n182 & ~pi047;
  assign n184 = ~n183 & ~pi048;
  assign n185 = ~n184 & ~pi049;
  assign n186 = ~n185 & ~pi050;
  assign n187 = ~n186 & ~pi051;
  assign n188 = ~n187 & ~pi052;
  assign n189 = ~n188 & ~pi053;
  assign n190 = ~n189 & ~pi054;
  assign n191 = ~n190 & ~pi055;
  assign n192 = ~n191 & ~pi056;
  assign n193 = ~n192 & ~pi057;
  assign n194 = ~n193 & ~pi058;
  assign n195 = ~n194 & ~pi059;
  assign n196 = ~n195 & ~pi060;
  assign n197 = ~n196 & ~pi061;
  assign n198 = ~n197 & ~pi062;
  assign n199 = ~n198 & ~pi063;
  assign n200 = ~n199 & ~pi064;
  assign n201 = ~n200 & ~pi065;
  assign n202 = ~n201 & ~pi066;
  assign n203 = ~n202 & ~pi067;
  assign n204 = ~n203 & ~pi068;
  assign n205 = ~n204 & ~pi069;
  assign n206 = ~n205 & ~pi070;
  assign n207 = ~n206 & ~pi071;
  assign n208 = ~n207 & ~pi072;
  assign n209 = ~n208 & ~pi073;
  assign n210 = ~n209 & ~pi074;
  assign n211 = ~n210 & ~pi075;
  assign n212 = ~n211 & ~pi076;
  assign n213 = ~n212 & ~pi077;
  assign n214 = ~n213 & ~pi078;
  assign n215 = ~n214 & ~pi079;
  assign n216 = ~n215 & ~pi080;
  assign n217 = ~n216 & ~pi081;
  assign n218 = ~n217 & ~pi082;
  assign n219 = ~n218 & ~pi083;
  assign n220 = ~n219 & ~pi084;
  assign n221 = ~n220 & ~pi085;
  assign n222 = ~n221 & ~pi086;
  assign n223 = ~n222 & ~pi087;
  assign n224 = ~n223 & ~pi088;
  assign n225 = ~n224 & ~pi089;
  assign n226 = ~n225 & ~pi090;
  assign n227 = ~n226 & ~pi091;
  assign n228 = ~n227 & ~pi092;
  assign n229 = ~n228 & ~pi093;
  assign n230 = ~n229 & ~pi094;
  assign n231 = ~n230 & ~pi095;
  assign n232 = ~n231 & ~pi096;
  assign n233 = ~n232 & ~pi097;
  assign n234 = ~n233 & ~pi098;
  assign n235 = ~n234 & ~pi099;
  assign n236 = ~n235 & ~pi100;
  assign n237 = ~n236 & ~pi101;
  assign n238 = ~n237 & ~pi102;
  assign n239 = ~n238 & ~pi103;
  assign n240 = ~n239 & ~pi104;
  assign n241 = ~n240 & ~pi105;
  assign n242 = ~n241 & ~pi106;
  assign n243 = ~n242 & ~pi107;
  assign n244 = ~n243 & ~pi108;
  assign n245 = ~n244 & ~pi109;
  assign n246 = ~n245 & ~pi110;
  assign n247 = ~n246 & ~pi111;
  assign n248 = ~n247 & ~pi112;
  assign n249 = ~n248 & ~pi113;
  assign n250 = ~n249 & ~pi114;
  assign n251 = ~n250 & ~pi115;
  assign n252 = ~n251 & ~pi116;
  assign n253 = ~n252 & ~pi117;
  assign n254 = ~n253 & ~pi118;
  assign n255 = ~n254 & ~pi119;
  assign n256 = ~n255 & ~pi120;
  assign n257 = ~n256 & ~pi121;
  assign n258 = ~n257 & ~pi122;
  assign n259 = ~n258 & ~pi123;
  assign n260 = ~n259 & ~pi124;
  assign n261 = ~n260 & ~pi125;
  assign n262 = ~n261 & ~pi126;
  assign po0 = n262 | pi127;
  assign n264 = ~pi126 & ~pi127;
  assign n265 = ~pi124 & ~pi125;
  assign n266 = ~pi122 & ~pi123;
  assign n267 = ~pi120 & ~pi121;
  assign n268 = n266 & n267;
  assign n269 = ~pi118 & ~pi119;
  assign n270 = ~pi116 & ~pi117;
  assign n271 = n269 & n270;
  assign n272 = n268 & n271;
  assign n273 = ~pi114 & ~pi115;
  assign n274 = n264 & n265;
  assign n275 = ~pi112 & ~pi113;
  assign n276 = n273 & n275;
  assign n277 = n272 & n276;
  assign n278 = n277 & n274;
  assign n279 = ~pi110 & ~pi111;
  assign n280 = ~pi108 & ~pi109;
  assign n281 = ~pi106 & ~pi107;
  assign n282 = ~pi104 & ~pi105;
  assign n283 = ~pi102 & ~pi103;
  assign n284 = ~pi100 & ~pi101;
  assign n285 = ~pi098 & ~pi099;
  assign n286 = ~pi096 & ~pi097;
  assign n287 = ~pi094 & ~pi095;
  assign n288 = ~pi092 & ~pi093;
  assign n289 = ~pi090 & ~pi091;
  assign n290 = ~pi088 & ~pi089;
  assign n291 = ~pi084 & ~pi085;
  assign n292 = ~pi086 & ~pi087;
  assign n293 = n291 & n292;
  assign n294 = n289 & n290;
  assign n295 = n287 & n288;
  assign n296 = n294 & n295;
  assign n297 = ~pi082 & ~pi083;
  assign n298 = ~pi080 & ~pi081;
  assign n299 = n297 & n298;
  assign n300 = n296 & n299;
  assign n301 = n300 & n293;
  assign n302 = ~pi078 & ~pi079;
  assign n303 = ~pi076 & ~pi077;
  assign n304 = ~pi074 & ~pi075;
  assign n305 = ~pi072 & ~pi073;
  assign n306 = ~pi070 & ~pi071;
  assign n307 = ~pi068 & ~pi069;
  assign n308 = ~pi066 & ~pi067;
  assign n309 = n304 & n305;
  assign n310 = n302 & n303;
  assign n311 = n309 & n310;
  assign n312 = n306 & n307;
  assign n313 = ~pi064 & ~pi065;
  assign n314 = n308 & n313;
  assign n315 = n312 & n314;
  assign n316 = n311 & n315;
  assign n317 = ~pi062 & ~pi063;
  assign n318 = ~pi060 & ~pi061;
  assign n319 = n317 & n318;
  assign n320 = ~pi058 & ~pi059;
  assign n321 = ~pi056 & ~pi057;
  assign n322 = n320 & n321;
  assign n323 = n319 & n322;
  assign n324 = ~pi054 & ~pi055;
  assign n325 = ~pi052 & ~pi053;
  assign n326 = n324 & n325;
  assign n327 = ~pi050 & ~pi051;
  assign n328 = ~pi048 & ~pi049;
  assign n329 = n327 & n328;
  assign n330 = n326 & n329;
  assign n331 = n323 & n330;
  assign n332 = ~pi046 & ~pi047;
  assign n333 = ~pi044 & ~pi045;
  assign n334 = n332 & n333;
  assign n335 = ~pi042 & ~pi043;
  assign n336 = ~pi040 & ~pi041;
  assign n337 = n335 & n336;
  assign n338 = n334 & n337;
  assign n339 = ~pi038 & ~pi039;
  assign n340 = ~pi036 & ~pi037;
  assign n341 = ~pi034 & ~pi035;
  assign n342 = n339 & n340;
  assign n343 = ~pi032 & ~pi033;
  assign n344 = n341 & n343;
  assign n345 = n342 & n344;
  assign n346 = n338 & n345;
  assign n347 = n331 & n346;
  assign n348 = ~pi018 & ~pi019;
  assign n349 = ~pi016 & ~pi017;
  assign n350 = n348 & n349;
  assign n351 = ~pi030 & ~pi031;
  assign n352 = ~pi028 & ~pi029;
  assign n353 = n351 & n352;
  assign n354 = ~pi026 & ~pi027;
  assign n355 = ~pi024 & ~pi025;
  assign n356 = n354 & n355;
  assign n357 = n353 & n356;
  assign n358 = ~pi022 & ~pi023;
  assign n359 = ~pi020 & ~pi021;
  assign n360 = n358 & n359;
  assign n361 = n357 & n360;
  assign n362 = n361 & n350;
  assign n363 = ~pi014 & ~pi015;
  assign n364 = ~pi012 & ~pi013;
  assign n365 = ~pi010 & ~pi011;
  assign n366 = n281 & n282;
  assign n367 = n279 & n280;
  assign n368 = n366 & n367;
  assign n369 = n285 & n286;
  assign n370 = n283 & n284;
  assign n371 = n369 & n370;
  assign n372 = n368 & n371;
  assign n373 = ~n362 & n346;
  assign n374 = ~n373 & n331;
  assign n375 = ~n374 & n316;
  assign n376 = ~n375 & n301;
  assign n377 = ~n376 & n372;
  assign n378 = n363 & n364;
  assign n379 = ~pi008 & ~pi009;
  assign n380 = n365 & n379;
  assign n381 = n378 & n380;
  assign n382 = ~n377 & ~n381;
  assign n383 = ~pi004 & ~pi005;
  assign n384 = ~pi002 & ~pi003;
  assign n385 = n383 & ~n384;
  assign n386 = ~pi006 & ~pi007;
  assign n387 = ~n385 & n386;
  assign n388 = ~n382 & ~n387;
  assign n389 = ~n388 & n365;
  assign n390 = ~n389 & n364;
  assign n391 = ~n390 & n363;
  assign n392 = ~n391 & n362;
  assign n393 = n356 & ~n358;
  assign n394 = ~n393 & n354;
  assign n395 = ~n394 & n353;
  assign n396 = n361 & ~n348;
  assign n397 = ~n396 & n351;
  assign n398 = n397 & ~n395;
  assign n399 = ~n392 & n398;
  assign n400 = ~n399 & n347;
  assign n401 = ~n400 & n341;
  assign n402 = ~n401 & n342;
  assign n403 = ~n402 & n339;
  assign n404 = ~n403 & n338;
  assign n405 = n333 & ~n335;
  assign n406 = ~n405 & n332;
  assign n407 = ~n404 & n406;
  assign n408 = ~n407 & n331;
  assign n409 = n325 & ~n327;
  assign n410 = ~n409 & n324;
  assign n411 = ~n408 & n410;
  assign n412 = ~n411 & n323;
  assign n413 = n318 & ~n320;
  assign n414 = ~n413 & n317;
  assign n415 = ~n412 & n414;
  assign n416 = ~n415 & n316;
  assign n417 = ~n416 & n308;
  assign n418 = ~n417 & n307;
  assign n419 = ~n418 & n306;
  assign n420 = ~n419 & n309;
  assign n421 = ~n420 & n304;
  assign n422 = ~n421 & n303;
  assign n423 = ~n422 & n302;
  assign n424 = ~n423 & n301;
  assign n425 = n291 & ~n297;
  assign n426 = ~n425 & n292;
  assign n427 = ~n424 & n426;
  assign n428 = ~n427 & n294;
  assign n429 = ~n428 & n289;
  assign n430 = ~n429 & n288;
  assign n431 = ~n430 & n287;
  assign n432 = ~n431 & n286;
  assign n433 = ~n432 & n285;
  assign n434 = ~n433 & n284;
  assign n435 = ~n434 & n283;
  assign n436 = ~n435 & n366;
  assign n437 = ~n436 & n281;
  assign n438 = ~n437 & n280;
  assign n439 = ~n438 & n279;
  assign n440 = ~n439 & n278;
  assign n441 = ~n440 & n273;
  assign n442 = ~n441 & n272;
  assign n443 = n267 & ~n269;
  assign n444 = ~n443 & n266;
  assign n445 = ~n442 & n444;
  assign n446 = ~n445 & n265;
  assign po1 = n446 | ~n264;
  assign n448 = n383 & n386;
  assign n449 = ~n382 & ~n448;
  assign n450 = ~n449 & n378;
  assign n451 = ~n450 & n350;
  assign n452 = ~n451 & n360;
  assign n453 = ~n452 & n356;
  assign n454 = ~n453 & n353;
  assign n455 = ~n454 & n344;
  assign n456 = ~n455 & n342;
  assign n457 = ~n456 & n337;
  assign n458 = ~n457 & n334;
  assign n459 = ~n458 & n329;
  assign n460 = ~n459 & n326;
  assign n461 = ~n460 & n322;
  assign n462 = ~n461 & n319;
  assign n463 = ~n462 & n314;
  assign n464 = ~n463 & n312;
  assign n465 = ~n464 & n309;
  assign n466 = ~n465 & n310;
  assign n467 = ~n466 & n300;
  assign n468 = ~n467 & n293;
  assign n469 = ~n468 & n294;
  assign n470 = ~n469 & n295;
  assign n471 = ~n470 & n369;
  assign n472 = ~n471 & n370;
  assign n473 = ~n472 & n366;
  assign n474 = ~n473 & n367;
  assign n475 = ~n474 & n277;
  assign n476 = ~n475 & n271;
  assign n477 = ~n476 & n268;
  assign po2 = n477 | ~n274;
  assign n479 = n268 & n274;
  assign n480 = ~n382 & n357;
  assign n481 = ~n480 & n347;
  assign n482 = n330 & ~n338;
  assign n483 = ~n482 & n323;
  assign n484 = ~n481 & n483;
  assign n485 = n301 & n316;
  assign n486 = ~n484 & n485;
  assign n487 = n301 & ~n311;
  assign n488 = ~n487 & n296;
  assign n489 = ~n486 & n488;
  assign n490 = ~n489 & n371;
  assign n491 = ~n490 & n368;
  assign n492 = ~n491 & n277;
  assign po3 = n492 | ~n479;
  assign po4 = n377 | ~n278;
  assign n495 = n278 & n372;
  assign n496 = n485 & ~n347;
  assign po6 = ~n485 | ~n495;
  assign po5 = n496 | ~n495;
  assign n499 = ~pi000 & ~pi001;
  assign n500 = n347 & n499;
  assign n501 = ~po6 & n500;
  assign n502 = ~n375 & n501;
  assign n503 = ~n388 & n502;
  assign n504 = ~n481 & n503;
  assign po7 = n451 | ~n504;
endmodule


