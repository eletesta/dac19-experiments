module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128;
  wire n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073;
  assign n257 = x128 ^ x0;
  assign n259 = x0 & x128;
  assign n258 = x129 ^ x1;
  assign n260 = n259 ^ n258;
  assign n264 = x130 ^ x2;
  assign n261 = n259 ^ x129;
  assign n262 = n258 & ~n261;
  assign n263 = n262 ^ x1;
  assign n265 = n264 ^ n263;
  assign n269 = x131 ^ x3;
  assign n266 = n263 ^ x130;
  assign n267 = n264 & ~n266;
  assign n268 = n267 ^ x2;
  assign n270 = n269 ^ n268;
  assign n274 = x132 ^ x4;
  assign n271 = n268 ^ x131;
  assign n272 = n269 & ~n271;
  assign n273 = n272 ^ x3;
  assign n275 = n274 ^ n273;
  assign n277 = n269 & n274;
  assign n278 = n268 & n277;
  assign n279 = x3 & x131;
  assign n280 = n279 ^ x132;
  assign n281 = n274 & ~n280;
  assign n282 = n281 ^ x4;
  assign n283 = ~n278 & ~n282;
  assign n276 = x133 ^ x5;
  assign n284 = n283 ^ n276;
  assign n288 = x134 ^ x6;
  assign n285 = n283 ^ x133;
  assign n286 = n276 & n285;
  assign n287 = n286 ^ x5;
  assign n289 = n288 ^ n287;
  assign n291 = n276 & n288;
  assign n292 = ~n283 & n291;
  assign n293 = x5 & x133;
  assign n294 = n293 ^ x134;
  assign n295 = n288 & ~n294;
  assign n296 = n295 ^ x6;
  assign n297 = ~n292 & ~n296;
  assign n290 = x135 ^ x7;
  assign n298 = n297 ^ n290;
  assign n302 = x136 ^ x8;
  assign n299 = n297 ^ x135;
  assign n300 = n290 & n299;
  assign n301 = n300 ^ x7;
  assign n303 = n302 ^ n301;
  assign n305 = n290 & n302;
  assign n306 = ~n297 & n305;
  assign n307 = x7 & x135;
  assign n308 = n307 ^ x136;
  assign n309 = n302 & ~n308;
  assign n310 = n309 ^ x8;
  assign n311 = ~n306 & ~n310;
  assign n304 = x137 ^ x9;
  assign n312 = n311 ^ n304;
  assign n314 = x9 & x137;
  assign n315 = n304 & ~n311;
  assign n316 = ~n314 & ~n315;
  assign n313 = x138 ^ x10;
  assign n317 = n316 ^ n313;
  assign n319 = n313 & n315;
  assign n320 = n314 ^ x138;
  assign n321 = n313 & ~n320;
  assign n322 = n321 ^ x10;
  assign n323 = ~n319 & ~n322;
  assign n318 = x139 ^ x11;
  assign n324 = n323 ^ n318;
  assign n328 = x140 ^ x12;
  assign n325 = n323 ^ x139;
  assign n326 = n318 & n325;
  assign n327 = n326 ^ x11;
  assign n329 = n328 ^ n327;
  assign n331 = n318 & n328;
  assign n332 = ~n323 & n331;
  assign n333 = x11 & x139;
  assign n334 = n333 ^ x140;
  assign n335 = n328 & ~n334;
  assign n336 = n335 ^ x12;
  assign n337 = ~n332 & ~n336;
  assign n330 = x141 ^ x13;
  assign n338 = n337 ^ n330;
  assign n342 = x142 ^ x14;
  assign n339 = n337 ^ x141;
  assign n340 = n330 & n339;
  assign n341 = n340 ^ x13;
  assign n343 = n342 ^ n341;
  assign n345 = n330 & n342;
  assign n346 = ~n337 & n345;
  assign n347 = x13 & x141;
  assign n348 = n347 ^ x142;
  assign n349 = n342 & ~n348;
  assign n350 = n349 ^ x14;
  assign n351 = ~n346 & ~n350;
  assign n344 = x143 ^ x15;
  assign n352 = n351 ^ n344;
  assign n356 = x144 ^ x16;
  assign n353 = n351 ^ x143;
  assign n354 = n344 & n353;
  assign n355 = n354 ^ x15;
  assign n357 = n356 ^ n355;
  assign n359 = n344 & n356;
  assign n360 = ~n351 & n359;
  assign n361 = x15 & x143;
  assign n362 = n361 ^ x144;
  assign n363 = n356 & ~n362;
  assign n364 = n363 ^ x16;
  assign n365 = ~n360 & ~n364;
  assign n358 = x145 ^ x17;
  assign n366 = n365 ^ n358;
  assign n370 = x146 ^ x18;
  assign n367 = n365 ^ x145;
  assign n368 = n358 & n367;
  assign n369 = n368 ^ x17;
  assign n371 = n370 ^ n369;
  assign n373 = n358 & n370;
  assign n374 = ~n365 & n373;
  assign n375 = x17 & x145;
  assign n376 = n375 ^ x146;
  assign n377 = n370 & ~n376;
  assign n378 = n377 ^ x18;
  assign n379 = ~n374 & ~n378;
  assign n372 = x147 ^ x19;
  assign n380 = n379 ^ n372;
  assign n382 = x19 & x147;
  assign n383 = n372 & ~n379;
  assign n384 = ~n382 & ~n383;
  assign n381 = x148 ^ x20;
  assign n385 = n384 ^ n381;
  assign n387 = n381 & n383;
  assign n388 = n382 ^ x148;
  assign n389 = n381 & ~n388;
  assign n390 = n389 ^ x20;
  assign n391 = ~n387 & ~n390;
  assign n386 = x149 ^ x21;
  assign n392 = n391 ^ n386;
  assign n396 = x150 ^ x22;
  assign n393 = n391 ^ x149;
  assign n394 = n386 & n393;
  assign n395 = n394 ^ x21;
  assign n397 = n396 ^ n395;
  assign n399 = n386 & n396;
  assign n400 = ~n391 & n399;
  assign n401 = x21 & x149;
  assign n402 = n401 ^ x150;
  assign n403 = n396 & ~n402;
  assign n404 = n403 ^ x22;
  assign n405 = ~n400 & ~n404;
  assign n398 = x151 ^ x23;
  assign n406 = n405 ^ n398;
  assign n410 = x152 ^ x24;
  assign n407 = n405 ^ x151;
  assign n408 = n398 & n407;
  assign n409 = n408 ^ x23;
  assign n411 = n410 ^ n409;
  assign n413 = n398 & n410;
  assign n414 = ~n405 & n413;
  assign n415 = x23 & x151;
  assign n416 = n415 ^ x152;
  assign n417 = n410 & ~n416;
  assign n418 = n417 ^ x24;
  assign n419 = ~n414 & ~n418;
  assign n412 = x153 ^ x25;
  assign n420 = n419 ^ n412;
  assign n424 = x154 ^ x26;
  assign n421 = n419 ^ x153;
  assign n422 = n412 & n421;
  assign n423 = n422 ^ x25;
  assign n425 = n424 ^ n423;
  assign n427 = n412 & n424;
  assign n428 = ~n419 & n427;
  assign n429 = x25 & x153;
  assign n430 = n429 ^ x154;
  assign n431 = n424 & ~n430;
  assign n432 = n431 ^ x26;
  assign n433 = ~n428 & ~n432;
  assign n426 = x155 ^ x27;
  assign n434 = n433 ^ n426;
  assign n438 = x156 ^ x28;
  assign n435 = n433 ^ x155;
  assign n436 = n426 & n435;
  assign n437 = n436 ^ x27;
  assign n439 = n438 ^ n437;
  assign n441 = n426 & n438;
  assign n442 = ~n433 & n441;
  assign n443 = x27 & x155;
  assign n444 = n443 ^ x156;
  assign n445 = n438 & ~n444;
  assign n446 = n445 ^ x28;
  assign n447 = ~n442 & ~n446;
  assign n440 = x157 ^ x29;
  assign n448 = n447 ^ n440;
  assign n450 = x29 & x157;
  assign n451 = n440 & ~n447;
  assign n452 = ~n450 & ~n451;
  assign n449 = x158 ^ x30;
  assign n453 = n452 ^ n449;
  assign n455 = n449 & n451;
  assign n456 = n450 ^ x158;
  assign n457 = n449 & ~n456;
  assign n458 = n457 ^ x30;
  assign n459 = ~n455 & ~n458;
  assign n454 = x159 ^ x31;
  assign n460 = n459 ^ n454;
  assign n464 = x160 ^ x32;
  assign n461 = n459 ^ x159;
  assign n462 = n454 & n461;
  assign n463 = n462 ^ x31;
  assign n465 = n464 ^ n463;
  assign n467 = n454 & n464;
  assign n468 = ~n459 & n467;
  assign n469 = x31 & x159;
  assign n470 = n469 ^ x160;
  assign n471 = n464 & ~n470;
  assign n472 = n471 ^ x32;
  assign n473 = ~n468 & ~n472;
  assign n466 = x161 ^ x33;
  assign n474 = n473 ^ n466;
  assign n478 = x162 ^ x34;
  assign n475 = n473 ^ x161;
  assign n476 = n466 & n475;
  assign n477 = n476 ^ x33;
  assign n479 = n478 ^ n477;
  assign n481 = n466 & n478;
  assign n482 = ~n473 & n481;
  assign n483 = x33 & x161;
  assign n484 = n483 ^ x162;
  assign n485 = n478 & ~n484;
  assign n486 = n485 ^ x34;
  assign n487 = ~n482 & ~n486;
  assign n480 = x163 ^ x35;
  assign n488 = n487 ^ n480;
  assign n492 = x164 ^ x36;
  assign n489 = n487 ^ x163;
  assign n490 = n480 & n489;
  assign n491 = n490 ^ x35;
  assign n493 = n492 ^ n491;
  assign n495 = n480 & n492;
  assign n496 = ~n487 & n495;
  assign n497 = x35 & x163;
  assign n498 = n497 ^ x164;
  assign n499 = n492 & ~n498;
  assign n500 = n499 ^ x36;
  assign n501 = ~n496 & ~n500;
  assign n494 = x165 ^ x37;
  assign n502 = n501 ^ n494;
  assign n506 = x166 ^ x38;
  assign n503 = n501 ^ x165;
  assign n504 = n494 & n503;
  assign n505 = n504 ^ x37;
  assign n507 = n506 ^ n505;
  assign n509 = n494 & n506;
  assign n510 = ~n501 & n509;
  assign n511 = x37 & x165;
  assign n512 = n511 ^ x166;
  assign n513 = n506 & ~n512;
  assign n514 = n513 ^ x38;
  assign n515 = ~n510 & ~n514;
  assign n508 = x167 ^ x39;
  assign n516 = n515 ^ n508;
  assign n518 = x39 & x167;
  assign n519 = n508 & ~n515;
  assign n520 = ~n518 & ~n519;
  assign n517 = x168 ^ x40;
  assign n521 = n520 ^ n517;
  assign n523 = n517 & n519;
  assign n524 = n518 ^ x168;
  assign n525 = n517 & ~n524;
  assign n526 = n525 ^ x40;
  assign n527 = ~n523 & ~n526;
  assign n522 = x169 ^ x41;
  assign n528 = n527 ^ n522;
  assign n532 = x170 ^ x42;
  assign n529 = n527 ^ x169;
  assign n530 = n522 & n529;
  assign n531 = n530 ^ x41;
  assign n533 = n532 ^ n531;
  assign n535 = n522 & n532;
  assign n536 = ~n527 & n535;
  assign n537 = x41 & x169;
  assign n538 = n537 ^ x170;
  assign n539 = n532 & ~n538;
  assign n540 = n539 ^ x42;
  assign n541 = ~n536 & ~n540;
  assign n534 = x171 ^ x43;
  assign n542 = n541 ^ n534;
  assign n546 = x172 ^ x44;
  assign n543 = n541 ^ x171;
  assign n544 = n534 & n543;
  assign n545 = n544 ^ x43;
  assign n547 = n546 ^ n545;
  assign n549 = n534 & n546;
  assign n550 = ~n541 & n549;
  assign n551 = x43 & x171;
  assign n552 = n551 ^ x172;
  assign n553 = n546 & ~n552;
  assign n554 = n553 ^ x44;
  assign n555 = ~n550 & ~n554;
  assign n548 = x173 ^ x45;
  assign n556 = n555 ^ n548;
  assign n560 = x174 ^ x46;
  assign n557 = n555 ^ x173;
  assign n558 = n548 & n557;
  assign n559 = n558 ^ x45;
  assign n561 = n560 ^ n559;
  assign n563 = n548 & n560;
  assign n564 = ~n555 & n563;
  assign n565 = x45 & x173;
  assign n566 = n565 ^ x174;
  assign n567 = n560 & ~n566;
  assign n568 = n567 ^ x46;
  assign n569 = ~n564 & ~n568;
  assign n562 = x175 ^ x47;
  assign n570 = n569 ^ n562;
  assign n574 = x176 ^ x48;
  assign n571 = n569 ^ x175;
  assign n572 = n562 & n571;
  assign n573 = n572 ^ x47;
  assign n575 = n574 ^ n573;
  assign n577 = n562 & n574;
  assign n578 = ~n569 & n577;
  assign n579 = x47 & x175;
  assign n580 = n579 ^ x176;
  assign n581 = n574 & ~n580;
  assign n582 = n581 ^ x48;
  assign n583 = ~n578 & ~n582;
  assign n576 = x177 ^ x49;
  assign n584 = n583 ^ n576;
  assign n586 = x49 & x177;
  assign n587 = n576 & ~n583;
  assign n588 = ~n586 & ~n587;
  assign n585 = x178 ^ x50;
  assign n589 = n588 ^ n585;
  assign n591 = n585 & n587;
  assign n592 = n586 ^ x178;
  assign n593 = n585 & ~n592;
  assign n594 = n593 ^ x50;
  assign n595 = ~n591 & ~n594;
  assign n590 = x179 ^ x51;
  assign n596 = n595 ^ n590;
  assign n600 = x180 ^ x52;
  assign n597 = n595 ^ x179;
  assign n598 = n590 & n597;
  assign n599 = n598 ^ x51;
  assign n601 = n600 ^ n599;
  assign n603 = n590 & n600;
  assign n604 = ~n595 & n603;
  assign n605 = x51 & x179;
  assign n606 = n605 ^ x180;
  assign n607 = n600 & ~n606;
  assign n608 = n607 ^ x52;
  assign n609 = ~n604 & ~n608;
  assign n602 = x181 ^ x53;
  assign n610 = n609 ^ n602;
  assign n614 = x182 ^ x54;
  assign n611 = n609 ^ x181;
  assign n612 = n602 & n611;
  assign n613 = n612 ^ x53;
  assign n615 = n614 ^ n613;
  assign n617 = n602 & n614;
  assign n618 = ~n609 & n617;
  assign n619 = x53 & x181;
  assign n620 = n619 ^ x182;
  assign n621 = n614 & ~n620;
  assign n622 = n621 ^ x54;
  assign n623 = ~n618 & ~n622;
  assign n616 = x183 ^ x55;
  assign n624 = n623 ^ n616;
  assign n628 = x184 ^ x56;
  assign n625 = n623 ^ x183;
  assign n626 = n616 & n625;
  assign n627 = n626 ^ x55;
  assign n629 = n628 ^ n627;
  assign n631 = n616 & n628;
  assign n632 = ~n623 & n631;
  assign n633 = x55 & x183;
  assign n634 = n633 ^ x184;
  assign n635 = n628 & ~n634;
  assign n636 = n635 ^ x56;
  assign n637 = ~n632 & ~n636;
  assign n630 = x185 ^ x57;
  assign n638 = n637 ^ n630;
  assign n642 = x186 ^ x58;
  assign n639 = n637 ^ x185;
  assign n640 = n630 & n639;
  assign n641 = n640 ^ x57;
  assign n643 = n642 ^ n641;
  assign n645 = n630 & n642;
  assign n646 = ~n637 & n645;
  assign n647 = x57 & x185;
  assign n648 = n647 ^ x186;
  assign n649 = n642 & ~n648;
  assign n650 = n649 ^ x58;
  assign n651 = ~n646 & ~n650;
  assign n644 = x187 ^ x59;
  assign n652 = n651 ^ n644;
  assign n654 = x59 & x187;
  assign n655 = n644 & ~n651;
  assign n656 = ~n654 & ~n655;
  assign n653 = x188 ^ x60;
  assign n657 = n656 ^ n653;
  assign n659 = n653 & n655;
  assign n660 = n654 ^ x188;
  assign n661 = n653 & ~n660;
  assign n662 = n661 ^ x60;
  assign n663 = ~n659 & ~n662;
  assign n658 = x189 ^ x61;
  assign n664 = n663 ^ n658;
  assign n668 = x190 ^ x62;
  assign n665 = n663 ^ x189;
  assign n666 = n658 & n665;
  assign n667 = n666 ^ x61;
  assign n669 = n668 ^ n667;
  assign n671 = n658 & n668;
  assign n672 = ~n663 & n671;
  assign n673 = x61 & x189;
  assign n674 = n673 ^ x190;
  assign n675 = n668 & ~n674;
  assign n676 = n675 ^ x62;
  assign n677 = ~n672 & ~n676;
  assign n670 = x191 ^ x63;
  assign n678 = n677 ^ n670;
  assign n682 = x192 ^ x64;
  assign n679 = n677 ^ x191;
  assign n680 = n670 & n679;
  assign n681 = n680 ^ x63;
  assign n683 = n682 ^ n681;
  assign n685 = n670 & n682;
  assign n686 = ~n677 & n685;
  assign n687 = x63 & x191;
  assign n688 = n687 ^ x192;
  assign n689 = n682 & ~n688;
  assign n690 = n689 ^ x64;
  assign n691 = ~n686 & ~n690;
  assign n684 = x193 ^ x65;
  assign n692 = n691 ^ n684;
  assign n696 = x194 ^ x66;
  assign n693 = n691 ^ x193;
  assign n694 = n684 & n693;
  assign n695 = n694 ^ x65;
  assign n697 = n696 ^ n695;
  assign n699 = n684 & n696;
  assign n700 = ~n691 & n699;
  assign n701 = x65 & x193;
  assign n702 = n701 ^ x194;
  assign n703 = n696 & ~n702;
  assign n704 = n703 ^ x66;
  assign n705 = ~n700 & ~n704;
  assign n698 = x195 ^ x67;
  assign n706 = n705 ^ n698;
  assign n710 = x196 ^ x68;
  assign n707 = n705 ^ x195;
  assign n708 = n698 & n707;
  assign n709 = n708 ^ x67;
  assign n711 = n710 ^ n709;
  assign n713 = n698 & n710;
  assign n714 = ~n705 & n713;
  assign n715 = x67 & x195;
  assign n716 = n715 ^ x196;
  assign n717 = n710 & ~n716;
  assign n718 = n717 ^ x68;
  assign n719 = ~n714 & ~n718;
  assign n712 = x197 ^ x69;
  assign n720 = n719 ^ n712;
  assign n722 = x69 & x197;
  assign n723 = n712 & ~n719;
  assign n724 = ~n722 & ~n723;
  assign n721 = x198 ^ x70;
  assign n725 = n724 ^ n721;
  assign n727 = n721 & n723;
  assign n728 = n722 ^ x198;
  assign n729 = n721 & ~n728;
  assign n730 = n729 ^ x70;
  assign n731 = ~n727 & ~n730;
  assign n726 = x199 ^ x71;
  assign n732 = n731 ^ n726;
  assign n736 = x200 ^ x72;
  assign n733 = n731 ^ x199;
  assign n734 = n726 & n733;
  assign n735 = n734 ^ x71;
  assign n737 = n736 ^ n735;
  assign n739 = n726 & n736;
  assign n740 = ~n731 & n739;
  assign n741 = x71 & x199;
  assign n742 = n741 ^ x200;
  assign n743 = n736 & ~n742;
  assign n744 = n743 ^ x72;
  assign n745 = ~n740 & ~n744;
  assign n738 = x201 ^ x73;
  assign n746 = n745 ^ n738;
  assign n750 = x202 ^ x74;
  assign n747 = n745 ^ x201;
  assign n748 = n738 & n747;
  assign n749 = n748 ^ x73;
  assign n751 = n750 ^ n749;
  assign n753 = n738 & n750;
  assign n754 = ~n745 & n753;
  assign n755 = x73 & x201;
  assign n756 = n755 ^ x202;
  assign n757 = n750 & ~n756;
  assign n758 = n757 ^ x74;
  assign n759 = ~n754 & ~n758;
  assign n752 = x203 ^ x75;
  assign n760 = n759 ^ n752;
  assign n764 = x204 ^ x76;
  assign n761 = n759 ^ x203;
  assign n762 = n752 & n761;
  assign n763 = n762 ^ x75;
  assign n765 = n764 ^ n763;
  assign n767 = n752 & n764;
  assign n768 = ~n759 & n767;
  assign n769 = x75 & x203;
  assign n770 = n769 ^ x204;
  assign n771 = n764 & ~n770;
  assign n772 = n771 ^ x76;
  assign n773 = ~n768 & ~n772;
  assign n766 = x205 ^ x77;
  assign n774 = n773 ^ n766;
  assign n778 = x206 ^ x78;
  assign n775 = n773 ^ x205;
  assign n776 = n766 & n775;
  assign n777 = n776 ^ x77;
  assign n779 = n778 ^ n777;
  assign n781 = n766 & n778;
  assign n782 = ~n773 & n781;
  assign n783 = x77 & x205;
  assign n784 = n783 ^ x206;
  assign n785 = n778 & ~n784;
  assign n786 = n785 ^ x78;
  assign n787 = ~n782 & ~n786;
  assign n780 = x207 ^ x79;
  assign n788 = n787 ^ n780;
  assign n790 = x79 & x207;
  assign n791 = n780 & ~n787;
  assign n792 = ~n790 & ~n791;
  assign n789 = x208 ^ x80;
  assign n793 = n792 ^ n789;
  assign n795 = n789 & n791;
  assign n796 = n790 ^ x208;
  assign n797 = n789 & ~n796;
  assign n798 = n797 ^ x80;
  assign n799 = ~n795 & ~n798;
  assign n794 = x209 ^ x81;
  assign n800 = n799 ^ n794;
  assign n804 = x210 ^ x82;
  assign n801 = n799 ^ x209;
  assign n802 = n794 & n801;
  assign n803 = n802 ^ x81;
  assign n805 = n804 ^ n803;
  assign n807 = n794 & n804;
  assign n808 = ~n799 & n807;
  assign n809 = x81 & x209;
  assign n810 = n809 ^ x210;
  assign n811 = n804 & ~n810;
  assign n812 = n811 ^ x82;
  assign n813 = ~n808 & ~n812;
  assign n806 = x211 ^ x83;
  assign n814 = n813 ^ n806;
  assign n818 = x212 ^ x84;
  assign n815 = n813 ^ x211;
  assign n816 = n806 & n815;
  assign n817 = n816 ^ x83;
  assign n819 = n818 ^ n817;
  assign n821 = n806 & n818;
  assign n822 = ~n813 & n821;
  assign n823 = x83 & x211;
  assign n824 = n823 ^ x212;
  assign n825 = n818 & ~n824;
  assign n826 = n825 ^ x84;
  assign n827 = ~n822 & ~n826;
  assign n820 = x213 ^ x85;
  assign n828 = n827 ^ n820;
  assign n832 = x214 ^ x86;
  assign n829 = n827 ^ x213;
  assign n830 = n820 & n829;
  assign n831 = n830 ^ x85;
  assign n833 = n832 ^ n831;
  assign n835 = n820 & n832;
  assign n836 = ~n827 & n835;
  assign n837 = x85 & x213;
  assign n838 = n837 ^ x214;
  assign n839 = n832 & ~n838;
  assign n840 = n839 ^ x86;
  assign n841 = ~n836 & ~n840;
  assign n834 = x215 ^ x87;
  assign n842 = n841 ^ n834;
  assign n846 = x216 ^ x88;
  assign n843 = n841 ^ x215;
  assign n844 = n834 & n843;
  assign n845 = n844 ^ x87;
  assign n847 = n846 ^ n845;
  assign n849 = n834 & n846;
  assign n850 = ~n841 & n849;
  assign n851 = x87 & x215;
  assign n852 = n851 ^ x216;
  assign n853 = n846 & ~n852;
  assign n854 = n853 ^ x88;
  assign n855 = ~n850 & ~n854;
  assign n848 = x217 ^ x89;
  assign n856 = n855 ^ n848;
  assign n858 = x89 & x217;
  assign n859 = n848 & ~n855;
  assign n860 = ~n858 & ~n859;
  assign n857 = x218 ^ x90;
  assign n861 = n860 ^ n857;
  assign n863 = n857 & n859;
  assign n864 = n858 ^ x218;
  assign n865 = n857 & ~n864;
  assign n866 = n865 ^ x90;
  assign n867 = ~n863 & ~n866;
  assign n862 = x219 ^ x91;
  assign n868 = n867 ^ n862;
  assign n870 = x91 & x219;
  assign n871 = n862 & ~n867;
  assign n872 = ~n870 & ~n871;
  assign n869 = x220 ^ x92;
  assign n873 = n872 ^ n869;
  assign n875 = n869 & n871;
  assign n876 = n870 ^ x220;
  assign n877 = n869 & ~n876;
  assign n878 = n877 ^ x92;
  assign n879 = ~n875 & ~n878;
  assign n874 = x221 ^ x93;
  assign n880 = n879 ^ n874;
  assign n884 = x222 ^ x94;
  assign n881 = n879 ^ x221;
  assign n882 = n874 & n881;
  assign n883 = n882 ^ x93;
  assign n885 = n884 ^ n883;
  assign n889 = x223 ^ x95;
  assign n886 = n883 ^ x222;
  assign n887 = n884 & ~n886;
  assign n888 = n887 ^ x94;
  assign n890 = n889 ^ n888;
  assign n894 = x224 ^ x96;
  assign n891 = n888 ^ x223;
  assign n892 = n889 & ~n891;
  assign n893 = n892 ^ x95;
  assign n895 = n894 ^ n893;
  assign n899 = x225 ^ x97;
  assign n896 = n893 ^ x224;
  assign n897 = n894 & ~n896;
  assign n898 = n897 ^ x96;
  assign n900 = n899 ^ n898;
  assign n904 = x226 ^ x98;
  assign n901 = n898 ^ x225;
  assign n902 = n899 & ~n901;
  assign n903 = n902 ^ x97;
  assign n905 = n904 ^ n903;
  assign n907 = n899 & n904;
  assign n908 = n898 & n907;
  assign n909 = x97 & x225;
  assign n910 = n909 ^ x226;
  assign n911 = n904 & ~n910;
  assign n912 = n911 ^ x98;
  assign n913 = ~n908 & ~n912;
  assign n906 = x227 ^ x99;
  assign n914 = n913 ^ n906;
  assign n918 = x228 ^ x100;
  assign n915 = n913 ^ x227;
  assign n916 = n906 & n915;
  assign n917 = n916 ^ x99;
  assign n919 = n918 ^ n917;
  assign n921 = n906 & n918;
  assign n922 = ~n913 & n921;
  assign n923 = x99 & x227;
  assign n924 = n923 ^ x228;
  assign n925 = n918 & ~n924;
  assign n926 = n925 ^ x100;
  assign n927 = ~n922 & ~n926;
  assign n920 = x229 ^ x101;
  assign n928 = n927 ^ n920;
  assign n932 = x230 ^ x102;
  assign n929 = n927 ^ x229;
  assign n930 = n920 & n929;
  assign n931 = n930 ^ x101;
  assign n933 = n932 ^ n931;
  assign n935 = n920 & n932;
  assign n936 = ~n927 & n935;
  assign n937 = x101 & x229;
  assign n938 = n937 ^ x230;
  assign n939 = n932 & ~n938;
  assign n940 = n939 ^ x102;
  assign n941 = ~n936 & ~n940;
  assign n934 = x231 ^ x103;
  assign n942 = n941 ^ n934;
  assign n946 = x232 ^ x104;
  assign n943 = n941 ^ x231;
  assign n944 = n934 & n943;
  assign n945 = n944 ^ x103;
  assign n947 = n946 ^ n945;
  assign n951 = x233 ^ x105;
  assign n948 = n945 ^ x232;
  assign n949 = n946 & ~n948;
  assign n950 = n949 ^ x104;
  assign n952 = n951 ^ n950;
  assign n956 = x234 ^ x106;
  assign n953 = n950 ^ x233;
  assign n954 = n951 & ~n953;
  assign n955 = n954 ^ x105;
  assign n957 = n956 ^ n955;
  assign n959 = n951 & n956;
  assign n960 = n950 & n959;
  assign n961 = x105 & x233;
  assign n962 = n961 ^ x234;
  assign n963 = n956 & ~n962;
  assign n964 = n963 ^ x106;
  assign n965 = ~n960 & ~n964;
  assign n958 = x235 ^ x107;
  assign n966 = n965 ^ n958;
  assign n970 = x236 ^ x108;
  assign n967 = n965 ^ x235;
  assign n968 = n958 & n967;
  assign n969 = n968 ^ x107;
  assign n971 = n970 ^ n969;
  assign n975 = x237 ^ x109;
  assign n972 = n969 ^ x236;
  assign n973 = n970 & ~n972;
  assign n974 = n973 ^ x108;
  assign n976 = n975 ^ n974;
  assign n980 = x238 ^ x110;
  assign n977 = n974 ^ x237;
  assign n978 = n975 & ~n977;
  assign n979 = n978 ^ x109;
  assign n981 = n980 ^ n979;
  assign n983 = n975 & n980;
  assign n984 = n974 & n983;
  assign n985 = x109 & x237;
  assign n986 = n985 ^ x238;
  assign n987 = n980 & ~n986;
  assign n988 = n987 ^ x110;
  assign n989 = ~n984 & ~n988;
  assign n982 = x239 ^ x111;
  assign n990 = n989 ^ n982;
  assign n994 = x240 ^ x112;
  assign n991 = n989 ^ x239;
  assign n992 = n982 & n991;
  assign n993 = n992 ^ x111;
  assign n995 = n994 ^ n993;
  assign n999 = x241 ^ x113;
  assign n996 = n993 ^ x240;
  assign n997 = n994 & ~n996;
  assign n998 = n997 ^ x112;
  assign n1000 = n999 ^ n998;
  assign n1004 = x242 ^ x114;
  assign n1001 = n998 ^ x241;
  assign n1002 = n999 & ~n1001;
  assign n1003 = n1002 ^ x113;
  assign n1005 = n1004 ^ n1003;
  assign n1009 = x243 ^ x115;
  assign n1006 = n1003 ^ x242;
  assign n1007 = n1004 & ~n1006;
  assign n1008 = n1007 ^ x114;
  assign n1010 = n1009 ^ n1008;
  assign n1014 = x244 ^ x116;
  assign n1011 = n1008 ^ x243;
  assign n1012 = n1009 & ~n1011;
  assign n1013 = n1012 ^ x115;
  assign n1015 = n1014 ^ n1013;
  assign n1019 = x245 ^ x117;
  assign n1016 = n1013 ^ x244;
  assign n1017 = n1014 & ~n1016;
  assign n1018 = n1017 ^ x116;
  assign n1020 = n1019 ^ n1018;
  assign n1024 = x246 ^ x118;
  assign n1021 = n1018 ^ x245;
  assign n1022 = n1019 & ~n1021;
  assign n1023 = n1022 ^ x117;
  assign n1025 = n1024 ^ n1023;
  assign n1029 = x247 ^ x119;
  assign n1026 = n1023 ^ x246;
  assign n1027 = n1024 & ~n1026;
  assign n1028 = n1027 ^ x118;
  assign n1030 = n1029 ^ n1028;
  assign n1034 = x248 ^ x120;
  assign n1031 = n1028 ^ x247;
  assign n1032 = n1029 & ~n1031;
  assign n1033 = n1032 ^ x119;
  assign n1035 = n1034 ^ n1033;
  assign n1039 = x249 ^ x121;
  assign n1036 = n1033 ^ x248;
  assign n1037 = n1034 & ~n1036;
  assign n1038 = n1037 ^ x120;
  assign n1040 = n1039 ^ n1038;
  assign n1044 = x250 ^ x122;
  assign n1041 = n1038 ^ x249;
  assign n1042 = n1039 & ~n1041;
  assign n1043 = n1042 ^ x121;
  assign n1045 = n1044 ^ n1043;
  assign n1049 = x251 ^ x123;
  assign n1046 = n1043 ^ x250;
  assign n1047 = n1044 & ~n1046;
  assign n1048 = n1047 ^ x122;
  assign n1050 = n1049 ^ n1048;
  assign n1054 = x252 ^ x124;
  assign n1051 = n1048 ^ x251;
  assign n1052 = n1049 & ~n1051;
  assign n1053 = n1052 ^ x123;
  assign n1055 = n1054 ^ n1053;
  assign n1059 = x253 ^ x125;
  assign n1056 = n1053 ^ x252;
  assign n1057 = n1054 & ~n1056;
  assign n1058 = n1057 ^ x124;
  assign n1060 = n1059 ^ n1058;
  assign n1064 = x254 ^ x126;
  assign n1061 = n1058 ^ x253;
  assign n1062 = n1059 & ~n1061;
  assign n1063 = n1062 ^ x125;
  assign n1065 = n1064 ^ n1063;
  assign n1069 = x255 ^ x127;
  assign n1066 = n1063 ^ x254;
  assign n1067 = n1064 & ~n1066;
  assign n1068 = n1067 ^ x126;
  assign n1070 = n1069 ^ n1068;
  assign n1071 = n1068 ^ x255;
  assign n1072 = n1069 & ~n1071;
  assign n1073 = n1072 ^ x127;
  assign y0 = n257;
  assign y1 = n260;
  assign y2 = n265;
  assign y3 = n270;
  assign y4 = n275;
  assign y5 = ~n284;
  assign y6 = n289;
  assign y7 = ~n298;
  assign y8 = n303;
  assign y9 = ~n312;
  assign y10 = ~n317;
  assign y11 = ~n324;
  assign y12 = n329;
  assign y13 = ~n338;
  assign y14 = n343;
  assign y15 = ~n352;
  assign y16 = n357;
  assign y17 = ~n366;
  assign y18 = n371;
  assign y19 = ~n380;
  assign y20 = ~n385;
  assign y21 = ~n392;
  assign y22 = n397;
  assign y23 = ~n406;
  assign y24 = n411;
  assign y25 = ~n420;
  assign y26 = n425;
  assign y27 = ~n434;
  assign y28 = n439;
  assign y29 = ~n448;
  assign y30 = ~n453;
  assign y31 = ~n460;
  assign y32 = n465;
  assign y33 = ~n474;
  assign y34 = n479;
  assign y35 = ~n488;
  assign y36 = n493;
  assign y37 = ~n502;
  assign y38 = n507;
  assign y39 = ~n516;
  assign y40 = ~n521;
  assign y41 = ~n528;
  assign y42 = n533;
  assign y43 = ~n542;
  assign y44 = n547;
  assign y45 = ~n556;
  assign y46 = n561;
  assign y47 = ~n570;
  assign y48 = n575;
  assign y49 = ~n584;
  assign y50 = ~n589;
  assign y51 = ~n596;
  assign y52 = n601;
  assign y53 = ~n610;
  assign y54 = n615;
  assign y55 = ~n624;
  assign y56 = n629;
  assign y57 = ~n638;
  assign y58 = n643;
  assign y59 = ~n652;
  assign y60 = ~n657;
  assign y61 = ~n664;
  assign y62 = n669;
  assign y63 = ~n678;
  assign y64 = n683;
  assign y65 = ~n692;
  assign y66 = n697;
  assign y67 = ~n706;
  assign y68 = n711;
  assign y69 = ~n720;
  assign y70 = ~n725;
  assign y71 = ~n732;
  assign y72 = n737;
  assign y73 = ~n746;
  assign y74 = n751;
  assign y75 = ~n760;
  assign y76 = n765;
  assign y77 = ~n774;
  assign y78 = n779;
  assign y79 = ~n788;
  assign y80 = ~n793;
  assign y81 = ~n800;
  assign y82 = n805;
  assign y83 = ~n814;
  assign y84 = n819;
  assign y85 = ~n828;
  assign y86 = n833;
  assign y87 = ~n842;
  assign y88 = n847;
  assign y89 = ~n856;
  assign y90 = ~n861;
  assign y91 = ~n868;
  assign y92 = ~n873;
  assign y93 = ~n880;
  assign y94 = n885;
  assign y95 = n890;
  assign y96 = n895;
  assign y97 = n900;
  assign y98 = n905;
  assign y99 = ~n914;
  assign y100 = n919;
  assign y101 = ~n928;
  assign y102 = n933;
  assign y103 = ~n942;
  assign y104 = n947;
  assign y105 = n952;
  assign y106 = n957;
  assign y107 = ~n966;
  assign y108 = n971;
  assign y109 = n976;
  assign y110 = n981;
  assign y111 = ~n990;
  assign y112 = n995;
  assign y113 = n1000;
  assign y114 = n1005;
  assign y115 = n1010;
  assign y116 = n1015;
  assign y117 = n1020;
  assign y118 = n1025;
  assign y119 = n1030;
  assign y120 = n1035;
  assign y121 = n1040;
  assign y122 = n1045;
  assign y123 = n1050;
  assign y124 = n1055;
  assign y125 = n1060;
  assign y126 = n1065;
  assign y127 = n1070;
  assign y128 = n1073;
endmodule
