module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24;
  wire n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790;
  assign n25 = ~x0 & ~x1;
  assign n26 = ~x2 & n25;
  assign n27 = ~x3 & n26;
  assign n28 = ~x4 & n27;
  assign n29 = ~x5 & n28;
  assign n30 = ~x6 & ~x7;
  assign n31 = n29 & n30;
  assign n32 = ~x8 & n31;
  assign n33 = ~x9 & n32;
  assign n34 = ~x10 & n33;
  assign n35 = ~x11 & n34;
  assign n36 = ~x12 & ~x13;
  assign n37 = ~x14 & n36;
  assign n38 = n35 & n37;
  assign n49 = ~x22 & ~n38;
  assign n50 = n49 ^ x15;
  assign n39 = ~x15 & n38;
  assign n40 = ~x22 & ~n39;
  assign n41 = ~x18 & ~x19;
  assign n42 = ~x16 & ~x17;
  assign n43 = n41 & n42;
  assign n44 = ~n40 & n43;
  assign n45 = ~x22 & ~n44;
  assign n46 = n45 ^ x20;
  assign n52 = x21 & ~x22;
  assign n53 = x20 & n52;
  assign n54 = ~x20 & ~x21;
  assign n55 = ~n53 & ~n54;
  assign n56 = ~n46 & n55;
  assign n83 = ~n50 & n56;
  assign n70 = n39 ^ x16;
  assign n71 = x17 & ~n70;
  assign n86 = x18 & x19;
  assign n87 = ~x22 & n86;
  assign n88 = n71 & n87;
  assign n75 = x16 & ~x17;
  assign n89 = x22 & n41;
  assign n90 = n75 & n89;
  assign n91 = ~n88 & ~n90;
  assign n198 = n83 & ~n91;
  assign n47 = x22 ^ x21;
  assign n48 = n46 & n47;
  assign n51 = n48 & ~n50;
  assign n72 = x19 & ~x22;
  assign n103 = n42 & n86;
  assign n104 = n39 ^ x18;
  assign n105 = n104 ^ x22;
  assign n106 = n42 ^ n39;
  assign n107 = n106 ^ n42;
  assign n108 = x16 & x17;
  assign n109 = n108 ^ n42;
  assign n110 = ~n107 & n109;
  assign n111 = n110 ^ n42;
  assign n112 = n111 ^ n104;
  assign n113 = n105 & ~n112;
  assign n114 = n113 ^ n110;
  assign n115 = n114 ^ n42;
  assign n116 = n115 ^ x22;
  assign n117 = ~n104 & ~n116;
  assign n118 = n117 ^ n104;
  assign n119 = ~n103 & n118;
  assign n120 = ~n72 & ~n119;
  assign n352 = n51 & n120;
  assign n1976 = ~n198 & ~n352;
  assign n139 = n48 & n50;
  assign n59 = x18 & ~x19;
  assign n60 = ~x22 & n59;
  assign n122 = ~x17 & ~n70;
  assign n178 = n60 & n122;
  assign n66 = ~x18 & x19;
  assign n67 = x22 & n66;
  assign n179 = n67 & n108;
  assign n180 = ~n178 & ~n179;
  assign n252 = n139 & ~n180;
  assign n128 = ~x22 & n41;
  assign n163 = n71 & n128;
  assign n130 = x22 & n86;
  assign n164 = n75 & n130;
  assign n165 = ~n163 & ~n164;
  assign n324 = n83 & ~n165;
  assign n1977 = ~n252 & ~n324;
  assign n1978 = n1976 & n1977;
  assign n100 = x21 ^ x20;
  assign n101 = n47 & ~n100;
  assign n102 = n50 & n101;
  assign n61 = x17 ^ x16;
  assign n62 = n39 ^ x17;
  assign n63 = n61 & ~n62;
  assign n135 = n63 & n87;
  assign n65 = ~x16 & x17;
  assign n136 = n65 & n89;
  assign n137 = ~n135 & ~n136;
  assign n138 = n102 & ~n137;
  assign n73 = ~x18 & n72;
  assign n74 = n71 & n73;
  assign n76 = x22 & n59;
  assign n77 = n75 & n76;
  assign n78 = ~n74 & ~n77;
  assign n288 = n51 & ~n78;
  assign n289 = ~n138 & ~n288;
  assign n57 = n50 & n56;
  assign n145 = ~n39 & n108;
  assign n146 = n87 & n145;
  assign n147 = ~n44 & ~n146;
  assign n308 = n57 & ~n147;
  assign n771 = n51 & ~n165;
  assign n888 = ~n308 & ~n771;
  assign n1979 = n289 & n888;
  assign n1980 = n1978 & n1979;
  assign n148 = n73 & n122;
  assign n149 = n76 & n108;
  assign n150 = ~n148 & ~n149;
  assign n154 = x19 & ~n118;
  assign n155 = n42 & n76;
  assign n156 = ~n154 & ~n155;
  assign n493 = n150 & n156;
  assign n494 = ~n56 & n493;
  assign n174 = n46 & ~n47;
  assign n227 = n60 & n71;
  assign n228 = n67 & n75;
  assign n229 = ~n227 & ~n228;
  assign n246 = n60 & n145;
  assign n247 = n42 & n66;
  assign n248 = ~n40 & n247;
  assign n249 = ~n246 & ~n248;
  assign n495 = n229 & n249;
  assign n496 = ~n174 & n495;
  assign n497 = ~n494 & ~n496;
  assign n2075 = ~n91 & n101;
  assign n2076 = n147 & ~n2075;
  assign n393 = n51 & ~n180;
  assign n2367 = ~n165 & n174;
  assign n2368 = ~n393 & ~n2367;
  assign n2369 = n2076 & n2368;
  assign n2370 = ~n497 & n2369;
  assign n84 = ~n47 & n50;
  assign n85 = n46 & n84;
  assign n95 = n63 & n73;
  assign n96 = n65 & n76;
  assign n97 = ~n95 & ~n96;
  assign n299 = n85 & ~n97;
  assign n166 = n122 & n128;
  assign n167 = n108 & n130;
  assign n168 = ~n166 & ~n167;
  assign n309 = n57 & ~n168;
  assign n503 = ~n299 & ~n309;
  assign n123 = n87 & n122;
  assign n124 = n89 & n108;
  assign n125 = ~n123 & ~n124;
  assign n296 = n102 & ~n125;
  assign n356 = ~n97 & n139;
  assign n808 = ~n296 & ~n356;
  assign n2371 = n503 & n808;
  assign n2372 = n2370 & n2371;
  assign n129 = n63 & n128;
  assign n131 = n65 & n130;
  assign n132 = ~n129 & ~n131;
  assign n175 = ~n50 & n174;
  assign n418 = ~n132 & n175;
  assign n226 = n57 & ~n91;
  assign n162 = ~n50 & n101;
  assign n592 = ~n125 & n162;
  assign n758 = ~n226 & ~n592;
  assign n2373 = ~n418 & n758;
  assign n231 = ~n156 & n162;
  assign n282 = ~n137 & n162;
  assign n2257 = ~n231 & ~n282;
  assign n414 = n120 & n139;
  assign n585 = n85 & ~n229;
  assign n2374 = ~n414 & ~n585;
  assign n2375 = n2257 & n2374;
  assign n2376 = n2373 & n2375;
  assign n2377 = n2372 & n2376;
  assign n2378 = n1980 & n2377;
  assign n234 = ~n57 & n147;
  assign n406 = n78 & n156;
  assign n407 = ~n139 & n406;
  assign n408 = ~n234 & ~n407;
  assign n169 = n165 & n168;
  assign n170 = n132 & n169;
  assign n514 = ~n120 & n132;
  assign n515 = n50 & ~n514;
  assign n522 = n170 & ~n515;
  assign n523 = n101 & ~n522;
  assign n524 = n51 & ~n147;
  assign n525 = n56 & ~n406;
  assign n526 = ~n524 & ~n525;
  assign n527 = ~n523 & n526;
  assign n528 = ~n408 & n527;
  assign n64 = n60 & n63;
  assign n68 = n65 & n67;
  assign n69 = ~n64 & ~n68;
  assign n191 = ~n69 & n175;
  assign n192 = n175 & ~n180;
  assign n193 = ~n191 & ~n192;
  assign n239 = ~n69 & n85;
  assign n479 = ~n125 & n174;
  assign n480 = ~n239 & ~n479;
  assign n276 = ~n120 & n165;
  assign n481 = n57 & ~n276;
  assign n482 = n480 & ~n481;
  assign n483 = n193 & n482;
  assign n283 = n139 & ~n150;
  assign n362 = n139 & ~n168;
  assign n975 = ~n283 & ~n362;
  assign n432 = ~n78 & n139;
  assign n265 = n97 & n150;
  assign n2073 = n51 & ~n265;
  assign n2074 = ~n432 & ~n2073;
  assign n2379 = n975 & n2074;
  assign n209 = n83 & n120;
  assign n638 = ~n91 & n175;
  assign n2380 = ~n209 & ~n638;
  assign n2381 = n2379 & n2380;
  assign n2382 = n483 & n2381;
  assign n2383 = n528 & n2382;
  assign n2384 = n2378 & n2383;
  assign n243 = n162 & ~n165;
  assign n244 = n83 & ~n147;
  assign n245 = ~n243 & ~n244;
  assign n250 = n175 & ~n249;
  assign n251 = n245 & ~n250;
  assign n297 = ~n69 & n83;
  assign n298 = n51 & ~n125;
  assign n300 = ~n298 & ~n299;
  assign n301 = ~n297 & n300;
  assign n322 = n251 & n301;
  assign n323 = n162 & ~n168;
  assign n325 = ~n125 & n139;
  assign n326 = ~n324 & ~n325;
  assign n327 = ~n323 & n326;
  assign n328 = n46 & n50;
  assign n329 = ~n165 & n328;
  assign n330 = n47 & n329;
  assign n331 = n78 & n125;
  assign n332 = ~n120 & n331;
  assign n333 = n83 & ~n332;
  assign n334 = ~n330 & ~n333;
  assign n335 = n327 & n334;
  assign n336 = n322 & n335;
  assign n210 = ~n91 & n102;
  assign n158 = n91 & n147;
  assign n337 = n85 & ~n158;
  assign n338 = ~n210 & ~n337;
  assign n339 = n132 & n338;
  assign n340 = n84 & ~n339;
  assign n341 = n83 & ~n249;
  assign n342 = ~n340 & ~n341;
  assign n343 = n336 & n342;
  assign n344 = ~n78 & n162;
  assign n345 = n51 & ~n249;
  assign n346 = ~n344 & ~n345;
  assign n347 = ~n69 & n102;
  assign n348 = n139 & ~n229;
  assign n349 = ~n347 & ~n348;
  assign n350 = n346 & n349;
  assign n221 = ~n83 & ~n102;
  assign n222 = ~n156 & ~n221;
  assign n351 = n83 & ~n150;
  assign n353 = ~n351 & ~n352;
  assign n354 = ~n222 & n353;
  assign n355 = n350 & n354;
  assign n357 = ~n78 & n102;
  assign n271 = ~n50 & ~n229;
  assign n358 = n174 & n271;
  assign n359 = ~n357 & ~n358;
  assign n360 = ~n356 & n359;
  assign n361 = n355 & n360;
  assign n363 = n83 & ~n180;
  assign n364 = ~n362 & ~n363;
  assign n238 = ~n69 & n162;
  assign n365 = n180 & n229;
  assign n366 = n85 & ~n365;
  assign n367 = ~n238 & ~n366;
  assign n368 = n364 & n367;
  assign n159 = n125 & n137;
  assign n369 = n156 & n159;
  assign n370 = n276 & n369;
  assign n371 = n175 & ~n370;
  assign n372 = n368 & ~n371;
  assign n373 = n361 & n372;
  assign n374 = n83 & ~n137;
  assign n375 = ~n137 & n175;
  assign n376 = ~n374 & ~n375;
  assign n377 = ~n97 & n102;
  assign n378 = n376 & ~n377;
  assign n379 = ~n198 & ~n309;
  assign n380 = n102 & ~n168;
  assign n79 = n69 & n78;
  assign n381 = ~n79 & n85;
  assign n382 = ~n380 & ~n381;
  assign n383 = n379 & n382;
  assign n384 = n378 & n383;
  assign n385 = n83 & ~n97;
  assign n386 = n48 & ~n91;
  assign n387 = ~n385 & ~n386;
  assign n388 = ~n132 & n139;
  assign n389 = ~n288 & ~n388;
  assign n390 = n387 & n389;
  assign n230 = n102 & ~n229;
  assign n290 = n56 & n271;
  assign n391 = ~n230 & ~n290;
  assign n392 = ~n221 & ~n276;
  assign n394 = n85 & ~n168;
  assign n395 = ~n150 & n162;
  assign n396 = ~n97 & n162;
  assign n397 = ~n395 & ~n396;
  assign n398 = ~n394 & n397;
  assign n399 = ~n393 & n398;
  assign n400 = ~n392 & n399;
  assign n401 = n391 & n400;
  assign n402 = n390 & n401;
  assign n403 = n384 & n402;
  assign n404 = n373 & n403;
  assign n405 = n343 & n404;
  assign n58 = ~n51 & ~n57;
  assign n80 = ~n50 & n69;
  assign n81 = ~n79 & ~n80;
  assign n82 = ~n58 & n81;
  assign n207 = n83 & ~n132;
  assign n558 = n162 & ~n249;
  assign n559 = ~n207 & ~n558;
  assign n560 = ~n82 & n559;
  assign n253 = n97 & n229;
  assign n254 = n175 & ~n253;
  assign n431 = n57 & ~n132;
  assign n577 = ~n254 & ~n431;
  assign n578 = n193 & n577;
  assign n579 = n389 & n578;
  assign n2092 = ~n132 & ~n579;
  assign n663 = n57 & ~n125;
  assign n664 = ~n432 & ~n663;
  assign n202 = n51 & ~n137;
  assign n800 = n51 & ~n156;
  assign n980 = ~n202 & ~n800;
  assign n151 = n147 & n150;
  assign n981 = n51 & ~n151;
  assign n982 = n980 & ~n981;
  assign n983 = n664 & n982;
  assign n240 = ~n238 & ~n239;
  assign n2093 = ~n323 & ~n374;
  assign n2094 = n240 & n2093;
  assign n656 = ~n132 & n162;
  assign n2095 = n102 & ~n156;
  assign n2096 = ~n656 & ~n2095;
  assign n2097 = ~n230 & n2096;
  assign n2098 = ~n363 & n2097;
  assign n2099 = n2094 & n2098;
  assign n2100 = n983 & n2099;
  assign n2101 = ~n2092 & n2100;
  assign n2102 = n560 & n2101;
  assign n581 = ~n85 & n150;
  assign n582 = ~n102 & n132;
  assign n583 = ~n581 & ~n582;
  assign n255 = n51 & ~n168;
  assign n747 = ~n255 & ~n297;
  assign n2103 = ~n583 & n747;
  assign n2104 = n2102 & n2103;
  assign n273 = n50 & ~n137;
  assign n274 = n56 & n273;
  assign n759 = ~n274 & ~n357;
  assign n606 = n102 & ~n180;
  assign n766 = ~n290 & ~n606;
  assign n912 = n56 & ~n156;
  assign n913 = n766 & ~n912;
  assign n914 = n759 & n913;
  assign n915 = n139 & ~n249;
  assign n916 = ~n356 & ~n915;
  assign n459 = n84 & ~n150;
  assign n917 = ~n120 & ~n459;
  assign n918 = n46 & ~n917;
  assign n919 = n916 & ~n918;
  assign n920 = n914 & n919;
  assign n1023 = ~n83 & ~n139;
  assign n1024 = ~n168 & ~n1023;
  assign n1025 = ~n137 & n174;
  assign n1026 = n50 & n1025;
  assign n1027 = ~n418 & ~n1026;
  assign n1028 = ~n1024 & n1027;
  assign n938 = n57 & ~n150;
  assign n939 = ~n78 & n85;
  assign n940 = ~n938 & ~n939;
  assign n303 = n57 & ~n97;
  assign n1029 = n125 & n249;
  assign n1030 = n51 & ~n1029;
  assign n1031 = ~n303 & ~n1030;
  assign n1032 = n940 & n1031;
  assign n1033 = n1028 & n1032;
  assign n767 = n57 & ~n229;
  assign n926 = ~n147 & n162;
  assign n927 = ~n767 & ~n926;
  assign n2247 = ~n375 & n927;
  assign n2248 = n1033 & n2247;
  assign n2309 = n920 & n2248;
  assign n121 = n102 & n120;
  assign n126 = n83 & ~n125;
  assign n127 = ~n121 & ~n126;
  assign n410 = ~n78 & n175;
  assign n2186 = ~n410 & ~n585;
  assign n2310 = n127 & n2186;
  assign n2108 = n78 & n265;
  assign n2109 = n83 & ~n2108;
  assign n2110 = ~n309 & ~n2109;
  assign n281 = n102 & ~n147;
  assign n2311 = ~n191 & ~n281;
  assign n2312 = n2110 & n2311;
  assign n2313 = n2310 & n2312;
  assign n624 = n85 & n120;
  assign n2314 = n175 & ~n1029;
  assign n2315 = ~n624 & ~n2314;
  assign n468 = n57 & ~n249;
  assign n1040 = n51 & ~n91;
  assign n2316 = ~n468 & ~n1040;
  assign n2317 = n2315 & n2316;
  assign n756 = ~n91 & n162;
  assign n2318 = ~n341 & ~n756;
  assign n627 = n162 & ~n180;
  assign n2319 = ~n344 & ~n627;
  assign n2320 = n2318 & n2319;
  assign n2321 = n2317 & n2320;
  assign n2322 = n2313 & n2321;
  assign n2323 = n2309 & n2322;
  assign n2324 = n2104 & n2323;
  assign n268 = n83 & ~n168;
  assign n484 = n132 & ~n174;
  assign n485 = ~n268 & n484;
  assign n486 = ~n56 & ~n120;
  assign n487 = n85 & ~n180;
  assign n488 = n486 & ~n487;
  assign n489 = ~n485 & ~n488;
  assign n490 = n83 & ~n276;
  assign n491 = ~n489 & ~n490;
  assign n492 = n483 & n491;
  assign n498 = n150 & n180;
  assign n499 = n69 & n498;
  assign n500 = n56 & ~n499;
  assign n501 = ~n303 & ~n500;
  assign n502 = ~n497 & n501;
  assign n504 = ~n174 & n503;
  assign n505 = n502 & n504;
  assign n506 = n492 & n505;
  assign n92 = n85 & ~n91;
  assign n93 = ~n83 & ~n92;
  assign n94 = ~n82 & n93;
  assign n98 = n80 & n97;
  assign n99 = ~n94 & ~n98;
  assign n133 = n58 & ~n132;
  assign n134 = n127 & ~n133;
  assign n140 = ~n91 & n139;
  assign n141 = ~n138 & ~n140;
  assign n142 = n134 & n141;
  assign n143 = ~n99 & n142;
  assign n144 = ~n51 & n143;
  assign n152 = ~n85 & n151;
  assign n153 = ~n144 & ~n152;
  assign n157 = n132 & n156;
  assign n160 = n158 & n159;
  assign n161 = n56 & n160;
  assign n171 = n162 & n170;
  assign n172 = ~n161 & ~n171;
  assign n173 = n157 & n172;
  assign n176 = n78 & ~n175;
  assign n177 = ~n173 & ~n176;
  assign n181 = n156 & n180;
  assign n182 = n137 & n181;
  assign n183 = n85 & ~n182;
  assign n184 = n132 & n150;
  assign n185 = ~n83 & n184;
  assign n186 = n78 & ~n102;
  assign n187 = n97 & n186;
  assign n188 = ~n185 & ~n187;
  assign n189 = ~n183 & ~n188;
  assign n190 = ~n125 & n175;
  assign n194 = ~n190 & n193;
  assign n195 = n189 & n194;
  assign n196 = ~n177 & n195;
  assign n197 = ~n153 & n196;
  assign n634 = ~n283 & ~n558;
  assign n284 = n51 & ~n69;
  assign n635 = ~n284 & ~n394;
  assign n636 = n634 & n635;
  assign n637 = n197 & n636;
  assign n411 = n46 & ~n50;
  assign n639 = ~n249 & n411;
  assign n640 = ~n638 & ~n639;
  assign n641 = ~n308 & ~n357;
  assign n642 = n640 & n641;
  assign n643 = n57 & ~n156;
  assign n644 = ~n231 & ~n643;
  assign n645 = n127 & n644;
  assign n646 = n642 & n645;
  assign n647 = ~n151 & n174;
  assign n648 = ~n175 & ~n647;
  assign n649 = ~n348 & n648;
  assign n650 = ~n50 & n78;
  assign n651 = ~n649 & ~n650;
  assign n652 = ~n139 & n156;
  assign n424 = ~n102 & n249;
  assign n653 = n147 & n424;
  assign n654 = ~n652 & ~n653;
  assign n655 = n174 & ~n253;
  assign n446 = ~n50 & ~n97;
  assign n657 = ~n446 & ~n656;
  assign n658 = ~n655 & n657;
  assign n659 = ~n654 & n658;
  assign n660 = ~n651 & n659;
  assign n661 = n646 & n660;
  assign n662 = n637 & n661;
  assign n438 = n85 & ~n249;
  assign n665 = ~n150 & n175;
  assign n666 = ~n438 & ~n665;
  assign n667 = ~n395 & n666;
  assign n668 = n664 & n667;
  assign n669 = n147 & ~n175;
  assign n670 = ~n486 & ~n669;
  assign n671 = ~n243 & ~n670;
  assign n672 = n668 & n671;
  assign n261 = n168 & n180;
  assign n262 = n175 & ~n261;
  assign n263 = n102 & ~n150;
  assign n264 = ~n262 & ~n263;
  assign n266 = n139 & ~n265;
  assign n267 = n264 & ~n266;
  assign n269 = ~n147 & n175;
  assign n270 = ~n268 & ~n269;
  assign n272 = n48 & n271;
  assign n275 = ~n272 & ~n274;
  assign n277 = n85 & ~n276;
  assign n278 = n275 & ~n277;
  assign n279 = n270 & n278;
  assign n280 = n267 & n279;
  assign n673 = n280 & n527;
  assign n674 = n672 & n673;
  assign n675 = n85 & ~n125;
  assign n467 = ~n165 & n175;
  assign n676 = ~n226 & ~n467;
  assign n677 = ~n675 & n676;
  assign n678 = n384 & n677;
  assign n679 = n674 & n678;
  assign n680 = n662 & n679;
  assign n561 = n334 & n560;
  assign n562 = ~n168 & n174;
  assign n563 = ~n50 & n562;
  assign n564 = ~n347 & ~n563;
  assign n565 = ~n272 & n564;
  assign n566 = n139 & ~n156;
  assign n567 = ~n345 & ~n566;
  assign n568 = n565 & n567;
  assign n569 = n561 & n568;
  assign n570 = n125 & n181;
  assign n571 = n57 & ~n570;
  assign n572 = ~n299 & ~n571;
  assign n531 = n120 & n162;
  assign n573 = ~n362 & ~n531;
  assign n574 = ~n250 & n573;
  assign n575 = n572 & n574;
  assign n576 = n569 & n575;
  assign n429 = n51 & ~n132;
  assign n580 = ~n429 & ~n467;
  assign n584 = n580 & ~n583;
  assign n586 = ~n102 & n150;
  assign n587 = ~n585 & n586;
  assign n588 = n97 & ~n174;
  assign n589 = ~n587 & ~n588;
  assign n590 = n584 & ~n589;
  assign n591 = n579 & n590;
  assign n593 = ~n395 & ~n592;
  assign n594 = ~n255 & n593;
  assign n454 = n57 & n120;
  assign n595 = n51 & ~n157;
  assign n596 = ~n454 & ~n595;
  assign n597 = ~n249 & n328;
  assign n598 = ~n524 & ~n597;
  assign n599 = n596 & n598;
  assign n600 = n594 & n599;
  assign n601 = n591 & n600;
  assign n602 = n576 & n601;
  assign n603 = ~n78 & n174;
  assign n604 = ~n138 & ~n396;
  assign n605 = ~n603 & n604;
  assign n607 = ~n323 & ~n606;
  assign n608 = n605 & n607;
  assign n609 = ~n296 & ~n380;
  assign n610 = ~n325 & n609;
  assign n611 = ~n282 & ~n418;
  assign n510 = n69 & n168;
  assign n612 = n180 & n510;
  assign n613 = n85 & ~n612;
  assign n614 = n165 & ~n446;
  assign n615 = n56 & ~n614;
  assign n616 = ~n613 & ~n615;
  assign n617 = n611 & n616;
  assign n618 = n610 & n617;
  assign n619 = n608 & n618;
  assign n620 = n85 & ~n165;
  assign n621 = n120 & n175;
  assign n622 = ~n348 & ~n621;
  assign n623 = ~n620 & n622;
  assign n625 = n139 & ~n147;
  assign n626 = ~n624 & ~n625;
  assign n628 = ~n83 & ~n627;
  assign n629 = ~n181 & ~n628;
  assign n630 = n626 & ~n629;
  assign n631 = n623 & n630;
  assign n632 = n619 & n631;
  assign n633 = n602 & n632;
  assign n694 = n680 ^ n633;
  assign n507 = n56 & n506;
  assign n508 = n83 & ~n160;
  assign n509 = ~n429 & ~n508;
  assign n511 = n139 & ~n510;
  assign n512 = n509 & ~n511;
  assign n513 = ~n352 & n512;
  assign n516 = n165 & n180;
  assign n517 = ~n515 & n516;
  assign n518 = n48 & ~n517;
  assign n519 = ~n255 & ~n518;
  assign n520 = n513 & n519;
  assign n521 = ~n507 & n520;
  assign n529 = n69 & n365;
  assign n530 = n101 & ~n529;
  assign n470 = n102 & ~n249;
  assign n532 = ~n470 & ~n531;
  assign n533 = ~n530 & n532;
  assign n534 = n528 & n533;
  assign n535 = n521 & n534;
  assign n695 = n680 ^ n535;
  assign n537 = ~x22 & ~n35;
  assign n541 = x12 & ~x22;
  assign n542 = ~n537 & ~n541;
  assign n549 = x13 & ~x22;
  assign n550 = n542 & ~n549;
  assign n551 = n550 ^ x14;
  assign n696 = n680 ^ n551;
  assign n697 = n695 & n696;
  assign n698 = n697 ^ n680;
  assign n699 = ~n694 & ~n698;
  assign n700 = n699 ^ n535;
  assign n536 = ~n48 & n535;
  assign n538 = n537 ^ x12;
  assign n539 = ~n506 & ~n538;
  assign n540 = n536 & ~n539;
  assign n543 = n542 ^ x13;
  assign n544 = n506 & n521;
  assign n545 = n543 & n544;
  assign n546 = ~n521 & ~n538;
  assign n547 = ~n545 & ~n546;
  assign n548 = ~n540 & n547;
  assign n552 = n551 ^ n543;
  assign n553 = n521 & n552;
  assign n554 = n553 ^ n543;
  assign n555 = ~n536 & ~n554;
  assign n556 = ~n506 & n543;
  assign n557 = ~n555 & ~n556;
  assign n708 = ~n548 & n557;
  assign n681 = ~n633 & ~n680;
  assign n682 = ~n535 & ~n681;
  assign n683 = ~x22 & ~n34;
  assign n684 = n683 ^ x11;
  assign n685 = n684 ^ n538;
  assign n686 = ~n506 & n685;
  assign n687 = ~n682 & ~n686;
  assign n707 = n543 & ~n687;
  assign n709 = n708 ^ n707;
  assign n710 = n700 & n709;
  assign n711 = n710 ^ n708;
  assign n712 = ~n506 & n711;
  assign n688 = n687 ^ n557;
  assign n701 = ~n548 & n700;
  assign n702 = ~n688 & n701;
  assign n704 = n557 & ~n687;
  assign n1942 = ~n702 & ~n704;
  assign n1943 = ~n712 & n1942;
  assign n1937 = ~n521 & ~n551;
  assign n1938 = ~n538 & ~n684;
  assign n1939 = n1938 ^ n552;
  assign n1940 = ~n506 & n1939;
  assign n1941 = ~n1937 & ~n1940;
  assign n1944 = n1943 ^ n1941;
  assign n859 = n700 ^ n548;
  assign n849 = ~x22 & ~n33;
  assign n850 = n849 ^ x10;
  assign n731 = ~x22 & ~n32;
  assign n732 = n731 ^ x9;
  assign n851 = n850 ^ n732;
  assign n739 = ~n230 & ~n324;
  assign n740 = ~n431 & n739;
  assign n741 = n623 & n740;
  assign n471 = n125 & n229;
  assign n742 = n58 & n471;
  assign n743 = ~n85 & ~n120;
  assign n744 = ~n298 & n743;
  assign n745 = ~n742 & ~n744;
  assign n746 = n741 & ~n745;
  assign n748 = n376 & n747;
  assign n749 = ~n239 & ~n656;
  assign n750 = n573 & n749;
  assign n751 = n748 & n750;
  assign n752 = n746 & n751;
  assign n753 = ~n120 & n150;
  assign n754 = n137 & n753;
  assign n755 = n139 & ~n754;
  assign n757 = n389 & ~n756;
  assign n760 = ~n238 & n759;
  assign n761 = n758 & n760;
  assign n762 = n757 & n761;
  assign n763 = ~n755 & n762;
  assign n764 = ~n202 & ~n210;
  assign n765 = n626 & n764;
  assign n469 = ~n467 & ~n468;
  assign n768 = n766 & ~n767;
  assign n769 = n469 & n768;
  assign n770 = n765 & n769;
  assign n211 = n125 & n165;
  assign n772 = n102 & ~n211;
  assign n773 = ~n207 & ~n772;
  assign n774 = ~n771 & n773;
  assign n291 = n57 & ~n165;
  assign n775 = ~n562 & ~n566;
  assign n776 = ~n291 & n775;
  assign n777 = n774 & n776;
  assign n778 = n770 & n777;
  assign n779 = n763 & n778;
  assign n780 = n752 & n779;
  assign n781 = n637 & n780;
  assign n430 = ~n341 & ~n429;
  assign n782 = ~n222 & n430;
  assign n783 = ~n357 & ~n362;
  assign n784 = n782 & n783;
  assign n423 = n97 & ~n139;
  assign n425 = ~n423 & ~n424;
  assign n785 = ~n243 & ~n425;
  assign n786 = n162 & ~n229;
  assign n787 = ~n288 & ~n786;
  assign n788 = ~n190 & n787;
  assign n789 = n785 & n788;
  assign n790 = n784 & n789;
  assign n791 = ~n209 & ~n385;
  assign n792 = ~n297 & n791;
  assign n793 = n667 & n792;
  assign n794 = n790 & n793;
  assign n458 = ~n252 & ~n380;
  assign n460 = ~n48 & n180;
  assign n461 = ~n101 & n125;
  assign n462 = ~n50 & ~n461;
  assign n463 = ~n460 & n462;
  assign n464 = ~n459 & ~n463;
  assign n465 = n458 & n464;
  assign n795 = ~n102 & ~n175;
  assign n796 = ~n158 & ~n795;
  assign n797 = ~n238 & ~n531;
  assign n798 = ~n771 & n797;
  assign n799 = ~n796 & n798;
  assign n801 = ~n675 & ~n800;
  assign n802 = n799 & n801;
  assign n803 = n465 & n802;
  assign n804 = ~n198 & ~n291;
  assign n805 = n132 & ~n274;
  assign n806 = n804 & n805;
  assign n807 = n56 & ~n806;
  assign n809 = n91 & n156;
  assign n810 = n175 & ~n809;
  assign n811 = ~n288 & ~n810;
  assign n812 = n85 & ~n147;
  assign n813 = n85 & ~n156;
  assign n814 = ~n812 & ~n813;
  assign n815 = n811 & n814;
  assign n816 = n808 & n815;
  assign n817 = ~n807 & n816;
  assign n818 = n803 & n817;
  assign n819 = n794 & n818;
  assign n820 = ~n162 & ~n175;
  assign n821 = ~n249 & ~n820;
  assign n822 = n102 & ~n132;
  assign n823 = n51 & ~n253;
  assign n824 = ~n822 & ~n823;
  assign n825 = ~n821 & n824;
  assign n826 = ~n140 & n825;
  assign n409 = ~n138 & ~n408;
  assign n827 = ~n358 & ~n755;
  assign n828 = n409 & n827;
  assign n829 = n826 & n828;
  assign n830 = n57 & ~n365;
  assign n831 = ~n284 & ~n830;
  assign n832 = ~n210 & ~n656;
  assign n833 = n831 & n832;
  assign n834 = n829 & n833;
  assign n835 = n819 & n834;
  assign n852 = ~n781 & ~n835;
  assign n853 = ~n633 & ~n852;
  assign n854 = n853 ^ n850;
  assign n855 = n851 & n854;
  assign n856 = n855 ^ n732;
  assign n857 = n856 ^ n684;
  assign n858 = ~n506 & n857;
  assign n860 = n859 ^ n858;
  assign n721 = n535 & n681;
  assign n722 = n633 & n680;
  assign n723 = ~n535 & n722;
  assign n724 = ~n721 & ~n723;
  assign n725 = n543 ^ n535;
  assign n726 = ~n724 & n725;
  assign n727 = n551 ^ n535;
  assign n728 = n694 & n727;
  assign n729 = ~n726 & ~n728;
  assign n715 = n521 & ~n536;
  assign n716 = n538 & n715;
  assign n717 = n521 ^ n506;
  assign n718 = n684 & n717;
  assign n719 = n718 ^ n506;
  assign n720 = ~n716 & n719;
  assign n730 = n729 ^ n720;
  assign n734 = n538 ^ n535;
  assign n735 = ~n724 & ~n734;
  assign n736 = n694 & n725;
  assign n737 = ~n735 & ~n736;
  assign n733 = ~n506 & n732;
  assign n738 = n737 ^ n733;
  assign n836 = n835 ^ n781;
  assign n837 = n781 ^ n633;
  assign n838 = n781 ^ n551;
  assign n839 = n837 & n838;
  assign n840 = n839 ^ n781;
  assign n841 = ~n836 & ~n840;
  assign n842 = n841 ^ n633;
  assign n843 = n842 ^ n733;
  assign n844 = n738 & ~n843;
  assign n845 = n844 ^ n737;
  assign n846 = n845 ^ n729;
  assign n847 = ~n730 & n846;
  assign n848 = n847 ^ n845;
  assign n861 = n860 ^ n848;
  assign n862 = n684 & ~n859;
  assign n863 = n861 & n862;
  assign n864 = ~n848 & n856;
  assign n865 = ~n863 & ~n864;
  assign n866 = ~n506 & ~n865;
  assign n867 = ~n848 & ~n858;
  assign n868 = ~n506 & ~n684;
  assign n869 = n856 & n868;
  assign n870 = ~n867 & ~n869;
  assign n871 = n859 & ~n870;
  assign n872 = ~n866 & ~n871;
  assign n689 = n506 & n688;
  assign n690 = ~n557 & n687;
  assign n691 = ~n684 & n690;
  assign n692 = ~n689 & ~n691;
  assign n693 = n548 & ~n692;
  assign n703 = ~n693 & ~n702;
  assign n705 = ~n689 & ~n704;
  assign n706 = ~n700 & ~n705;
  assign n713 = ~n706 & ~n712;
  assign n714 = n703 & n713;
  assign n873 = n872 ^ n714;
  assign n874 = ~n48 & ~n99;
  assign n875 = n69 & n156;
  assign n876 = ~n411 & ~n875;
  assign n877 = n180 & ~n876;
  assign n878 = ~n874 & ~n877;
  assign n879 = ~n822 & ~n878;
  assign n880 = n56 & ~n160;
  assign n881 = ~n51 & ~n880;
  assign n882 = ~n137 & ~n881;
  assign n883 = ~n281 & ~n470;
  assign n884 = ~n812 & n883;
  assign n885 = ~n283 & n884;
  assign n886 = ~n620 & n885;
  assign n887 = ~n882 & n886;
  assign n889 = ~n138 & ~n395;
  assign n890 = n888 & n889;
  assign n447 = n174 & n446;
  assign n891 = ~n230 & ~n273;
  assign n892 = ~n447 & n891;
  assign n893 = ~n209 & n892;
  assign n894 = n608 & n893;
  assign n895 = n890 & n894;
  assign n896 = n887 & n895;
  assign n897 = n879 & n896;
  assign n898 = n390 & n565;
  assign n899 = ~n324 & ~n394;
  assign n900 = ~n438 & ~n810;
  assign n901 = n899 & n900;
  assign n902 = n898 & n901;
  assign n903 = ~n282 & ~n362;
  assign n904 = n125 & n132;
  assign n905 = n83 & ~n904;
  assign n906 = n903 & ~n905;
  assign n907 = ~n308 & ~n351;
  assign n908 = ~n243 & ~n624;
  assign n909 = n907 & n908;
  assign n910 = n906 & n909;
  assign n911 = n902 & n910;
  assign n921 = ~n190 & ~n813;
  assign n922 = n495 & n904;
  assign n923 = n57 & ~n922;
  assign n924 = ~n231 & ~n923;
  assign n925 = n921 & n924;
  assign n928 = n925 & n927;
  assign n929 = n920 & n928;
  assign n930 = n911 & n929;
  assign n931 = n897 & n930;
  assign n932 = n85 & ~n157;
  assign n933 = ~n558 & ~n932;
  assign n934 = n666 & n933;
  assign n935 = n102 & ~n165;
  assign n936 = ~n191 & ~n935;
  assign n937 = n934 & n936;
  assign n941 = ~n418 & ~n562;
  assign n942 = n940 & n941;
  assign n943 = ~n298 & ~n344;
  assign n944 = ~n244 & ~n348;
  assign n945 = n943 & n944;
  assign n946 = n942 & n945;
  assign n947 = n937 & n946;
  assign n232 = ~n230 & ~n231;
  assign n233 = ~n226 & n232;
  assign n948 = ~n274 & ~n767;
  assign n419 = ~n120 & n168;
  assign n949 = n97 & n419;
  assign n950 = n85 & ~n949;
  assign n951 = n948 & ~n950;
  assign n952 = n233 & n951;
  assign n953 = n947 & n952;
  assign n954 = n879 & n953;
  assign n955 = n83 & ~n253;
  assign n956 = n338 & ~n955;
  assign n957 = n270 & n956;
  assign n958 = ~n363 & ~n531;
  assign n959 = n957 & n958;
  assign n960 = n151 & n181;
  assign n961 = ~n57 & n960;
  assign n962 = n181 & n186;
  assign n963 = ~n46 & n50;
  assign n964 = ~n962 & n963;
  assign n965 = ~n961 & n964;
  assign n966 = ~n238 & ~n431;
  assign n967 = ~n158 & n162;
  assign n968 = ~n395 & ~n967;
  assign n969 = n165 & n249;
  assign n970 = n56 & ~n969;
  assign n971 = n968 & ~n970;
  assign n972 = n966 & n971;
  assign n973 = ~n965 & n972;
  assign n974 = n959 & n973;
  assign n976 = n276 & n975;
  assign n977 = ~n48 & ~n162;
  assign n978 = ~n976 & ~n977;
  assign n979 = n974 & ~n978;
  assign n984 = n175 & ~n962;
  assign n985 = ~n675 & ~n984;
  assign n235 = n69 & n132;
  assign n986 = n91 & n235;
  assign n987 = n51 & ~n986;
  assign n988 = ~n254 & ~n987;
  assign n989 = n985 & n988;
  assign n990 = n983 & n989;
  assign n991 = n979 & n990;
  assign n992 = n954 & n991;
  assign n993 = ~n931 & ~n992;
  assign n199 = n78 & ~n198;
  assign n200 = ~n83 & ~n162;
  assign n201 = ~n199 & ~n200;
  assign n203 = ~n121 & ~n202;
  assign n204 = ~n201 & n203;
  assign n205 = ~n48 & ~n57;
  assign n206 = ~n180 & ~n205;
  assign n208 = ~n206 & ~n207;
  assign n212 = n162 & ~n211;
  assign n213 = ~n210 & ~n212;
  assign n214 = n137 & n168;
  assign n215 = n139 & ~n214;
  assign n216 = n213 & ~n215;
  assign n217 = ~n209 & n216;
  assign n218 = n208 & n217;
  assign n219 = n204 & n218;
  assign n220 = ~n83 & n219;
  assign n223 = ~n102 & ~n120;
  assign n224 = ~n222 & n223;
  assign n225 = ~n220 & ~n224;
  assign n236 = ~n85 & n235;
  assign n237 = ~n234 & ~n236;
  assign n994 = ~n470 & ~n786;
  assign n995 = ~n374 & n994;
  assign n996 = ~n255 & n995;
  assign n997 = n610 & n996;
  assign n998 = n85 & ~n211;
  assign n999 = ~n271 & ~n998;
  assign n1000 = ~n288 & n999;
  assign n1001 = ~n351 & n1000;
  assign n1002 = ~n85 & n249;
  assign n1003 = n69 & n150;
  assign n1004 = ~n56 & n1003;
  assign n1005 = ~n1002 & ~n1004;
  assign n1006 = ~n284 & ~n1005;
  assign n1007 = n125 & n168;
  assign n1008 = n162 & ~n1007;
  assign n1009 = n1006 & ~n1008;
  assign n1010 = n1001 & n1009;
  assign n1011 = n997 & n1010;
  assign n1012 = ~n237 & n1011;
  assign n1013 = ~n225 & n1012;
  assign n1014 = ~n352 & ~n606;
  assign n1015 = ~n454 & n1014;
  assign n1016 = n267 & n1015;
  assign n1017 = ~n140 & n958;
  assign n1018 = ~n297 & ~n638;
  assign n1019 = ~n281 & ~n531;
  assign n1020 = n1018 & n1019;
  assign n1021 = n1017 & n1020;
  assign n1022 = n1016 & n1021;
  assign n1034 = n580 & n890;
  assign n1035 = n1033 & n1034;
  assign n1036 = n1022 & n1035;
  assign n1037 = ~n57 & ~n282;
  assign n1038 = ~n182 & ~n1037;
  assign n1039 = n503 & ~n1038;
  assign n1041 = ~n566 & ~n1040;
  assign n1042 = n933 & n1041;
  assign n1043 = n1039 & n1042;
  assign n1044 = ~n756 & n927;
  assign n1045 = ~n394 & ~n822;
  assign n1046 = ~n393 & n1045;
  assign n1047 = n1044 & n1046;
  assign n1048 = n1043 & n1047;
  assign n1049 = n1036 & n1048;
  assign n1050 = n1013 & n1049;
  assign n1051 = n993 & n1050;
  assign n1052 = n931 & n992;
  assign n1053 = ~n1050 & n1052;
  assign n1054 = ~n1051 & ~n1053;
  assign n1055 = ~x22 & ~n28;
  assign n1056 = n1055 ^ x5;
  assign n1057 = n1056 ^ n1050;
  assign n1058 = ~n1054 & ~n1057;
  assign n1059 = n992 ^ n931;
  assign n1060 = ~x22 & ~n29;
  assign n1061 = n1060 ^ x6;
  assign n1062 = n1061 ^ n1050;
  assign n1063 = n1059 & ~n1062;
  assign n1064 = ~n1058 & ~n1063;
  assign n1065 = n343 & ~n756;
  assign n1066 = ~n939 & n948;
  assign n453 = ~n226 & ~n282;
  assign n1067 = n364 & n453;
  assign n1068 = n1066 & n1067;
  assign n1069 = n594 & n1068;
  assign n1070 = n102 & ~n753;
  assign n1071 = ~n272 & ~n1070;
  assign n1072 = ~n284 & n1071;
  assign n1073 = n147 ^ n57;
  assign n1074 = n147 ^ n125;
  assign n1075 = n1074 ^ n125;
  assign n1076 = n977 ^ n125;
  assign n1077 = ~n1075 & ~n1076;
  assign n1078 = n1077 ^ n125;
  assign n1079 = ~n1073 & n1078;
  assign n1080 = n1079 ^ n57;
  assign n1081 = n1072 & ~n1080;
  assign n1082 = n1069 & n1081;
  assign n1083 = n78 & ~n120;
  assign n1084 = ~n50 & ~n1083;
  assign n1085 = ~n101 & ~n1084;
  assign n1086 = ~n50 & ~n174;
  assign n1087 = ~n1083 & ~n1086;
  assign n1088 = n156 & ~n1087;
  assign n1089 = ~n1085 & ~n1088;
  assign n1090 = n139 & ~n406;
  assign n1091 = ~n656 & ~n1090;
  assign n1092 = ~n1089 & n1091;
  assign n1093 = n483 & n1092;
  assign n1094 = n1082 & n1093;
  assign n1095 = n1065 & n1094;
  assign n1099 = x6 & ~x22;
  assign n1100 = ~n1060 & ~n1099;
  assign n1101 = n1100 ^ x7;
  assign n1096 = ~x22 & ~n31;
  assign n1097 = n1096 ^ x8;
  assign n1098 = n1097 ^ n931;
  assign n1102 = n1101 ^ n1098;
  assign n1103 = n1102 ^ n1098;
  assign n1104 = n1098 ^ n1097;
  assign n1105 = n1103 & ~n1104;
  assign n1106 = n1105 ^ n1098;
  assign n1107 = n1095 & ~n1106;
  assign n1108 = n1107 ^ n1098;
  assign n1109 = ~n1064 & ~n1108;
  assign n1110 = ~n198 & ~n375;
  assign n1111 = ~n625 & ~n771;
  assign n1112 = n1110 & n1111;
  assign n1113 = ~n207 & ~n230;
  assign n1114 = n503 & n1113;
  assign n1115 = n1112 & n1114;
  assign n1116 = n901 & n1115;
  assign n420 = n175 & ~n419;
  assign n421 = ~n418 & ~n420;
  assign n1117 = ~n329 & n421;
  assign n1118 = ~n395 & n1117;
  assign n1119 = ~n624 & ~n821;
  assign n1120 = n996 & n1119;
  assign n1121 = n1118 & n1120;
  assign n1122 = n1116 & n1121;
  assign n1123 = ~n254 & ~n272;
  assign n1124 = ~n290 & ~n323;
  assign n1125 = ~n524 & n1124;
  assign n1126 = n1123 & n1125;
  assign n1127 = n189 & n1126;
  assign n1128 = ~n180 & n1086;
  assign n1129 = ~n356 & ~n1128;
  assign n1130 = ~n643 & n1129;
  assign n1131 = n1127 & n1130;
  assign n1132 = n102 & ~n510;
  assign n1133 = ~n298 & ~n1132;
  assign n1134 = ~n341 & ~n467;
  assign n1135 = n1133 & n1134;
  assign n1136 = n907 & n966;
  assign n1137 = n1135 & n1136;
  assign n1138 = n125 & n365;
  assign n1139 = n139 & ~n1138;
  assign n1140 = ~n663 & ~n1139;
  assign n1141 = n51 & ~n493;
  assign n1142 = n85 & ~n132;
  assign n1143 = ~n1141 & ~n1142;
  assign n1144 = n1140 & n1143;
  assign n1145 = n792 & n1144;
  assign n1146 = n1137 & n1145;
  assign n1147 = n1131 & n1146;
  assign n1148 = n1122 & n1147;
  assign n1149 = ~n1050 & ~n1148;
  assign n1150 = ~n835 & ~n1149;
  assign n1151 = ~x22 & ~n26;
  assign n1152 = n1151 ^ x3;
  assign n1153 = n1148 ^ n1050;
  assign n1154 = n1152 & n1153;
  assign n1155 = n1150 & ~n1154;
  assign n1156 = ~x22 & ~n27;
  assign n1157 = n1156 ^ x4;
  assign n1158 = n1157 ^ n835;
  assign n1159 = n1153 & ~n1158;
  assign n1160 = n835 & n1149;
  assign n1161 = n1160 ^ n1152;
  assign n1162 = n1161 ^ n1160;
  assign n1163 = n1050 & n1148;
  assign n1164 = ~n835 & n1163;
  assign n1165 = n1164 ^ n1160;
  assign n1166 = ~n1162 & n1165;
  assign n1167 = n1166 ^ n1160;
  assign n1168 = ~n1159 & ~n1167;
  assign n1169 = n1155 & ~n1168;
  assign n1170 = n1109 & n1169;
  assign n1171 = n836 & n1152;
  assign n1172 = n1108 ^ n1064;
  assign n1173 = ~n1155 & n1168;
  assign n1174 = n1173 ^ n1108;
  assign n1175 = n1172 & ~n1174;
  assign n1176 = n1175 ^ n1064;
  assign n1177 = n1171 & ~n1176;
  assign n1178 = ~n1170 & ~n1177;
  assign n1184 = ~n1054 & ~n1062;
  assign n1185 = n1101 ^ n1050;
  assign n1186 = n1059 & n1185;
  assign n1187 = ~n1184 & ~n1186;
  assign n1179 = ~n1160 & ~n1164;
  assign n1180 = ~n1158 & ~n1179;
  assign n1181 = n1056 ^ n835;
  assign n1182 = n1153 & ~n1181;
  assign n1183 = ~n1180 & ~n1182;
  assign n1188 = n1187 ^ n1183;
  assign n1189 = n931 ^ n732;
  assign n1190 = n1189 ^ n1097;
  assign n1191 = n1190 ^ n1189;
  assign n1192 = n1189 ^ n732;
  assign n1193 = ~n1191 & ~n1192;
  assign n1194 = n1193 ^ n1189;
  assign n1195 = n1095 & ~n1194;
  assign n1196 = n1195 ^ n1189;
  assign n1197 = n1196 ^ n1183;
  assign n1198 = n1188 & ~n1197;
  assign n1199 = n1198 ^ n1187;
  assign n1200 = n1178 & n1199;
  assign n1202 = n1097 ^ n1050;
  assign n1254 = ~n1054 & ~n1202;
  assign n1255 = n1050 ^ n732;
  assign n1256 = n1059 & ~n1255;
  assign n1257 = ~n1254 & ~n1256;
  assign n1246 = n931 ^ n684;
  assign n1247 = n1246 ^ n850;
  assign n1248 = n1247 ^ n1246;
  assign n1249 = n1246 ^ n684;
  assign n1250 = ~n1248 & ~n1249;
  assign n1251 = n1250 ^ n1246;
  assign n1252 = n1095 & ~n1251;
  assign n1253 = n1252 ^ n1246;
  assign n1258 = n1257 ^ n1253;
  assign n1206 = n1061 ^ n835;
  assign n1242 = ~n1179 & ~n1206;
  assign n1243 = n1101 ^ n835;
  assign n1244 = n1153 & n1243;
  assign n1245 = ~n1242 & ~n1244;
  assign n1259 = n1258 ^ n1245;
  assign n1213 = n781 & n835;
  assign n1214 = ~n633 & n1213;
  assign n1231 = n853 & ~n1152;
  assign n1232 = ~n1214 & ~n1231;
  assign n1233 = n931 ^ n850;
  assign n1234 = n1233 ^ n732;
  assign n1235 = n1234 ^ n1233;
  assign n1236 = n1233 ^ n850;
  assign n1237 = ~n1235 & ~n1236;
  assign n1238 = n1237 ^ n1233;
  assign n1239 = n1095 & ~n1238;
  assign n1240 = n1239 ^ n1233;
  assign n1241 = ~n1232 & ~n1240;
  assign n1260 = n1259 ^ n1241;
  assign n1210 = n1157 ^ n633;
  assign n1212 = n633 & n852;
  assign n1225 = ~n1212 & ~n1214;
  assign n1226 = ~n1210 & ~n1225;
  assign n1227 = n1056 ^ n633;
  assign n1228 = n836 & ~n1227;
  assign n1229 = ~n1226 & ~n1228;
  assign n1224 = n694 & n1152;
  assign n1230 = n1229 ^ n1224;
  assign n1261 = n1260 ^ n1230;
  assign n1205 = ~n1179 & ~n1181;
  assign n1207 = n1153 & ~n1206;
  assign n1208 = ~n1205 & ~n1207;
  assign n1201 = ~n1054 & n1185;
  assign n1203 = n1059 & ~n1202;
  assign n1204 = ~n1201 & ~n1203;
  assign n1209 = n1208 ^ n1204;
  assign n1211 = n836 & ~n1210;
  assign n1215 = n1214 ^ n1212;
  assign n1216 = n1214 ^ n1152;
  assign n1217 = n1216 ^ n1214;
  assign n1218 = n1215 & n1217;
  assign n1219 = n1218 ^ n1214;
  assign n1220 = ~n1211 & ~n1219;
  assign n1221 = n1220 ^ n1204;
  assign n1222 = n1209 & ~n1221;
  assign n1223 = n1222 ^ n1208;
  assign n1262 = n1261 ^ n1223;
  assign n1263 = ~n1200 & ~n1262;
  assign n1268 = n1196 ^ n1188;
  assign n1264 = n1176 ^ n1171;
  assign n1265 = n1264 ^ n1109;
  assign n1266 = ~n1169 & n1265;
  assign n1267 = n1266 ^ n1109;
  assign n1269 = n1268 ^ n1267;
  assign n1270 = n1056 & n1095;
  assign n1272 = n1061 & n1095;
  assign n1271 = n1061 ^ n931;
  assign n1273 = n1272 ^ n1271;
  assign n1274 = ~n1270 & ~n1273;
  assign n1283 = n1157 ^ n1050;
  assign n1284 = ~n1054 & ~n1283;
  assign n1285 = ~n1057 & n1059;
  assign n1286 = ~n1284 & ~n1285;
  assign n1275 = n1101 ^ n931;
  assign n1276 = n1275 ^ n1061;
  assign n1277 = n1276 ^ n1275;
  assign n1278 = n1275 ^ n1101;
  assign n1279 = ~n1277 & ~n1278;
  assign n1280 = n1279 ^ n1275;
  assign n1281 = n1095 & n1280;
  assign n1282 = n1281 ^ n1275;
  assign n1287 = n1286 ^ n1282;
  assign n1288 = ~n993 & ~n1050;
  assign n1289 = ~n1052 & n1152;
  assign n1290 = n1288 & ~n1289;
  assign n1291 = ~n1154 & ~n1290;
  assign n1292 = ~n1287 & ~n1291;
  assign n1293 = ~n1274 & ~n1292;
  assign n1294 = n1059 & ~n1283;
  assign n1295 = n1053 ^ n1051;
  assign n1296 = n1152 ^ n1053;
  assign n1297 = n1296 ^ n1053;
  assign n1298 = n1295 & n1297;
  assign n1299 = n1298 ^ n1053;
  assign n1300 = ~n1294 & ~n1299;
  assign n1301 = n1287 & n1300;
  assign n1302 = ~n1290 & n1301;
  assign n1303 = ~n1293 & ~n1302;
  assign n1304 = ~n1287 & ~n1300;
  assign n1305 = ~n1154 & ~n1304;
  assign n1306 = n1303 & ~n1305;
  assign n1308 = ~n992 & n1152;
  assign n1307 = n1056 & ~n1095;
  assign n1309 = n1308 ^ n1307;
  assign n1310 = n1152 ^ n1095;
  assign n1311 = n1095 ^ n931;
  assign n1312 = ~n1095 & n1311;
  assign n1313 = n1312 ^ n1095;
  assign n1314 = ~n1310 & ~n1313;
  assign n1315 = n1314 ^ n1312;
  assign n1316 = n1315 ^ n1095;
  assign n1317 = n1316 ^ n931;
  assign n1318 = n1157 & n1317;
  assign n1319 = n1318 ^ n931;
  assign n1320 = n1319 ^ n1307;
  assign n1321 = n1320 ^ n1319;
  assign n1322 = n1319 ^ n931;
  assign n1323 = n1321 & ~n1322;
  assign n1324 = n1323 ^ n1319;
  assign n1325 = ~n1309 & ~n1324;
  assign n1326 = ~n1306 & ~n1325;
  assign n1327 = ~n1301 & ~n1305;
  assign n1328 = ~n1274 & ~n1327;
  assign n1329 = n1282 & ~n1286;
  assign n1330 = n1168 ^ n1155;
  assign n1331 = n1330 ^ n1172;
  assign n1332 = ~n1329 & n1331;
  assign n1333 = n1287 & n1291;
  assign n1334 = ~n1332 & ~n1333;
  assign n1335 = ~n1328 & n1334;
  assign n1336 = ~n1326 & n1335;
  assign n1337 = n1336 ^ n1268;
  assign n1338 = n1337 ^ n1268;
  assign n1339 = n1274 & n1290;
  assign n1340 = n1339 ^ n1282;
  assign n1341 = ~n1287 & ~n1340;
  assign n1342 = n1341 ^ n1286;
  assign n1343 = ~n1331 & ~n1342;
  assign n1344 = n1343 ^ n1268;
  assign n1345 = n1344 ^ n1268;
  assign n1346 = ~n1338 & ~n1345;
  assign n1347 = n1346 ^ n1268;
  assign n1348 = n1269 & ~n1347;
  assign n1349 = n1348 ^ n1267;
  assign n1350 = ~n1263 & n1349;
  assign n1351 = ~n1178 & ~n1199;
  assign n1352 = n1262 & ~n1351;
  assign n1353 = n1240 ^ n1232;
  assign n1354 = n1220 ^ n1209;
  assign n1355 = ~n1353 & n1354;
  assign n1356 = ~n1352 & ~n1355;
  assign n1357 = ~n1350 & n1356;
  assign n1358 = n1353 & ~n1354;
  assign n1359 = n1358 ^ n1262;
  assign n1360 = n1358 ^ n1200;
  assign n1361 = n1360 ^ n1358;
  assign n1362 = n1349 & ~n1351;
  assign n1363 = n1362 ^ n1358;
  assign n1364 = n1363 ^ n1358;
  assign n1365 = ~n1361 & ~n1364;
  assign n1366 = n1365 ^ n1358;
  assign n1367 = ~n1359 & ~n1366;
  assign n1368 = n1367 ^ n1262;
  assign n1369 = ~n1357 & n1368;
  assign n1379 = ~n1225 & ~n1227;
  assign n1380 = n1061 ^ n633;
  assign n1381 = n836 & ~n1380;
  assign n1382 = ~n1379 & ~n1381;
  assign n1374 = ~n1179 & n1243;
  assign n1375 = n1097 ^ n835;
  assign n1376 = n1153 & ~n1375;
  assign n1377 = ~n1374 & ~n1376;
  assign n1370 = ~n1054 & ~n1255;
  assign n1371 = n1050 ^ n850;
  assign n1372 = n1059 & ~n1371;
  assign n1373 = ~n1370 & ~n1372;
  assign n1378 = n1377 ^ n1373;
  assign n1383 = n1382 ^ n1378;
  assign n1384 = n1369 & n1383;
  assign n1421 = n1253 ^ n1245;
  assign n1422 = n1258 & ~n1421;
  assign n1423 = n1422 ^ n1257;
  assign n1390 = n931 ^ n538;
  assign n1391 = n1390 ^ n684;
  assign n1392 = n1391 ^ n1390;
  assign n1393 = n1390 ^ n538;
  assign n1394 = ~n1392 & ~n1393;
  assign n1395 = n1394 ^ n1390;
  assign n1396 = n1095 & ~n1395;
  assign n1397 = n1396 ^ n1390;
  assign n1389 = n682 & ~n1224;
  assign n1419 = n1397 ^ n1389;
  assign n1411 = n1157 ^ n535;
  assign n1412 = n694 & ~n1411;
  assign n1413 = n1152 ^ n721;
  assign n1414 = n1413 ^ n721;
  assign n1415 = n723 ^ n721;
  assign n1416 = ~n1414 & n1415;
  assign n1417 = n1416 ^ n721;
  assign n1418 = ~n1412 & ~n1417;
  assign n1420 = n1419 ^ n1418;
  assign n1447 = n1423 ^ n1420;
  assign n1440 = ~n724 & ~n1411;
  assign n1441 = n1056 ^ n535;
  assign n1442 = n694 & ~n1441;
  assign n1443 = ~n1440 & ~n1442;
  assign n1435 = ~n1054 & ~n1371;
  assign n1436 = n1050 ^ n684;
  assign n1437 = n1059 & ~n1436;
  assign n1438 = ~n1435 & ~n1437;
  assign n1427 = n931 ^ n543;
  assign n1428 = n1427 ^ n538;
  assign n1429 = n1428 ^ n1427;
  assign n1430 = n1427 ^ n543;
  assign n1431 = ~n1429 & ~n1430;
  assign n1432 = n1431 ^ n1427;
  assign n1433 = n1095 & n1432;
  assign n1434 = n1433 ^ n1427;
  assign n1439 = n1438 ^ n1434;
  assign n1444 = n1443 ^ n1439;
  assign n1424 = n1423 ^ n1418;
  assign n1425 = ~n1420 & n1424;
  assign n1426 = n1425 ^ n1423;
  assign n1445 = n1444 ^ n1426;
  assign n1403 = ~n1225 & ~n1380;
  assign n1404 = n1101 ^ n633;
  assign n1405 = n836 & n1404;
  assign n1406 = ~n1403 & ~n1405;
  assign n1399 = ~n1179 & ~n1375;
  assign n1400 = n835 ^ n732;
  assign n1401 = n1153 & ~n1400;
  assign n1402 = ~n1399 & ~n1401;
  assign n1407 = n1406 ^ n1402;
  assign n1398 = n1389 & ~n1397;
  assign n1408 = n1407 ^ n1398;
  assign n1388 = n715 & n1152;
  assign n1409 = n1408 ^ n1388;
  assign n1385 = n1382 ^ n1377;
  assign n1386 = ~n1378 & n1385;
  assign n1387 = n1386 ^ n1382;
  assign n1410 = n1409 ^ n1387;
  assign n1446 = n1445 ^ n1410;
  assign n1448 = n1447 ^ n1446;
  assign n1449 = n1223 & n1259;
  assign n1450 = n1241 ^ n1229;
  assign n1451 = n1230 & ~n1450;
  assign n1452 = n1451 ^ n1241;
  assign n1453 = n1449 & ~n1452;
  assign n1454 = ~n1223 & ~n1259;
  assign n1455 = ~n1224 & n1229;
  assign n1456 = ~n1241 & n1455;
  assign n1457 = ~n1454 & n1456;
  assign n1458 = ~n1453 & ~n1457;
  assign n1459 = n1458 ^ n1446;
  assign n1460 = n1459 ^ n1458;
  assign n1461 = n1452 & n1454;
  assign n1462 = n1224 & ~n1229;
  assign n1463 = n1241 & n1462;
  assign n1464 = ~n1449 & n1463;
  assign n1465 = ~n1461 & ~n1464;
  assign n1466 = n1465 ^ n1458;
  assign n1467 = ~n1460 & n1466;
  assign n1468 = n1467 ^ n1458;
  assign n1469 = ~n1448 & n1468;
  assign n1470 = n1469 ^ n1447;
  assign n1471 = ~n1384 & ~n1470;
  assign n1472 = ~n1447 & n1458;
  assign n1473 = n1465 & ~n1472;
  assign n1474 = n1473 ^ n1446;
  assign n1475 = n1473 ^ n1383;
  assign n1476 = n1475 ^ n1473;
  assign n1477 = n1473 ^ n1369;
  assign n1478 = n1477 ^ n1473;
  assign n1479 = ~n1476 & ~n1478;
  assign n1480 = n1479 ^ n1473;
  assign n1481 = ~n1474 & n1480;
  assign n1482 = n1481 ^ n1446;
  assign n1483 = ~n1471 & ~n1482;
  assign n1505 = ~n1054 & ~n1436;
  assign n1506 = n1050 ^ n538;
  assign n1507 = n1059 & ~n1506;
  assign n1508 = ~n1505 & ~n1507;
  assign n1495 = n931 ^ n551;
  assign n1496 = n1495 ^ n543;
  assign n1497 = n1496 ^ n1495;
  assign n1498 = n1495 ^ n551;
  assign n1499 = n1497 & ~n1498;
  assign n1500 = n1499 ^ n1495;
  assign n1501 = n1095 & n1500;
  assign n1502 = n1501 ^ n1495;
  assign n1503 = n1502 ^ n506;
  assign n1484 = n506 & n536;
  assign n1485 = n1152 ^ n506;
  assign n1486 = n1485 ^ n521;
  assign n1487 = n1486 ^ n1485;
  assign n1488 = n1485 ^ n1157;
  assign n1489 = n1488 ^ n1485;
  assign n1490 = n1487 & n1489;
  assign n1491 = n1490 ^ n1485;
  assign n1492 = ~n717 & ~n1491;
  assign n1493 = n1492 ^ n1485;
  assign n1494 = ~n1484 & ~n1493;
  assign n1504 = n1503 ^ n1494;
  assign n1509 = n1508 ^ n1504;
  assign n1510 = n1444 ^ n1410;
  assign n1511 = ~n1445 & n1510;
  assign n1512 = n1511 ^ n1426;
  assign n1513 = ~n1509 & n1512;
  assign n1576 = ~n506 & n1502;
  assign n1569 = ~n506 & ~n1157;
  assign n1570 = n536 & ~n1569;
  assign n1571 = n506 & ~n1056;
  assign n1572 = n1571 ^ n1157;
  assign n1573 = n521 & ~n1572;
  assign n1574 = n1573 ^ n1157;
  assign n1575 = ~n1570 & n1574;
  assign n1577 = n1576 ^ n1575;
  assign n1521 = ~n1225 & n1404;
  assign n1522 = n1097 ^ n633;
  assign n1523 = n836 & ~n1522;
  assign n1524 = ~n1521 & ~n1523;
  assign n1517 = ~n1179 & ~n1400;
  assign n1518 = n850 ^ n835;
  assign n1519 = n1153 & ~n1518;
  assign n1520 = ~n1517 & ~n1519;
  assign n1525 = n1524 ^ n1520;
  assign n1526 = ~n724 & ~n1441;
  assign n1527 = n1061 ^ n535;
  assign n1528 = n694 & ~n1527;
  assign n1529 = ~n1526 & ~n1528;
  assign n1566 = n1529 ^ n1524;
  assign n1567 = ~n1525 & n1566;
  assign n1568 = n1567 ^ n1529;
  assign n1578 = n1577 ^ n1568;
  assign n1559 = ~n1054 & ~n1506;
  assign n1560 = n1050 ^ n543;
  assign n1561 = n1059 & n1560;
  assign n1562 = ~n1559 & ~n1561;
  assign n1557 = ~n506 & n1152;
  assign n1555 = ~n551 & n1095;
  assign n1556 = ~n931 & ~n1555;
  assign n1558 = n1557 ^ n1556;
  assign n1563 = n1562 ^ n1558;
  assign n1552 = n1508 ^ n1503;
  assign n1553 = n1504 & n1552;
  assign n1554 = n1553 ^ n1508;
  assign n1564 = n1563 ^ n1554;
  assign n1547 = ~n724 & ~n1527;
  assign n1548 = n1101 ^ n535;
  assign n1549 = n694 & n1548;
  assign n1550 = ~n1547 & ~n1549;
  assign n1542 = ~n1225 & ~n1522;
  assign n1543 = n732 ^ n633;
  assign n1544 = n836 & ~n1543;
  assign n1545 = ~n1542 & ~n1544;
  assign n1538 = ~n1179 & ~n1518;
  assign n1539 = n835 ^ n684;
  assign n1540 = n1153 & ~n1539;
  assign n1541 = ~n1538 & ~n1540;
  assign n1546 = n1545 ^ n1541;
  assign n1551 = n1550 ^ n1546;
  assign n1565 = n1564 ^ n1551;
  assign n1579 = n1578 ^ n1565;
  assign n1530 = n1529 ^ n1525;
  assign n1514 = n1402 ^ n1398;
  assign n1515 = n1407 & n1514;
  assign n1516 = n1515 ^ n1406;
  assign n1531 = n1530 ^ n1516;
  assign n1532 = n1443 ^ n1438;
  assign n1533 = n1439 & n1532;
  assign n1534 = n1533 ^ n1443;
  assign n1535 = n1534 ^ n1530;
  assign n1536 = n1531 & ~n1535;
  assign n1537 = n1536 ^ n1516;
  assign n1580 = n1579 ^ n1537;
  assign n1581 = ~n1513 & ~n1580;
  assign n1582 = n1483 & ~n1581;
  assign n1583 = n1509 & ~n1512;
  assign n1584 = n1580 & ~n1583;
  assign n1585 = n1534 ^ n1531;
  assign n1586 = n1388 ^ n1387;
  assign n1587 = n1409 & n1586;
  assign n1588 = n1587 ^ n1408;
  assign n1589 = n1585 & ~n1588;
  assign n1590 = ~n1584 & ~n1589;
  assign n1591 = ~n1582 & n1590;
  assign n1592 = ~n1585 & n1588;
  assign n1593 = n1592 ^ n1580;
  assign n1594 = n1512 ^ n1483;
  assign n1595 = n1512 ^ n1509;
  assign n1596 = n1594 & n1595;
  assign n1597 = n1596 ^ n1483;
  assign n1598 = n1597 ^ n1580;
  assign n1599 = ~n1593 & n1598;
  assign n1600 = n1599 ^ n1580;
  assign n1601 = ~n1591 & n1600;
  assign n1602 = n1563 ^ n1551;
  assign n1603 = n1564 & ~n1602;
  assign n1604 = n1603 ^ n1554;
  assign n1605 = n1601 & n1604;
  assign n1650 = n715 & n1061;
  assign n1651 = n717 & n1056;
  assign n1652 = n1651 ^ n506;
  assign n1653 = ~n1650 & n1652;
  assign n1646 = n1562 ^ n1557;
  assign n1647 = n1562 ^ n1556;
  assign n1648 = ~n1646 & n1647;
  assign n1649 = n1648 ^ n1557;
  assign n1654 = n1653 ^ n1649;
  assign n1643 = n1550 ^ n1545;
  assign n1644 = ~n1546 & n1643;
  assign n1645 = n1644 ^ n1550;
  assign n1655 = n1654 ^ n1645;
  assign n1636 = ~n724 & n1548;
  assign n1637 = n1097 ^ n535;
  assign n1638 = n694 & ~n1637;
  assign n1639 = ~n1636 & ~n1638;
  assign n1631 = ~n1225 & ~n1543;
  assign n1632 = n850 ^ n633;
  assign n1633 = n836 & ~n1632;
  assign n1634 = ~n1631 & ~n1633;
  assign n1627 = ~n1179 & ~n1539;
  assign n1628 = n835 ^ n538;
  assign n1629 = n1153 & ~n1628;
  assign n1630 = ~n1627 & ~n1629;
  assign n1635 = n1634 ^ n1630;
  assign n1640 = n1639 ^ n1635;
  assign n1610 = ~n1051 & ~n1052;
  assign n1611 = ~n543 & ~n1610;
  assign n1612 = n1050 ^ n931;
  assign n1613 = n1612 ^ n551;
  assign n1614 = n1613 ^ n992;
  assign n1615 = n1614 ^ n1050;
  assign n1616 = n1615 ^ n551;
  assign n1617 = n992 ^ n551;
  assign n1618 = n1617 ^ n551;
  assign n1619 = n1050 ^ n551;
  assign n1620 = n1619 ^ n551;
  assign n1621 = ~n1618 & ~n1620;
  assign n1622 = n1621 ^ n551;
  assign n1623 = ~n1616 & ~n1622;
  assign n1624 = n1623 ^ n1613;
  assign n1625 = ~n1611 & ~n1624;
  assign n1609 = ~n506 & n1157;
  assign n1626 = n1625 ^ n1609;
  assign n1641 = n1640 ^ n1626;
  assign n1606 = n1576 ^ n1568;
  assign n1607 = ~n1577 & ~n1606;
  assign n1608 = n1607 ^ n1568;
  assign n1642 = n1641 ^ n1608;
  assign n1656 = n1655 ^ n1642;
  assign n1657 = n1578 ^ n1537;
  assign n1658 = ~n1579 & n1657;
  assign n1659 = n1658 ^ n1537;
  assign n1660 = n1659 ^ n1655;
  assign n1661 = ~n1656 & ~n1660;
  assign n1662 = n1661 ^ n1659;
  assign n1663 = ~n1605 & ~n1662;
  assign n1706 = ~n724 & ~n1637;
  assign n1707 = n732 ^ n535;
  assign n1708 = n694 & ~n1707;
  assign n1709 = ~n1706 & ~n1708;
  assign n1701 = ~n1225 & ~n1632;
  assign n1702 = n684 ^ n633;
  assign n1703 = n836 & ~n1702;
  assign n1704 = ~n1701 & ~n1703;
  assign n1697 = ~n1179 & ~n1628;
  assign n1698 = n835 ^ n543;
  assign n1699 = n1153 & n1698;
  assign n1700 = ~n1697 & ~n1699;
  assign n1705 = n1704 ^ n1700;
  assign n1710 = n1709 ^ n1705;
  assign n1673 = n992 & ~n1050;
  assign n1691 = ~n931 & n1673;
  assign n1692 = n931 & n1050;
  assign n1693 = ~n1691 & ~n1692;
  assign n1694 = ~n551 & ~n1610;
  assign n1695 = n1693 & ~n1694;
  assign n1690 = ~n506 & n1056;
  assign n1696 = n1695 ^ n1690;
  assign n1711 = n1710 ^ n1696;
  assign n1687 = n1653 ^ n1645;
  assign n1688 = ~n1654 & ~n1687;
  assign n1689 = n1688 ^ n1649;
  assign n1712 = n1711 ^ n1689;
  assign n1681 = n715 & ~n1101;
  assign n1682 = n717 & n1061;
  assign n1683 = n1682 ^ n506;
  assign n1684 = ~n1681 & n1683;
  assign n1678 = n1639 ^ n1634;
  assign n1679 = ~n1635 & n1678;
  assign n1680 = n1679 ^ n1639;
  assign n1685 = n1684 ^ n1680;
  assign n1667 = n1609 ^ n931;
  assign n1668 = ~n992 & ~n1667;
  assign n1669 = n1668 ^ n931;
  assign n1670 = ~n1626 & ~n1669;
  assign n1671 = ~n543 & n1051;
  assign n1672 = ~n1609 & ~n1671;
  assign n1674 = n543 & n1673;
  assign n1675 = n931 & ~n1674;
  assign n1676 = ~n1672 & ~n1675;
  assign n1677 = ~n1670 & ~n1676;
  assign n1686 = n1685 ^ n1677;
  assign n1713 = n1712 ^ n1686;
  assign n1664 = n1640 ^ n1608;
  assign n1665 = n1641 & n1664;
  assign n1666 = n1665 ^ n1608;
  assign n1714 = n1713 ^ n1666;
  assign n1715 = ~n1663 & n1714;
  assign n1716 = ~n1601 & ~n1604;
  assign n1717 = n1655 & ~n1659;
  assign n1718 = n1642 & n1717;
  assign n1719 = ~n1655 & n1659;
  assign n1720 = ~n1642 & n1719;
  assign n1721 = ~n1718 & ~n1720;
  assign n1722 = n1714 & n1721;
  assign n1723 = n1722 ^ n1720;
  assign n1724 = ~n1716 & n1723;
  assign n1725 = n1605 & n1662;
  assign n1726 = ~n1724 & ~n1725;
  assign n1727 = ~n1715 & n1726;
  assign n1744 = ~n724 & ~n1707;
  assign n1745 = n850 ^ n535;
  assign n1746 = n694 & ~n1745;
  assign n1747 = ~n1744 & ~n1746;
  assign n1739 = ~n1179 & n1698;
  assign n1740 = n835 ^ n551;
  assign n1741 = n1153 & n1740;
  assign n1742 = ~n1739 & ~n1741;
  assign n1734 = n544 & ~n1097;
  assign n1735 = n717 & n1101;
  assign n1736 = n1735 ^ n506;
  assign n1737 = ~n1734 & n1736;
  assign n1738 = ~n1484 & n1737;
  assign n1743 = n1742 ^ n1738;
  assign n1748 = n1747 ^ n1743;
  assign n1731 = n1709 ^ n1704;
  assign n1732 = ~n1705 & n1731;
  assign n1733 = n1732 ^ n1709;
  assign n1749 = n1748 ^ n1733;
  assign n1728 = n1684 ^ n1677;
  assign n1729 = n1685 & ~n1728;
  assign n1730 = n1729 ^ n1680;
  assign n1750 = n1749 ^ n1730;
  assign n1751 = ~n1727 & ~n1750;
  assign n1761 = n931 & ~n1695;
  assign n1762 = ~n1690 & ~n1694;
  assign n1763 = ~n1761 & ~n1762;
  assign n1764 = ~n1691 & n1763;
  assign n1765 = ~n1692 & ~n1764;
  assign n1756 = ~n1225 & ~n1702;
  assign n1757 = n633 ^ n538;
  assign n1758 = n836 & ~n1757;
  assign n1759 = ~n1756 & ~n1758;
  assign n1755 = ~n506 & n1061;
  assign n1760 = n1759 ^ n1755;
  assign n1766 = n1765 ^ n1760;
  assign n1752 = n1710 ^ n1689;
  assign n1753 = n1711 & ~n1752;
  assign n1754 = n1753 ^ n1689;
  assign n1767 = n1766 ^ n1754;
  assign n1768 = n1712 ^ n1666;
  assign n1769 = ~n1713 & n1768;
  assign n1770 = n1769 ^ n1666;
  assign n1771 = n1770 ^ n1754;
  assign n1772 = n1767 & ~n1771;
  assign n1773 = n1772 ^ n1770;
  assign n1774 = ~n1751 & ~n1773;
  assign n1810 = ~n1755 & n1764;
  assign n1811 = n1755 ^ n1692;
  assign n1812 = ~n1763 & n1811;
  assign n1813 = ~n1759 & ~n1812;
  assign n1814 = ~n1810 & ~n1813;
  assign n1815 = ~n1755 & n1759;
  assign n1816 = n1691 & ~n1815;
  assign n1817 = n1814 & ~n1816;
  assign n1803 = ~n724 & ~n1745;
  assign n1804 = n684 ^ n535;
  assign n1805 = n694 & ~n1804;
  assign n1806 = ~n1803 & ~n1805;
  assign n1800 = ~n1692 & ~n1755;
  assign n1801 = ~n1691 & ~n1800;
  assign n1794 = ~n506 & ~n1097;
  assign n1795 = n536 & ~n1794;
  assign n1796 = n544 & ~n732;
  assign n1797 = ~n521 & ~n1097;
  assign n1798 = ~n1796 & ~n1797;
  assign n1799 = ~n1795 & n1798;
  assign n1802 = n1801 ^ n1799;
  assign n1807 = n1806 ^ n1802;
  assign n1789 = ~n1225 & ~n1757;
  assign n1790 = n633 ^ n543;
  assign n1791 = n836 & n1790;
  assign n1792 = ~n1789 & ~n1791;
  assign n1787 = ~n506 & ~n1101;
  assign n1781 = n1148 ^ n835;
  assign n1782 = n1148 ^ n551;
  assign n1783 = n1781 & n1782;
  assign n1784 = n1783 ^ n1148;
  assign n1785 = ~n1153 & ~n1784;
  assign n1786 = n1785 ^ n835;
  assign n1788 = n1787 ^ n1786;
  assign n1793 = n1792 ^ n1788;
  assign n1808 = n1807 ^ n1793;
  assign n1778 = n1747 ^ n1742;
  assign n1779 = n1743 & n1778;
  assign n1780 = n1779 ^ n1747;
  assign n1809 = n1808 ^ n1780;
  assign n1818 = n1817 ^ n1809;
  assign n1775 = n1733 ^ n1730;
  assign n1776 = n1749 & n1775;
  assign n1777 = n1776 ^ n1730;
  assign n1819 = n1818 ^ n1777;
  assign n1820 = ~n1774 & n1819;
  assign n1821 = n1727 & n1750;
  assign n1822 = n1754 & ~n1766;
  assign n1823 = ~n1770 & n1822;
  assign n1824 = ~n1754 & n1766;
  assign n1825 = n1770 & n1824;
  assign n1826 = ~n1819 & ~n1825;
  assign n1827 = ~n1823 & ~n1826;
  assign n1828 = ~n1821 & n1827;
  assign n1829 = n1751 & n1773;
  assign n1830 = ~n1828 & ~n1829;
  assign n1831 = ~n1820 & n1830;
  assign n1867 = n521 & ~n850;
  assign n1868 = ~n536 & n850;
  assign n1869 = ~n1867 & ~n1868;
  assign n1870 = n544 & ~n684;
  assign n1871 = ~n1484 & ~n1870;
  assign n1872 = ~n1869 & n1871;
  assign n1836 = n1101 ^ n1097;
  assign n1863 = n1150 ^ n1101;
  assign n1864 = ~n1836 & n1863;
  assign n1865 = n1864 ^ n1101;
  assign n1866 = ~n506 & ~n1865;
  assign n1873 = n1872 ^ n1866;
  assign n1852 = ~n1225 & n1790;
  assign n1853 = n633 ^ n551;
  assign n1854 = n836 & n1853;
  assign n1855 = ~n1852 & ~n1854;
  assign n1847 = n521 & n851;
  assign n1848 = n1847 ^ n732;
  assign n1849 = ~n536 & n1848;
  assign n1850 = ~n506 & ~n732;
  assign n1851 = ~n1849 & ~n1850;
  assign n1856 = n1855 ^ n1851;
  assign n1857 = ~n724 & ~n1804;
  assign n1858 = n694 & ~n734;
  assign n1859 = ~n1857 & ~n1858;
  assign n1860 = n1859 ^ n1855;
  assign n1861 = ~n1856 & n1860;
  assign n1862 = n1861 ^ n1859;
  assign n1874 = n1873 ^ n1862;
  assign n1846 = n842 ^ n738;
  assign n1875 = n1874 ^ n1846;
  assign n1837 = ~n506 & ~n1836;
  assign n1838 = n1837 ^ n1150;
  assign n1832 = n1792 ^ n1787;
  assign n1833 = n1792 ^ n1786;
  assign n1834 = n1832 & ~n1833;
  assign n1835 = n1834 ^ n1787;
  assign n1839 = n1838 ^ n1835;
  assign n1840 = n1806 ^ n1801;
  assign n1841 = ~n1802 & ~n1840;
  assign n1842 = n1841 ^ n1806;
  assign n1843 = n1842 ^ n1835;
  assign n1844 = ~n1839 & n1843;
  assign n1845 = n1844 ^ n1842;
  assign n1876 = n1875 ^ n1845;
  assign n1877 = n1842 ^ n1839;
  assign n1878 = n1817 ^ n1777;
  assign n1879 = ~n1818 & n1878;
  assign n1880 = n1879 ^ n1777;
  assign n1881 = ~n1877 & ~n1880;
  assign n1882 = n1876 & ~n1881;
  assign n1883 = n1831 & ~n1882;
  assign n1884 = n1859 ^ n1856;
  assign n1885 = n1793 ^ n1780;
  assign n1886 = n1808 & ~n1885;
  assign n1887 = n1886 ^ n1807;
  assign n1888 = ~n1884 & ~n1887;
  assign n1889 = n1877 & n1880;
  assign n1890 = ~n1876 & ~n1889;
  assign n1891 = ~n1888 & ~n1890;
  assign n1892 = ~n1883 & n1891;
  assign n1893 = n1884 & n1887;
  assign n1894 = n1893 ^ n1876;
  assign n1895 = n1881 ^ n1876;
  assign n1896 = n1895 ^ n1876;
  assign n1897 = n1831 & ~n1889;
  assign n1898 = n1897 ^ n1876;
  assign n1899 = n1898 ^ n1876;
  assign n1900 = ~n1896 & ~n1899;
  assign n1901 = n1900 ^ n1876;
  assign n1902 = n1894 & ~n1901;
  assign n1903 = n1902 ^ n1893;
  assign n1904 = ~n1892 & ~n1903;
  assign n1905 = ~n506 & n851;
  assign n1906 = n1905 ^ n853;
  assign n1907 = n845 ^ n730;
  assign n1908 = n1866 ^ n1862;
  assign n1909 = ~n1873 & ~n1908;
  assign n1910 = n1909 ^ n1862;
  assign n1911 = n1907 & n1910;
  assign n1912 = n1906 & n1911;
  assign n1913 = n1874 ^ n1845;
  assign n1914 = ~n1875 & n1913;
  assign n1915 = n1914 ^ n1845;
  assign n1916 = ~n1912 & ~n1915;
  assign n1917 = n1910 ^ n1907;
  assign n1918 = n1910 ^ n1906;
  assign n1919 = n1917 & ~n1918;
  assign n1920 = n1919 ^ n1907;
  assign n1921 = ~n1916 & n1920;
  assign n1922 = ~n1907 & ~n1910;
  assign n1923 = ~n1906 & n1922;
  assign n1924 = ~n1915 & n1923;
  assign n1925 = n861 & ~n1924;
  assign n1926 = ~n1921 & ~n1925;
  assign n1927 = ~n1904 & ~n1926;
  assign n1928 = n1915 & ~n1923;
  assign n1929 = ~n1920 & ~n1928;
  assign n1930 = n1912 & n1915;
  assign n1931 = ~n861 & ~n1930;
  assign n1932 = ~n1929 & ~n1931;
  assign n1933 = ~n1927 & ~n1932;
  assign n1934 = n1933 ^ n872;
  assign n1935 = ~n873 & ~n1934;
  assign n1936 = n1935 ^ n1933;
  assign n1945 = n1944 ^ n1936;
  assign n412 = ~n174 & ~n411;
  assign n413 = ~n147 & ~n412;
  assign n415 = ~n413 & ~n414;
  assign n416 = ~n410 & n415;
  assign n417 = n409 & n416;
  assign n422 = n387 & n421;
  assign n426 = ~n263 & ~n425;
  assign n427 = n422 & n426;
  assign n428 = n417 & n427;
  assign n433 = ~n431 & ~n432;
  assign n434 = n430 & n433;
  assign n435 = ~n330 & ~n396;
  assign n436 = n434 & n435;
  assign n437 = n428 & n436;
  assign n439 = ~n375 & ~n438;
  assign n440 = ~n283 & n439;
  assign n441 = ~n323 & ~n351;
  assign n442 = ~n222 & n441;
  assign n443 = n440 & n442;
  assign n444 = n219 & n443;
  assign n445 = n437 & n444;
  assign n448 = ~n255 & ~n447;
  assign n449 = n78 & n150;
  assign n450 = n51 & ~n449;
  assign n451 = n391 & ~n450;
  assign n452 = n448 & n451;
  assign n455 = ~n348 & ~n454;
  assign n456 = n453 & n455;
  assign n457 = n452 & n456;
  assign n466 = n193 & ~n303;
  assign n472 = n85 & ~n471;
  assign n473 = ~n470 & ~n472;
  assign n474 = n469 & n473;
  assign n475 = n466 & n474;
  assign n476 = n465 & n475;
  assign n477 = n457 & n476;
  assign n478 = n445 & n477;
  assign n1946 = n1945 ^ n478;
  assign n2285 = n1933 ^ n873;
  assign n1985 = ~n1924 & ~n1930;
  assign n1986 = n1929 ^ n1921;
  assign n1987 = ~n1904 & n1986;
  assign n1988 = n1987 ^ n1929;
  assign n1989 = n1985 & ~n1988;
  assign n1990 = n1989 ^ n861;
  assign n1947 = ~n85 & n221;
  assign n1948 = ~n78 & ~n1947;
  assign n1949 = n434 & ~n1948;
  assign n1950 = n57 & ~n169;
  assign n1951 = n473 & ~n1950;
  assign n1952 = n139 & ~n159;
  assign n1953 = n1951 & ~n1952;
  assign n1954 = n560 & n1953;
  assign n1955 = n1949 & n1954;
  assign n1956 = ~n274 & ~n375;
  assign n1957 = n270 & n1956;
  assign n1958 = n1045 & n1957;
  assign n1959 = n1955 & n1958;
  assign n1960 = ~n356 & ~n786;
  assign n1961 = ~n938 & n1960;
  assign n1962 = ~n396 & ~n468;
  assign n1963 = n48 & n446;
  assign n1964 = n1962 & ~n1963;
  assign n1965 = ~n583 & ~n1026;
  assign n1966 = n1964 & n1965;
  assign n1967 = n1961 & n1966;
  assign n1968 = n102 & ~n522;
  assign n1969 = n671 & ~n1968;
  assign n1970 = n1967 & n1969;
  assign n1971 = n575 & n1970;
  assign n1972 = n567 & ~n767;
  assign n1973 = ~n210 & ~n487;
  assign n1974 = n1972 & n1973;
  assign n1975 = n565 & n1974;
  assign n1981 = ~n651 & n1980;
  assign n1982 = n1975 & n1981;
  assign n1983 = n1971 & n1982;
  assign n1984 = n1959 & n1983;
  assign n1991 = n1990 ^ n1984;
  assign n2023 = n1917 ^ n1906;
  assign n2024 = n2023 ^ n1915;
  assign n2025 = n2024 ^ n1904;
  assign n1992 = n102 & ~n181;
  assign n1993 = ~n192 & ~n1992;
  assign n1994 = n1959 & n1993;
  assign n302 = ~n296 & n301;
  assign n1995 = n56 & ~n125;
  assign n1996 = ~n620 & ~n1995;
  assign n1997 = n927 & n1996;
  assign n1998 = n302 & n1997;
  assign n1999 = ~n252 & ~n395;
  assign n2000 = ~n57 & n1999;
  assign n2001 = ~n498 & ~n2000;
  assign n2002 = ~n810 & ~n2001;
  assign n2003 = n1998 & n2002;
  assign n2004 = ~n50 & ~n809;
  assign n2005 = n614 & ~n2004;
  assign n2006 = ~n48 & ~n231;
  assign n2007 = ~n2005 & ~n2006;
  assign n2008 = ~n363 & ~n2007;
  assign n2009 = n101 & ~n168;
  assign n2010 = n175 ^ n120;
  assign n2011 = n175 ^ n139;
  assign n2012 = n2011 ^ n139;
  assign n2013 = n922 ^ n139;
  assign n2014 = n2012 & n2013;
  assign n2015 = n2014 ^ n139;
  assign n2016 = n2010 & ~n2015;
  assign n2017 = n2016 ^ n120;
  assign n2018 = ~n2009 & ~n2017;
  assign n2019 = n2008 & n2018;
  assign n2020 = n457 & n2019;
  assign n2021 = n2003 & n2020;
  assign n2022 = n1994 & n2021;
  assign n2026 = n2025 ^ n2022;
  assign n241 = ~n237 & n240;
  assign n242 = n233 & n241;
  assign n256 = ~n254 & ~n255;
  assign n257 = ~n252 & n256;
  assign n258 = n251 & n257;
  assign n259 = n242 & n258;
  assign n260 = ~n225 & n259;
  assign n2047 = ~n162 & ~n328;
  assign n2048 = ~n180 & ~n2047;
  assign n2049 = ~n150 & n411;
  assign n2050 = ~n2048 & ~n2049;
  assign n2051 = ~n767 & n2050;
  assign n2052 = ~n284 & ~n325;
  assign n2053 = ~n625 & n2052;
  assign n2054 = n2051 & n2053;
  assign n2055 = ~n92 & ~n375;
  assign n2056 = ~n675 & n2055;
  assign n2057 = ~n120 & n249;
  assign n2058 = ~n175 & n2057;
  assign n2059 = ~n652 & ~n2058;
  assign n2060 = ~n344 & ~n656;
  assign n2061 = ~n786 & n2060;
  assign n2062 = ~n330 & n2061;
  assign n2063 = ~n2059 & n2062;
  assign n2064 = n2056 & n2063;
  assign n2065 = n2054 & n2064;
  assign n2066 = ~n79 & n963;
  assign n2067 = ~n438 & ~n2066;
  assign n2068 = ~n388 & n2067;
  assign n2069 = n2065 & n2068;
  assign n2070 = n1036 & n2069;
  assign n2071 = n260 & n2070;
  assign n2027 = n1880 ^ n1877;
  assign n2028 = n1877 & n1893;
  assign n2029 = ~n1877 & n1888;
  assign n2030 = ~n2028 & ~n2029;
  assign n2031 = ~n2027 & ~n2030;
  assign n2032 = ~n1880 & ~n2028;
  assign n2033 = n1887 ^ n1884;
  assign n2034 = n1887 ^ n1877;
  assign n2035 = ~n2033 & n2034;
  assign n2036 = n2035 ^ n1877;
  assign n2037 = ~n2032 & n2036;
  assign n2038 = n2037 ^ n1831;
  assign n2039 = n2038 ^ n2037;
  assign n2040 = ~n1880 & ~n2036;
  assign n2041 = ~n2029 & ~n2040;
  assign n2042 = n2041 ^ n2037;
  assign n2043 = n2039 & ~n2042;
  assign n2044 = n2043 ^ n2037;
  assign n2045 = ~n2031 & ~n2044;
  assign n2046 = n2045 ^ n1876;
  assign n2072 = n2071 ^ n2046;
  assign n2089 = n2033 ^ n2027;
  assign n2090 = n2089 ^ n1831;
  assign n2077 = ~n221 & ~n2076;
  assign n2078 = n2074 & ~n2077;
  assign n2079 = n996 & n2078;
  assign n2080 = n361 & n2079;
  assign n2081 = n175 & ~n498;
  assign n2082 = ~n566 & ~n2081;
  assign n2083 = n940 & n2082;
  assign n2084 = n1009 & n2083;
  assign n2085 = n1117 & n2084;
  assign n2086 = n2080 & n2085;
  assign n2087 = n143 & n1116;
  assign n2088 = n2086 & n2087;
  assign n2091 = n2090 ^ n2088;
  assign n2130 = n1750 ^ n1727;
  assign n2132 = ~n1823 & ~n1825;
  assign n2131 = n1773 ^ n1750;
  assign n2133 = n2132 ^ n2131;
  assign n2134 = ~n2130 & ~n2133;
  assign n2135 = n2134 ^ n2132;
  assign n2136 = n2135 ^ n1819;
  assign n2105 = ~n190 & ~n272;
  assign n2106 = ~n92 & ~n296;
  assign n2107 = n2105 & n2106;
  assign n2111 = ~n643 & n2110;
  assign n2112 = n2107 & n2111;
  assign n2113 = ~n330 & ~n606;
  assign n2114 = ~n396 & n2113;
  assign n2115 = n2112 & n2114;
  assign n2116 = n1034 & n2115;
  assign n2117 = ~n282 & ~n822;
  assign n2118 = ~n268 & n2117;
  assign n2119 = ~n324 & ~n938;
  assign n2120 = n2118 & n2119;
  assign n2121 = ~n69 & n139;
  assign n2122 = ~n254 & ~n2121;
  assign n2123 = n2120 & n2122;
  assign n2124 = ~n562 & ~n939;
  assign n2125 = ~n206 & n2124;
  assign n2126 = n785 & n2125;
  assign n2127 = n2123 & n2126;
  assign n2128 = n2116 & n2127;
  assign n2129 = n2104 & n2128;
  assign n2137 = n2136 ^ n2129;
  assign n2166 = n1770 ^ n1767;
  assign n2167 = n2166 ^ n2130;
  assign n2138 = n175 & ~n493;
  assign n2139 = ~n299 & ~n2138;
  assign n2140 = ~n613 & n2139;
  assign n2141 = n346 & n2140;
  assign n2142 = n391 & n888;
  assign n2143 = n1961 & n2142;
  assign n2144 = n2141 & n2143;
  assign n2145 = n757 & n2114;
  assign n2146 = ~n1029 & ~n2047;
  assign n2147 = ~n468 & ~n2146;
  assign n2148 = n2145 & n2147;
  assign n2149 = ~n175 & n406;
  assign n2150 = ~n83 & n147;
  assign n2151 = ~n2149 & ~n2150;
  assign n2152 = ~n915 & ~n2151;
  assign n2153 = n139 & ~n875;
  assign n2154 = n57 & ~n1007;
  assign n2155 = ~n2153 & ~n2154;
  assign n2156 = ~n323 & n2155;
  assign n2157 = n2152 & n2156;
  assign n2158 = n120 & n963;
  assign n2159 = ~n656 & ~n2158;
  assign n2160 = ~n207 & n2159;
  assign n2161 = n421 & n2160;
  assign n2162 = n2157 & n2161;
  assign n2163 = n2148 & n2162;
  assign n2164 = n2144 & n2163;
  assign n2165 = n834 & n2164;
  assign n2168 = n2167 ^ n2165;
  assign n2201 = n1604 ^ n1601;
  assign n2233 = n1662 ^ n1604;
  assign n2234 = n2233 ^ n1721;
  assign n2235 = ~n2201 & n2234;
  assign n2236 = n2235 ^ n1721;
  assign n2237 = n2236 ^ n1714;
  assign n2200 = n1659 ^ n1656;
  assign n2202 = n2201 ^ n2200;
  assign n2169 = n174 & ~n180;
  assign n2170 = n1962 & ~n2169;
  assign n2171 = n448 & n2170;
  assign n2172 = ~n432 & ~n620;
  assign n2173 = n83 & ~n214;
  assign n2174 = ~n377 & ~n2173;
  assign n2175 = n2172 & n2174;
  assign n2176 = ~n56 & n156;
  assign n2177 = ~n50 & n125;
  assign n2178 = ~n48 & n2177;
  assign n2179 = ~n2176 & ~n2178;
  assign n2180 = n50 & n91;
  assign n2181 = n2179 & ~n2180;
  assign n2182 = n101 & ~n150;
  assign n2183 = ~n2181 & ~n2182;
  assign n2184 = n2175 & n2183;
  assign n2185 = n2171 & n2184;
  assign n2187 = ~n786 & ~n822;
  assign n2188 = ~n981 & n2187;
  assign n2189 = n2186 & n2188;
  assign n2190 = ~n198 & ~n250;
  assign n2191 = n2113 & n2190;
  assign n2192 = n2189 & n2191;
  assign n2193 = ~n767 & ~n2121;
  assign n2194 = n57 & ~n510;
  assign n2195 = n2193 & ~n2194;
  assign n2196 = n774 & n2195;
  assign n2197 = n2192 & n2196;
  assign n2198 = n2185 & n2197;
  assign n2199 = n361 & n2198;
  assign n2203 = n2202 ^ n2199;
  assign n2204 = ~n1483 & n1583;
  assign n2205 = n1483 & n1513;
  assign n2206 = n1588 ^ n1585;
  assign n2207 = ~n2205 & ~n2206;
  assign n2208 = ~n2204 & n2207;
  assign n2209 = n1597 ^ n1592;
  assign n2210 = n2209 ^ n1592;
  assign n2211 = n1592 ^ n1589;
  assign n2212 = ~n2210 & n2211;
  assign n2213 = n2212 ^ n1592;
  assign n2214 = ~n2208 & ~n2213;
  assign n2215 = n2214 ^ n1580;
  assign n2216 = ~n58 & ~n897;
  assign n2217 = n101 & ~n156;
  assign n2218 = n56 & ~n211;
  assign n2219 = ~n2217 & ~n2218;
  assign n2220 = ~n363 & n2219;
  assign n2221 = n804 & n2220;
  assign n2222 = n275 & n908;
  assign n2223 = n2221 & n2222;
  assign n2224 = n833 & n1020;
  assign n2225 = n2223 & n2224;
  assign n2226 = n2144 & n2225;
  assign n2227 = n437 & n2226;
  assign n2228 = ~n2216 & n2227;
  assign n2229 = n2215 & n2228;
  assign n2230 = n2229 ^ n2199;
  assign n2231 = ~n2203 & ~n2230;
  assign n2232 = n2231 ^ n2202;
  assign n2238 = n2237 ^ n2232;
  assign n2239 = ~n363 & n634;
  assign n2240 = ~n138 & ~n341;
  assign n2241 = ~n250 & ~n812;
  assign n2242 = n2240 & n2241;
  assign n2243 = n2239 & n2242;
  assign n292 = ~n290 & ~n291;
  assign n2244 = n292 & n901;
  assign n2245 = n2243 & n2244;
  assign n2246 = n2157 & n2245;
  assign n2249 = n591 & n2248;
  assign n2250 = n2246 & n2249;
  assign n2251 = n1999 & n2113;
  assign n2252 = ~n243 & ~n296;
  assign n2253 = ~n1132 & n2252;
  assign n2254 = n980 & n2253;
  assign n2255 = n2251 & n2254;
  assign n2256 = ~n352 & ~n935;
  assign n2258 = ~n1040 & n2257;
  assign n2259 = n2256 & n2258;
  assign n2260 = n2255 & n2259;
  assign n2261 = n2079 & n2097;
  assign n2262 = n2260 & n2261;
  assign n2263 = n2250 & n2262;
  assign n2264 = n2263 ^ n2232;
  assign n2265 = n2238 & n2264;
  assign n2266 = n2265 ^ n2237;
  assign n2267 = n2266 ^ n2167;
  assign n2268 = ~n2168 & ~n2267;
  assign n2269 = n2268 ^ n2266;
  assign n2270 = n2269 ^ n2129;
  assign n2271 = ~n2137 & n2270;
  assign n2272 = n2271 ^ n2136;
  assign n2273 = n2272 ^ n2090;
  assign n2274 = ~n2091 & ~n2273;
  assign n2275 = n2274 ^ n2272;
  assign n2276 = n2275 ^ n2046;
  assign n2277 = n2072 & n2276;
  assign n2278 = n2277 ^ n2275;
  assign n2279 = n2278 ^ n2025;
  assign n2280 = ~n2026 & ~n2279;
  assign n2281 = n2280 ^ n2278;
  assign n2282 = n2281 ^ n1990;
  assign n2283 = n1991 & n2282;
  assign n2284 = n2283 ^ n2281;
  assign n2286 = n2285 ^ n2284;
  assign n2287 = ~n296 & ~n303;
  assign n2288 = ~n524 & n2287;
  assign n2289 = ~n226 & n1027;
  assign n2290 = n2288 & n2289;
  assign n2291 = n120 & ~n977;
  assign n2292 = ~n627 & ~n822;
  assign n2293 = ~n2291 & n2292;
  assign n2294 = n270 & n2293;
  assign n2295 = n2290 & n2294;
  assign n2296 = n580 & n764;
  assign n2297 = n831 & n2296;
  assign n2298 = n659 & n2297;
  assign n2299 = n2295 & n2298;
  assign n2300 = n911 & n2299;
  assign n2301 = ~n620 & n1145;
  assign n2302 = n2300 & n2301;
  assign n2303 = n2302 ^ n2285;
  assign n2304 = ~n2286 & ~n2303;
  assign n2305 = n2304 ^ n2284;
  assign n2306 = n2305 ^ n1945;
  assign n2307 = ~n1946 & ~n2306;
  assign n2308 = n2307 ^ n2305;
  assign n2325 = n2324 ^ n2308;
  assign n2326 = n543 & n1938;
  assign n2327 = ~n551 & ~n2326;
  assign n2328 = ~n506 & n2327;
  assign n2329 = ~n1937 & ~n2328;
  assign n2330 = n1943 & ~n2329;
  assign n2331 = n521 & ~n551;
  assign n2332 = ~n543 & ~n1938;
  assign n2333 = ~n506 & n2332;
  assign n2334 = n2331 & n2333;
  assign n2335 = ~n2330 & ~n2334;
  assign n2336 = n1936 & ~n2335;
  assign n2337 = n2336 ^ n2324;
  assign n2338 = ~n2325 & ~n2337;
  assign n2339 = n2338 ^ n2308;
  assign n2340 = n405 & ~n2339;
  assign n304 = n137 & ~n175;
  assign n305 = n78 & ~n139;
  assign n306 = ~n304 & ~n305;
  assign n307 = ~n303 & ~n306;
  assign n310 = ~n308 & ~n309;
  assign n311 = n307 & n310;
  assign n2341 = n435 & ~n583;
  assign n2342 = n936 & n2172;
  assign n2343 = n2341 & n2342;
  assign n2344 = ~n299 & ~n454;
  assign n2345 = ~n487 & n2344;
  assign n2346 = n2343 & n2345;
  assign n2347 = n311 & n2346;
  assign n2348 = n794 & n2347;
  assign n2349 = ~n121 & ~n1040;
  assign n2350 = ~n269 & n2349;
  assign n2351 = ~n207 & ~n244;
  assign n2352 = ~n252 & n2060;
  assign n2353 = n2351 & n2352;
  assign n2354 = n2350 & n2353;
  assign n2355 = n137 & n249;
  assign n2356 = ~n881 & ~n2355;
  assign n2357 = n2354 & ~n2356;
  assign n2358 = ~n393 & ~n563;
  assign n2359 = n57 & ~n875;
  assign n2360 = ~n92 & ~n2359;
  assign n2361 = n2358 & n2360;
  assign n2362 = n474 & n2361;
  assign n2363 = n2357 & n2362;
  assign n2364 = n826 & n2363;
  assign n2365 = n2348 & n2364;
  assign n2366 = n2340 & n2365;
  assign n2420 = n2384 ^ n2366;
  assign n317 = x22 ^ x2;
  assign n3265 = n2420 ^ n317;
  assign n3266 = x1 & n3265;
  assign n318 = ~x1 & x2;
  assign n3235 = n2365 ^ n2340;
  assign n3267 = n318 & n3235;
  assign n3268 = ~x0 & ~n3267;
  assign n3269 = ~n3266 & n3268;
  assign n2386 = n91 & n369;
  assign n2387 = n48 & ~n2386;
  assign n2388 = n528 & ~n2387;
  assign n2389 = n97 & n406;
  assign n2390 = ~n56 & ~n175;
  assign n2391 = ~n2389 & ~n2390;
  assign n2392 = ~n585 & ~n813;
  assign n2393 = ~n2391 & n2392;
  assign n2394 = n51 & ~n514;
  assign n2395 = ~n351 & ~n2394;
  assign n2396 = n940 & n2395;
  assign n2397 = n2393 & n2396;
  assign n2398 = n519 & n2397;
  assign n2399 = n492 & n2398;
  assign n2400 = n2388 & n2399;
  assign n2385 = n2366 & n2384;
  assign n2417 = n2400 ^ n2385;
  assign n3273 = n2417 ^ x22;
  assign n320 = x2 ^ x1;
  assign n2434 = n2305 ^ n1946;
  assign n2435 = n2286 & n2302;
  assign n2436 = n2284 & ~n2285;
  assign n2437 = ~n1946 & ~n2436;
  assign n2438 = ~n2435 & ~n2437;
  assign n2439 = n2281 ^ n1991;
  assign n2440 = n2278 ^ n2026;
  assign n2441 = n2275 ^ n2072;
  assign n2442 = n2272 ^ n2091;
  assign n2443 = n2269 ^ n2137;
  assign n2444 = n2266 ^ n2168;
  assign n2445 = n2263 ^ n2237;
  assign n2446 = n2445 ^ n2232;
  assign n2447 = n2229 ^ n2203;
  assign n2448 = ~n2446 & n2447;
  assign n2449 = ~n2444 & ~n2448;
  assign n2450 = ~n2443 & ~n2449;
  assign n2451 = ~n2442 & ~n2450;
  assign n2452 = ~n2441 & ~n2451;
  assign n2453 = ~n2440 & ~n2452;
  assign n2454 = ~n2439 & ~n2453;
  assign n2455 = ~n2438 & ~n2454;
  assign n2456 = n2434 & ~n2455;
  assign n2457 = n2329 & ~n2333;
  assign n2458 = n2457 ^ n1936;
  assign n2459 = n1944 & n2458;
  assign n2460 = n2459 ^ n2336;
  assign n2461 = n2325 & ~n2460;
  assign n2462 = n2461 ^ n2336;
  assign n2463 = ~n2456 & ~n2462;
  assign n2464 = ~n405 & n2339;
  assign n2465 = ~n2463 & n2464;
  assign n2466 = n2365 & ~n2465;
  assign n2467 = n2340 & n2463;
  assign n2468 = ~n2384 & ~n2467;
  assign n2469 = ~n2466 & n2468;
  assign n2472 = ~n2340 & ~n2365;
  assign n2488 = ~n2308 & n2324;
  assign n2489 = n2459 & n2488;
  assign n2473 = n2302 ^ n2286;
  assign n2474 = n2228 ^ n2215;
  assign n2475 = n2447 & ~n2474;
  assign n2476 = n2446 & ~n2475;
  assign n2477 = n2444 & ~n2476;
  assign n2478 = n2443 & ~n2477;
  assign n2479 = n2442 & ~n2478;
  assign n2480 = n2441 & ~n2479;
  assign n2481 = n2440 & ~n2480;
  assign n2482 = n2439 & ~n2481;
  assign n2483 = n2473 & ~n2482;
  assign n2484 = ~n2434 & ~n2483;
  assign n2490 = ~n2339 & n2484;
  assign n2491 = ~n2489 & ~n2490;
  assign n2485 = n2308 & ~n2324;
  assign n2486 = ~n2459 & n2485;
  assign n2487 = ~n2484 & n2486;
  assign n2492 = n2491 ^ n2487;
  assign n2493 = n2492 ^ n2491;
  assign n2494 = n2491 ^ n2339;
  assign n2495 = n2494 ^ n2491;
  assign n2496 = ~n2493 & n2495;
  assign n2497 = n2496 ^ n2491;
  assign n2498 = n405 & ~n2497;
  assign n2499 = n2498 ^ n2491;
  assign n2500 = n2472 & n2499;
  assign n2501 = n2384 & ~n2500;
  assign n3270 = ~n2469 & ~n2501;
  assign n3271 = n320 & ~n3270;
  assign n3272 = n3271 ^ x1;
  assign n3274 = n3273 ^ n3272;
  assign n3275 = x0 & ~n3274;
  assign n3276 = ~n3269 & ~n3275;
  assign n3019 = n1056 & ~n1157;
  assign n3154 = n1157 & n2462;
  assign n3155 = ~n3019 & ~n3154;
  assign n319 = n317 & ~n318;
  assign n2428 = ~n26 & ~n319;
  assign n2509 = x0 & ~x22;
  assign n2510 = x2 & n2509;
  assign n2511 = n2428 & ~n2510;
  assign n2821 = ~n1152 & ~n2511;
  assign n2830 = ~n1157 & n2821;
  assign n3156 = ~n2434 & n2830;
  assign n3157 = n3156 ^ n2821;
  assign n3158 = ~n3155 & n3157;
  assign n2819 = n1152 & n2511;
  assign n2820 = ~n1157 & n2819;
  assign n3159 = n2462 & n2820;
  assign n2831 = ~n1056 & n1157;
  assign n2832 = n2819 & n2831;
  assign n3160 = n2434 & n2832;
  assign n3161 = ~n3159 & ~n3160;
  assign n3162 = ~n3158 & n3161;
  assign n3163 = n1056 & ~n3162;
  assign n2846 = ~n2456 & ~n2484;
  assign n3164 = n2462 ^ n2434;
  assign n3165 = ~n2846 & n3164;
  assign n2845 = n2511 ^ n1152;
  assign n3166 = n2339 ^ n405;
  assign n3167 = n3166 ^ n1157;
  assign n3168 = n2845 & ~n3167;
  assign n3169 = n3165 & n3168;
  assign n3170 = ~n3163 & ~n3169;
  assign n2895 = n1056 & n2845;
  assign n3171 = ~n3165 & n3166;
  assign n3172 = n2895 & n3171;
  assign n3173 = n3170 & ~n3172;
  assign n3174 = ~n1056 & n3162;
  assign n3175 = ~n3165 & ~n3166;
  assign n3176 = n2845 & ~n3175;
  assign n3177 = n3174 & ~n3176;
  assign n3178 = n3173 & ~n3177;
  assign n2598 = n1061 ^ n1056;
  assign n2893 = ~n2454 & ~n2482;
  assign n2894 = n2473 & ~n2893;
  assign n3137 = n2598 & n2894;
  assign n2603 = n1056 & n1061;
  assign n2602 = ~n1056 & ~n1061;
  assign n2604 = n2603 ^ n2602;
  assign n2605 = ~n1101 & n2604;
  assign n2606 = n2605 ^ n2603;
  assign n3138 = ~n2439 & n2606;
  assign n2608 = n1101 & n2604;
  assign n2609 = n2608 ^ n2603;
  assign n2610 = ~n1836 & n2609;
  assign n3139 = n2440 & n2610;
  assign n3140 = ~n3138 & ~n3139;
  assign n3141 = ~n3137 & n3140;
  assign n3142 = n1097 & ~n3141;
  assign n2910 = ~n2473 & ~n2893;
  assign n3143 = n2598 & ~n2910;
  assign n3144 = ~n1097 & n3140;
  assign n3145 = ~n3143 & n3144;
  assign n3146 = n2473 ^ n1101;
  assign n3147 = n2598 & n2893;
  assign n3148 = n3146 & n3147;
  assign n3149 = ~n3145 & ~n3148;
  assign n3150 = ~n3142 & n3149;
  assign n2522 = n1097 ^ n732;
  assign n2632 = ~n2451 & ~n2479;
  assign n3115 = n2522 & n2632;
  assign n3116 = n2441 ^ n850;
  assign n3117 = n3115 & n3116;
  assign n2524 = n732 & n1097;
  assign n2525 = ~n850 & ~n2524;
  assign n2526 = ~n732 & ~n1097;
  assign n2527 = n850 & ~n2526;
  assign n2528 = ~n2525 & ~n2527;
  assign n3118 = n2442 & n2528;
  assign n2519 = n850 ^ n684;
  assign n2530 = n2526 ^ n2524;
  assign n2531 = n2524 ^ n850;
  assign n2532 = n2531 ^ n2524;
  assign n2533 = n2530 & ~n2532;
  assign n2534 = n2533 ^ n2524;
  assign n2535 = n2519 & n2534;
  assign n3119 = ~n2443 & n2535;
  assign n3120 = ~n3118 & ~n3119;
  assign n3121 = n3120 ^ n684;
  assign n2640 = n2441 & ~n2632;
  assign n3122 = n2522 & ~n2640;
  assign n3123 = n3122 ^ n684;
  assign n2633 = ~n2441 & ~n2632;
  assign n2777 = n684 & n2522;
  assign n3124 = n2633 & n2777;
  assign n3125 = n3124 ^ n684;
  assign n3126 = ~n684 & n3125;
  assign n3127 = n3126 ^ n684;
  assign n3128 = ~n3123 & ~n3127;
  assign n3129 = n3128 ^ n3126;
  assign n3130 = n3129 ^ n684;
  assign n3131 = n3130 ^ n3124;
  assign n3132 = n3121 & n3131;
  assign n3133 = n3132 ^ n3124;
  assign n3134 = ~n3117 & ~n3133;
  assign n2569 = n538 & n684;
  assign n2751 = n543 & ~n2474;
  assign n2752 = n2569 & ~n2751;
  assign n2539 = ~n2203 & n2474;
  assign n2572 = ~n543 & ~n2474;
  assign n2753 = ~n551 & n1938;
  assign n2754 = ~n2572 & n2753;
  assign n2755 = ~n2539 & ~n2754;
  assign n2756 = ~n2752 & n2755;
  assign n2518 = n2203 & n2474;
  assign n2758 = n552 & n2518;
  assign n2759 = n2758 ^ n2446;
  assign n2760 = n685 & ~n2759;
  assign n2761 = n543 & n2569;
  assign n2762 = ~n543 & n1938;
  assign n2763 = ~n2761 & ~n2762;
  assign n2764 = n2447 & ~n2763;
  assign n2765 = n551 & n2569;
  assign n2766 = ~n2753 & ~n2765;
  assign n2767 = n552 & ~n2766;
  assign n2768 = ~n2474 & n2767;
  assign n2769 = ~n2764 & ~n2768;
  assign n2770 = ~n2760 & n2769;
  assign n3088 = ~n2756 & n2770;
  assign n3089 = n3088 ^ n2474;
  assign n3090 = n3088 ^ n551;
  assign n3091 = n3090 ^ n551;
  assign n2553 = ~n2448 & ~n2476;
  assign n3092 = n552 & n2553;
  assign n3093 = n3092 ^ n2444;
  assign n3094 = n685 & ~n3093;
  assign n3098 = n543 & ~n551;
  assign n3099 = n2447 & n3098;
  assign n3100 = n1938 & ~n3099;
  assign n3095 = ~n543 & n551;
  assign n3096 = n2447 & n3095;
  assign n3097 = n2569 & ~n3096;
  assign n3101 = n3100 ^ n3097;
  assign n3102 = n2446 ^ n543;
  assign n3103 = n3102 ^ n543;
  assign n3104 = n3097 ^ n543;
  assign n3105 = n3103 & ~n3104;
  assign n3106 = n3105 ^ n543;
  assign n3107 = n3101 & ~n3106;
  assign n3108 = n3107 ^ n3100;
  assign n3109 = ~n3094 & ~n3108;
  assign n3110 = n3109 ^ n551;
  assign n3111 = n3091 & n3110;
  assign n3112 = n3111 ^ n551;
  assign n3113 = n3089 & ~n3112;
  assign n3114 = n3113 ^ n3109;
  assign n3135 = n3134 ^ n3114;
  assign n2722 = ~n2450 & ~n2478;
  assign n2772 = ~n2443 & n2528;
  assign n2773 = n2444 & n2535;
  assign n2774 = ~n2772 & ~n2773;
  assign n2775 = ~n684 & n2774;
  assign n2776 = n2722 & n2775;
  assign n2778 = ~n2776 & ~n2777;
  assign n2779 = ~n850 & n2722;
  assign n2780 = n2442 & ~n2779;
  assign n2781 = ~n2778 & n2780;
  assign n2782 = n2774 ^ n684;
  assign n2730 = ~n2442 & ~n2722;
  assign n2783 = n2522 & ~n2730;
  assign n2784 = n2783 ^ n684;
  assign n2785 = ~n850 & n2522;
  assign n2786 = ~n2442 & n2785;
  assign n2787 = n2722 & n2786;
  assign n2788 = n2787 ^ n684;
  assign n2789 = ~n684 & n2788;
  assign n2790 = n2789 ^ n684;
  assign n2791 = ~n2784 & ~n2790;
  assign n2792 = n2791 ^ n2789;
  assign n2793 = n2792 ^ n684;
  assign n2794 = n2793 ^ n2787;
  assign n2795 = n2782 & n2794;
  assign n2796 = n2795 ^ n2787;
  assign n2797 = ~n2781 & ~n2796;
  assign n2757 = ~n551 & n2756;
  assign n2771 = n2770 ^ n2757;
  assign n2798 = n2797 ^ n2771;
  assign n2576 = ~n2449 & ~n2477;
  assign n2577 = ~n2443 & n2522;
  assign n2578 = ~n2576 & n2577;
  assign n2579 = n2444 & n2528;
  assign n2580 = ~n2446 & n2535;
  assign n2581 = ~n2579 & ~n2580;
  assign n2582 = ~n2578 & n2581;
  assign n2583 = ~n684 & ~n2582;
  assign n2584 = n2522 & n2576;
  assign n2585 = n2443 ^ n850;
  assign n2586 = n2585 ^ n2577;
  assign n2587 = n2586 ^ n2585;
  assign n2588 = n684 & n2581;
  assign n2589 = n2588 ^ n2585;
  assign n2590 = n2589 ^ n2585;
  assign n2591 = ~n2587 & n2590;
  assign n2592 = n2591 ^ n2585;
  assign n2593 = ~n2584 & ~n2592;
  assign n2594 = n2593 ^ n2585;
  assign n2595 = ~n2583 & n2594;
  assign n2568 = n685 & n2447;
  assign n2570 = n2569 ^ n543;
  assign n2571 = ~n2474 & ~n2570;
  assign n2573 = n2572 ^ n2571;
  assign n2574 = ~n2568 & ~n2573;
  assign n2575 = n2574 ^ n2572;
  assign n2596 = n2595 ^ n2575;
  assign n2517 = n685 & ~n2474;
  assign n2520 = n2518 & n2519;
  assign n2521 = n2520 ^ n2446;
  assign n2523 = ~n2521 & n2522;
  assign n2529 = n2447 & n2528;
  assign n2536 = ~n2474 & n2535;
  assign n2537 = ~n2529 & ~n2536;
  assign n2538 = ~n2523 & n2537;
  assign n2540 = ~n2474 & n2524;
  assign n2541 = ~n850 & n2540;
  assign n2542 = n2541 ^ n2524;
  assign n2543 = ~n2539 & ~n2542;
  assign n2544 = n850 & ~n2474;
  assign n2545 = n2526 & ~n2544;
  assign n2546 = n2543 & ~n2545;
  assign n2547 = n684 & ~n2546;
  assign n2548 = n2538 & n2547;
  assign n2549 = ~n2517 & ~n2548;
  assign n2550 = ~n2446 & n2528;
  assign n2551 = n2447 & n2535;
  assign n2552 = ~n2550 & ~n2551;
  assign n2554 = n850 & n2553;
  assign n2555 = n2554 ^ n2444;
  assign n2556 = n2522 & n2555;
  assign n2557 = n2556 ^ n684;
  assign n2558 = n2557 ^ n2556;
  assign n2559 = ~n850 & n2553;
  assign n2560 = n2559 ^ n2444;
  assign n2561 = n2522 & n2560;
  assign n2562 = n2561 ^ n2556;
  assign n2563 = n2558 & n2562;
  assign n2564 = n2563 ^ n2556;
  assign n2565 = n2552 & ~n2564;
  assign n2566 = n2565 ^ n684;
  assign n2567 = ~n2549 & ~n2566;
  assign n2748 = n2575 ^ n2567;
  assign n2749 = n2596 & n2748;
  assign n2750 = n2749 ^ n2595;
  assign n3085 = n2771 ^ n2750;
  assign n3086 = ~n2798 & ~n3085;
  assign n3087 = n3086 ^ n2797;
  assign n3136 = n3135 ^ n3087;
  assign n3151 = n3150 ^ n3136;
  assign n2800 = ~n2453 & ~n2481;
  assign n2801 = ~n2439 & ~n2800;
  assign n2802 = n2598 & n2801;
  assign n2803 = n2440 & n2606;
  assign n2804 = ~n2441 & n2610;
  assign n2805 = ~n2803 & ~n2804;
  assign n2806 = ~n2802 & n2805;
  assign n2807 = n1097 & ~n2806;
  assign n2808 = n2439 & ~n2800;
  assign n2809 = n2598 & ~n2808;
  assign n2810 = ~n1097 & n2805;
  assign n2811 = ~n2809 & n2810;
  assign n2812 = n2598 & n2800;
  assign n2813 = n2439 ^ n1101;
  assign n2814 = n2812 & ~n2813;
  assign n2815 = ~n2811 & ~n2814;
  assign n2816 = ~n2807 & n2815;
  assign n2799 = n2798 ^ n2750;
  assign n2817 = n2816 ^ n2799;
  assign n2599 = ~n2452 & ~n2480;
  assign n2600 = n2440 & ~n2599;
  assign n2601 = n2598 & n2600;
  assign n2607 = ~n2441 & n2606;
  assign n2611 = n2442 & n2610;
  assign n2612 = ~n2607 & ~n2611;
  assign n2613 = ~n2601 & n2612;
  assign n2614 = ~n1097 & ~n2613;
  assign n2615 = ~n2440 & ~n2599;
  assign n2616 = n2598 & ~n2615;
  assign n2617 = n1097 & n2612;
  assign n2618 = ~n2616 & n2617;
  assign n2619 = n2598 & n2599;
  assign n2620 = n2440 ^ n1101;
  assign n2621 = n2619 & ~n2620;
  assign n2622 = ~n2618 & ~n2621;
  assign n2623 = ~n2614 & n2622;
  assign n2597 = n2596 ^ n2567;
  assign n2624 = n2623 ^ n2597;
  assign n2634 = n2598 & n2633;
  assign n2635 = n2442 & n2606;
  assign n2636 = ~n2443 & n2610;
  assign n2637 = ~n2635 & ~n2636;
  assign n2638 = ~n2634 & n2637;
  assign n2639 = ~n1097 & ~n2638;
  assign n2641 = n2598 & ~n2640;
  assign n2642 = n1097 & n2637;
  assign n2643 = ~n2641 & n2642;
  assign n2644 = n2598 & n2632;
  assign n2645 = n2441 ^ n1101;
  assign n2646 = n2644 & n2645;
  assign n2647 = ~n2643 & ~n2646;
  assign n2648 = ~n2639 & n2647;
  assign n2628 = n2566 ^ n2517;
  assign n2625 = n684 & n2552;
  assign n2626 = ~n2561 & n2625;
  assign n2627 = ~n2517 & n2626;
  assign n2629 = n2628 ^ n2627;
  assign n2630 = n2548 & n2629;
  assign n2631 = n2630 ^ n2628;
  assign n2649 = n2648 ^ n2631;
  assign n2719 = n684 & n2546;
  assign n2720 = n2719 ^ n2538;
  assign n2659 = ~n1836 & n2518;
  assign n2660 = n2659 ^ n2446;
  assign n2661 = n2598 & ~n2660;
  assign n2662 = n2447 & n2606;
  assign n2663 = ~n2474 & n2610;
  assign n2664 = ~n2662 & ~n2663;
  assign n2665 = ~n2661 & n2664;
  assign n2666 = n2447 & n2598;
  assign n2667 = n2474 & ~n2666;
  assign n2668 = ~n2609 & ~n2667;
  assign n2669 = n1097 & ~n2668;
  assign n2670 = n2665 & n2669;
  assign n2671 = ~n2474 & n2522;
  assign n2672 = ~n2670 & ~n2671;
  assign n2673 = ~n2446 & n2606;
  assign n2674 = n2447 & n2610;
  assign n2675 = ~n2673 & ~n2674;
  assign n2676 = n2675 ^ n1097;
  assign n2677 = ~n2444 & ~n2553;
  assign n2678 = n2598 & ~n2677;
  assign n2679 = n2678 ^ n2675;
  assign n2680 = ~n1097 & ~n2553;
  assign n2681 = n2598 & ~n2680;
  assign n2682 = n1101 & n2553;
  assign n2683 = n2682 ^ n2444;
  assign n2684 = n2681 & n2683;
  assign n2685 = n2684 ^ n2675;
  assign n2686 = n2675 & ~n2685;
  assign n2687 = n2686 ^ n2675;
  assign n2688 = n2679 & n2687;
  assign n2689 = n2688 ^ n2686;
  assign n2690 = n2689 ^ n2675;
  assign n2691 = n2690 ^ n2684;
  assign n2692 = n2676 & ~n2691;
  assign n2693 = n2692 ^ n2684;
  assign n2694 = ~n2672 & ~n2693;
  assign n2650 = n2474 ^ n2447;
  assign n2651 = n2650 ^ n2447;
  assign n2652 = n2447 ^ n732;
  assign n2653 = n2652 ^ n2447;
  assign n2654 = ~n2651 & n2653;
  assign n2655 = n2654 ^ n2447;
  assign n2656 = ~n2522 & n2655;
  assign n2657 = n2656 ^ n2447;
  assign n2658 = n2657 ^ n2544;
  assign n2695 = n2694 ^ n2658;
  assign n2696 = n2576 ^ n2443;
  assign n2697 = ~n1101 & n2598;
  assign n2698 = ~n2696 & n2697;
  assign n2699 = n1097 & ~n1101;
  assign n2700 = n2444 & n2606;
  assign n2701 = ~n2446 & n2610;
  assign n2702 = ~n2700 & ~n2701;
  assign n2703 = ~n2699 & n2702;
  assign n2704 = n1101 & n2598;
  assign n2705 = ~n2443 & n2704;
  assign n2706 = n2703 & ~n2705;
  assign n2707 = ~n2698 & n2706;
  assign n2708 = n2443 & n2702;
  assign n2709 = n1097 & ~n2708;
  assign n2710 = ~n2707 & ~n2709;
  assign n2711 = n2598 & ~n2696;
  assign n2712 = n1097 & ~n2697;
  assign n2713 = n2702 & n2712;
  assign n2714 = ~n2711 & n2713;
  assign n2715 = ~n2710 & ~n2714;
  assign n2716 = n2715 ^ n2658;
  assign n2717 = n2695 & n2716;
  assign n2718 = n2717 ^ n2694;
  assign n2721 = n2720 ^ n2718;
  assign n2723 = n2442 & ~n2722;
  assign n2724 = n2598 & n2723;
  assign n2725 = ~n2443 & n2606;
  assign n2726 = n2444 & n2610;
  assign n2727 = ~n2725 & ~n2726;
  assign n2728 = ~n2724 & n2727;
  assign n2729 = n1097 & ~n2728;
  assign n2731 = n2598 & ~n2730;
  assign n2732 = ~n1097 & n2727;
  assign n2733 = ~n2731 & n2732;
  assign n2734 = n2598 & n2722;
  assign n2735 = n2442 ^ n1101;
  assign n2736 = n2734 & n2735;
  assign n2737 = ~n2733 & ~n2736;
  assign n2738 = ~n2729 & n2737;
  assign n2739 = n2738 ^ n2720;
  assign n2740 = n2721 & ~n2739;
  assign n2741 = n2740 ^ n2738;
  assign n2742 = n2741 ^ n2648;
  assign n2743 = ~n2649 & ~n2742;
  assign n2744 = n2743 ^ n2741;
  assign n2745 = n2744 ^ n2623;
  assign n2746 = n2624 & ~n2745;
  assign n2747 = n2746 ^ n2744;
  assign n3082 = n2799 ^ n2747;
  assign n3083 = n2817 & ~n3082;
  assign n3084 = n3083 ^ n2816;
  assign n3152 = n3151 ^ n3084;
  assign n2825 = ~n2820 & ~n2821;
  assign n2826 = ~n1056 & ~n2825;
  assign n2822 = n1157 & n2821;
  assign n2823 = ~n2820 & ~n2822;
  assign n2824 = n1056 & ~n2823;
  assign n2827 = n2826 ^ n2824;
  assign n2828 = n2434 & n2827;
  assign n2829 = n2828 ^ n2826;
  assign n2833 = n2832 ^ n2830;
  assign n2834 = n2830 ^ n1056;
  assign n2835 = n2830 ^ n2473;
  assign n2836 = n2830 & ~n2835;
  assign n2837 = n2836 ^ n2830;
  assign n2838 = ~n2834 & n2837;
  assign n2839 = n2838 ^ n2836;
  assign n2840 = n2839 ^ n2830;
  assign n2841 = n2840 ^ n2473;
  assign n2842 = n2833 & ~n2841;
  assign n2843 = n2842 ^ n2830;
  assign n2844 = ~n2829 & ~n2843;
  assign n2847 = n1157 ^ n1056;
  assign n2848 = n2846 & n2847;
  assign n2849 = n2848 ^ n1056;
  assign n2850 = n2849 ^ n2462;
  assign n2851 = n2845 & ~n2850;
  assign n2852 = n2844 & ~n2851;
  assign n2818 = n2817 ^ n2747;
  assign n2853 = n2852 ^ n2818;
  assign n2890 = n2744 ^ n2624;
  assign n2854 = n2473 ^ n2439;
  assign n2855 = n2854 ^ n2473;
  assign n2856 = n2473 ^ n1056;
  assign n2857 = n2856 ^ n2473;
  assign n2858 = ~n2855 & n2857;
  assign n2859 = n2858 ^ n2473;
  assign n2860 = ~n1157 & n2859;
  assign n2861 = n2860 ^ n2473;
  assign n2862 = n2821 & n2861;
  assign n2863 = n2473 & n2820;
  assign n2864 = ~n2439 & n2832;
  assign n2865 = ~n2863 & ~n2864;
  assign n2866 = ~n2862 & n2865;
  assign n2867 = n2866 ^ n1056;
  assign n2868 = n2482 ^ n2454;
  assign n2869 = ~n2473 & n2868;
  assign n2870 = n2869 ^ n2482;
  assign n2871 = ~n2434 & ~n2870;
  assign n2872 = n2845 & ~n2871;
  assign n2873 = n2872 ^ n1056;
  assign n2874 = ~n1056 & n2845;
  assign n2875 = n2434 & ~n2870;
  assign n2876 = n2874 & n2875;
  assign n2877 = n2434 ^ n1157;
  assign n2878 = n2845 & n2870;
  assign n2879 = n2877 & n2878;
  assign n2880 = ~n2876 & ~n2879;
  assign n2881 = n2880 ^ n1056;
  assign n2882 = n1056 & n2881;
  assign n2883 = n2882 ^ n1056;
  assign n2884 = n2873 & n2883;
  assign n2885 = n2884 ^ n2882;
  assign n2886 = n2885 ^ n1056;
  assign n2887 = n2886 ^ n2880;
  assign n2888 = ~n2867 & n2887;
  assign n2889 = n2888 ^ n2880;
  assign n2891 = n2890 ^ n2889;
  assign n2896 = n2894 & n2895;
  assign n2897 = ~n2439 & ~n2823;
  assign n2898 = n1157 & ~n2819;
  assign n2899 = ~n1157 & ~n2821;
  assign n2900 = ~n2898 & ~n2899;
  assign n2901 = n2847 & n2900;
  assign n2902 = n2440 & n2901;
  assign n2903 = ~n2897 & ~n2902;
  assign n2904 = n1056 & ~n2903;
  assign n2905 = ~n2896 & ~n2904;
  assign n2906 = n2473 ^ n1157;
  assign n2907 = n2845 & n2893;
  assign n2908 = ~n2906 & n2907;
  assign n2909 = n2905 & ~n2908;
  assign n2911 = n2845 & ~n2910;
  assign n2912 = ~n1056 & n2903;
  assign n2913 = ~n2911 & n2912;
  assign n2914 = n2909 & ~n2913;
  assign n2892 = n2741 ^ n2649;
  assign n2915 = n2914 ^ n2892;
  assign n2917 = ~n2808 & n2845;
  assign n2918 = n2440 & ~n2823;
  assign n2919 = ~n2441 & n2901;
  assign n2920 = ~n2918 & ~n2919;
  assign n2921 = n1056 & n2920;
  assign n2922 = ~n2917 & n2921;
  assign n2923 = n2800 & n2845;
  assign n2924 = n2439 ^ n1157;
  assign n2925 = n2923 & ~n2924;
  assign n2926 = ~n2922 & ~n2925;
  assign n2927 = n2801 & n2874;
  assign n2928 = ~n1056 & ~n2920;
  assign n2929 = ~n2927 & ~n2928;
  assign n2930 = n2926 & n2929;
  assign n2916 = n2738 ^ n2721;
  assign n2931 = n2930 ^ n2916;
  assign n2933 = n2599 & n2845;
  assign n2934 = n2440 ^ n1157;
  assign n2935 = n2933 & ~n2934;
  assign n2936 = ~n2441 & ~n2823;
  assign n2937 = n2442 & n2901;
  assign n2938 = ~n2936 & ~n2937;
  assign n2939 = n2938 ^ n1056;
  assign n2940 = ~n2615 & n2845;
  assign n2941 = n2940 ^ n2938;
  assign n2942 = n2600 & n2895;
  assign n2943 = n2942 ^ n2940;
  assign n2944 = n2940 & ~n2943;
  assign n2945 = n2944 ^ n2940;
  assign n2946 = n2941 & n2945;
  assign n2947 = n2946 ^ n2944;
  assign n2948 = n2947 ^ n2940;
  assign n2949 = n2948 ^ n2942;
  assign n2950 = n2939 & ~n2949;
  assign n2951 = n2950 ^ n2942;
  assign n2952 = ~n2935 & ~n2951;
  assign n2932 = n2715 ^ n2695;
  assign n2953 = n2952 ^ n2932;
  assign n2957 = n2442 & ~n2823;
  assign n2958 = ~n2443 & n2901;
  assign n2959 = ~n2957 & ~n2958;
  assign n2960 = n1056 & n2959;
  assign n2961 = n2632 & n2960;
  assign n2962 = ~n2874 & ~n2961;
  assign n2963 = n1157 & n2632;
  assign n2964 = ~n2441 & ~n2963;
  assign n2965 = ~n2962 & n2964;
  assign n2966 = n2959 ^ n1056;
  assign n2967 = ~n2640 & n2845;
  assign n2968 = n2967 ^ n1056;
  assign n2969 = n2441 & n2632;
  assign n2970 = n1157 & n2845;
  assign n2971 = n2969 & n2970;
  assign n2972 = n2971 ^ n1056;
  assign n2973 = n1056 & ~n2972;
  assign n2974 = n2973 ^ n1056;
  assign n2975 = n2968 & n2974;
  assign n2976 = n2975 ^ n2973;
  assign n2977 = n2976 ^ n1056;
  assign n2978 = n2977 ^ n2971;
  assign n2979 = ~n2966 & ~n2978;
  assign n2980 = n2979 ^ n2971;
  assign n2981 = ~n2965 & ~n2980;
  assign n2954 = n2693 ^ n2672;
  assign n2955 = n2670 & n2671;
  assign n2956 = ~n2954 & ~n2955;
  assign n2982 = n2981 ^ n2956;
  assign n2985 = n2723 & n2874;
  assign n2986 = ~n2443 & ~n2823;
  assign n2987 = n2444 & n2901;
  assign n2988 = ~n2986 & ~n2987;
  assign n2989 = ~n1056 & ~n2988;
  assign n2990 = ~n2985 & ~n2989;
  assign n2991 = n2442 ^ n1157;
  assign n2992 = n2722 & n2845;
  assign n2993 = n2991 & n2992;
  assign n2994 = n2990 & ~n2993;
  assign n2995 = ~n2730 & n2845;
  assign n2996 = n1056 & n2988;
  assign n2997 = ~n2995 & n2996;
  assign n2998 = n2994 & ~n2997;
  assign n2983 = n1097 & n2668;
  assign n2984 = n2983 ^ n2665;
  assign n2999 = n2998 ^ n2984;
  assign n3008 = n2553 & n2847;
  assign n3009 = n3008 ^ n2444;
  assign n3010 = n2845 & n3009;
  assign n3011 = ~n2446 & ~n2823;
  assign n3012 = n2447 & n2901;
  assign n3013 = ~n3011 & ~n3012;
  assign n3014 = ~n3010 & n3013;
  assign n3017 = ~n2539 & ~n2900;
  assign n3018 = n1056 & ~n3017;
  assign n3024 = n2518 & n2847;
  assign n3025 = n3024 ^ n2446;
  assign n3020 = n3019 ^ n2831;
  assign n3021 = n1152 & n3020;
  assign n3022 = n3021 ^ n3019;
  assign n3023 = ~n2474 & n3022;
  assign n3026 = n3025 ^ n3023;
  assign n3027 = n3026 ^ n3025;
  assign n3028 = n1157 ^ n1152;
  assign n3029 = n2447 & n3028;
  assign n3030 = n3029 ^ n3025;
  assign n3031 = n3030 ^ n3025;
  assign n3032 = ~n3027 & ~n3031;
  assign n3033 = n3032 ^ n3025;
  assign n3034 = ~n2845 & n3033;
  assign n3035 = n3034 ^ n3025;
  assign n3036 = n3018 & n3035;
  assign n3015 = ~n1056 & n1061;
  assign n3016 = ~n2474 & n3015;
  assign n3037 = n3036 ^ n3016;
  assign n3038 = n3037 ^ n3016;
  assign n3039 = n1056 & ~n1061;
  assign n3040 = ~n2474 & n3039;
  assign n3041 = n3040 ^ n3016;
  assign n3042 = n3041 ^ n3016;
  assign n3043 = ~n3038 & ~n3042;
  assign n3044 = n3043 ^ n3016;
  assign n3045 = n3014 & ~n3044;
  assign n3046 = n3045 ^ n3016;
  assign n3000 = n2666 ^ n1101;
  assign n3001 = n3000 ^ n1101;
  assign n3002 = n2603 ^ n1101;
  assign n3003 = n3002 ^ n1101;
  assign n3004 = ~n3001 & n3003;
  assign n3005 = n3004 ^ n1101;
  assign n3006 = ~n2474 & ~n3005;
  assign n3007 = n3006 ^ n2666;
  assign n3047 = n3046 ^ n3007;
  assign n3052 = n2576 & n2847;
  assign n3053 = n3052 ^ n1056;
  assign n3054 = n3053 ^ n2443;
  assign n3048 = n2444 & n3028;
  assign n3049 = ~n2446 & n3022;
  assign n3050 = ~n3048 & ~n3049;
  assign n3051 = n3050 ^ n1056;
  assign n3055 = n3054 ^ n3051;
  assign n3056 = ~n2845 & n3055;
  assign n3057 = n3056 ^ n3054;
  assign n3058 = n3057 ^ n3007;
  assign n3059 = n3047 & n3058;
  assign n3060 = n3059 ^ n3046;
  assign n3061 = n3060 ^ n2984;
  assign n3062 = n2999 & n3061;
  assign n3063 = n3062 ^ n2998;
  assign n3064 = n3063 ^ n2956;
  assign n3065 = n2982 & ~n3064;
  assign n3066 = n3065 ^ n2981;
  assign n3067 = n3066 ^ n2932;
  assign n3068 = ~n2953 & ~n3067;
  assign n3069 = n3068 ^ n2952;
  assign n3070 = n3069 ^ n2916;
  assign n3071 = n2931 & n3070;
  assign n3072 = n3071 ^ n2930;
  assign n3073 = n3072 ^ n2892;
  assign n3074 = n2915 & n3073;
  assign n3075 = n3074 ^ n2914;
  assign n3076 = n3075 ^ n2889;
  assign n3077 = ~n2891 & ~n3076;
  assign n3078 = n3077 ^ n3075;
  assign n3079 = n3078 ^ n2818;
  assign n3080 = n2853 & ~n3079;
  assign n3081 = n3080 ^ n2852;
  assign n3153 = n3152 ^ n3081;
  assign n3264 = n3178 ^ n3153;
  assign n3277 = n3276 ^ n3264;
  assign n3290 = n3078 ^ n2853;
  assign n3278 = x1 & ~n3235;
  assign n3279 = n318 & n3166;
  assign n3280 = ~x0 & ~n3279;
  assign n3281 = ~n3278 & n3280;
  assign n3282 = ~n2463 & ~n2472;
  assign n3283 = n2499 & ~n3282;
  assign n3284 = ~n2466 & ~n3283;
  assign n3285 = n320 & n3284;
  assign n3286 = n3285 ^ n2420;
  assign n3287 = x0 & n3286;
  assign n3288 = ~n3281 & ~n3287;
  assign n3289 = n3288 ^ n2511;
  assign n3641 = n3290 ^ n3289;
  assign n3294 = n3289 & n3290;
  assign n3642 = n3641 ^ n3294;
  assign n2425 = x1 & ~x2;
  assign n2426 = x0 & x22;
  assign n2427 = n2425 & n2426;
  assign n3236 = ~n2486 & ~n2489;
  assign n3237 = n3236 ^ n405;
  assign n3238 = ~n3165 & n3237;
  assign n3239 = n3238 ^ n3235;
  assign n3496 = n2427 & ~n3239;
  assign n3418 = ~n25 & n319;
  assign n2416 = ~x0 & x1;
  assign n3497 = ~n320 & ~n2416;
  assign n3498 = ~n3235 & n3497;
  assign n3499 = n318 & ~n2462;
  assign n3500 = x1 ^ x0;
  assign n3501 = x1 & ~n3500;
  assign n3502 = n3501 ^ x1;
  assign n3503 = n3166 ^ x1;
  assign n3504 = n3502 & ~n3503;
  assign n3505 = n3504 ^ n3501;
  assign n3506 = n3505 ^ x1;
  assign n3507 = n3506 ^ x0;
  assign n3508 = ~n3499 & ~n3507;
  assign n3509 = ~n3498 & ~n3508;
  assign n3510 = n3418 & ~n3509;
  assign n3511 = ~n3496 & ~n3510;
  assign n3512 = n2428 & n3509;
  assign n2429 = x22 ^ x1;
  assign n2430 = x0 & n2429;
  assign n3414 = n2510 ^ n2430;
  assign n3513 = n3239 ^ n2430;
  assign n3514 = n3513 ^ n2430;
  assign n3515 = n3414 & n3514;
  assign n3516 = n3515 ^ n2430;
  assign n3517 = n3512 & ~n3516;
  assign n3518 = n3511 & ~n3517;
  assign n3296 = n2462 ^ n317;
  assign n3297 = x1 & ~n3296;
  assign n3298 = n318 & ~n2434;
  assign n3299 = ~x0 & ~n3298;
  assign n3300 = ~n3297 & n3299;
  assign n3302 = n320 & n3165;
  assign n3301 = n3166 ^ n2511;
  assign n3303 = n3302 ^ n3301;
  assign n3304 = x0 & ~n3303;
  assign n3305 = ~n3300 & ~n3304;
  assign n3295 = n3072 ^ n2915;
  assign n3306 = n3305 ^ n3295;
  assign n3308 = x1 & n2434;
  assign n3309 = n318 & n2473;
  assign n3310 = ~x0 & ~n3309;
  assign n3311 = ~n3308 & n3310;
  assign n3312 = n320 & n2846;
  assign n3313 = n3312 ^ n2462;
  assign n3314 = x0 & ~n3313;
  assign n3315 = ~n3311 & ~n3314;
  assign n3316 = n3315 ^ n2511;
  assign n3307 = n3069 ^ n2931;
  assign n3317 = n3316 ^ n3307;
  assign n3319 = n320 & n2870;
  assign n3320 = n3319 ^ n2434;
  assign n3321 = x0 & n3320;
  assign n3322 = n2416 & n2473;
  assign n2419 = ~x0 & n318;
  assign n3323 = n2419 & ~n2439;
  assign n3324 = ~n3322 & ~n3323;
  assign n3325 = ~n3321 & n3324;
  assign n3326 = n3325 ^ n2511;
  assign n3318 = n3066 ^ n2953;
  assign n3327 = n3326 ^ n3318;
  assign n3328 = n3060 ^ n2999;
  assign n3330 = n320 & n2599;
  assign n3331 = n3330 ^ n2440;
  assign n3332 = x0 & n3331;
  assign n3333 = n2416 & ~n2441;
  assign n3334 = n2419 & n2442;
  assign n3335 = ~n3333 & ~n3334;
  assign n3336 = ~n3332 & n3335;
  assign n3337 = n3336 ^ n2511;
  assign n3329 = n3057 ^ n3047;
  assign n3338 = n3337 ^ n3329;
  assign n321 = x0 & ~n320;
  assign n3346 = n321 & ~n2441;
  assign n3347 = n2416 & n2442;
  assign n3348 = n2419 & ~n2443;
  assign n3349 = ~n3347 & ~n3348;
  assign n3350 = ~n3346 & n3349;
  assign n3351 = n2511 & n3350;
  assign n3352 = n2632 ^ n2441;
  assign n3353 = n2430 & ~n3352;
  assign n3354 = n3351 & ~n3353;
  assign n3355 = n319 & ~n3350;
  assign n3356 = n318 & n2509;
  assign n3357 = ~n2427 & ~n3356;
  assign n3358 = ~n3352 & ~n3357;
  assign n3359 = ~n3355 & ~n3358;
  assign n3360 = ~n3354 & n3359;
  assign n3341 = n3014 & ~n3036;
  assign n3342 = n3341 ^ n1061;
  assign n3339 = n1056 & ~n3036;
  assign n3340 = n3339 ^ n3014;
  assign n3343 = n3342 ^ n3340;
  assign n3344 = n2474 & n3343;
  assign n3345 = n3344 ^ n3342;
  assign n3361 = n3360 ^ n3345;
  assign n3372 = n2447 & n2845;
  assign n3426 = n2474 & ~n3372;
  assign n3427 = n1056 & ~n2900;
  assign n3428 = ~n3426 & n3427;
  assign n3429 = n3428 ^ n3035;
  assign n3384 = n320 & n2553;
  assign n3385 = n3384 ^ n2444;
  assign n3386 = x0 & n3385;
  assign n3387 = n2416 & ~n2446;
  assign n3388 = n2419 & n2447;
  assign n3389 = ~n3387 & ~n3388;
  assign n3390 = ~n3386 & n3389;
  assign n3393 = n2446 ^ n1152;
  assign n3394 = n3393 ^ n1152;
  assign n3395 = n2203 ^ n1152;
  assign n3396 = n3395 ^ n1152;
  assign n3397 = n3394 & ~n3396;
  assign n3398 = n3397 ^ n1152;
  assign n3399 = n2474 & ~n3398;
  assign n3400 = n3399 ^ n1152;
  assign n3401 = n2511 & ~n3400;
  assign n3391 = n1152 & ~n2511;
  assign n3392 = ~n2474 & n3391;
  assign n3402 = n3401 ^ n3392;
  assign n3403 = ~n3390 & n3402;
  assign n3404 = n3403 ^ n3401;
  assign n3362 = n3028 ^ n1157;
  assign n3363 = n3362 ^ n2511;
  assign n3364 = n2511 ^ n1157;
  assign n3365 = n3364 ^ n2511;
  assign n3366 = n2511 ^ n2447;
  assign n3367 = n3366 ^ n2511;
  assign n3368 = n3365 & n3367;
  assign n3369 = n3368 ^ n2511;
  assign n3370 = n3363 & ~n3369;
  assign n3371 = n3370 ^ n3028;
  assign n3373 = n3372 ^ n3371;
  assign n3374 = n3372 ^ n1157;
  assign n3375 = n3372 ^ n2474;
  assign n3376 = n3372 & ~n3375;
  assign n3377 = n3376 ^ n3372;
  assign n3378 = ~n3374 & n3377;
  assign n3379 = n3378 ^ n3376;
  assign n3380 = n3379 ^ n3372;
  assign n3381 = n3380 ^ n2474;
  assign n3382 = n3373 & ~n3381;
  assign n3383 = n3382 ^ n3372;
  assign n3405 = n3404 ^ n3383;
  assign n3406 = x0 & n2443;
  assign n3407 = n2416 & ~n2444;
  assign n3408 = n318 & n2446;
  assign n3409 = x0 & n320;
  assign n3410 = ~n3408 & ~n3409;
  assign n3411 = ~n3407 & n3410;
  assign n3412 = ~n3406 & n3411;
  assign n3413 = n2428 & ~n3412;
  assign n3415 = ~n2696 & n3414;
  assign n3416 = n3415 ^ n2510;
  assign n3417 = n3413 & ~n3416;
  assign n3419 = n3412 & n3418;
  assign n3420 = n2427 & ~n2696;
  assign n3421 = ~n3419 & ~n3420;
  assign n3422 = ~n3417 & n3421;
  assign n3423 = n3422 ^ n3383;
  assign n3424 = n3405 & n3423;
  assign n3425 = n3424 ^ n3404;
  assign n3430 = n3429 ^ n3425;
  assign n3431 = n321 & n2442;
  assign n3432 = n2416 & ~n2443;
  assign n3433 = n2419 & n2444;
  assign n3434 = ~n3432 & ~n3433;
  assign n3435 = ~n3431 & n3434;
  assign n3436 = n2511 & n3435;
  assign n3437 = n2722 ^ n2442;
  assign n3438 = n3409 & n3437;
  assign n3439 = n3436 & ~n3438;
  assign n3440 = n319 & ~n3435;
  assign n3441 = ~n3357 & n3437;
  assign n3442 = ~n3440 & ~n3441;
  assign n3443 = ~n3439 & n3442;
  assign n3444 = n3443 ^ n3429;
  assign n3445 = ~n3430 & ~n3444;
  assign n3446 = n3445 ^ n3425;
  assign n3447 = n3446 ^ n3345;
  assign n3448 = n3361 & n3447;
  assign n3449 = n3448 ^ n3360;
  assign n3450 = n3449 ^ n3329;
  assign n3451 = n3338 & ~n3450;
  assign n3452 = n3451 ^ n3337;
  assign n3453 = n3328 & ~n3452;
  assign n3455 = n320 & n2800;
  assign n3456 = n3455 ^ n2439;
  assign n3454 = n318 & ~n2441;
  assign n3457 = n3456 ^ n3454;
  assign n3458 = n3457 ^ n3456;
  assign n3459 = x1 & n2440;
  assign n3460 = n3459 ^ n3456;
  assign n3461 = n3460 ^ n3456;
  assign n3462 = ~n3458 & ~n3461;
  assign n3463 = n3462 ^ n3456;
  assign n3464 = ~x0 & n3463;
  assign n3465 = n3464 ^ n3456;
  assign n3466 = n3465 ^ n2511;
  assign n3467 = n3063 ^ n2982;
  assign n3468 = n320 & n2893;
  assign n3469 = n3468 ^ n2473;
  assign n3470 = x0 & n3469;
  assign n3471 = n2416 & ~n2439;
  assign n3472 = n2419 & n2440;
  assign n3473 = ~n3471 & ~n3472;
  assign n3474 = ~n3470 & n3473;
  assign n3475 = n3474 ^ n3465;
  assign n3476 = ~n3467 & n3475;
  assign n3477 = n3466 & n3476;
  assign n3478 = n3477 ^ n3466;
  assign n3479 = ~n3453 & n3478;
  assign n3480 = n3474 ^ n2511;
  assign n3481 = n3480 ^ n3467;
  assign n3482 = ~n3328 & n3452;
  assign n3483 = n3482 ^ n3480;
  assign n3484 = n3481 & ~n3483;
  assign n3485 = n3484 ^ n3467;
  assign n3486 = ~n3479 & ~n3485;
  assign n3487 = n3486 ^ n3318;
  assign n3488 = ~n3327 & ~n3487;
  assign n3489 = n3488 ^ n3326;
  assign n3490 = n3489 ^ n3307;
  assign n3491 = n3317 & n3490;
  assign n3492 = n3491 ^ n3316;
  assign n3493 = n3492 ^ n3295;
  assign n3494 = ~n3306 & n3493;
  assign n3495 = n3494 ^ n3305;
  assign n3519 = n3518 ^ n3495;
  assign n3520 = n3075 ^ n2891;
  assign n3521 = n3520 ^ n3518;
  assign n3522 = ~n3519 & n3521;
  assign n3523 = n3522 ^ n3495;
  assign n3643 = ~n351 & ~n467;
  assign n3644 = ~n395 & n3643;
  assign n3645 = n2288 & n3644;
  assign n3646 = n2054 & n3645;
  assign n3647 = ~n272 & ~n935;
  assign n3648 = n3646 & n3647;
  assign n3649 = ~n269 & n3648;
  assign n3650 = ~n356 & ~n374;
  assign n3651 = ~n191 & n3650;
  assign n3652 = n84 & ~n159;
  assign n3653 = n2113 & ~n3652;
  assign n3654 = n3651 & n3653;
  assign n3655 = n2123 & n3654;
  assign n3656 = n127 & ~n209;
  assign n3657 = n2239 & n3656;
  assign n3658 = n3655 & n3657;
  assign n3659 = n85 & ~n184;
  assign n3660 = n2317 & ~n3659;
  assign n3661 = n762 & n3660;
  assign n3662 = n3658 & n3661;
  assign n3663 = n3649 & n3662;
  assign n3664 = n3523 & ~n3663;
  assign n3665 = ~n57 & ~n380;
  assign n3666 = ~n2095 & n3665;
  assign n3667 = n168 & n186;
  assign n3668 = ~n3666 & ~n3667;
  assign n3669 = n952 & ~n3668;
  assign n285 = ~n283 & ~n284;
  assign n286 = ~n282 & n285;
  assign n3670 = ~n140 & ~n786;
  assign n3671 = n286 & n3670;
  assign n3672 = n2094 & n3671;
  assign n3673 = n3669 & n3672;
  assign n3674 = ~n324 & ~n915;
  assign n3675 = n774 & n3674;
  assign n3676 = n3673 & n3675;
  assign n3677 = ~n198 & ~n388;
  assign n3678 = n2349 & n3677;
  assign n3679 = n907 & n3678;
  assign n3680 = n150 & ~n162;
  assign n3681 = ~n139 & n3680;
  assign n3682 = ~n743 & ~n3681;
  assign n3683 = ~n810 & ~n3682;
  assign n3684 = n3679 & n3683;
  assign n3685 = n2171 & n3684;
  assign n3686 = ~n191 & ~n656;
  assign n3687 = n57 & ~n184;
  assign n3688 = ~n358 & ~n3687;
  assign n3689 = n3686 & n3688;
  assign n3690 = n292 & n596;
  assign n3691 = n3689 & n3690;
  assign n3692 = ~n210 & ~n345;
  assign n3693 = n102 & ~n498;
  assign n3694 = ~n1963 & ~n3693;
  assign n3695 = n3692 & n3694;
  assign n3696 = n3691 & n3695;
  assign n3697 = n3685 & n3696;
  assign n3698 = n3676 & n3697;
  assign n3699 = n3664 & ~n3698;
  assign n3700 = n3699 ^ n3641;
  assign n3701 = n3700 ^ n3699;
  assign n3702 = n3699 ^ n3523;
  assign n3703 = n3701 & n3702;
  assign n3704 = n3703 ^ n3699;
  assign n3705 = n3642 & n3704;
  assign n3706 = n3705 ^ n3294;
  assign n3707 = n3277 & ~n3706;
  assign n3708 = ~n3294 & n3698;
  assign n3709 = ~n3277 & ~n3708;
  assign n3291 = ~n3289 & ~n3290;
  assign n3710 = n3291 & ~n3664;
  assign n3711 = n3709 & ~n3710;
  assign n3524 = ~n3294 & ~n3523;
  assign n3712 = n3524 & n3663;
  assign n3713 = n3711 & ~n3712;
  assign n3714 = ~n3707 & ~n3713;
  assign n3715 = n3641 & ~n3663;
  assign n3716 = ~n3664 & n3698;
  assign n3717 = ~n3715 & n3716;
  assign n3718 = ~n3714 & ~n3717;
  assign n3719 = ~n147 & ~n260;
  assign n3720 = ~n291 & ~n2121;
  assign n3721 = ~n438 & ~n487;
  assign n3722 = n3720 & n3721;
  assign n3723 = n1113 & n3722;
  assign n3724 = n2052 & n2380;
  assign n3725 = n102 & ~n369;
  assign n3726 = ~n675 & ~n3725;
  assign n3727 = ~n78 & n84;
  assign n3728 = ~n822 & ~n3727;
  assign n3729 = ~n299 & n3728;
  assign n3730 = n3726 & n3729;
  assign n3731 = n3724 & n3730;
  assign n3732 = n3723 & n3731;
  assign n3733 = n783 & n3732;
  assign n3734 = ~n3719 & n3733;
  assign n3735 = ~n352 & n591;
  assign n3736 = ~n190 & ~n454;
  assign n3737 = n57 & ~n180;
  assign n3738 = ~n771 & ~n3737;
  assign n3739 = n3736 & n3738;
  assign n3740 = n2361 & n3739;
  assign n3741 = n631 & n3740;
  assign n3742 = n307 & n2318;
  assign n3743 = ~n418 & n749;
  assign n3744 = n379 & n3743;
  assign n3745 = n1972 & n3744;
  assign n3746 = n3742 & n3745;
  assign n3747 = n3741 & n3746;
  assign n3748 = n3735 & n3747;
  assign n3749 = n3734 & n3748;
  assign n3750 = n3718 & ~n3749;
  assign n3292 = n3291 ^ n3264;
  assign n3293 = n3292 ^ n3264;
  assign n3525 = n3524 ^ n3264;
  assign n3526 = n3525 ^ n3264;
  assign n3527 = ~n3293 & ~n3526;
  assign n3528 = n3527 ^ n3264;
  assign n3529 = n3277 & ~n3528;
  assign n3530 = n3529 ^ n3276;
  assign n3240 = ~n2847 & n3235;
  assign n3241 = n3240 ^ n1056;
  assign n3242 = n2845 & n3241;
  assign n3243 = ~n3239 & n3242;
  assign n3244 = ~n3235 & n3238;
  assign n3245 = n2970 & n3244;
  assign n3246 = ~n3243 & ~n3245;
  assign n3247 = n3235 & ~n3238;
  assign n3248 = n2874 & ~n3247;
  assign n3249 = ~n2823 & n3166;
  assign n3250 = n2819 & n3154;
  assign n3251 = n3250 ^ n1056;
  assign n3252 = n3251 ^ n3250;
  assign n3253 = n2462 & n2830;
  assign n3254 = n3253 ^ n3250;
  assign n3255 = n3252 & n3254;
  assign n3256 = n3255 ^ n3250;
  assign n3257 = ~n3249 & ~n3256;
  assign n3258 = n3257 ^ n1056;
  assign n3259 = ~n3248 & n3258;
  assign n3260 = n3246 & ~n3259;
  assign n3219 = n2598 & n2875;
  assign n3220 = n2473 & n2606;
  assign n3221 = ~n2439 & n2610;
  assign n3222 = ~n3220 & ~n3221;
  assign n3223 = ~n3219 & n3222;
  assign n3224 = n1097 & ~n3223;
  assign n3225 = n2598 & ~n2871;
  assign n3226 = ~n1097 & n3222;
  assign n3227 = ~n3225 & n3226;
  assign n3228 = n2598 & n2870;
  assign n3229 = n2434 ^ n1101;
  assign n3230 = n3228 & n3229;
  assign n3231 = ~n3227 & ~n3230;
  assign n3232 = ~n3224 & n3231;
  assign n3203 = n2522 & n2600;
  assign n3204 = ~n2441 & n2528;
  assign n3205 = n2442 & n2535;
  assign n3206 = ~n3204 & ~n3205;
  assign n3207 = ~n3203 & n3206;
  assign n3208 = ~n684 & ~n3207;
  assign n3209 = n2522 & ~n2615;
  assign n3210 = n684 & n3206;
  assign n3211 = ~n3209 & n3210;
  assign n3212 = n2522 & n2599;
  assign n3213 = n2440 ^ n850;
  assign n3214 = n3212 & n3213;
  assign n3215 = ~n3211 & ~n3214;
  assign n3216 = ~n3208 & n3215;
  assign n3195 = ~n551 & ~n2474;
  assign n3196 = ~n3088 & ~n3195;
  assign n3197 = ~n3109 & ~n3196;
  assign n3198 = ~n2447 & ~n3197;
  assign n3199 = ~n551 & n3198;
  assign n3200 = n2447 & n3197;
  assign n3201 = ~n3199 & ~n3200;
  assign n3188 = n552 & n2576;
  assign n3189 = n3188 ^ n2443;
  assign n3190 = n685 & ~n3189;
  assign n3191 = n2444 & ~n2763;
  assign n3192 = ~n2446 & n2767;
  assign n3193 = ~n3191 & ~n3192;
  assign n3194 = ~n3190 & n3193;
  assign n3202 = n3201 ^ n3194;
  assign n3217 = n3216 ^ n3202;
  assign n3185 = n3114 ^ n3087;
  assign n3186 = n3135 & ~n3185;
  assign n3187 = n3186 ^ n3134;
  assign n3218 = n3217 ^ n3187;
  assign n3233 = n3232 ^ n3218;
  assign n3182 = n3136 ^ n3084;
  assign n3183 = n3151 & ~n3182;
  assign n3184 = n3183 ^ n3150;
  assign n3234 = n3233 ^ n3184;
  assign n3261 = n3260 ^ n3234;
  assign n3179 = n3178 ^ n3081;
  assign n3180 = ~n3153 & n3179;
  assign n3181 = n3180 ^ n3178;
  assign n3262 = n3261 ^ n3181;
  assign n2401 = n2385 & n2400;
  assign n2402 = ~n288 & n2388;
  assign n2403 = n78 & n1029;
  assign n2404 = n174 & ~n2403;
  assign n2405 = ~n299 & ~n2404;
  assign n2406 = ~n385 & n2405;
  assign n2407 = n265 & n495;
  assign n2408 = ~n81 & n2407;
  assign n2409 = n48 & ~n2408;
  assign n2410 = n2122 & ~n2409;
  assign n2411 = n2406 & n2410;
  assign n2412 = n502 & n2411;
  assign n2413 = n2402 & n2412;
  assign n2414 = ~n2401 & ~n2413;
  assign n2415 = n321 & n2414;
  assign n2418 = n2416 & ~n2417;
  assign n2421 = n2419 & ~n2420;
  assign n2422 = ~n2418 & ~n2421;
  assign n2423 = ~n2415 & n2422;
  assign n2424 = n319 & ~n2423;
  assign n2470 = ~n2385 & n2400;
  assign n2471 = ~n2469 & n2470;
  assign n2502 = n2501 ^ n2385;
  assign n2503 = n2400 & ~n2502;
  assign n2504 = n2503 ^ n2501;
  assign n2505 = ~n2471 & n2504;
  assign n2506 = n2505 ^ n2414;
  assign n2431 = n2428 & ~n2430;
  assign n2432 = n2423 & n2431;
  assign n2433 = ~n2427 & ~n2432;
  assign n2507 = n2506 ^ n2433;
  assign n2508 = n2507 ^ n2433;
  assign n2512 = n2423 & n2511;
  assign n2513 = n2512 ^ n2433;
  assign n2514 = ~n2508 & ~n2513;
  assign n2515 = n2514 ^ n2433;
  assign n2516 = ~n2424 & n2515;
  assign n3263 = n3262 ^ n2516;
  assign n3751 = n3530 ^ n3263;
  assign n3752 = n3750 & n3751;
  assign n3753 = ~n3718 & n3749;
  assign n3754 = ~n3751 & n3753;
  assign n3755 = ~n3752 & ~n3754;
  assign n3612 = x1 & n2414;
  assign n3613 = n318 & ~n2417;
  assign n3614 = ~x0 & ~n3613;
  assign n3615 = ~n3612 & n3614;
  assign n3630 = n2413 & n2504;
  assign n3631 = n2414 & ~n2471;
  assign n3632 = ~n3630 & ~n3631;
  assign n3633 = n320 & n3632;
  assign n3616 = n253 & n753;
  assign n3617 = n57 & ~n3616;
  assign n3618 = ~n138 & ~n347;
  assign n3619 = n101 & ~n125;
  assign n3620 = n3618 & ~n3619;
  assign n3621 = ~n3617 & n3620;
  assign n3622 = ~n297 & ~n786;
  assign n3623 = n3621 & n3622;
  assign n3624 = ~n638 & ~n1025;
  assign n3625 = n172 & n3624;
  assign n3626 = n101 & ~n2408;
  assign n3627 = n3625 & ~n3626;
  assign n3628 = n3623 & n3627;
  assign n3629 = n974 & n3628;
  assign n3634 = n3633 ^ n3629;
  assign n3635 = x0 & n3634;
  assign n3636 = ~n3615 & ~n3635;
  assign n3637 = n3636 ^ n2511;
  assign n3593 = n2462 & ~n2846;
  assign n3594 = n2598 & n3593;
  assign n3595 = n2434 & n2606;
  assign n3596 = n2473 & n2610;
  assign n3597 = ~n3595 & ~n3596;
  assign n3598 = ~n3594 & n3597;
  assign n3599 = n1097 & ~n3598;
  assign n3600 = ~n2462 & ~n2846;
  assign n3601 = n2598 & ~n3600;
  assign n3602 = ~n1097 & n3597;
  assign n3603 = ~n3601 & n3602;
  assign n3604 = n2598 & n2846;
  assign n3605 = n2462 ^ n1101;
  assign n3606 = n3604 & n3605;
  assign n3607 = ~n3603 & ~n3606;
  assign n3608 = ~n3599 & n3607;
  assign n3576 = n2522 & n2801;
  assign n3577 = n2440 & n2528;
  assign n3578 = ~n2441 & n2535;
  assign n3579 = ~n3577 & ~n3578;
  assign n3580 = ~n3576 & n3579;
  assign n3581 = ~n684 & ~n3580;
  assign n3582 = n2522 & ~n2808;
  assign n3583 = n684 & n3579;
  assign n3584 = ~n3582 & n3583;
  assign n3585 = n2522 & n2800;
  assign n3586 = n2439 ^ n850;
  assign n3587 = n3585 & ~n3586;
  assign n3588 = ~n3584 & ~n3587;
  assign n3589 = ~n3581 & n3588;
  assign n3569 = n3197 ^ n2447;
  assign n3570 = n3197 ^ n3194;
  assign n3571 = n3569 & ~n3570;
  assign n3572 = n3571 ^ n2447;
  assign n3573 = n3572 ^ n2446;
  assign n3574 = ~n551 & n3573;
  assign n3562 = n552 & n2722;
  assign n3563 = n3562 ^ n2442;
  assign n3564 = n685 & n3563;
  assign n3565 = ~n2443 & ~n2763;
  assign n3566 = n2444 & n2767;
  assign n3567 = ~n3565 & ~n3566;
  assign n3568 = ~n3564 & n3567;
  assign n3575 = n3574 ^ n3568;
  assign n3590 = n3589 ^ n3575;
  assign n3559 = n3202 ^ n3187;
  assign n3560 = ~n3217 & ~n3559;
  assign n3561 = n3560 ^ n3216;
  assign n3591 = n3590 ^ n3561;
  assign n3556 = n3232 ^ n3184;
  assign n3557 = n3233 & n3556;
  assign n3558 = n3557 ^ n3184;
  assign n3592 = n3591 ^ n3558;
  assign n3609 = n3608 ^ n3592;
  assign n3553 = n3260 ^ n3181;
  assign n3554 = n3261 & n3553;
  assign n3555 = n3554 ^ n3181;
  assign n3610 = n3609 ^ n3555;
  assign n3534 = n2847 & n3284;
  assign n3535 = n3534 ^ n1056;
  assign n3536 = n3535 ^ n2420;
  assign n3537 = n2845 & n3536;
  assign n3538 = n2826 & n3235;
  assign n3539 = n3166 ^ n2830;
  assign n3540 = n2830 & ~n3539;
  assign n3541 = n3540 ^ n2830;
  assign n3542 = ~n2834 & n3541;
  assign n3543 = n3542 ^ n3540;
  assign n3544 = n3543 ^ n2830;
  assign n3545 = n3544 ^ n3166;
  assign n3546 = n2833 & ~n3545;
  assign n3547 = n3546 ^ n2830;
  assign n3548 = ~n3538 & ~n3547;
  assign n3549 = n1056 & ~n3235;
  assign n3550 = ~n2823 & n3549;
  assign n3551 = n3548 & ~n3550;
  assign n3552 = ~n3537 & n3551;
  assign n3611 = n3610 ^ n3552;
  assign n3638 = n3637 ^ n3611;
  assign n3531 = n3530 ^ n2516;
  assign n3532 = ~n3263 & ~n3531;
  assign n3533 = n3532 ^ n3530;
  assign n3639 = n3638 ^ n3533;
  assign n287 = ~n281 & n286;
  assign n293 = ~n207 & n292;
  assign n294 = n289 & n293;
  assign n295 = n287 & n294;
  assign n312 = n302 & n311;
  assign n313 = n295 & n312;
  assign n314 = n280 & n313;
  assign n315 = n260 & n314;
  assign n316 = n197 & n315;
  assign n3640 = n3639 ^ n316;
  assign n3756 = n3755 ^ n3640;
  assign n3907 = x23 ^ x22;
  assign n3908 = n3907 ^ n316;
  assign n3909 = n3640 & n3908;
  assign n3910 = n3909 ^ n3639;
  assign n3911 = n3754 & n3910;
  assign n3912 = n316 & n3639;
  assign n3913 = ~n3907 & n3912;
  assign n3914 = n3913 ^ n3910;
  assign n3915 = ~n3752 & ~n3914;
  assign n3916 = n3915 ^ n3910;
  assign n3917 = ~n3911 & n3916;
  assign n3918 = ~n316 & ~n3639;
  assign n3919 = ~n3754 & n3918;
  assign n3920 = n3907 & n3919;
  assign n3921 = n3917 & ~n3920;
  assign n3877 = n318 & n2414;
  assign n3878 = x1 & ~n3629;
  assign n3879 = ~x0 & ~n3878;
  assign n3880 = ~n3877 & n3879;
  assign n3896 = ~n3629 & ~n3630;
  assign n3897 = n3629 & ~n3631;
  assign n3898 = ~n3896 & ~n3897;
  assign n3899 = n320 & n3898;
  assign n3772 = ~n298 & ~n393;
  assign n3773 = ~n356 & n3772;
  assign n3881 = n162 & ~n949;
  assign n3882 = n3773 & ~n3881;
  assign n3883 = n1081 & n3882;
  assign n3884 = n141 & n346;
  assign n3885 = n3883 & n3884;
  assign n3886 = n471 & n493;
  assign n3887 = n139 & ~n3886;
  assign n3888 = n512 & ~n3887;
  assign n3889 = ~n558 & n2292;
  assign n3890 = ~n771 & n3889;
  assign n3891 = ~n425 & n3890;
  assign n3892 = n3888 & n3891;
  assign n3893 = n763 & n3892;
  assign n3894 = n3885 & n3893;
  assign n3895 = n2262 & n3894;
  assign n3900 = n3899 ^ n3895;
  assign n3901 = x0 & n3900;
  assign n3902 = ~n3880 & ~n3901;
  assign n3903 = n3902 ^ n2511;
  assign n3859 = ~n2417 & ~n3270;
  assign n3860 = n2895 & n3859;
  assign n3861 = ~n2420 & ~n2823;
  assign n3862 = n2901 & ~n3235;
  assign n3863 = ~n3861 & ~n3862;
  assign n3864 = n1056 & ~n3863;
  assign n3865 = ~n3860 & ~n3864;
  assign n3866 = n2845 & n3270;
  assign n3867 = n2417 ^ n1157;
  assign n3868 = n3866 & n3867;
  assign n3869 = n3865 & ~n3868;
  assign n3870 = n2417 & ~n3270;
  assign n3871 = n2845 & ~n3870;
  assign n3872 = ~n1056 & n3863;
  assign n3873 = ~n3871 & n3872;
  assign n3874 = n3869 & ~n3873;
  assign n3843 = n2598 & n3171;
  assign n3844 = n2462 & n2606;
  assign n3845 = n2434 & n2610;
  assign n3846 = ~n3844 & ~n3845;
  assign n3847 = ~n3843 & n3846;
  assign n3848 = ~n1097 & ~n3847;
  assign n3849 = n2598 & ~n3175;
  assign n3850 = n1097 & n3846;
  assign n3851 = ~n3849 & n3850;
  assign n3852 = n3166 ^ n1101;
  assign n3853 = n2598 & ~n3852;
  assign n3854 = n3165 & n3853;
  assign n3855 = ~n3851 & ~n3854;
  assign n3856 = ~n3848 & n3855;
  assign n3821 = n2473 ^ n850;
  assign n3822 = n2522 & n2893;
  assign n3823 = ~n3821 & n3822;
  assign n3824 = ~n2439 & n2528;
  assign n3825 = n2440 & n2535;
  assign n3826 = ~n3824 & ~n3825;
  assign n3827 = n3826 ^ n684;
  assign n3828 = n2522 & ~n2910;
  assign n3829 = n3828 ^ n3826;
  assign n3830 = n2777 & n2894;
  assign n3831 = n3830 ^ n3828;
  assign n3832 = n3828 & ~n3831;
  assign n3833 = n3832 ^ n3828;
  assign n3834 = n3829 & n3833;
  assign n3835 = n3834 ^ n3832;
  assign n3836 = n3835 ^ n3828;
  assign n3837 = n3836 ^ n3830;
  assign n3838 = n3827 & ~n3837;
  assign n3839 = n3838 ^ n3830;
  assign n3840 = ~n3823 & ~n3839;
  assign n3814 = n3568 ^ n2446;
  assign n3815 = ~n3573 & ~n3814;
  assign n3816 = n3815 ^ n2446;
  assign n3817 = ~n551 & ~n3816;
  assign n3818 = n3817 ^ n2444;
  assign n3819 = ~n551 & ~n3818;
  assign n3792 = n552 & n2632;
  assign n3793 = n3792 ^ n2441;
  assign n3794 = n685 & n3793;
  assign n3795 = n2443 ^ n2442;
  assign n3796 = n3795 ^ n2442;
  assign n3797 = n2442 ^ n551;
  assign n3798 = n3797 ^ n2442;
  assign n3799 = ~n3796 & n3798;
  assign n3800 = n3799 ^ n2442;
  assign n3801 = n684 & n3800;
  assign n3802 = n3801 ^ n2442;
  assign n3803 = ~n543 & n3802;
  assign n3804 = n543 & n2442;
  assign n3805 = n3804 ^ n538;
  assign n3806 = n3805 ^ n3804;
  assign n3807 = ~n2443 & n3098;
  assign n3808 = n3807 ^ n3804;
  assign n3809 = ~n3806 & n3808;
  assign n3810 = n3809 ^ n3804;
  assign n3811 = ~n685 & ~n3810;
  assign n3812 = ~n3803 & n3811;
  assign n3813 = ~n3794 & ~n3812;
  assign n3820 = n3819 ^ n3813;
  assign n3841 = n3840 ^ n3820;
  assign n3789 = n3575 ^ n3561;
  assign n3790 = n3590 & ~n3789;
  assign n3791 = n3790 ^ n3589;
  assign n3842 = n3841 ^ n3791;
  assign n3857 = n3856 ^ n3842;
  assign n3786 = n3608 ^ n3558;
  assign n3787 = n3592 & n3786;
  assign n3788 = n3787 ^ n3608;
  assign n3858 = n3857 ^ n3788;
  assign n3875 = n3874 ^ n3858;
  assign n3783 = n3609 ^ n3552;
  assign n3784 = ~n3610 & n3783;
  assign n3785 = n3784 ^ n3555;
  assign n3876 = n3875 ^ n3785;
  assign n3904 = n3903 ^ n3876;
  assign n3780 = n3637 ^ n3533;
  assign n3781 = n3638 & n3780;
  assign n3782 = n3781 ^ n3533;
  assign n3905 = n3904 ^ n3782;
  assign n3757 = ~n566 & ~n786;
  assign n3758 = n85 & ~n514;
  assign n3759 = ~n643 & ~n3758;
  assign n3760 = n3757 & n3759;
  assign n3761 = n307 & n3760;
  assign n3762 = n57 & ~n2355;
  assign n3763 = ~n344 & ~n3762;
  assign n3764 = n3643 & n3763;
  assign n3765 = n3761 & n3764;
  assign n3766 = n2019 & n3765;
  assign n3767 = n270 & ~n425;
  assign n3768 = ~n388 & ~n665;
  assign n3769 = n3767 & n3768;
  assign n3770 = n3766 & n3769;
  assign n3771 = n3732 & n3770;
  assign n3774 = n2392 & n3773;
  assign n3775 = n3742 & n3774;
  assign n3776 = ~n809 & ~n3775;
  assign n3777 = ~n432 & ~n447;
  assign n3778 = ~n3776 & n3777;
  assign n3779 = n3771 & n3778;
  assign n3906 = n3905 ^ n3779;
  assign n3922 = n3921 ^ n3906;
  assign n3940 = ~n3906 & ~n3912;
  assign n3941 = n3752 & ~n3940;
  assign n3923 = n3749 ^ n3718;
  assign n3924 = n3751 ^ n3749;
  assign n3925 = ~n3923 & n3924;
  assign n3926 = n3925 ^ n3718;
  assign n3942 = n3640 & ~n3754;
  assign n3943 = ~n3926 & n3942;
  assign n3944 = ~n3941 & ~n3943;
  assign n3945 = n3752 & n3918;
  assign n3946 = n3906 & ~n3945;
  assign n3947 = ~n3944 & ~n3946;
  assign n3927 = ~n3912 & n3926;
  assign n3928 = ~n3752 & n3927;
  assign n3929 = ~n3906 & ~n3918;
  assign n3930 = ~n3928 & n3929;
  assign n3931 = n3906 ^ n3754;
  assign n3932 = n3918 ^ n3912;
  assign n3933 = n3918 ^ n3906;
  assign n3934 = n3933 ^ n3918;
  assign n3935 = n3932 & n3934;
  assign n3936 = n3935 ^ n3918;
  assign n3937 = ~n3931 & ~n3936;
  assign n3938 = n3937 ^ n3754;
  assign n3939 = ~n3930 & n3938;
  assign n3948 = n3947 ^ n3939;
  assign n4051 = n3895 ^ n317;
  assign n4052 = x1 & n4051;
  assign n4053 = n318 & n3629;
  assign n4054 = ~x0 & ~n4053;
  assign n4055 = ~n4052 & n4054;
  assign n4056 = n3897 ^ n3896;
  assign n4057 = ~n3895 & n4056;
  assign n4058 = n4057 ^ n3896;
  assign n4059 = n4058 ^ n2429;
  assign n4060 = n4059 ^ n2429;
  assign n4061 = n2429 ^ n317;
  assign n4062 = ~n4060 & n4061;
  assign n4063 = n4062 ^ n2429;
  assign n4064 = x0 & n4063;
  assign n4065 = ~n4055 & ~n4064;
  assign n4021 = n1157 & ~n2417;
  assign n4022 = ~n2420 & n3019;
  assign n4023 = ~n4021 & ~n4022;
  assign n4024 = n2821 & ~n4023;
  assign n4025 = ~n2417 & n2820;
  assign n4026 = ~n2420 & n2832;
  assign n4027 = ~n4025 & ~n4026;
  assign n4028 = ~n4024 & n4027;
  assign n4029 = n1056 & n4028;
  assign n4030 = n2505 & n4029;
  assign n4031 = ~n2874 & ~n4030;
  assign n4032 = n1157 & n2505;
  assign n4033 = n2414 & ~n4032;
  assign n4034 = ~n4031 & n4033;
  assign n4035 = n4028 ^ n1056;
  assign n4036 = ~n2414 & ~n2505;
  assign n4037 = n2845 & ~n4036;
  assign n4038 = n4037 ^ n1056;
  assign n4039 = ~n2414 & n2505;
  assign n4040 = n2970 & n4039;
  assign n4041 = n4040 ^ n1056;
  assign n4042 = n1056 & ~n4041;
  assign n4043 = n4042 ^ n1056;
  assign n4044 = n4038 & n4043;
  assign n4045 = n4044 ^ n4042;
  assign n4046 = n4045 ^ n1056;
  assign n4047 = n4046 ^ n4040;
  assign n4048 = ~n4035 & ~n4047;
  assign n4049 = n4048 ^ n4040;
  assign n4050 = ~n4034 & ~n4049;
  assign n4066 = n4065 ^ n4050;
  assign n3996 = n3166 ^ n1097;
  assign n3997 = n2602 & n3996;
  assign n3998 = ~n1101 & ~n2603;
  assign n3999 = ~n1101 & ~n2462;
  assign n4000 = ~n1097 & n3999;
  assign n4001 = ~n3998 & ~n4000;
  assign n4002 = ~n3997 & ~n4001;
  assign n4003 = ~n1097 & n2603;
  assign n4004 = n3166 & n4003;
  assign n4005 = n1097 & n2602;
  assign n4006 = ~n2462 & n4005;
  assign n4007 = n1101 & ~n4006;
  assign n4008 = ~n4004 & n4007;
  assign n4009 = ~n4002 & ~n4008;
  assign n4010 = n1097 & ~n3166;
  assign n4011 = n2603 & n4010;
  assign n4012 = ~n4009 & ~n4011;
  assign n4013 = ~n1836 & n3238;
  assign n4014 = n4013 ^ n1097;
  assign n4015 = n4014 ^ n3235;
  assign n4016 = n2598 & ~n4015;
  assign n4017 = n4012 & ~n4016;
  assign n3974 = n2434 ^ n850;
  assign n3975 = n2522 & n2870;
  assign n3976 = ~n3974 & n3975;
  assign n3977 = n2473 & n2528;
  assign n3978 = ~n2439 & n2535;
  assign n3979 = ~n3977 & ~n3978;
  assign n3980 = n3979 ^ n684;
  assign n3981 = n2522 & ~n2871;
  assign n3982 = n3981 ^ n684;
  assign n3983 = n2777 & n2875;
  assign n3984 = n3983 ^ n684;
  assign n3985 = ~n684 & n3984;
  assign n3986 = n3985 ^ n684;
  assign n3987 = ~n3982 & ~n3986;
  assign n3988 = n3987 ^ n3985;
  assign n3989 = n3988 ^ n684;
  assign n3990 = n3989 ^ n3983;
  assign n3991 = n3980 & n3990;
  assign n3992 = n3991 ^ n3983;
  assign n3993 = ~n3976 & ~n3992;
  assign n3968 = n3817 ^ n3813;
  assign n3969 = n3818 & n3968;
  assign n3970 = n3969 ^ n2444;
  assign n3971 = n3970 ^ n2443;
  assign n3972 = ~n551 & n3971;
  assign n3961 = n552 & n2599;
  assign n3962 = n3961 ^ n2440;
  assign n3963 = n685 & n3962;
  assign n3964 = ~n2441 & ~n2763;
  assign n3965 = n2442 & n2767;
  assign n3966 = ~n3964 & ~n3965;
  assign n3967 = ~n3963 & n3966;
  assign n3973 = n3972 ^ n3967;
  assign n3994 = n3993 ^ n3973;
  assign n3958 = n3820 ^ n3791;
  assign n3959 = n3841 & n3958;
  assign n3960 = n3959 ^ n3840;
  assign n3995 = n3994 ^ n3960;
  assign n4018 = n4017 ^ n3995;
  assign n3955 = n3842 ^ n3788;
  assign n3956 = n3857 & n3955;
  assign n3957 = n3956 ^ n3856;
  assign n4019 = n4018 ^ n3957;
  assign n3952 = n3874 ^ n3785;
  assign n3953 = ~n3875 & n3952;
  assign n3954 = n3953 ^ n3785;
  assign n4020 = n4019 ^ n3954;
  assign n4067 = n4066 ^ n4020;
  assign n3949 = n3903 ^ n3782;
  assign n3950 = ~n3904 & n3949;
  assign n3951 = n3950 ^ n3782;
  assign n4068 = n4067 ^ n3951;
  assign n4069 = n184 & n249;
  assign n4070 = n139 & ~n4069;
  assign n4071 = ~n1963 & ~n4070;
  assign n4072 = ~n226 & ~n938;
  assign n4073 = n4071 & n4072;
  assign n4074 = ~n309 & ~n344;
  assign n4075 = n640 & n4074;
  assign n4076 = n4073 & n4075;
  assign n4077 = ~n377 & ~n429;
  assign n4078 = n156 & n235;
  assign n4079 = n175 & ~n4078;
  assign n4080 = ~n281 & ~n438;
  assign n4081 = ~n4079 & n4080;
  assign n4082 = n4077 & n4081;
  assign n4083 = n4076 & n4082;
  assign n4084 = n752 & n4083;
  assign n4085 = n3649 & n4084;
  assign n4086 = ~n4068 & n4085;
  assign n4087 = n3927 ^ n3779;
  assign n4088 = n4087 ^ n3779;
  assign n4089 = n3918 ^ n3779;
  assign n4090 = n4089 ^ n3779;
  assign n4091 = ~n4088 & ~n4090;
  assign n4092 = n4091 ^ n3779;
  assign n4093 = ~n3906 & ~n4092;
  assign n4094 = n4093 ^ n3905;
  assign n4095 = n4086 & ~n4094;
  assign n4096 = n4094 ^ n4068;
  assign n4097 = n4085 ^ n4068;
  assign n4098 = n4096 & n4097;
  assign n4099 = n4098 ^ n4094;
  assign n4100 = ~n4095 & ~n4099;
  assign n4101 = n4068 & ~n4085;
  assign n4102 = n4094 & n4101;
  assign n4103 = ~n4100 & ~n4102;
  assign n4104 = n4103 ^ n3947;
  assign n4105 = n4104 ^ n3939;
  assign n4106 = n4105 ^ n4104;
  assign n4107 = n4104 ^ n3907;
  assign n4108 = ~n4106 & n4107;
  assign n4109 = n4108 ^ n4104;
  assign n4110 = ~n3948 & n4109;
  assign n4111 = n4110 ^ n4104;
  assign n4268 = n3907 & ~n3939;
  assign n4269 = n4099 & n4268;
  assign n4270 = n3939 & n4095;
  assign n4271 = ~n4269 & ~n4270;
  assign n4272 = ~n3907 & ~n3947;
  assign n4273 = n4102 & ~n4272;
  assign n4274 = n4271 & ~n4273;
  assign n4275 = ~n3907 & ~n4099;
  assign n4276 = n3947 & ~n4095;
  assign n4277 = n4275 & ~n4276;
  assign n4278 = n4274 & ~n4277;
  assign n4248 = n3954 & ~n4019;
  assign n4249 = n4065 ^ n3951;
  assign n4250 = n4066 & n4249;
  assign n4251 = n4250 ^ n3951;
  assign n4252 = n4248 & n4251;
  assign n4253 = n4050 & ~n4065;
  assign n4254 = ~n4248 & n4253;
  assign n4255 = ~n3951 & n4254;
  assign n4258 = ~n3954 & n4019;
  assign n4256 = ~n4050 & n4065;
  assign n4257 = n3951 & n4256;
  assign n4259 = n4258 ^ n4257;
  assign n4260 = n4259 ^ n4257;
  assign n4261 = n4257 ^ n4251;
  assign n4262 = n4260 & ~n4261;
  assign n4263 = n4262 ^ n4257;
  assign n4264 = ~n4255 & ~n4263;
  assign n4265 = ~n4252 & n4264;
  assign n4223 = ~n3895 & ~n3897;
  assign n4224 = x1 & n4223;
  assign n4225 = x2 & n3897;
  assign n4226 = ~n4224 & ~n4225;
  assign n4227 = n2426 & ~n4226;
  assign n4228 = ~x2 & ~x22;
  assign n4229 = n2416 & n4228;
  assign n4230 = x2 & x22;
  assign n4231 = n4230 ^ n3895;
  assign n4232 = n4230 ^ n2419;
  assign n4233 = n4232 ^ n2419;
  assign n4234 = n2419 ^ x1;
  assign n4235 = n4233 & ~n4234;
  assign n4236 = n4235 ^ n2419;
  assign n4237 = n4231 & ~n4236;
  assign n4238 = n4237 ^ n3895;
  assign n4239 = ~n4229 & ~n4238;
  assign n4240 = ~n4227 & n4239;
  assign n4241 = n4223 ^ x2;
  assign n4242 = n4241 ^ x2;
  assign n4243 = n320 & n4242;
  assign n4244 = n4243 ^ x2;
  assign n4245 = n2509 & ~n4244;
  assign n4246 = n4240 & ~n4245;
  assign n4191 = n2414 & n2820;
  assign n4192 = ~n2417 & n2832;
  assign n4193 = ~n4191 & ~n4192;
  assign n4194 = ~n1056 & ~n1157;
  assign n4195 = n2821 & ~n4194;
  assign n4196 = n3867 ^ n2417;
  assign n4197 = n2417 ^ n2414;
  assign n4198 = n4196 & ~n4197;
  assign n4199 = n4198 ^ n2417;
  assign n4200 = n4195 & ~n4199;
  assign n4201 = n4193 & ~n4200;
  assign n4202 = ~n1056 & n4201;
  assign n4203 = n2895 & n3632;
  assign n4204 = ~n4202 & ~n4203;
  assign n4205 = n1157 & n3632;
  assign n4206 = n3629 & ~n4205;
  assign n4207 = ~n4204 & n4206;
  assign n4208 = n2970 & ~n3629;
  assign n4209 = n3632 & n4208;
  assign n4210 = n1056 & ~n4201;
  assign n4211 = ~n4209 & ~n4210;
  assign n4212 = ~n4207 & n4211;
  assign n4213 = n2845 ^ n1056;
  assign n4214 = ~n3629 & ~n3632;
  assign n4215 = n4214 ^ n4201;
  assign n4216 = n4214 ^ n2845;
  assign n4217 = n4216 ^ n4214;
  assign n4218 = n4215 & ~n4217;
  assign n4219 = n4218 ^ n4214;
  assign n4220 = ~n4213 & n4219;
  assign n4221 = n4212 & ~n4220;
  assign n4166 = ~n1836 & n3284;
  assign n4167 = n4166 ^ n1097;
  assign n4168 = n4167 ^ n2420;
  assign n4169 = n2598 & n4168;
  assign n4170 = ~n1097 & n2602;
  assign n4171 = n3235 & n4170;
  assign n4172 = n4010 ^ n1061;
  assign n4173 = n4172 ^ n4010;
  assign n4174 = n3235 ^ n1097;
  assign n4175 = n4174 ^ n4010;
  assign n4176 = n4173 & ~n4175;
  assign n4177 = n4176 ^ n4010;
  assign n4178 = ~n2598 & ~n4177;
  assign n4179 = n4178 ^ n1101;
  assign n4180 = n4179 ^ n4178;
  assign n4181 = ~n3235 & n4005;
  assign n4182 = ~n3166 & n4003;
  assign n4183 = ~n4181 & ~n4182;
  assign n4184 = n4183 ^ n4178;
  assign n4185 = ~n4180 & ~n4184;
  assign n4186 = n4185 ^ n4178;
  assign n4187 = ~n4171 & ~n4186;
  assign n4188 = ~n4169 & n4187;
  assign n4147 = n2522 & n3593;
  assign n4148 = n2434 & n2528;
  assign n4149 = n2473 & n2535;
  assign n4150 = ~n4148 & ~n4149;
  assign n4151 = ~n4147 & n4150;
  assign n4152 = ~n684 & ~n4151;
  assign n4153 = n2522 & ~n3600;
  assign n4154 = n684 & n4150;
  assign n4155 = ~n4153 & n4154;
  assign n4156 = n2785 ^ n2462;
  assign n4157 = n4156 ^ n2785;
  assign n4158 = ~n2524 & n2527;
  assign n4159 = n4158 ^ n2785;
  assign n4160 = ~n4157 & n4159;
  assign n4161 = n4160 ^ n2785;
  assign n4162 = n2846 & n4161;
  assign n4163 = ~n4155 & ~n4162;
  assign n4164 = ~n4152 & n4163;
  assign n4137 = n3967 ^ n2443;
  assign n4138 = ~n3971 & ~n4137;
  assign n4139 = n4138 ^ n2443;
  assign n4140 = ~n551 & ~n4139;
  assign n4141 = ~n2442 & ~n4140;
  assign n4142 = ~n551 & n4141;
  assign n4143 = n2442 & n4140;
  assign n4144 = ~n4142 & ~n4143;
  assign n4130 = n552 & n2800;
  assign n4131 = n4130 ^ n2439;
  assign n4132 = n685 & ~n4131;
  assign n4133 = n2440 & ~n2763;
  assign n4134 = ~n2441 & n2767;
  assign n4135 = ~n4133 & ~n4134;
  assign n4136 = ~n4132 & n4135;
  assign n4145 = n4144 ^ n4136;
  assign n4127 = n3973 ^ n3960;
  assign n4128 = ~n3994 & n4127;
  assign n4129 = n4128 ^ n3993;
  assign n4146 = n4145 ^ n4129;
  assign n4165 = n4164 ^ n4146;
  assign n4189 = n4188 ^ n4165;
  assign n4124 = n4017 ^ n3957;
  assign n4125 = ~n4018 & n4124;
  assign n4126 = n4125 ^ n3957;
  assign n4190 = n4189 ^ n4126;
  assign n4222 = n4221 ^ n4190;
  assign n4247 = n4246 ^ n4222;
  assign n4266 = n4265 ^ n4247;
  assign n4112 = n353 & n3768;
  assign n4113 = ~n138 & ~n303;
  assign n4114 = n4112 & n4113;
  assign n4115 = ~n374 & ~n624;
  assign n4116 = ~n1026 & n4115;
  assign n4117 = n1046 & n4116;
  assign n4118 = n4114 & n4117;
  assign n4119 = n457 & n4118;
  assign n4120 = n560 & n3695;
  assign n4121 = n802 & n4120;
  assign n4122 = n4119 & n4121;
  assign n4123 = n1065 & n4122;
  assign n4267 = n4266 ^ n4123;
  assign n4279 = n4278 ^ n4267;
  assign n4286 = n4123 & n4266;
  assign n4287 = n4099 & ~n4286;
  assign n4288 = ~n4123 & ~n4266;
  assign n4289 = n3939 & ~n4102;
  assign n4290 = ~n4288 & n4289;
  assign n4291 = n4287 & n4290;
  assign n4292 = ~n4267 & n4270;
  assign n4293 = ~n4291 & ~n4292;
  assign n4280 = n4102 ^ n4100;
  assign n4281 = n4267 ^ n4102;
  assign n4282 = n4281 ^ n4102;
  assign n4283 = n4280 & n4282;
  assign n4284 = n4283 ^ n4102;
  assign n4285 = n3947 & n4284;
  assign n4294 = n4293 ^ n4285;
  assign n4295 = ~n4287 & ~n4288;
  assign n4383 = n4247 & ~n4257;
  assign n4384 = ~n4255 & ~n4258;
  assign n4385 = ~n4383 & n4384;
  assign n4386 = n4247 & ~n4248;
  assign n4387 = n4251 & ~n4386;
  assign n4388 = ~n4385 & ~n4387;
  assign n4378 = ~n4190 & ~n4221;
  assign n4379 = ~n4246 & ~n4378;
  assign n4380 = n4190 & n4221;
  assign n4381 = ~n4379 & ~n4380;
  assign n4356 = n3895 & ~n3898;
  assign n4357 = n2845 & ~n4356;
  assign n4358 = n1157 & ~n2414;
  assign n4359 = n2820 & ~n3629;
  assign n4360 = ~n2832 & ~n4359;
  assign n4361 = ~n4358 & ~n4360;
  assign n4362 = n2822 & ~n3629;
  assign n4363 = ~n4361 & ~n4362;
  assign n4364 = n2414 & n2830;
  assign n4365 = n1056 & ~n4364;
  assign n4366 = n4363 & n4365;
  assign n4367 = ~n4357 & n4366;
  assign n4368 = ~n3895 & ~n3898;
  assign n4369 = n2874 & n4368;
  assign n4370 = n3895 ^ n1157;
  assign n4371 = n2845 & ~n4370;
  assign n4372 = n3898 & n4371;
  assign n4373 = ~n1056 & ~n4363;
  assign n4374 = ~n4372 & ~n4373;
  assign n4375 = ~n4369 & n4374;
  assign n4376 = ~n4367 & n4375;
  assign n4340 = n2598 & n3859;
  assign n4341 = ~n2420 & n2606;
  assign n4342 = n2610 & ~n3235;
  assign n4343 = ~n4341 & ~n4342;
  assign n4344 = ~n4340 & n4343;
  assign n4345 = n1097 & ~n4344;
  assign n4346 = n2598 & ~n3870;
  assign n4347 = ~n1097 & n4343;
  assign n4348 = ~n4346 & n4347;
  assign n4349 = n2598 & n3270;
  assign n4350 = n2417 ^ n1101;
  assign n4351 = n4349 & ~n4350;
  assign n4352 = ~n4348 & ~n4351;
  assign n4353 = ~n4345 & n4352;
  assign n4323 = n3166 ^ n850;
  assign n4324 = n2522 & ~n4323;
  assign n4325 = n3165 & n4324;
  assign n4326 = n2462 & n2528;
  assign n4327 = n2434 & n2535;
  assign n4328 = ~n4326 & ~n4327;
  assign n4329 = n684 & ~n4328;
  assign n4330 = ~n4325 & ~n4329;
  assign n4331 = n2777 & n3171;
  assign n4332 = n4330 & ~n4331;
  assign n4333 = n2522 & ~n3175;
  assign n4334 = ~n684 & n4328;
  assign n4335 = ~n4333 & n4334;
  assign n4336 = n4332 & ~n4335;
  assign n4308 = n685 & n2894;
  assign n4309 = ~n2439 & ~n2763;
  assign n4310 = n2440 & n2767;
  assign n4311 = ~n4309 & ~n4310;
  assign n4312 = ~n4308 & n4311;
  assign n4313 = ~n551 & ~n4312;
  assign n4314 = n685 & ~n2910;
  assign n4315 = n551 & n4311;
  assign n4316 = ~n4314 & n4315;
  assign n4317 = n2473 ^ n543;
  assign n4318 = n685 & n2893;
  assign n4319 = n4317 & n4318;
  assign n4320 = ~n4316 & ~n4319;
  assign n4321 = ~n4313 & n4320;
  assign n4322 = n4321 ^ n2511;
  assign n4337 = n4336 ^ n4322;
  assign n4302 = n4140 ^ n2442;
  assign n4303 = n4140 ^ n4136;
  assign n4304 = n4302 & ~n4303;
  assign n4305 = n4304 ^ n2442;
  assign n4306 = n4305 ^ n2441;
  assign n4307 = ~n551 & ~n4306;
  assign n4338 = n4337 ^ n4307;
  assign n4299 = n4164 ^ n4129;
  assign n4300 = ~n4146 & ~n4299;
  assign n4301 = n4300 ^ n4164;
  assign n4339 = n4338 ^ n4301;
  assign n4354 = n4353 ^ n4339;
  assign n4296 = n4165 ^ n4126;
  assign n4297 = ~n4189 & ~n4296;
  assign n4298 = n4297 ^ n4188;
  assign n4355 = n4354 ^ n4298;
  assign n4377 = n4376 ^ n4355;
  assign n4382 = n4381 ^ n4377;
  assign n4389 = n4388 ^ n4382;
  assign n4390 = n759 & n1041;
  assign n4391 = ~n92 & n2311;
  assign n4392 = n4390 & n4391;
  assign n4393 = n162 & ~n369;
  assign n4394 = n671 & ~n4393;
  assign n4395 = n4392 & n4394;
  assign n4396 = n1137 & n4395;
  assign n4397 = n2185 & n4396;
  assign n4398 = n834 & n4397;
  assign n4399 = ~n4389 & n4398;
  assign n4400 = ~n4295 & ~n4399;
  assign n4401 = n4389 & ~n4398;
  assign n4402 = ~n4400 & ~n4401;
  assign n4403 = ~n4295 & n4401;
  assign n4404 = ~n4402 & ~n4403;
  assign n4405 = n4295 & n4399;
  assign n4406 = ~n4404 & ~n4405;
  assign n4407 = n4406 ^ n4285;
  assign n4408 = n4407 ^ n4293;
  assign n4409 = n4408 ^ n4407;
  assign n4410 = n4407 ^ n3907;
  assign n4411 = n4409 & ~n4410;
  assign n4412 = n4411 ^ n4407;
  assign n4413 = n4294 & ~n4412;
  assign n4414 = n4413 ^ n4407;
  assign n4565 = ~n4376 & ~n4381;
  assign n4566 = n4388 & ~n4565;
  assign n4567 = ~n4298 & n4354;
  assign n4568 = n4298 & ~n4354;
  assign n4569 = n4376 & ~n4568;
  assign n4570 = n4381 & n4569;
  assign n4571 = ~n4567 & ~n4570;
  assign n4572 = n4566 & ~n4571;
  assign n4573 = ~n4567 & ~n4569;
  assign n4574 = ~n4376 & n4568;
  assign n4575 = n4573 & ~n4574;
  assign n4576 = ~n4381 & n4575;
  assign n4577 = n4576 ^ n4574;
  assign n4578 = ~n4388 & n4577;
  assign n4579 = n4376 & n4567;
  assign n4580 = n4579 ^ n4574;
  assign n4581 = n4381 & n4580;
  assign n4582 = n4581 ^ n4574;
  assign n4583 = ~n4578 & ~n4582;
  assign n4584 = ~n4572 & n4583;
  assign n4547 = ~n2823 & ~n3895;
  assign n4548 = n2832 & ~n3629;
  assign n4549 = ~n4547 & ~n4548;
  assign n4550 = ~n1056 & ~n4549;
  assign n4551 = n1056 & ~n4547;
  assign n4552 = ~n1157 & ~n2511;
  assign n4553 = ~n3629 & n4552;
  assign n4554 = n4551 & ~n4553;
  assign n4555 = ~n2845 & ~n4554;
  assign n4556 = ~n2819 & n2899;
  assign n4557 = n4556 ^ n4058;
  assign n4558 = n4557 ^ n4556;
  assign n4559 = n4556 ^ n4551;
  assign n4560 = ~n4558 & ~n4559;
  assign n4561 = n4560 ^ n4556;
  assign n4562 = ~n4555 & ~n4561;
  assign n4563 = ~n4550 & ~n4562;
  assign n4530 = n2414 & ~n2505;
  assign n4531 = n2598 & n4530;
  assign n4532 = ~n2417 & n2606;
  assign n4533 = ~n2420 & n2610;
  assign n4534 = ~n4532 & ~n4533;
  assign n4535 = ~n4531 & n4534;
  assign n4536 = ~n1097 & ~n4535;
  assign n4537 = n2598 & ~n4036;
  assign n4538 = n1097 & n4534;
  assign n4539 = ~n4537 & n4538;
  assign n4540 = n2414 ^ n1101;
  assign n4541 = n2598 & ~n4540;
  assign n4542 = n2505 & n4541;
  assign n4543 = ~n4539 & ~n4542;
  assign n4544 = ~n4536 & n4543;
  assign n4489 = ~n551 & ~n2441;
  assign n4519 = n4322 & n4336;
  assign n4520 = ~n4489 & n4519;
  assign n4521 = n4322 ^ n2441;
  assign n4522 = n4305 & ~n4521;
  assign n4523 = ~n4336 & ~n4522;
  assign n4524 = ~n2441 & ~n4322;
  assign n4525 = ~n4305 & ~n4524;
  assign n4526 = ~n551 & ~n4525;
  assign n4527 = ~n4523 & n4526;
  assign n4528 = ~n4520 & ~n4527;
  assign n4495 = n2528 & n3166;
  assign n4496 = n2462 & n2535;
  assign n4497 = ~n4495 & ~n4496;
  assign n4498 = n684 & n4497;
  assign n4499 = n3235 ^ n850;
  assign n4500 = n4499 ^ n3235;
  assign n4501 = n3239 ^ n3235;
  assign n4502 = ~n4500 & n4501;
  assign n4503 = n4502 ^ n3235;
  assign n4504 = n2522 & ~n4503;
  assign n4505 = n4498 & ~n4504;
  assign n4506 = n850 & n3238;
  assign n4507 = ~n684 & ~n3235;
  assign n4508 = n2522 & n4507;
  assign n4509 = ~n4506 & n4508;
  assign n4510 = ~n684 & ~n4497;
  assign n4511 = ~n684 & n850;
  assign n4512 = n2522 & n4511;
  assign n4513 = n3235 & n4512;
  assign n4514 = n3238 & n4513;
  assign n4515 = ~n4510 & ~n4514;
  assign n4516 = ~n4509 & n4515;
  assign n4517 = ~n4505 & n4516;
  assign n4479 = ~n2511 & n4321;
  assign n4480 = ~n2441 & n4479;
  assign n4481 = ~n551 & n2440;
  assign n4482 = ~n4480 & n4481;
  assign n4483 = n2511 & ~n4321;
  assign n4484 = n2441 & n4483;
  assign n4485 = n4482 & ~n4484;
  assign n4486 = n551 & n4483;
  assign n4487 = ~n4485 & ~n4486;
  assign n4488 = ~n2440 & n4484;
  assign n4490 = ~n2440 & n4489;
  assign n4491 = n4479 & n4490;
  assign n4492 = ~n4488 & ~n4491;
  assign n4493 = n4487 & n4492;
  assign n4449 = n2473 ^ n551;
  assign n4450 = n4449 ^ n2473;
  assign n4451 = ~n2855 & n4450;
  assign n4452 = n4451 ^ n2473;
  assign n4453 = ~n543 & n4452;
  assign n4454 = n4453 ^ n2473;
  assign n4455 = n2569 & n4454;
  assign n4456 = ~n543 & ~n2473;
  assign n4457 = ~n2439 & n2753;
  assign n4458 = ~n2762 & ~n4457;
  assign n4459 = ~n4456 & ~n4458;
  assign n4460 = ~n4455 & ~n4459;
  assign n4461 = n4460 ^ n551;
  assign n4462 = n685 & ~n2871;
  assign n4463 = n4462 ^ n551;
  assign n4464 = n551 & n685;
  assign n4465 = n2875 & n4464;
  assign n4466 = n2434 ^ n543;
  assign n4467 = n685 & n2870;
  assign n4468 = ~n4466 & n4467;
  assign n4469 = ~n4465 & ~n4468;
  assign n4470 = n4469 ^ n551;
  assign n4471 = ~n551 & ~n4470;
  assign n4472 = n4471 ^ n551;
  assign n4473 = ~n4463 & ~n4472;
  assign n4474 = n4473 ^ n4471;
  assign n4475 = n4474 ^ n551;
  assign n4476 = n4475 ^ n4469;
  assign n4477 = n4461 & ~n4476;
  assign n4478 = n4477 ^ n4469;
  assign n4494 = n4493 ^ n4478;
  assign n4518 = n4517 ^ n4494;
  assign n4529 = n4528 ^ n4518;
  assign n4545 = n4544 ^ n4529;
  assign n4446 = n4353 ^ n4338;
  assign n4447 = n4339 & n4446;
  assign n4448 = n4447 ^ n4353;
  assign n4546 = n4545 ^ n4448;
  assign n4564 = n4563 ^ n4546;
  assign n4585 = n4584 ^ n4564;
  assign n4430 = ~n51 & n137;
  assign n4431 = ~n85 & n156;
  assign n4432 = ~n4430 & ~n4431;
  assign n4433 = ~n243 & ~n4432;
  assign n4434 = ~n174 & n229;
  assign n4435 = ~n324 & n4434;
  assign n4436 = ~n486 & ~n4435;
  assign n4437 = n4433 & ~n4436;
  assign n4438 = n2068 & n4437;
  assign n4439 = ~n296 & n940;
  assign n4440 = n240 & n3736;
  assign n4441 = n4439 & n4440;
  assign n4442 = n4438 & n4441;
  assign n4443 = n3892 & n4442;
  assign n4444 = n3778 & n4443;
  assign n4445 = n2363 & n4444;
  assign n4586 = n4585 ^ n4445;
  assign n4415 = n3907 & n4293;
  assign n4416 = n4415 ^ n4402;
  assign n4417 = ~n3907 & ~n4285;
  assign n4418 = ~n4405 & ~n4417;
  assign n4419 = n4418 ^ n4402;
  assign n4420 = n4403 & ~n4417;
  assign n4421 = n4420 ^ n4402;
  assign n4422 = n4402 & ~n4421;
  assign n4423 = n4422 ^ n4402;
  assign n4424 = n4419 & n4423;
  assign n4425 = n4424 ^ n4422;
  assign n4426 = n4425 ^ n4402;
  assign n4427 = n4426 ^ n4420;
  assign n4428 = n4416 & ~n4427;
  assign n4429 = n4428 ^ n4420;
  assign n4587 = n4586 ^ n4429;
  assign n4713 = n4405 ^ n4404;
  assign n4714 = n4586 & n4713;
  assign n4715 = n4714 ^ n4404;
  assign n4716 = ~n4293 & n4715;
  assign n4717 = n3907 & ~n4716;
  assign n4718 = n4400 & ~n4586;
  assign n4719 = n4285 & ~n4405;
  assign n4720 = ~n4718 & n4719;
  assign n4721 = n4586 ^ n4295;
  assign n4722 = ~n4401 & n4721;
  assign n4723 = n4722 ^ n4295;
  assign n4724 = n4720 & ~n4723;
  assign n4725 = ~n4717 & ~n4724;
  assign n4698 = n4564 & ~n4570;
  assign n4699 = n4388 & ~n4698;
  assign n4700 = ~n4564 & ~n4565;
  assign n4701 = ~n4567 & ~n4700;
  assign n4702 = ~n4699 & n4701;
  assign n4703 = ~n4564 & ~n4568;
  assign n4704 = n4388 ^ n4381;
  assign n4705 = n4388 ^ n4376;
  assign n4706 = n4704 & n4705;
  assign n4707 = n4706 ^ n4388;
  assign n4708 = ~n4703 & ~n4707;
  assign n4709 = ~n4702 & ~n4708;
  assign n4683 = n3897 ^ n1056;
  assign n4684 = n4683 ^ n1056;
  assign n4685 = ~n1157 & ~n3895;
  assign n4686 = n4685 ^ n1056;
  assign n4687 = ~n4684 & ~n4686;
  assign n4688 = n4687 ^ n1056;
  assign n4689 = ~n2819 & ~n4688;
  assign n4690 = n2821 ^ n1157;
  assign n4691 = n2821 ^ n1056;
  assign n4692 = n4690 & ~n4691;
  assign n4693 = ~n3895 & n4692;
  assign n4694 = n4693 ^ n1056;
  assign n4695 = ~n4689 & n4694;
  assign n4680 = n4563 ^ n4545;
  assign n4681 = n4546 & n4680;
  assign n4682 = n4681 ^ n4563;
  assign n4696 = n4695 ^ n4682;
  assign n4663 = n2598 & n4214;
  assign n4664 = n2414 & n2606;
  assign n4665 = ~n2417 & n2610;
  assign n4666 = ~n4664 & ~n4665;
  assign n4667 = ~n4663 & n4666;
  assign n4668 = ~n1097 & ~n4667;
  assign n4669 = n3629 & ~n3632;
  assign n4670 = n2598 & ~n4669;
  assign n4671 = n1097 & n4666;
  assign n4672 = ~n4670 & n4671;
  assign n4673 = n3629 ^ n1101;
  assign n4674 = n2598 & n4673;
  assign n4675 = n3632 & n4674;
  assign n4676 = ~n4672 & ~n4675;
  assign n4677 = ~n4668 & n4676;
  assign n4646 = ~n2420 & n2522;
  assign n4647 = ~n3284 & n4646;
  assign n4648 = n2528 & ~n3235;
  assign n4649 = n2535 & n3166;
  assign n4650 = ~n4648 & ~n4649;
  assign n4651 = ~n4647 & n4650;
  assign n4652 = ~n684 & ~n4651;
  assign n4653 = n2522 & n3284;
  assign n4655 = n684 & n4650;
  assign n4656 = ~n4646 & n4655;
  assign n4654 = n2420 ^ n850;
  assign n4657 = n4656 ^ n4654;
  assign n4658 = n4653 & ~n4657;
  assign n4659 = n4658 ^ n4656;
  assign n4660 = ~n4652 & ~n4659;
  assign n4632 = n4480 & n4481;
  assign n4633 = ~n4488 & ~n4632;
  assign n4634 = n2439 & ~n4633;
  assign n4635 = n2440 & ~n2441;
  assign n4636 = n4321 & n4635;
  assign n4637 = ~n551 & ~n2439;
  assign n4638 = ~n4636 & n4637;
  assign n4639 = ~n4488 & n4638;
  assign n4640 = n2511 & n4481;
  assign n4641 = ~n2439 & n4640;
  assign n4642 = ~n4486 & ~n4641;
  assign n4643 = ~n4639 & n4642;
  assign n4644 = ~n4634 & n4643;
  assign n4615 = ~n551 & n2434;
  assign n4616 = n2762 & n4615;
  assign n4617 = n2765 & n4456;
  assign n4618 = ~n551 & ~n2473;
  assign n4619 = n2326 & ~n4618;
  assign n4620 = ~n4617 & ~n4619;
  assign n4621 = ~n4616 & n4620;
  assign n4622 = n2434 ^ n551;
  assign n4623 = n551 & n1938;
  assign n4624 = ~n2761 & ~n4623;
  assign n4625 = n4622 & ~n4624;
  assign n4626 = n4621 & ~n4625;
  assign n4627 = n552 & ~n2846;
  assign n4628 = n4627 ^ n543;
  assign n4629 = n4628 ^ n2462;
  assign n4630 = n685 & n4629;
  assign n4631 = n4626 & ~n4630;
  assign n4645 = n4644 ^ n4631;
  assign n4661 = n4660 ^ n4645;
  assign n4612 = n4517 ^ n4493;
  assign n4613 = ~n4494 & n4612;
  assign n4614 = n4613 ^ n4517;
  assign n4662 = n4661 ^ n4614;
  assign n4678 = n4677 ^ n4662;
  assign n4609 = n4544 ^ n4528;
  assign n4610 = ~n4529 & n4609;
  assign n4611 = n4610 ^ n4544;
  assign n4679 = n4678 ^ n4611;
  assign n4697 = n4696 ^ n4679;
  assign n4710 = n4709 ^ n4697;
  assign n4591 = ~n50 & ~n151;
  assign n4592 = n249 & ~n4591;
  assign n4593 = ~n205 & ~n4592;
  assign n4594 = n3768 & ~n4593;
  assign n4595 = n3773 & n4594;
  assign n4596 = n240 & ~n583;
  assign n4597 = n448 & n4596;
  assign n4598 = n2259 & n4597;
  assign n4599 = n4595 & n4598;
  assign n4600 = ~n191 & ~n625;
  assign n4601 = n349 & n4600;
  assign n4602 = n458 & n4601;
  assign n4603 = ~n250 & ~n288;
  assign n4604 = n2392 & n4603;
  assign n4605 = n4602 & n4604;
  assign n4606 = n4599 & n4605;
  assign n4607 = n2175 & n4606;
  assign n4608 = n3734 & n4607;
  assign n4711 = n4710 ^ n4608;
  assign n4588 = n4585 ^ n4402;
  assign n4589 = n4586 & ~n4588;
  assign n4590 = n4589 ^ n4402;
  assign n4712 = n4711 ^ n4590;
  assign n4726 = n4725 ^ n4712;
  assign n4838 = n4716 & ~n4724;
  assign n4839 = n4712 & n4838;
  assign n4840 = ~n4712 & n4724;
  assign n4841 = ~n3907 & ~n4840;
  assign n4842 = ~n4839 & ~n4841;
  assign n4826 = ~n150 & ~n3684;
  assign n4827 = ~n91 & n328;
  assign n4828 = n791 & ~n4827;
  assign n4829 = ~n365 & ~n820;
  assign n4830 = n4828 & ~n4829;
  assign n4831 = n2373 & n4433;
  assign n4832 = n4830 & n4831;
  assign n4833 = n4599 & n4832;
  assign n4834 = ~n4826 & n4833;
  assign n4835 = n1994 & n4834;
  assign n4794 = n2462 & ~n2763;
  assign n4795 = n2434 & n2767;
  assign n4796 = ~n4794 & ~n4795;
  assign n4797 = n552 & n3165;
  assign n4798 = n4797 ^ n3166;
  assign n4799 = n685 & n4798;
  assign n4800 = n4796 & ~n4799;
  assign n4801 = ~n2439 & ~n2511;
  assign n4802 = n4636 & n4801;
  assign n4803 = ~n2473 & n4802;
  assign n4804 = n551 & ~n4483;
  assign n4805 = ~n4803 & ~n4804;
  assign n4806 = n4800 & ~n4805;
  assign n4807 = ~n4481 & ~n4489;
  assign n4808 = ~n4637 & n4807;
  assign n4809 = ~n4321 & n4808;
  assign n4810 = n2511 & n4809;
  assign n4811 = n2473 & ~n4810;
  assign n4812 = n4811 ^ n4800;
  assign n4813 = n4812 ^ n4811;
  assign n4814 = ~n4618 & ~n4810;
  assign n4815 = n4814 ^ n4811;
  assign n4816 = ~n4813 & ~n4815;
  assign n4817 = n4816 ^ n4811;
  assign n4818 = ~n4802 & n4817;
  assign n4819 = ~n4806 & ~n4818;
  assign n4820 = n4819 ^ n1056;
  assign n4791 = n4660 ^ n4644;
  assign n4792 = n4645 & n4791;
  assign n4793 = n4792 ^ n4660;
  assign n4821 = n4820 ^ n4793;
  assign n4765 = ~n2420 & n2528;
  assign n4766 = n2535 & ~n3235;
  assign n4767 = ~n4765 & ~n4766;
  assign n4768 = ~n684 & n4767;
  assign n4769 = n3270 & n4768;
  assign n4770 = ~n2777 & ~n4769;
  assign n4771 = ~n850 & n3270;
  assign n4772 = ~n2417 & ~n4771;
  assign n4773 = ~n4770 & n4772;
  assign n4774 = n4767 ^ n684;
  assign n4775 = n2522 & ~n3870;
  assign n4776 = n4775 ^ n684;
  assign n4777 = n2366 & ~n2499;
  assign n4778 = ~n3270 & ~n4777;
  assign n4779 = n2417 & n2785;
  assign n4780 = ~n4778 & n4779;
  assign n4781 = n4780 ^ n684;
  assign n4782 = ~n684 & n4781;
  assign n4783 = n4782 ^ n684;
  assign n4784 = ~n4776 & ~n4783;
  assign n4785 = n4784 ^ n4782;
  assign n4786 = n4785 ^ n684;
  assign n4787 = n4786 ^ n4780;
  assign n4788 = n4774 & n4787;
  assign n4789 = n4788 ^ n4780;
  assign n4790 = ~n4773 & ~n4789;
  assign n4822 = n4821 ^ n4790;
  assign n4762 = n4677 ^ n4661;
  assign n4763 = n4662 & ~n4762;
  assign n4764 = n4763 ^ n4677;
  assign n4823 = n4822 ^ n4764;
  assign n4748 = n2598 & n4368;
  assign n4749 = n2414 & n2610;
  assign n4750 = n2606 & ~n3629;
  assign n4751 = ~n4749 & ~n4750;
  assign n4752 = ~n4748 & n4751;
  assign n4753 = n1097 & ~n4752;
  assign n4754 = n2598 & ~n4356;
  assign n4755 = ~n1097 & n4751;
  assign n4756 = ~n4754 & n4755;
  assign n4757 = n3895 ^ n1101;
  assign n4758 = n2598 & ~n4757;
  assign n4759 = n3898 & n4758;
  assign n4760 = ~n4756 & ~n4759;
  assign n4761 = ~n4753 & n4760;
  assign n4824 = n4823 ^ n4761;
  assign n4730 = n4611 & ~n4678;
  assign n4731 = ~n4695 & n4730;
  assign n4732 = ~n4611 & n4678;
  assign n4733 = n4695 & n4732;
  assign n4734 = ~n4731 & ~n4733;
  assign n4735 = n4696 & ~n4734;
  assign n4736 = ~n4695 & ~n4732;
  assign n4737 = ~n4730 & ~n4736;
  assign n4738 = ~n4682 & ~n4731;
  assign n4739 = ~n4737 & ~n4738;
  assign n4740 = n4739 ^ n4709;
  assign n4741 = n4740 ^ n4739;
  assign n4742 = ~n4682 & n4737;
  assign n4743 = ~n4733 & ~n4742;
  assign n4744 = n4743 ^ n4739;
  assign n4745 = ~n4741 & ~n4744;
  assign n4746 = n4745 ^ n4739;
  assign n4747 = ~n4735 & ~n4746;
  assign n4825 = n4824 ^ n4747;
  assign n4836 = n4835 ^ n4825;
  assign n4727 = n4710 ^ n4590;
  assign n4728 = ~n4711 & n4727;
  assign n4729 = n4728 ^ n4590;
  assign n4837 = n4836 ^ n4729;
  assign n4843 = n4842 ^ n4837;
  assign n4946 = ~n4732 & ~n4824;
  assign n4947 = n4709 ^ n4682;
  assign n4948 = n4696 & n4947;
  assign n4949 = n4948 ^ n4709;
  assign n4950 = ~n4946 & ~n4949;
  assign n4951 = n4682 & n4736;
  assign n4952 = n4824 & ~n4951;
  assign n4953 = n4709 & ~n4952;
  assign n4954 = ~n4682 & n4695;
  assign n4955 = ~n4824 & ~n4954;
  assign n4956 = ~n4730 & ~n4955;
  assign n4957 = ~n4953 & n4956;
  assign n4958 = ~n4950 & ~n4957;
  assign n4924 = ~n850 & n2414;
  assign n4925 = ~n4530 & ~n4924;
  assign n4926 = n2522 & ~n4925;
  assign n4927 = ~n2417 & n2528;
  assign n4928 = ~n2420 & n2535;
  assign n4929 = ~n4927 & ~n4928;
  assign n4930 = ~n4926 & n4929;
  assign n4931 = ~n684 & ~n4930;
  assign n4932 = n684 & n4929;
  assign n4933 = n2414 ^ n850;
  assign n4934 = n4933 ^ n2414;
  assign n4935 = n2506 ^ n2414;
  assign n4936 = ~n4934 & n4935;
  assign n4937 = n4936 ^ n2414;
  assign n4938 = n2522 & n4937;
  assign n4939 = n4932 & ~n4938;
  assign n4940 = n4039 & n4512;
  assign n4941 = ~n4939 & ~n4940;
  assign n4942 = ~n4931 & n4941;
  assign n4907 = n685 & ~n3235;
  assign n4908 = ~n3238 & n4907;
  assign n4909 = ~n2763 & n3166;
  assign n4910 = n2462 & n2767;
  assign n4911 = ~n4909 & ~n4910;
  assign n4912 = ~n4908 & n4911;
  assign n4913 = ~n551 & ~n4912;
  assign n4914 = n3235 ^ n543;
  assign n4915 = n685 & ~n4914;
  assign n4916 = n3238 & n4915;
  assign n4917 = ~n4913 & ~n4916;
  assign n4918 = n685 & ~n3247;
  assign n4919 = n551 & n4911;
  assign n4920 = ~n4918 & n4919;
  assign n4921 = n4917 & ~n4920;
  assign n4897 = n2511 ^ n1056;
  assign n4898 = n2511 ^ n551;
  assign n4899 = n4898 ^ n2511;
  assign n4900 = n2511 ^ n2473;
  assign n4901 = n4900 ^ n2511;
  assign n4902 = ~n4899 & n4901;
  assign n4903 = n4902 ^ n2511;
  assign n4904 = n4897 & n4903;
  assign n4905 = n4904 ^ n1056;
  assign n4906 = n4905 ^ n4615;
  assign n4922 = n4921 ^ n4906;
  assign n4871 = n4636 & n4637;
  assign n4872 = n2511 & ~n4809;
  assign n4873 = ~n4871 & ~n4872;
  assign n4874 = n551 & ~n4800;
  assign n4875 = ~n4873 & n4874;
  assign n4876 = n2473 & ~n2511;
  assign n4877 = n4800 & ~n4876;
  assign n4878 = n2473 & ~n4873;
  assign n4879 = ~n4877 & ~n4878;
  assign n4880 = ~n551 & ~n4879;
  assign n4881 = ~n4871 & ~n4874;
  assign n4882 = ~n2511 & ~n4881;
  assign n4883 = ~n4880 & ~n4882;
  assign n4884 = n4883 ^ n1056;
  assign n4885 = n4884 ^ n4883;
  assign n4886 = ~n2473 & ~n4873;
  assign n4887 = ~n4874 & ~n4886;
  assign n4888 = n2511 & ~n4887;
  assign n4889 = ~n551 & n4876;
  assign n4890 = n4873 & ~n4889;
  assign n4891 = n4800 & ~n4890;
  assign n4892 = ~n4888 & ~n4891;
  assign n4893 = n4892 ^ n4883;
  assign n4894 = ~n4885 & n4893;
  assign n4895 = n4894 ^ n4883;
  assign n4896 = ~n4875 & n4895;
  assign n4923 = n4922 ^ n4896;
  assign n4943 = n4942 ^ n4923;
  assign n4868 = n4822 ^ n4761;
  assign n4869 = n4823 & n4868;
  assign n4870 = n4869 ^ n4764;
  assign n4944 = n4943 ^ n4870;
  assign n4851 = n2606 & ~n3895;
  assign n4852 = n2610 & ~n3629;
  assign n4853 = ~n4851 & ~n4852;
  assign n4854 = n4853 ^ n1097;
  assign n4855 = n4854 ^ n1101;
  assign n4856 = n4854 ^ n4853;
  assign n4857 = n2598 & n4058;
  assign n4858 = n4857 ^ n4853;
  assign n4859 = ~n4853 & ~n4858;
  assign n4860 = n4859 ^ n4853;
  assign n4861 = ~n4856 & ~n4860;
  assign n4862 = n4861 ^ n4859;
  assign n4863 = n4862 ^ n4853;
  assign n4864 = n4863 ^ n4857;
  assign n4865 = n4855 & ~n4864;
  assign n4866 = n4865 ^ n4854;
  assign n4848 = n4820 ^ n4790;
  assign n4849 = ~n4821 & ~n4848;
  assign n4850 = n4849 ^ n4793;
  assign n4867 = n4866 ^ n4850;
  assign n4945 = n4944 ^ n4867;
  assign n4959 = n4958 ^ n4945;
  assign n4960 = n57 & ~n516;
  assign n4961 = n641 & ~n4960;
  assign n4962 = n78 & n369;
  assign n4963 = n85 & ~n4962;
  assign n4964 = n4961 & ~n4963;
  assign n4965 = n416 & n4964;
  assign n4966 = n3735 & n4965;
  assign n4967 = n349 & n664;
  assign n4968 = n2240 & n2352;
  assign n4969 = n4967 & n4968;
  assign n4970 = ~n156 & n175;
  assign n4971 = n56 & ~n97;
  assign n4972 = ~n4970 & ~n4971;
  assign n4973 = ~n2121 & n4972;
  assign n4974 = n1130 & n4973;
  assign n4975 = n4969 & n4974;
  assign n4976 = n4966 & n4975;
  assign n4977 = n3676 & n4976;
  assign n4978 = ~n4959 & n4977;
  assign n4979 = n4825 ^ n4729;
  assign n4980 = n4836 & ~n4979;
  assign n4981 = n4980 ^ n4729;
  assign n4982 = ~n4978 & ~n4981;
  assign n4983 = n4959 & ~n4977;
  assign n4984 = n4982 & ~n4983;
  assign n4985 = n4977 ^ n4959;
  assign n4986 = n4981 & n4985;
  assign n4987 = ~n4984 & ~n4986;
  assign n4844 = ~n4837 & n4839;
  assign n4845 = n3907 & ~n4844;
  assign n4846 = n4837 & n4840;
  assign n4847 = ~n4845 & ~n4846;
  assign n4988 = n4987 ^ n4847;
  assign n5081 = n4977 ^ n4845;
  assign n5082 = ~n3907 & ~n4846;
  assign n5083 = n4959 & ~n5082;
  assign n5084 = n5083 ^ n4977;
  assign n5085 = ~n5081 & ~n5084;
  assign n5086 = n5085 ^ n4977;
  assign n5087 = ~n4981 & ~n5086;
  assign n5088 = n5082 ^ n4845;
  assign n5089 = n5081 ^ n4845;
  assign n5090 = n5088 & n5089;
  assign n5091 = n5090 ^ n4845;
  assign n5092 = n4985 & n5091;
  assign n5093 = ~n5087 & ~n5092;
  assign n5094 = ~n4845 & n4978;
  assign n5095 = ~n4983 & n5082;
  assign n5096 = ~n5094 & ~n5095;
  assign n5097 = n4981 & ~n5096;
  assign n5098 = n5093 & ~n5097;
  assign n5062 = n4870 & ~n4943;
  assign n5063 = ~n4850 & ~n4866;
  assign n5069 = n5062 & ~n5063;
  assign n5065 = ~n4870 & n4943;
  assign n5066 = n4850 & n4866;
  assign n5070 = ~n5065 & n5066;
  assign n5071 = ~n5069 & ~n5070;
  assign n5064 = ~n5062 & n5063;
  assign n5067 = n5065 & ~n5066;
  assign n5068 = ~n5064 & ~n5067;
  assign n5072 = n5071 ^ n5068;
  assign n5073 = ~n4958 & n5072;
  assign n5074 = n5073 ^ n5071;
  assign n5075 = n4943 ^ n4866;
  assign n5076 = ~n4867 & n5075;
  assign n5077 = n4944 & n5076;
  assign n5078 = n5074 & ~n5077;
  assign n5045 = n2522 & n4214;
  assign n5046 = n2414 & n2528;
  assign n5047 = ~n2417 & n2535;
  assign n5048 = ~n5046 & ~n5047;
  assign n5049 = ~n5045 & n5048;
  assign n5050 = ~n684 & ~n5049;
  assign n5051 = n2522 & ~n4669;
  assign n5052 = n684 & n5048;
  assign n5053 = ~n5051 & n5052;
  assign n5054 = n3629 ^ n850;
  assign n5055 = n2522 & ~n5054;
  assign n5056 = n3632 & n5055;
  assign n5057 = ~n5053 & ~n5056;
  assign n5058 = ~n5050 & n5057;
  assign n5041 = n4921 ^ n4615;
  assign n5042 = n4921 ^ n4905;
  assign n5043 = ~n5041 & n5042;
  assign n5044 = n5043 ^ n4615;
  assign n5059 = n5058 ^ n5044;
  assign n5026 = n3098 & n3166;
  assign n5027 = n1938 & ~n5026;
  assign n5028 = n2761 & ~n3235;
  assign n5029 = n5028 ^ n2569;
  assign n5030 = ~n5027 & ~n5029;
  assign n5031 = n551 & n684;
  assign n5032 = n3166 & n5031;
  assign n5033 = ~n4507 & ~n5032;
  assign n5034 = ~n543 & ~n5033;
  assign n5035 = ~n5030 & ~n5034;
  assign n5036 = n552 & n3284;
  assign n5037 = n5036 ^ n2420;
  assign n5038 = n685 & n5037;
  assign n5039 = ~n5035 & ~n5038;
  assign n5022 = n2434 & ~n2462;
  assign n5023 = ~n551 & ~n5022;
  assign n5024 = ~n2434 & n2462;
  assign n5025 = n5023 & ~n5024;
  assign n5040 = n5039 ^ n5025;
  assign n5060 = n5059 ^ n5040;
  assign n5018 = n4942 ^ n4896;
  assign n5019 = n4923 & n5018;
  assign n5020 = n5019 ^ n4942;
  assign n4998 = n3897 ^ n1097;
  assign n4999 = n4998 ^ n1097;
  assign n5000 = n1101 & ~n3895;
  assign n5001 = n5000 ^ n1097;
  assign n5002 = ~n4999 & ~n5001;
  assign n5003 = n5002 ^ n1097;
  assign n5004 = ~n2603 & ~n5003;
  assign n5005 = ~n1097 & n1101;
  assign n5006 = ~n2602 & ~n5005;
  assign n5007 = n5006 ^ n1097;
  assign n5008 = n3895 ^ n1097;
  assign n5009 = n5008 ^ n1097;
  assign n5010 = n5007 & ~n5009;
  assign n5011 = n5010 ^ n1097;
  assign n5012 = n5004 ^ n2699;
  assign n5013 = n5011 & ~n5012;
  assign n5014 = n5013 ^ n2699;
  assign n5015 = ~n5004 & n5014;
  assign n5016 = n5015 ^ n5004;
  assign n5017 = n5016 ^ n5004;
  assign n5021 = n5020 ^ n5017;
  assign n5061 = n5060 ^ n5021;
  assign n5079 = n5078 ^ n5061;
  assign n4989 = ~n524 & n2052;
  assign n4990 = ~n291 & ~n431;
  assign n4991 = n758 & n4990;
  assign n4992 = n4989 & n4991;
  assign n4993 = n3764 & n4992;
  assign n4994 = n793 & n4604;
  assign n4995 = n4993 & n4994;
  assign n4996 = n3741 & n4995;
  assign n4997 = n2262 & n4996;
  assign n5080 = n5079 ^ n4997;
  assign n5099 = n5098 ^ n5080;
  assign n5186 = n4846 & ~n4986;
  assign n5187 = n5080 ^ n4983;
  assign n5188 = n5187 ^ n4983;
  assign n5189 = n4983 ^ n4982;
  assign n5190 = ~n5188 & ~n5189;
  assign n5191 = n5190 ^ n4983;
  assign n5192 = n5186 & n5191;
  assign n5193 = ~n3907 & ~n5192;
  assign n5194 = ~n4978 & n5080;
  assign n5195 = n4844 & ~n5194;
  assign n5196 = n4981 ^ n4978;
  assign n5197 = n5196 ^ n4978;
  assign n5198 = n5080 ^ n4978;
  assign n5199 = n5197 & n5198;
  assign n5200 = n5199 ^ n4978;
  assign n5201 = ~n4983 & ~n5200;
  assign n5202 = n5201 ^ n4981;
  assign n5203 = n5195 & n5202;
  assign n5204 = ~n5193 & ~n5203;
  assign n5173 = ~n5061 & ~n5063;
  assign n5174 = ~n5069 & ~n5173;
  assign n5175 = ~n5061 & ~n5065;
  assign n5176 = ~n5070 & ~n5175;
  assign n5177 = n5174 & n5176;
  assign n5178 = n4958 & ~n5177;
  assign n5179 = n5066 & ~n5174;
  assign n5180 = ~n5064 & n5175;
  assign n5181 = ~n5179 & ~n5180;
  assign n5182 = ~n5178 & n5181;
  assign n5167 = n5017 & ~n5020;
  assign n5168 = n5060 & ~n5167;
  assign n5169 = ~n5017 & n5020;
  assign n5170 = ~n5168 & ~n5169;
  assign n5153 = n2522 & ~n4356;
  assign n5154 = n2414 & n2535;
  assign n5155 = n2528 & ~n3629;
  assign n5156 = ~n5154 & ~n5155;
  assign n5157 = ~n684 & n5156;
  assign n5158 = ~n5153 & n5157;
  assign n5159 = n2777 & n4368;
  assign n5160 = n3895 ^ n850;
  assign n5161 = n2522 & n5160;
  assign n5162 = n3898 & n5161;
  assign n5163 = n684 & ~n5156;
  assign n5164 = ~n5162 & ~n5163;
  assign n5165 = ~n5159 & n5164;
  assign n5166 = ~n5158 & n5165;
  assign n5171 = n5170 ^ n5166;
  assign n5147 = n3166 ^ n2434;
  assign n5148 = ~n551 & n5147;
  assign n5149 = n5148 ^ n1097;
  assign n5141 = n5039 ^ n551;
  assign n5142 = n5141 ^ n2462;
  assign n5143 = n5039 ^ n2434;
  assign n5144 = n3164 & n5143;
  assign n5145 = ~n5142 & n5144;
  assign n5146 = n5145 ^ n5141;
  assign n5150 = n5149 ^ n5146;
  assign n5119 = n552 & ~n3270;
  assign n5120 = n5119 ^ n543;
  assign n5121 = n5120 ^ n2417;
  assign n5122 = n685 & n5121;
  assign n5123 = ~n551 & n2569;
  assign n5124 = n2420 & n5123;
  assign n5125 = n2420 ^ n551;
  assign n5126 = n1938 & n5125;
  assign n5127 = n2765 & n3235;
  assign n5128 = n5127 ^ n2569;
  assign n5129 = ~n5126 & ~n5128;
  assign n5130 = n5129 ^ n543;
  assign n5131 = n5130 ^ n5129;
  assign n5132 = ~n2420 & n2765;
  assign n5133 = ~n551 & n3235;
  assign n5134 = n1938 & n5133;
  assign n5135 = ~n5132 & ~n5134;
  assign n5136 = n5135 ^ n5129;
  assign n5137 = n5131 & n5136;
  assign n5138 = n5137 ^ n5129;
  assign n5139 = ~n5124 & n5138;
  assign n5140 = ~n5122 & n5139;
  assign n5151 = n5150 ^ n5140;
  assign n5116 = n5044 ^ n5040;
  assign n5117 = n5059 & ~n5116;
  assign n5118 = n5117 ^ n5058;
  assign n5152 = n5151 ^ n5118;
  assign n5172 = n5171 ^ n5152;
  assign n5183 = n5182 ^ n5172;
  assign n5108 = n83 & ~n261;
  assign n5109 = n285 & ~n5108;
  assign n5110 = ~n408 & ~n2194;
  assign n5111 = n5109 & n5110;
  assign n5112 = n3775 & n5111;
  assign n5113 = n678 & n5112;
  assign n5114 = n911 & n3696;
  assign n5115 = n5113 & n5114;
  assign n5184 = n5183 ^ n5115;
  assign n5100 = n4997 ^ n4983;
  assign n5101 = n5100 ^ n4997;
  assign n5102 = n4997 ^ n4982;
  assign n5103 = n5102 ^ n4997;
  assign n5104 = ~n5101 & ~n5103;
  assign n5105 = n5104 ^ n4997;
  assign n5106 = ~n5080 & ~n5105;
  assign n5107 = n5106 ^ n5079;
  assign n5185 = n5184 ^ n5107;
  assign n5205 = n5204 ^ n5185;
  assign n5283 = ~n5185 & n5192;
  assign n5284 = ~n3907 & ~n5283;
  assign n5285 = n5185 & n5203;
  assign n5286 = ~n5284 & ~n5285;
  assign n5272 = n1017 & n3623;
  assign n5273 = n51 & ~n159;
  assign n5274 = n56 & ~n249;
  assign n5275 = ~n5273 & ~n5274;
  assign n5276 = ~n518 & n5275;
  assign n5277 = n966 & n1041;
  assign n5278 = n5276 & n5277;
  assign n5279 = n5272 & n5278;
  assign n5280 = n662 & n5279;
  assign n5254 = n685 & ~n4036;
  assign n5255 = ~n2417 & ~n2763;
  assign n5256 = ~n2420 & n2767;
  assign n5257 = ~n5255 & ~n5256;
  assign n5258 = ~n551 & n5257;
  assign n5259 = ~n5254 & n5258;
  assign n5260 = n4464 & n4530;
  assign n5261 = n2414 ^ n543;
  assign n5262 = n685 & ~n5261;
  assign n5263 = n2505 & n5262;
  assign n5264 = n551 & ~n5257;
  assign n5265 = ~n5263 & ~n5264;
  assign n5266 = ~n5260 & n5265;
  assign n5267 = ~n5259 & n5266;
  assign n5247 = n2434 ^ n1097;
  assign n5248 = ~n5147 & ~n5247;
  assign n5249 = n5248 ^ n1097;
  assign n5250 = n3235 & n5249;
  assign n5251 = ~n551 & ~n5250;
  assign n5252 = ~n3235 & ~n5249;
  assign n5253 = n5251 & ~n5252;
  assign n5268 = n5267 ^ n5253;
  assign n5244 = n5149 ^ n5140;
  assign n5245 = n5150 & ~n5244;
  assign n5246 = n5245 ^ n5146;
  assign n5269 = n5268 ^ n5246;
  assign n5228 = n2528 & ~n3895;
  assign n5229 = n2535 & ~n3629;
  assign n5230 = ~n5228 & ~n5229;
  assign n5231 = n5230 ^ n684;
  assign n5232 = n2522 & n4058;
  assign n5233 = n5232 ^ n684;
  assign n5234 = n4058 & n4158;
  assign n5235 = n5234 ^ n684;
  assign n5236 = n684 & ~n5235;
  assign n5237 = n5236 ^ n684;
  assign n5238 = n5233 & n5237;
  assign n5239 = n5238 ^ n5236;
  assign n5240 = n5239 ^ n684;
  assign n5241 = n5240 ^ n5234;
  assign n5242 = ~n5231 & ~n5241;
  assign n5243 = n5242 ^ n5234;
  assign n5270 = n5269 ^ n5243;
  assign n5209 = ~n5118 & ~n5151;
  assign n5210 = n5166 & n5209;
  assign n5211 = n5118 & n5151;
  assign n5212 = ~n5166 & n5211;
  assign n5213 = ~n5210 & ~n5212;
  assign n5214 = ~n5171 & ~n5213;
  assign n5215 = n5166 ^ n5118;
  assign n5216 = ~n5152 & ~n5215;
  assign n5217 = n5216 ^ n5166;
  assign n5218 = n5170 & n5217;
  assign n5219 = ~n5210 & ~n5218;
  assign n5220 = n5219 ^ n5182;
  assign n5221 = n5220 ^ n5219;
  assign n5222 = n5170 & ~n5212;
  assign n5223 = ~n5217 & ~n5222;
  assign n5224 = n5223 ^ n5219;
  assign n5225 = ~n5221 & ~n5224;
  assign n5226 = n5225 ^ n5219;
  assign n5227 = ~n5214 & n5226;
  assign n5271 = n5270 ^ n5227;
  assign n5281 = n5280 ^ n5271;
  assign n5206 = n5183 ^ n5107;
  assign n5207 = n5184 & n5206;
  assign n5208 = n5207 ^ n5107;
  assign n5282 = n5281 ^ n5208;
  assign n5287 = n5286 ^ n5282;
  assign n5378 = n5282 & n5283;
  assign n5379 = ~n3907 & ~n5378;
  assign n5380 = ~n5282 & n5285;
  assign n5381 = ~n5379 & ~n5380;
  assign n5364 = ~n652 & ~n1013;
  assign n5365 = ~n303 & ~n1040;
  assign n5366 = ~n454 & n5365;
  assign n5367 = ~n5364 & n5366;
  assign n5368 = n174 & ~n229;
  assign n5369 = ~n357 & ~n5368;
  assign n5370 = n2106 & n5369;
  assign n5371 = n1046 & n5370;
  assign n5372 = n4082 & n5371;
  assign n5373 = n1982 & n5372;
  assign n5374 = n2102 & n5373;
  assign n5375 = n5367 & n5374;
  assign n5335 = n5252 & ~n5267;
  assign n5336 = ~n2420 & ~n5335;
  assign n5337 = n5249 & n5267;
  assign n5338 = n5133 & n5337;
  assign n5339 = n5336 & ~n5338;
  assign n5340 = n5251 & ~n5335;
  assign n5341 = n3235 & ~n5267;
  assign n5342 = n2420 & ~n5341;
  assign n5343 = ~n5340 & n5342;
  assign n5344 = ~n5339 & ~n5343;
  assign n5345 = n551 & ~n5267;
  assign n5346 = ~n5344 & ~n5345;
  assign n5347 = n5268 ^ n5243;
  assign n5348 = ~n5269 & ~n5347;
  assign n5349 = n5348 ^ n5246;
  assign n5350 = ~n5346 & n5349;
  assign n5351 = ~n551 & ~n5252;
  assign n5352 = ~n5337 & n5351;
  assign n5353 = ~n5133 & n5267;
  assign n5354 = ~n2420 & ~n5353;
  assign n5355 = ~n5352 & n5354;
  assign n5356 = ~n551 & n5335;
  assign n5357 = ~n5251 & n5267;
  assign n5358 = n2420 & ~n5357;
  assign n5359 = ~n5356 & n5358;
  assign n5360 = ~n5355 & ~n5359;
  assign n5361 = ~n5349 & n5360;
  assign n5362 = ~n5350 & ~n5361;
  assign n5319 = ~n5166 & ~n5170;
  assign n5320 = ~n5209 & n5319;
  assign n5321 = ~n5270 & ~n5320;
  assign n5322 = ~n5182 & ~n5321;
  assign n5323 = n5166 & n5170;
  assign n5324 = n5270 & ~n5323;
  assign n5325 = ~n5211 & ~n5324;
  assign n5326 = ~n5322 & n5325;
  assign n5327 = ~n5209 & n5270;
  assign n5328 = n5182 ^ n5170;
  assign n5329 = n5182 ^ n5166;
  assign n5330 = n5328 & n5329;
  assign n5331 = n5330 ^ n5182;
  assign n5332 = ~n5327 & n5331;
  assign n5333 = ~n5326 & ~n5332;
  assign n5304 = n685 & ~n4669;
  assign n5305 = n2414 & ~n2763;
  assign n5306 = ~n2417 & n2767;
  assign n5307 = ~n5305 & ~n5306;
  assign n5308 = ~n551 & n5307;
  assign n5309 = ~n5304 & n5308;
  assign n5310 = n4214 & n4464;
  assign n5311 = n3629 ^ n543;
  assign n5312 = n685 & n5311;
  assign n5313 = n3632 & n5312;
  assign n5314 = n551 & ~n5307;
  assign n5315 = ~n5313 & ~n5314;
  assign n5316 = ~n5310 & n5315;
  assign n5317 = ~n5309 & n5316;
  assign n5291 = n3897 ^ n684;
  assign n5292 = n5291 ^ n684;
  assign n5293 = ~n850 & ~n3895;
  assign n5294 = n5293 ^ n684;
  assign n5295 = ~n5292 & ~n5294;
  assign n5296 = n5295 ^ n684;
  assign n5297 = ~n2524 & ~n5296;
  assign n5298 = n2526 ^ n684;
  assign n5299 = n2526 ^ n850;
  assign n5300 = ~n5298 & n5299;
  assign n5301 = ~n3895 & n5300;
  assign n5302 = n5301 ^ n684;
  assign n5303 = ~n5297 & n5302;
  assign n5318 = n5317 ^ n5303;
  assign n5334 = n5333 ^ n5318;
  assign n5363 = n5362 ^ n5334;
  assign n5376 = n5375 ^ n5363;
  assign n5288 = n5271 ^ n5208;
  assign n5289 = ~n5281 & ~n5288;
  assign n5290 = n5289 ^ n5208;
  assign n5377 = n5376 ^ n5290;
  assign n5382 = n5381 ^ n5377;
  assign n5473 = ~n5377 & n5378;
  assign n5474 = ~n3907 & ~n5473;
  assign n5475 = n5377 & n5380;
  assign n5476 = ~n5474 & ~n5475;
  assign n5402 = ~n5333 & ~n5350;
  assign n5403 = ~n5361 & n5402;
  assign n5436 = ~n551 & n5336;
  assign n5437 = ~n5357 & ~n5436;
  assign n5409 = n3895 ^ n543;
  assign n5410 = n3898 & n5409;
  assign n5411 = ~n4356 & ~n5410;
  assign n5412 = n2326 & n2414;
  assign n5413 = ~n2763 & ~n3629;
  assign n5414 = ~n551 & ~n5413;
  assign n5415 = ~n5412 & n5414;
  assign n5416 = ~n5411 & n5415;
  assign n5417 = n551 & ~n2414;
  assign n5418 = n2569 & ~n5417;
  assign n5419 = n3629 ^ n551;
  assign n5420 = n1938 & n5419;
  assign n5421 = ~n543 & ~n5420;
  assign n5422 = ~n5418 & n5421;
  assign n5423 = ~n2414 & n2753;
  assign n5424 = n2765 & ~n3629;
  assign n5425 = n543 & ~n5424;
  assign n5426 = ~n5423 & n5425;
  assign n5427 = ~n5422 & ~n5426;
  assign n5428 = ~n551 & n3629;
  assign n5429 = n2569 & n5428;
  assign n5430 = ~n5427 & ~n5429;
  assign n5431 = ~n5416 & n5430;
  assign n5432 = ~n4368 & ~n5410;
  assign n5433 = n4464 & ~n5432;
  assign n5434 = n5431 & ~n5433;
  assign n5404 = ~n2417 & ~n2420;
  assign n5405 = n2400 & n2420;
  assign n5406 = ~n551 & ~n5405;
  assign n5407 = ~n5404 & n5406;
  assign n5408 = n5407 ^ n684;
  assign n5435 = n5434 ^ n5408;
  assign n5438 = n5437 ^ n5435;
  assign n5439 = ~n5361 & ~n5438;
  assign n5440 = n5333 & ~n5439;
  assign n5441 = ~n5403 & ~n5440;
  assign n5442 = ~n5350 & n5438;
  assign n5443 = n5303 & ~n5317;
  assign n5444 = ~n5442 & ~n5443;
  assign n5445 = ~n5441 & n5444;
  assign n5446 = ~n5333 & ~n5438;
  assign n5447 = n5438 ^ n5361;
  assign n5448 = ~n5303 & n5317;
  assign n5449 = n5448 ^ n5443;
  assign n5450 = n5449 ^ n5443;
  assign n5451 = n5443 ^ n5438;
  assign n5452 = n5451 ^ n5443;
  assign n5453 = n5450 & n5452;
  assign n5454 = n5453 ^ n5443;
  assign n5455 = n5447 & n5454;
  assign n5456 = n5455 ^ n5443;
  assign n5457 = ~n5446 & n5456;
  assign n5458 = ~n5403 & n5457;
  assign n5459 = n5402 & ~n5438;
  assign n5460 = n5448 & n5459;
  assign n5461 = ~n5458 & ~n5460;
  assign n5462 = ~n5445 & n5461;
  assign n5463 = n5402 & n5443;
  assign n5464 = n5333 & ~n5362;
  assign n5465 = ~n5361 & n5438;
  assign n5466 = ~n5448 & ~n5465;
  assign n5467 = ~n5464 & n5466;
  assign n5468 = ~n5463 & ~n5467;
  assign n5469 = ~n5459 & ~n5468;
  assign n5470 = n5462 & ~n5469;
  assign n5386 = n914 & n3683;
  assign n5387 = ~n394 & ~n566;
  assign n5388 = ~n92 & ~n2154;
  assign n5389 = n5387 & n5388;
  assign n5390 = n5386 & n5389;
  assign n5391 = ~n200 & ~n1029;
  assign n5392 = n139 & ~n495;
  assign n5393 = ~n420 & ~n5392;
  assign n5394 = ~n5391 & n5393;
  assign n5395 = ~n356 & ~n583;
  assign n5396 = ~n2394 & n5395;
  assign n5397 = n5394 & n5396;
  assign n5398 = n5390 & n5397;
  assign n5399 = n219 & n5398;
  assign n5400 = n3648 & n5399;
  assign n5401 = n3778 & n5400;
  assign n5471 = n5470 ^ n5401;
  assign n5383 = n5363 ^ n5290;
  assign n5384 = n5376 & n5383;
  assign n5385 = n5384 ^ n5290;
  assign n5472 = n5471 ^ n5385;
  assign n5477 = n5476 ^ n5472;
  assign n5532 = n5472 & n5473;
  assign n5533 = ~n3907 & ~n5532;
  assign n5534 = ~n5472 & n5475;
  assign n5535 = ~n5533 & ~n5534;
  assign n5518 = ~n5442 & n5448;
  assign n5519 = ~n5439 & ~n5518;
  assign n5520 = ~n5333 & n5519;
  assign n5521 = n5442 & ~n5448;
  assign n5522 = ~n5438 & ~n5443;
  assign n5523 = n5438 & n5443;
  assign n5524 = ~n5361 & ~n5523;
  assign n5525 = ~n5522 & ~n5524;
  assign n5526 = ~n5521 & ~n5525;
  assign n5527 = ~n5520 & n5526;
  assign n5528 = ~n5463 & n5527;
  assign n5502 = n552 & n4058;
  assign n5503 = n685 & ~n5502;
  assign n5504 = n543 & ~n3895;
  assign n5505 = n3095 & ~n3629;
  assign n5506 = n2569 & ~n5505;
  assign n5507 = ~n5504 & n5506;
  assign n5508 = n5409 ^ n3895;
  assign n5509 = ~n551 & ~n3629;
  assign n5510 = n5509 ^ n3895;
  assign n5511 = n5508 & ~n5510;
  assign n5512 = n5511 ^ n3895;
  assign n5513 = n1938 & n5512;
  assign n5514 = ~n5507 & ~n5513;
  assign n5515 = ~n5503 & n5514;
  assign n5496 = ~n684 & ~n5405;
  assign n5497 = ~n5404 & ~n5496;
  assign n5498 = n2414 & n5497;
  assign n5499 = ~n551 & ~n5498;
  assign n5500 = ~n2414 & ~n5497;
  assign n5501 = n5499 & ~n5500;
  assign n5516 = n5515 ^ n5501;
  assign n5493 = n5437 ^ n5434;
  assign n5494 = ~n5435 & ~n5493;
  assign n5495 = n5494 ^ n5437;
  assign n5517 = n5516 ^ n5495;
  assign n5529 = n5528 ^ n5517;
  assign n5481 = ~n468 & ~n665;
  assign n5482 = n2106 & n5481;
  assign n5483 = n83 & ~n4962;
  assign n5484 = n5482 & ~n5483;
  assign n5485 = ~n239 & ~n1963;
  assign n5486 = n634 & n5485;
  assign n5487 = n2392 & n5486;
  assign n5488 = n5484 & n5487;
  assign n5489 = n901 & n5488;
  assign n5490 = n1069 & n5489;
  assign n5491 = n437 & n2301;
  assign n5492 = n5490 & n5491;
  assign n5530 = n5529 ^ n5492;
  assign n5478 = n5470 ^ n5385;
  assign n5479 = ~n5471 & ~n5478;
  assign n5480 = n5479 ^ n5385;
  assign n5531 = n5530 ^ n5480;
  assign n5536 = n5535 ^ n5531;
  assign n5608 = n5531 & n5534;
  assign n5609 = n3907 & ~n5608;
  assign n5610 = ~n5531 & n5532;
  assign n5611 = ~n5609 & ~n5610;
  assign n5593 = ~n250 & n1110;
  assign n5594 = n954 & n5593;
  assign n5595 = ~n207 & ~n210;
  assign n5596 = n5485 & n5595;
  assign n5597 = n57 & ~n331;
  assign n5598 = ~n524 & ~n5597;
  assign n5599 = ~n1132 & n5598;
  assign n5600 = n5596 & n5599;
  assign n5601 = n3656 & n5600;
  assign n5602 = n887 & n5601;
  assign n5603 = n2116 & n5602;
  assign n5604 = n5594 & n5603;
  assign n5605 = n5367 & n5604;
  assign n5540 = n5528 ^ n5495;
  assign n5541 = n5517 & ~n5540;
  assign n5542 = n5541 ^ n5528;
  assign n5548 = n685 & n3897;
  assign n5549 = n552 & n2763;
  assign n5550 = ~n3895 & n5549;
  assign n5551 = ~n5548 & n5550;
  assign n5552 = ~n2414 & ~n5551;
  assign n5569 = ~n3629 & n5552;
  assign n5570 = n5515 ^ n551;
  assign n5571 = n5570 ^ n5515;
  assign n5547 = n5497 & n5515;
  assign n5572 = n5547 ^ n5515;
  assign n5573 = ~n5571 & ~n5572;
  assign n5574 = n5573 ^ n5515;
  assign n5575 = n5569 & n5574;
  assign n5543 = n2414 & n5509;
  assign n5544 = n5501 & n5515;
  assign n5545 = n5544 ^ n5499;
  assign n5546 = n5543 & n5545;
  assign n5556 = ~n2414 & n3629;
  assign n5576 = n551 & ~n5515;
  assign n5577 = ~n5556 & ~n5576;
  assign n5578 = ~n5546 & n5577;
  assign n5579 = n5578 ^ n5551;
  assign n5580 = n5579 ^ n5578;
  assign n5558 = n551 & n5515;
  assign n5559 = ~n5545 & ~n5558;
  assign n5581 = ~n551 & ~n2414;
  assign n5582 = ~n5509 & ~n5581;
  assign n5583 = ~n5559 & n5582;
  assign n5584 = n5543 & ~n5545;
  assign n5585 = ~n5583 & ~n5584;
  assign n5586 = n5585 ^ n5578;
  assign n5587 = ~n5580 & n5586;
  assign n5588 = n5587 ^ n5578;
  assign n5589 = ~n5575 & n5588;
  assign n5553 = n5428 & n5552;
  assign n5554 = ~n5547 & n5553;
  assign n5555 = ~n5546 & ~n5554;
  assign n5557 = n5551 & ~n5556;
  assign n5560 = n5559 ^ n5557;
  assign n5561 = n5560 ^ n5557;
  assign n5562 = n3629 ^ n2414;
  assign n5563 = ~n551 & n5562;
  assign n5564 = ~n5551 & ~n5563;
  assign n5565 = n5564 ^ n5557;
  assign n5566 = n5561 & n5565;
  assign n5567 = n5566 ^ n5557;
  assign n5568 = n5555 & ~n5567;
  assign n5590 = n5589 ^ n5568;
  assign n5591 = ~n5542 & n5590;
  assign n5592 = n5591 ^ n5589;
  assign n5606 = n5605 ^ n5592;
  assign n5537 = n5529 ^ n5480;
  assign n5538 = n5530 & n5537;
  assign n5539 = n5538 ^ n5480;
  assign n5607 = n5606 ^ n5539;
  assign n5612 = n5611 ^ n5607;
  assign n5650 = ~n5607 & n5610;
  assign n5651 = ~n3907 & ~n5650;
  assign n5652 = n5607 & n5608;
  assign n5653 = ~n5651 & ~n5652;
  assign n5634 = n3629 & n5551;
  assign n5635 = n5634 ^ n5563;
  assign n5636 = n5634 ^ n5559;
  assign n5637 = ~n5634 & n5636;
  assign n5638 = n5637 ^ n5634;
  assign n5639 = ~n5635 & ~n5638;
  assign n5640 = n5639 ^ n5637;
  assign n5641 = n5640 ^ n5634;
  assign n5642 = n5641 ^ n5559;
  assign n5643 = ~n5557 & n5642;
  assign n5644 = n5542 & ~n5643;
  assign n5645 = n5559 & ~n5564;
  assign n5646 = ~n5644 & ~n5645;
  assign n5627 = n551 & ~n5551;
  assign n5628 = n543 & n3629;
  assign n5629 = n5423 & n5628;
  assign n5630 = n2414 & ~n5428;
  assign n5631 = n3895 & ~n5630;
  assign n5632 = ~n5629 & ~n5631;
  assign n5633 = ~n5627 & n5632;
  assign n5647 = n5646 ^ n5633;
  assign n5616 = ~n57 & n1983;
  assign n5617 = ~n2149 & ~n5616;
  assign n5618 = ~n380 & ~n1963;
  assign n5619 = ~n620 & n5618;
  assign n5620 = n3647 & n5619;
  assign n5621 = n2352 & n5620;
  assign n5622 = n3723 & n5621;
  assign n5623 = n5389 & n5622;
  assign n5624 = n3661 & n5623;
  assign n5625 = n1036 & n5624;
  assign n5626 = ~n5617 & n5625;
  assign n5648 = n5647 ^ n5626;
  assign n5613 = n5592 ^ n5539;
  assign n5614 = n5606 & n5613;
  assign n5615 = n5614 ^ n5539;
  assign n5649 = n5648 ^ n5615;
  assign n5654 = n5653 ^ n5649;
  assign n5670 = ~n5649 & n5652;
  assign n5671 = n3907 & ~n5670;
  assign n5672 = n5649 & n5650;
  assign n5673 = ~n5671 & ~n5672;
  assign n5658 = n466 & n815;
  assign n5659 = n5395 & n5658;
  assign n5660 = ~n238 & ~n358;
  assign n5661 = n2318 & n5660;
  assign n5662 = ~n120 & n582;
  assign n5663 = ~n652 & ~n5662;
  assign n5664 = n888 & ~n5663;
  assign n5665 = n5661 & n5664;
  assign n5666 = n5659 & n5665;
  assign n5667 = n632 & n5666;
  assign n5668 = n2363 & n5667;
  assign n5655 = n5647 ^ n5615;
  assign n5656 = ~n5648 & ~n5655;
  assign n5657 = n5656 ^ n5615;
  assign n5669 = n5668 ^ n5657;
  assign n5674 = n5673 ^ n5669;
  assign n5684 = n5672 ^ n5657;
  assign n5685 = n5669 & n5684;
  assign n5686 = n5685 ^ n5672;
  assign n5687 = ~n3907 & ~n5686;
  assign n5688 = ~n5657 & n5668;
  assign n5689 = n5670 & n5688;
  assign n5690 = n5657 & ~n5668;
  assign n5691 = n5671 & n5690;
  assign n5692 = ~n5689 & ~n5691;
  assign n5693 = ~n5687 & n5692;
  assign n5675 = n204 & n1118;
  assign n5676 = n640 & ~n1141;
  assign n5677 = n3721 & n4113;
  assign n5678 = n5676 & n5677;
  assign n5679 = n959 & n5678;
  assign n5680 = n5675 & n5679;
  assign n5681 = n591 & n5680;
  assign n5682 = n879 & n5681;
  assign n5683 = n3673 & n5682;
  assign n5694 = n5693 ^ n5683;
  assign n5706 = ~n5683 & ~n5690;
  assign n5707 = n5670 & ~n5706;
  assign n5708 = ~n5669 & n5672;
  assign n5709 = ~n5707 & ~n5708;
  assign n5710 = n5683 & ~n5689;
  assign n5711 = ~n5709 & ~n5710;
  assign n5712 = n3907 & ~n5711;
  assign n5704 = ~n5683 & n5686;
  assign n5695 = n139 & ~n2355;
  assign n5696 = n2096 & ~n5695;
  assign n5697 = n158 & n175;
  assign n5698 = ~n308 & ~n5697;
  assign n5699 = n5696 & n5698;
  assign n5700 = n4433 & n5699;
  assign n5701 = n372 & n5700;
  assign n5702 = n1011 & n5701;
  assign n5703 = n5594 & n5702;
  assign n5705 = n5704 ^ n5703;
  assign n5713 = n5712 ^ n5705;
  assign n5722 = ~n85 & ~n396;
  assign n5723 = ~n274 & n5722;
  assign n5724 = ~n226 & n5723;
  assign n5725 = n147 & n419;
  assign n5726 = ~n1023 & ~n5725;
  assign n5727 = n5724 & ~n5726;
  assign n5728 = n4440 & n5727;
  assign n5729 = ~n2387 & n5728;
  assign n5730 = n1122 & n5729;
  assign n5731 = n4966 & n5730;
  assign n5714 = n5711 ^ n5703;
  assign n5715 = n5714 ^ n5703;
  assign n5716 = n5703 ^ n3907;
  assign n5717 = n5716 ^ n5703;
  assign n5718 = n5715 & n5717;
  assign n5719 = n5718 ^ n5703;
  assign n5720 = n5705 & ~n5719;
  assign n5721 = n5720 ^ n3907;
  assign n5732 = n5731 ^ n5721;
  assign n5739 = ~n5703 & n5704;
  assign n5740 = n5712 & n5739;
  assign n5741 = ~n5731 & n5740;
  assign n5742 = n5704 ^ n3907;
  assign n5743 = ~n5703 & ~n5731;
  assign n5744 = n5743 ^ n5704;
  assign n5745 = n5744 ^ n5743;
  assign n5746 = n5703 & n5731;
  assign n5747 = n5746 ^ n5743;
  assign n5748 = ~n5745 & n5747;
  assign n5749 = n5748 ^ n5743;
  assign n5750 = n5742 & n5749;
  assign n5751 = n5750 ^ n3907;
  assign n5752 = ~n5712 & ~n5751;
  assign n5753 = ~n5741 & ~n5752;
  assign n5733 = ~n56 & n180;
  assign n5734 = ~n633 & ~n5733;
  assign n5735 = ~n347 & ~n531;
  assign n5736 = n506 & n5735;
  assign n5737 = n2402 & n5736;
  assign n5738 = ~n5734 & n5737;
  assign n5754 = n5753 ^ n5738;
  assign n5755 = n544 & ~n2409;
  assign n5756 = ~n5738 & n5743;
  assign n5757 = n5704 & n5756;
  assign n5760 = n5757 ^ n5704;
  assign n5761 = ~n5755 & ~n5760;
  assign n5762 = n5761 ^ n5704;
  assign n5758 = n5757 ^ n5755;
  assign n5759 = n5758 ^ n3907;
  assign n5763 = n5762 ^ n5759;
  assign n5764 = n5762 ^ n5758;
  assign n5765 = n5738 & n5746;
  assign n5766 = n5765 ^ n5756;
  assign n5767 = ~n5704 & n5766;
  assign n5768 = n5767 ^ n5756;
  assign n5769 = n5711 & n5768;
  assign n5770 = n5769 ^ n5758;
  assign n5771 = ~n5758 & ~n5770;
  assign n5772 = n5771 ^ n5758;
  assign n5773 = n5764 & ~n5772;
  assign n5774 = n5773 ^ n5771;
  assign n5775 = n5774 ^ n5758;
  assign n5776 = n5775 ^ n5769;
  assign n5777 = ~n5763 & ~n5776;
  assign n5778 = n5777 ^ n5759;
  assign n5779 = ~x21 & ~x22;
  assign n5780 = n544 & n5779;
  assign n5781 = ~n5755 & n5757;
  assign n5782 = n5712 ^ n3907;
  assign n5783 = n5781 & ~n5782;
  assign n5784 = n5783 ^ n3907;
  assign n5785 = ~n5780 & ~n5784;
  assign n5786 = n5755 & ~n5757;
  assign n5787 = ~n5779 & n5786;
  assign n5788 = n5769 & n5787;
  assign n5789 = ~n5785 & ~n5788;
  assign n5790 = n3907 & ~n5788;
  assign y0 = n3756;
  assign y1 = ~n3922;
  assign y2 = ~n4111;
  assign y3 = n4279;
  assign y4 = n4414;
  assign y5 = n4587;
  assign y6 = n4726;
  assign y7 = n4843;
  assign y8 = ~n4988;
  assign y9 = ~n5099;
  assign y10 = ~n5205;
  assign y11 = n5287;
  assign y12 = ~n5382;
  assign y13 = n5477;
  assign y14 = ~n5536;
  assign y15 = n5612;
  assign y16 = n5654;
  assign y17 = n5674;
  assign y18 = ~n5694;
  assign y19 = ~n5713;
  assign y20 = ~n5732;
  assign y21 = ~n5754;
  assign y22 = ~n5778;
  assign y23 = n5789;
  assign y24 = n5790;
endmodule
