module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, y0, y1, y2, y3, y4, y5, y6, y7);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127;
  output y0, y1, y2, y3, y4, y5, y6, y7;
  wire n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496;
  assign n129 = ~x2 & ~x3;
  assign n130 = x1 & n129;
  assign n131 = n130 ^ x3;
  assign n132 = ~x4 & n131;
  assign n133 = ~x5 & ~n132;
  assign n134 = ~x6 & ~n133;
  assign n135 = ~x7 & ~n134;
  assign n136 = ~x8 & ~n135;
  assign n137 = ~x9 & ~n136;
  assign n138 = ~x10 & ~n137;
  assign n139 = ~x11 & ~n138;
  assign n140 = ~x12 & ~n139;
  assign n141 = ~x13 & ~n140;
  assign n142 = ~x14 & ~n141;
  assign n143 = ~x15 & ~n142;
  assign n144 = ~x16 & ~n143;
  assign n145 = ~x17 & ~n144;
  assign n146 = ~x18 & ~n145;
  assign n147 = ~x19 & ~n146;
  assign n148 = ~x20 & ~n147;
  assign n149 = ~x21 & ~n148;
  assign n150 = ~x22 & ~n149;
  assign n151 = ~x23 & ~n150;
  assign n152 = ~x24 & ~n151;
  assign n153 = ~x25 & ~n152;
  assign n154 = ~x26 & ~n153;
  assign n155 = ~x27 & ~n154;
  assign n156 = ~x28 & ~n155;
  assign n157 = ~x29 & ~n156;
  assign n158 = ~x30 & ~n157;
  assign n159 = ~x31 & ~n158;
  assign n160 = ~x32 & ~n159;
  assign n161 = ~x33 & ~n160;
  assign n162 = ~x34 & ~n161;
  assign n163 = ~x35 & ~n162;
  assign n164 = ~x36 & ~n163;
  assign n165 = ~x37 & ~n164;
  assign n166 = ~x38 & ~n165;
  assign n167 = ~x39 & ~n166;
  assign n168 = ~x40 & ~n167;
  assign n169 = ~x41 & ~n168;
  assign n170 = ~x42 & ~n169;
  assign n171 = ~x43 & ~n170;
  assign n172 = ~x44 & ~n171;
  assign n173 = ~x45 & ~n172;
  assign n174 = ~x46 & ~n173;
  assign n175 = ~x47 & ~n174;
  assign n176 = ~x48 & ~n175;
  assign n177 = ~x49 & ~n176;
  assign n178 = ~x50 & ~n177;
  assign n179 = ~x51 & ~n178;
  assign n180 = ~x52 & ~n179;
  assign n181 = ~x53 & ~n180;
  assign n182 = ~x54 & ~n181;
  assign n183 = ~x55 & ~n182;
  assign n184 = ~x56 & ~n183;
  assign n185 = ~x57 & ~n184;
  assign n186 = ~x58 & ~n185;
  assign n187 = ~x59 & ~n186;
  assign n188 = ~x60 & ~n187;
  assign n189 = ~x61 & ~n188;
  assign n190 = ~x62 & ~n189;
  assign n191 = ~x63 & ~n190;
  assign n192 = ~x64 & ~n191;
  assign n193 = ~x65 & ~n192;
  assign n194 = ~x66 & ~n193;
  assign n195 = ~x67 & ~n194;
  assign n196 = ~x68 & ~n195;
  assign n197 = ~x69 & ~n196;
  assign n198 = ~x70 & ~n197;
  assign n199 = ~x71 & ~n198;
  assign n200 = ~x72 & ~n199;
  assign n201 = ~x73 & ~n200;
  assign n202 = ~x74 & ~n201;
  assign n203 = ~x75 & ~n202;
  assign n204 = ~x76 & ~n203;
  assign n205 = ~x77 & ~n204;
  assign n206 = ~x78 & ~n205;
  assign n207 = ~x79 & ~n206;
  assign n208 = ~x80 & ~n207;
  assign n209 = ~x81 & ~n208;
  assign n210 = ~x82 & ~n209;
  assign n211 = ~x83 & ~n210;
  assign n212 = ~x84 & ~n211;
  assign n213 = ~x85 & ~n212;
  assign n214 = ~x86 & ~n213;
  assign n215 = ~x87 & ~n214;
  assign n216 = ~x88 & ~n215;
  assign n217 = ~x89 & ~n216;
  assign n218 = ~x90 & ~n217;
  assign n219 = ~x91 & ~n218;
  assign n220 = ~x92 & ~n219;
  assign n221 = ~x93 & ~n220;
  assign n222 = ~x94 & ~n221;
  assign n223 = ~x95 & ~n222;
  assign n224 = ~x96 & ~n223;
  assign n225 = ~x97 & ~n224;
  assign n226 = ~x98 & ~n225;
  assign n227 = ~x99 & ~n226;
  assign n228 = ~x100 & ~n227;
  assign n229 = ~x101 & ~n228;
  assign n230 = ~x102 & ~n229;
  assign n231 = ~x103 & ~n230;
  assign n232 = ~x104 & ~n231;
  assign n233 = ~x105 & ~n232;
  assign n234 = ~x106 & ~n233;
  assign n235 = ~x107 & ~n234;
  assign n236 = ~x108 & ~n235;
  assign n237 = ~x109 & ~n236;
  assign n238 = ~x110 & ~n237;
  assign n239 = ~x111 & ~n238;
  assign n240 = ~x112 & ~n239;
  assign n241 = ~x113 & ~n240;
  assign n242 = ~x114 & ~n241;
  assign n243 = ~x115 & ~n242;
  assign n244 = ~x116 & ~n243;
  assign n245 = ~x117 & ~n244;
  assign n246 = ~x118 & ~n245;
  assign n247 = ~x119 & ~n246;
  assign n248 = ~x120 & ~n247;
  assign n249 = ~x121 & ~n248;
  assign n250 = ~x122 & ~n249;
  assign n251 = ~x123 & ~n250;
  assign n252 = ~x124 & ~n251;
  assign n253 = ~x125 & ~n252;
  assign n254 = ~x126 & ~n253;
  assign n255 = ~x127 & ~n254;
  assign n256 = ~x126 & ~x127;
  assign n257 = ~x124 & ~x125;
  assign n258 = ~x122 & ~x123;
  assign n259 = ~x120 & ~x121;
  assign n260 = n258 & n259;
  assign n261 = ~x118 & ~x119;
  assign n262 = ~x116 & ~x117;
  assign n263 = n261 & n262;
  assign n264 = n260 & n263;
  assign n265 = ~x114 & ~x115;
  assign n266 = n256 & n257;
  assign n267 = ~x112 & ~x113;
  assign n268 = n265 & n267;
  assign n269 = n264 & n268;
  assign n270 = n266 & n269;
  assign n271 = ~x110 & ~x111;
  assign n272 = ~x108 & ~x109;
  assign n273 = ~x106 & ~x107;
  assign n274 = ~x104 & ~x105;
  assign n275 = n273 & n274;
  assign n276 = ~x102 & ~x103;
  assign n277 = ~x100 & ~x101;
  assign n278 = ~x98 & ~x99;
  assign n279 = ~x96 & ~x97;
  assign n280 = ~x94 & ~x95;
  assign n281 = ~x92 & ~x93;
  assign n282 = ~x90 & ~x91;
  assign n283 = ~x88 & ~x89;
  assign n284 = n282 & n283;
  assign n285 = ~x84 & ~x85;
  assign n286 = ~x86 & ~x87;
  assign n287 = n285 & n286;
  assign n288 = n280 & n281;
  assign n289 = n284 & n288;
  assign n290 = ~x82 & ~x83;
  assign n291 = ~x80 & ~x81;
  assign n292 = n290 & n291;
  assign n293 = n289 & n292;
  assign n294 = n287 & n293;
  assign n295 = ~x78 & ~x79;
  assign n296 = ~x76 & ~x77;
  assign n297 = ~x74 & ~x75;
  assign n298 = ~x72 & ~x73;
  assign n299 = n297 & n298;
  assign n300 = ~x70 & ~x71;
  assign n301 = ~x68 & ~x69;
  assign n302 = ~x66 & ~x67;
  assign n303 = n295 & n296;
  assign n304 = n299 & n303;
  assign n305 = n300 & n301;
  assign n306 = ~x64 & ~x65;
  assign n307 = n302 & n306;
  assign n308 = n305 & n307;
  assign n309 = n304 & n308;
  assign n310 = ~x62 & ~x63;
  assign n311 = ~x60 & ~x61;
  assign n312 = n310 & n311;
  assign n313 = ~x58 & ~x59;
  assign n314 = ~x56 & ~x57;
  assign n315 = n313 & n314;
  assign n316 = n312 & n315;
  assign n317 = ~x54 & ~x55;
  assign n318 = ~x52 & ~x53;
  assign n319 = n317 & n318;
  assign n320 = ~x50 & ~x51;
  assign n321 = ~x48 & ~x49;
  assign n322 = n320 & n321;
  assign n323 = n319 & n322;
  assign n324 = n316 & n323;
  assign n325 = ~x46 & ~x47;
  assign n326 = ~x44 & ~x45;
  assign n327 = n325 & n326;
  assign n328 = ~x42 & ~x43;
  assign n329 = ~x40 & ~x41;
  assign n330 = n328 & n329;
  assign n331 = n327 & n330;
  assign n332 = ~x38 & ~x39;
  assign n333 = ~x36 & ~x37;
  assign n334 = n332 & n333;
  assign n335 = ~x34 & ~x35;
  assign n336 = ~x32 & ~x33;
  assign n337 = n335 & n336;
  assign n338 = n334 & n337;
  assign n339 = n331 & n338;
  assign n340 = n324 & n339;
  assign n341 = ~x18 & ~x19;
  assign n342 = ~x16 & ~x17;
  assign n343 = n341 & n342;
  assign n344 = ~x30 & ~x31;
  assign n345 = ~x28 & ~x29;
  assign n346 = n344 & n345;
  assign n347 = ~x26 & ~x27;
  assign n348 = ~x24 & ~x25;
  assign n349 = n347 & n348;
  assign n350 = n346 & n349;
  assign n351 = ~x22 & ~x23;
  assign n352 = ~x20 & ~x21;
  assign n353 = n351 & n352;
  assign n354 = n350 & n353;
  assign n355 = n343 & n354;
  assign n356 = ~x14 & ~x15;
  assign n357 = ~x12 & ~x13;
  assign n358 = ~x10 & ~x11;
  assign n359 = n271 & n272;
  assign n360 = n275 & n359;
  assign n361 = n278 & n279;
  assign n362 = n276 & n277;
  assign n363 = n361 & n362;
  assign n364 = n360 & n363;
  assign n365 = n339 & ~n355;
  assign n366 = n324 & ~n365;
  assign n367 = n309 & ~n366;
  assign n368 = n294 & ~n367;
  assign n369 = n364 & ~n368;
  assign n370 = n356 & n357;
  assign n371 = ~x8 & ~x9;
  assign n372 = n358 & n371;
  assign n373 = n370 & n372;
  assign n374 = ~n369 & ~n373;
  assign n375 = ~x4 & ~x5;
  assign n376 = ~n129 & n375;
  assign n377 = ~x6 & ~x7;
  assign n378 = ~n376 & n377;
  assign n379 = ~n374 & ~n378;
  assign n380 = n358 & ~n379;
  assign n381 = n357 & ~n380;
  assign n382 = n356 & ~n381;
  assign n383 = n355 & ~n382;
  assign n384 = n349 & ~n351;
  assign n385 = n347 & ~n384;
  assign n386 = n346 & ~n385;
  assign n387 = ~n341 & n354;
  assign n388 = n344 & ~n387;
  assign n389 = ~n386 & n388;
  assign n390 = ~n383 & n389;
  assign n391 = n340 & ~n390;
  assign n392 = n335 & ~n391;
  assign n393 = n334 & ~n392;
  assign n394 = n332 & ~n393;
  assign n395 = n331 & ~n394;
  assign n396 = n326 & ~n328;
  assign n397 = n325 & ~n396;
  assign n398 = ~n395 & n397;
  assign n399 = n324 & ~n398;
  assign n400 = n318 & ~n320;
  assign n401 = n317 & ~n400;
  assign n402 = ~n399 & n401;
  assign n403 = n316 & ~n402;
  assign n404 = n311 & ~n313;
  assign n405 = n310 & ~n404;
  assign n406 = ~n403 & n405;
  assign n407 = n309 & ~n406;
  assign n408 = n302 & ~n407;
  assign n409 = n301 & ~n408;
  assign n410 = n300 & ~n409;
  assign n411 = n299 & ~n410;
  assign n412 = n297 & ~n411;
  assign n413 = n296 & ~n412;
  assign n414 = n295 & ~n413;
  assign n415 = n294 & ~n414;
  assign n416 = n285 & ~n290;
  assign n417 = n286 & ~n416;
  assign n418 = ~n415 & n417;
  assign n419 = n284 & ~n418;
  assign n420 = n282 & ~n419;
  assign n421 = n281 & ~n420;
  assign n422 = n280 & ~n421;
  assign n423 = n279 & ~n422;
  assign n424 = n278 & ~n423;
  assign n425 = n277 & ~n424;
  assign n426 = n276 & ~n425;
  assign n427 = n275 & ~n426;
  assign n428 = n273 & ~n427;
  assign n429 = n272 & ~n428;
  assign n430 = n271 & ~n429;
  assign n431 = n270 & ~n430;
  assign n432 = n265 & ~n431;
  assign n433 = n264 & ~n432;
  assign n434 = n259 & ~n261;
  assign n435 = n258 & ~n434;
  assign n436 = ~n433 & n435;
  assign n437 = n257 & ~n436;
  assign n438 = n256 & ~n437;
  assign n439 = n375 & n377;
  assign n440 = ~n374 & ~n439;
  assign n441 = n370 & ~n440;
  assign n442 = n343 & ~n441;
  assign n443 = n353 & ~n442;
  assign n444 = n349 & ~n443;
  assign n445 = n346 & ~n444;
  assign n446 = n337 & ~n445;
  assign n447 = n334 & ~n446;
  assign n448 = n330 & ~n447;
  assign n449 = n327 & ~n448;
  assign n450 = n322 & ~n449;
  assign n451 = n319 & ~n450;
  assign n452 = n315 & ~n451;
  assign n453 = n312 & ~n452;
  assign n454 = n307 & ~n453;
  assign n455 = n305 & ~n454;
  assign n456 = n299 & ~n455;
  assign n457 = n303 & ~n456;
  assign n458 = n293 & ~n457;
  assign n459 = n287 & ~n458;
  assign n460 = n284 & ~n459;
  assign n461 = n288 & ~n460;
  assign n462 = n361 & ~n461;
  assign n463 = n362 & ~n462;
  assign n464 = n275 & ~n463;
  assign n465 = n359 & ~n464;
  assign n466 = n269 & ~n465;
  assign n467 = n263 & ~n466;
  assign n468 = n260 & ~n467;
  assign n469 = n266 & ~n468;
  assign n470 = n260 & n266;
  assign n471 = n350 & ~n374;
  assign n472 = n340 & ~n471;
  assign n473 = n323 & ~n331;
  assign n474 = n316 & ~n473;
  assign n475 = ~n472 & n474;
  assign n476 = n294 & n309;
  assign n477 = ~n475 & n476;
  assign n478 = n294 & ~n304;
  assign n479 = n289 & ~n478;
  assign n480 = ~n477 & n479;
  assign n481 = n363 & ~n480;
  assign n482 = n360 & ~n481;
  assign n483 = n269 & ~n482;
  assign n484 = n470 & ~n483;
  assign n485 = n270 & ~n369;
  assign n486 = n270 & n364;
  assign n487 = n476 & n486;
  assign n488 = ~n340 & n487;
  assign n489 = n488 ^ n486;
  assign n490 = ~x0 & ~x1;
  assign n491 = n340 & n490;
  assign n492 = n487 & n491;
  assign n493 = ~n367 & n492;
  assign n494 = ~n379 & n493;
  assign n495 = ~n472 & n494;
  assign n496 = ~n442 & n495;
  assign y0 = ~n255;
  assign y1 = ~n438;
  assign y2 = ~n469;
  assign y3 = ~n484;
  assign y4 = ~n485;
  assign y5 = ~n489;
  assign y6 = ~n487;
  assign y7 = ~n496;
endmodule
