module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127;
  wire n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592;
  assign n129 = ~x126 & ~x127;
  assign n130 = ~x125 & n129;
  assign n131 = ~x124 & n130;
  assign n132 = ~x123 & n131;
  assign n133 = x122 & n132;
  assign n134 = ~x122 & n132;
  assign n135 = ~x121 & n134;
  assign n136 = ~x118 & ~x119;
  assign n137 = ~x117 & n136;
  assign n138 = ~x116 & ~x120;
  assign n139 = n137 & n138;
  assign n140 = n135 & n139;
  assign n141 = ~x115 & n140;
  assign n142 = ~x111 & ~x112;
  assign n143 = ~x113 & ~x114;
  assign n144 = n142 & n143;
  assign n145 = n141 & n144;
  assign n146 = ~x110 & n145;
  assign n147 = ~x109 & n146;
  assign n148 = ~x104 & ~x105;
  assign n149 = ~x108 & n148;
  assign n150 = ~x106 & ~x107;
  assign n151 = n149 & n150;
  assign n152 = n147 & n151;
  assign n153 = ~x103 & n152;
  assign n154 = ~x102 & n153;
  assign n155 = ~x101 & n154;
  assign n156 = ~x97 & ~x98;
  assign n157 = ~x99 & ~x100;
  assign n158 = n156 & n157;
  assign n159 = ~x96 & n158;
  assign n160 = n155 & n159;
  assign n161 = ~x95 & n160;
  assign n162 = ~x94 & n161;
  assign n163 = ~x93 & n162;
  assign n164 = ~x92 & n163;
  assign n165 = ~x91 & n164;
  assign n166 = ~x90 & n165;
  assign n167 = ~x89 & n166;
  assign n168 = ~x88 & n167;
  assign n169 = ~x85 & ~x86;
  assign n170 = ~x84 & ~x87;
  assign n171 = n169 & n170;
  assign n172 = n168 & n171;
  assign n173 = ~x83 & n172;
  assign n174 = ~x82 & n173;
  assign n175 = ~x81 & n174;
  assign n176 = ~x80 & n175;
  assign n177 = ~x79 & n176;
  assign n178 = ~x78 & n177;
  assign n179 = ~x77 & n178;
  assign n180 = ~x76 & n179;
  assign n181 = ~x75 & n180;
  assign n182 = ~x74 & n181;
  assign n183 = ~x73 & n182;
  assign n184 = ~x72 & n183;
  assign n185 = ~x71 & n184;
  assign n186 = ~x70 & n185;
  assign n187 = ~x69 & n186;
  assign n188 = ~x68 & n187;
  assign n189 = ~x67 & n188;
  assign n190 = ~x63 & x65;
  assign n191 = ~x66 & ~n190;
  assign n192 = n189 & n191;
  assign n193 = ~x61 & x65;
  assign n194 = x62 & ~n193;
  assign n195 = ~n192 & n194;
  assign n196 = x61 & ~x65;
  assign n197 = x64 & ~n196;
  assign n198 = ~x62 & x65;
  assign n199 = ~n197 & ~n198;
  assign n200 = ~n195 & ~n199;
  assign n201 = x64 & ~n198;
  assign n202 = ~x64 & x65;
  assign n203 = ~x66 & ~n202;
  assign n204 = ~n201 & n203;
  assign n205 = n204 ^ x66;
  assign n206 = ~n200 & n205;
  assign n207 = n206 ^ x66;
  assign n208 = n189 & ~n207;
  assign n209 = x63 & ~n208;
  assign n210 = n189 & n209;
  assign n211 = x63 & n204;
  assign n212 = n200 & ~n211;
  assign n213 = ~x63 & x66;
  assign n214 = n189 & ~n213;
  assign n215 = ~n212 & n214;
  assign n216 = n215 ^ x61;
  assign n217 = ~x60 & x65;
  assign n218 = n216 & ~n217;
  assign n219 = x64 & ~x65;
  assign n220 = x60 & n219;
  assign n221 = n220 ^ x64;
  assign n222 = ~n218 & n221;
  assign n223 = x64 & n215;
  assign n224 = n193 & ~n223;
  assign n225 = ~n222 & ~n224;
  assign n226 = n225 ^ x66;
  assign n227 = x65 & n215;
  assign n228 = x64 & n192;
  assign n229 = x62 & ~n228;
  assign n230 = ~n227 & ~n229;
  assign n231 = n192 ^ x65;
  assign n232 = x64 & ~n231;
  assign n233 = n232 ^ x65;
  assign n234 = ~n196 & n233;
  assign n235 = n215 & n234;
  assign n236 = n192 & n193;
  assign n237 = ~n235 & ~n236;
  assign n238 = ~n230 & n237;
  assign n239 = n238 ^ n225;
  assign n240 = ~n226 & ~n239;
  assign n241 = n240 ^ x66;
  assign n242 = n210 & ~n241;
  assign n243 = ~x49 & x64;
  assign n244 = ~x63 & x67;
  assign n245 = n188 & ~n244;
  assign n246 = ~n241 & n245;
  assign n247 = ~n210 & ~n246;
  assign n248 = x65 & ~n247;
  assign n249 = n223 & ~n248;
  assign n250 = ~n219 & ~n227;
  assign n251 = ~x60 & ~n250;
  assign n252 = ~n202 & ~n251;
  assign n253 = x60 & ~n227;
  assign n254 = x65 & n253;
  assign n255 = n252 & ~n254;
  assign n256 = ~n247 & ~n255;
  assign n257 = ~n249 & ~n256;
  assign n258 = n257 ^ x61;
  assign n259 = n258 ^ x66;
  assign n260 = n247 ^ x60;
  assign n261 = ~x59 & x65;
  assign n262 = ~n260 & ~n261;
  assign n263 = x59 & ~x65;
  assign n264 = x64 & ~n263;
  assign n265 = ~n262 & n264;
  assign n266 = x64 & ~n247;
  assign n267 = n217 & ~n266;
  assign n268 = ~n265 & ~n267;
  assign n269 = n268 ^ n258;
  assign n270 = n259 & n269;
  assign n271 = n270 ^ x66;
  assign n272 = n271 ^ x67;
  assign n273 = ~n226 & ~n247;
  assign n274 = n273 ^ n238;
  assign n275 = n274 ^ n271;
  assign n276 = n272 & n275;
  assign n277 = n276 ^ x67;
  assign n278 = n277 ^ x68;
  assign n279 = n241 ^ x67;
  assign n280 = n188 & n279;
  assign n281 = n209 & ~n280;
  assign n282 = n281 ^ n277;
  assign n283 = n278 & n282;
  assign n284 = n283 ^ x68;
  assign n285 = n187 & ~n284;
  assign n286 = x64 & n285;
  assign n287 = n272 & n285;
  assign n288 = n287 ^ n274;
  assign n289 = x68 & ~n288;
  assign n290 = x59 & ~n248;
  assign n291 = n285 & ~n290;
  assign n292 = n266 & ~n291;
  assign n293 = n219 ^ x65;
  assign n294 = n247 & n293;
  assign n295 = n294 ^ x65;
  assign n296 = ~x59 & n295;
  assign n297 = ~n202 & ~n296;
  assign n298 = x65 & n290;
  assign n299 = n297 & ~n298;
  assign n300 = n285 & ~n299;
  assign n301 = ~n292 & ~n300;
  assign n302 = n301 ^ x60;
  assign n303 = n302 ^ x66;
  assign n304 = ~x65 & n285;
  assign n305 = ~x58 & ~n263;
  assign n306 = ~n304 & n305;
  assign n307 = x58 & ~x65;
  assign n308 = x59 & ~n307;
  assign n309 = n285 & n308;
  assign n310 = ~n306 & ~n309;
  assign n311 = x64 & ~n310;
  assign n312 = n261 & ~n286;
  assign n313 = ~n311 & ~n312;
  assign n314 = n313 ^ n302;
  assign n315 = n303 & n314;
  assign n316 = n315 ^ x66;
  assign n317 = n316 ^ x67;
  assign n318 = n268 ^ x66;
  assign n319 = n285 & ~n318;
  assign n320 = n319 ^ n258;
  assign n321 = n320 ^ n316;
  assign n322 = n317 & ~n321;
  assign n323 = n322 ^ x67;
  assign n324 = ~n289 & ~n323;
  assign n325 = ~x68 & n288;
  assign n326 = n278 & n281;
  assign n327 = n187 & n326;
  assign n328 = n327 ^ n281;
  assign n329 = ~x69 & n328;
  assign n330 = ~n325 & ~n329;
  assign n331 = ~n324 & n330;
  assign n332 = x69 & ~n281;
  assign n333 = n186 & ~n332;
  assign n334 = ~n331 & n333;
  assign n335 = x65 & n334;
  assign n336 = ~n286 & ~n335;
  assign n337 = x65 & n285;
  assign n338 = x58 & ~n337;
  assign n339 = ~n336 & n338;
  assign n340 = x65 ^ x64;
  assign n341 = n340 ^ x65;
  assign n342 = n285 ^ x65;
  assign n343 = n341 & ~n342;
  assign n344 = x58 & n343;
  assign n345 = n344 ^ n340;
  assign n346 = n334 & n345;
  assign n347 = n346 ^ n286;
  assign n348 = ~n339 & ~n347;
  assign n349 = n348 ^ x59;
  assign n350 = n349 ^ x66;
  assign n351 = ~x65 & n334;
  assign n352 = ~x57 & ~n307;
  assign n353 = ~n351 & n352;
  assign n354 = x57 & ~x65;
  assign n355 = x58 & ~n354;
  assign n356 = n334 & n355;
  assign n357 = ~n353 & ~n356;
  assign n358 = x64 & ~n357;
  assign n359 = x64 & n334;
  assign n360 = ~x58 & x65;
  assign n361 = ~n359 & n360;
  assign n362 = ~n358 & ~n361;
  assign n363 = n362 ^ n349;
  assign n364 = n350 & n363;
  assign n365 = n364 ^ x66;
  assign n366 = n365 ^ x67;
  assign n367 = n313 ^ x66;
  assign n368 = n334 & ~n367;
  assign n369 = n368 ^ n302;
  assign n370 = n369 ^ n365;
  assign n371 = n366 & ~n370;
  assign n372 = n371 ^ x67;
  assign n373 = n372 ^ x68;
  assign n374 = n317 & n334;
  assign n375 = n374 ^ n320;
  assign n376 = n375 ^ n372;
  assign n377 = n373 & ~n376;
  assign n378 = n377 ^ x68;
  assign n379 = n378 ^ x69;
  assign n380 = n328 & ~n334;
  assign n381 = ~n242 & ~n380;
  assign n382 = ~x70 & ~n381;
  assign n383 = n323 ^ x68;
  assign n384 = n334 & n383;
  assign n385 = n384 ^ n288;
  assign n386 = n385 ^ n378;
  assign n387 = n379 & n386;
  assign n388 = n387 ^ x69;
  assign n389 = ~n382 & n388;
  assign n390 = x70 & n381;
  assign n391 = n185 & ~n390;
  assign n392 = ~n389 & n391;
  assign n393 = n379 & n392;
  assign n394 = n393 ^ n385;
  assign n395 = ~x70 & n394;
  assign n396 = ~x65 & n392;
  assign n397 = ~x56 & ~n354;
  assign n398 = ~n396 & n397;
  assign n399 = x56 & ~x65;
  assign n400 = x57 & ~n399;
  assign n401 = n392 & n400;
  assign n402 = ~n398 & ~n401;
  assign n403 = x64 & ~n402;
  assign n404 = x64 & n392;
  assign n405 = ~x57 & x65;
  assign n406 = ~n404 & n405;
  assign n407 = ~n403 & ~n406;
  assign n408 = n407 ^ x66;
  assign n409 = x65 & n392;
  assign n410 = x57 & ~n335;
  assign n411 = n409 & n410;
  assign n412 = n293 & ~n334;
  assign n413 = n412 ^ x65;
  assign n414 = ~x57 & n413;
  assign n415 = ~n202 & ~n414;
  assign n416 = n392 & ~n415;
  assign n417 = ~n411 & ~n416;
  assign n418 = n392 & ~n410;
  assign n419 = n359 & ~n418;
  assign n420 = n417 & ~n419;
  assign n421 = n420 ^ x58;
  assign n422 = n421 ^ n407;
  assign n423 = ~n408 & n422;
  assign n424 = n423 ^ x66;
  assign n425 = n424 ^ x67;
  assign n426 = n362 ^ x66;
  assign n427 = n392 & ~n426;
  assign n428 = n427 ^ n349;
  assign n429 = n428 ^ n424;
  assign n430 = n425 & ~n429;
  assign n431 = n430 ^ x67;
  assign n432 = n431 ^ x68;
  assign n433 = n366 & n392;
  assign n434 = n433 ^ n369;
  assign n435 = n434 ^ n431;
  assign n436 = n432 & ~n435;
  assign n437 = n436 ^ x68;
  assign n438 = n437 ^ x69;
  assign n439 = n373 & n392;
  assign n440 = n439 ^ n375;
  assign n441 = n440 ^ n437;
  assign n442 = n438 & ~n441;
  assign n443 = n442 ^ x69;
  assign n444 = ~n395 & n443;
  assign n445 = x70 & ~n394;
  assign n446 = x71 & n381;
  assign n447 = ~n445 & ~n446;
  assign n448 = ~n444 & n447;
  assign n449 = x70 & ~x71;
  assign n450 = ~n381 & n449;
  assign n451 = n388 & n450;
  assign n452 = ~n448 & ~n451;
  assign n453 = n184 & ~n452;
  assign n454 = ~x65 & n453;
  assign n455 = ~x55 & ~n399;
  assign n456 = ~n454 & n455;
  assign n457 = x55 & ~x65;
  assign n458 = x56 & ~n457;
  assign n459 = n453 & n458;
  assign n460 = ~n456 & ~n459;
  assign n461 = x64 & ~n460;
  assign n462 = x64 & n453;
  assign n463 = ~x56 & x65;
  assign n464 = ~n462 & n463;
  assign n465 = ~n461 & ~n464;
  assign n466 = n465 ^ x66;
  assign n467 = x65 & n453;
  assign n468 = x56 & ~n409;
  assign n469 = n467 & n468;
  assign n470 = n293 & ~n392;
  assign n471 = n470 ^ x65;
  assign n472 = ~x56 & n471;
  assign n473 = ~n202 & ~n472;
  assign n474 = n453 & ~n473;
  assign n475 = ~n469 & ~n474;
  assign n476 = n453 & ~n468;
  assign n477 = n404 & ~n476;
  assign n478 = n475 & ~n477;
  assign n479 = n478 ^ x57;
  assign n480 = n479 ^ n465;
  assign n481 = ~n466 & n480;
  assign n482 = n481 ^ x66;
  assign n483 = n482 ^ x67;
  assign n484 = ~n408 & n453;
  assign n485 = n484 ^ n421;
  assign n486 = n485 ^ n482;
  assign n487 = n483 & ~n486;
  assign n488 = n487 ^ x67;
  assign n489 = n488 ^ x68;
  assign n490 = n425 & n453;
  assign n491 = n490 ^ n428;
  assign n492 = n491 ^ n488;
  assign n493 = n489 & ~n492;
  assign n494 = n493 ^ x68;
  assign n495 = n494 ^ x69;
  assign n496 = n443 ^ x70;
  assign n497 = n453 & n496;
  assign n498 = n497 ^ n394;
  assign n499 = ~x71 & n498;
  assign n500 = n432 & n453;
  assign n501 = n500 ^ n434;
  assign n502 = n501 ^ n494;
  assign n503 = n495 & ~n502;
  assign n504 = n503 ^ x69;
  assign n505 = n504 ^ x70;
  assign n506 = n438 & n453;
  assign n507 = n506 ^ n440;
  assign n508 = n507 ^ n504;
  assign n509 = n505 & ~n508;
  assign n510 = n509 ^ x70;
  assign n511 = ~n499 & n510;
  assign n512 = ~n381 & ~n392;
  assign n513 = ~n453 & n512;
  assign n514 = ~n242 & ~n513;
  assign n515 = ~x72 & ~n514;
  assign n516 = x72 & ~n512;
  assign n517 = n183 & ~n516;
  assign n518 = ~n515 & n517;
  assign n519 = x71 & ~n498;
  assign n520 = n518 & ~n519;
  assign n521 = ~n511 & n520;
  assign n522 = n452 & n512;
  assign n523 = ~n242 & ~n522;
  assign n524 = n184 & ~n523;
  assign n525 = ~n521 & ~n524;
  assign n526 = n495 & ~n525;
  assign n527 = n526 ^ n501;
  assign n528 = ~x70 & ~n527;
  assign n529 = x65 & ~n525;
  assign n530 = x55 & ~n467;
  assign n531 = n529 & n530;
  assign n532 = n293 & ~n453;
  assign n533 = n532 ^ x65;
  assign n534 = ~x55 & n533;
  assign n535 = ~n202 & ~n534;
  assign n536 = ~n525 & ~n535;
  assign n537 = ~n531 & ~n536;
  assign n538 = ~n525 & ~n530;
  assign n539 = n462 & ~n538;
  assign n540 = n537 & ~n539;
  assign n541 = n540 ^ x56;
  assign n542 = n541 ^ x66;
  assign n543 = x64 & ~n525;
  assign n544 = ~x55 & x65;
  assign n545 = ~n543 & n544;
  assign n546 = ~x65 & ~n525;
  assign n547 = ~x54 & x64;
  assign n548 = ~n457 & n547;
  assign n549 = ~n546 & n548;
  assign n550 = ~n545 & ~n549;
  assign n551 = x54 & n457;
  assign n552 = n551 ^ x55;
  assign n553 = n543 & n552;
  assign n554 = n550 & ~n553;
  assign n555 = n554 ^ n541;
  assign n556 = n542 & n555;
  assign n557 = n556 ^ x66;
  assign n558 = n557 ^ x67;
  assign n559 = ~n466 & ~n525;
  assign n560 = n559 ^ n479;
  assign n561 = n560 ^ n557;
  assign n562 = n558 & ~n561;
  assign n563 = n562 ^ x67;
  assign n564 = n563 ^ x68;
  assign n565 = n483 & ~n525;
  assign n566 = n565 ^ n485;
  assign n567 = n566 ^ n563;
  assign n568 = n564 & ~n567;
  assign n569 = n568 ^ x68;
  assign n570 = n569 ^ x69;
  assign n571 = n489 & ~n525;
  assign n572 = n571 ^ n491;
  assign n573 = n572 ^ n569;
  assign n574 = n570 & ~n573;
  assign n575 = n574 ^ x69;
  assign n576 = ~n528 & n575;
  assign n577 = n505 & ~n525;
  assign n578 = n577 ^ n507;
  assign n579 = x70 & x71;
  assign n580 = ~n578 & ~n579;
  assign n581 = n576 & ~n580;
  assign n582 = x71 & n527;
  assign n583 = n575 & n582;
  assign n584 = n578 ^ x71;
  assign n585 = x70 & n527;
  assign n586 = n585 ^ n578;
  assign n587 = n584 & ~n586;
  assign n588 = n587 ^ x71;
  assign n589 = ~n583 & ~n588;
  assign n590 = ~n581 & n589;
  assign n591 = n510 ^ x71;
  assign n592 = ~n525 & n591;
  assign n593 = n592 ^ n498;
  assign n594 = ~x72 & n593;
  assign n595 = ~n184 & ~n381;
  assign n596 = ~n521 & n595;
  assign n597 = ~x73 & n596;
  assign n598 = ~n594 & ~n597;
  assign n599 = ~n590 & n598;
  assign n600 = x72 & ~n597;
  assign n601 = ~n593 & n600;
  assign n602 = x73 & ~n596;
  assign n603 = n182 & ~n602;
  assign n604 = ~n601 & n603;
  assign n605 = ~n599 & n604;
  assign n606 = x65 & n605;
  assign n607 = x54 & ~n529;
  assign n608 = n606 & n607;
  assign n609 = n293 & n525;
  assign n610 = n609 ^ x65;
  assign n611 = ~x54 & n610;
  assign n612 = ~n202 & ~n611;
  assign n613 = n605 & ~n612;
  assign n614 = ~n608 & ~n613;
  assign n615 = n605 & ~n607;
  assign n616 = n543 & ~n615;
  assign n617 = n614 & ~n616;
  assign n618 = n617 ^ x55;
  assign n619 = n618 ^ x66;
  assign n620 = ~x53 & ~x54;
  assign n621 = ~n605 & n620;
  assign n622 = ~x53 & x65;
  assign n623 = ~n621 & ~n622;
  assign n624 = x64 & ~n623;
  assign n625 = x64 & n605;
  assign n627 = x53 & ~x65;
  assign n628 = x54 & ~n627;
  assign n626 = ~x54 & x65;
  assign n629 = n628 ^ n626;
  assign n630 = ~n625 & n629;
  assign n631 = n630 ^ n628;
  assign n632 = ~n624 & ~n631;
  assign n633 = n632 ^ n618;
  assign n634 = n619 & n633;
  assign n635 = n634 ^ x66;
  assign n636 = n635 ^ x67;
  assign n637 = n554 ^ x66;
  assign n638 = n605 & ~n637;
  assign n639 = n638 ^ n541;
  assign n640 = n639 ^ n635;
  assign n641 = n636 & ~n640;
  assign n642 = n641 ^ x67;
  assign n643 = n642 ^ x68;
  assign n644 = n558 & n605;
  assign n645 = n644 ^ n560;
  assign n646 = n645 ^ n642;
  assign n647 = n643 & ~n646;
  assign n648 = n647 ^ x68;
  assign n649 = n648 ^ x69;
  assign n650 = n564 & n605;
  assign n651 = n650 ^ n566;
  assign n652 = n651 ^ n648;
  assign n653 = n649 & ~n652;
  assign n654 = n653 ^ x69;
  assign n655 = n654 ^ x70;
  assign n656 = n570 & n605;
  assign n657 = n656 ^ n572;
  assign n658 = n657 ^ n654;
  assign n659 = n655 & ~n658;
  assign n660 = n659 ^ x70;
  assign n661 = n660 ^ x71;
  assign n662 = n575 ^ x70;
  assign n663 = n605 & n662;
  assign n664 = n663 ^ n527;
  assign n665 = n664 ^ n660;
  assign n666 = n661 & ~n665;
  assign n667 = n666 ^ x71;
  assign n668 = n667 ^ x72;
  assign n669 = ~n576 & ~n585;
  assign n670 = n669 ^ x71;
  assign n671 = n605 & ~n670;
  assign n672 = n671 ^ n578;
  assign n673 = n672 ^ n667;
  assign n674 = n668 & ~n673;
  assign n675 = n674 ^ x72;
  assign n676 = ~x73 & ~n675;
  assign n677 = n590 ^ x72;
  assign n678 = n605 & ~n677;
  assign n679 = n678 ^ n593;
  assign n680 = ~n676 & ~n679;
  assign n681 = x73 & n675;
  assign n682 = n596 & ~n605;
  assign n683 = ~n242 & ~n682;
  assign n684 = x74 & n683;
  assign n685 = n181 & ~n684;
  assign n686 = ~n681 & n685;
  assign n687 = ~n680 & n686;
  assign n688 = n182 & ~n683;
  assign n689 = ~n687 & ~n688;
  assign n690 = ~x65 & ~n689;
  assign n691 = ~x52 & x64;
  assign n692 = ~n627 & n691;
  assign n693 = ~n690 & n692;
  assign n694 = x64 & ~n689;
  assign n695 = x52 & ~x65;
  assign n696 = x53 & ~n695;
  assign n697 = n696 ^ n622;
  assign n698 = n694 & n697;
  assign n699 = n698 ^ n622;
  assign n700 = ~n693 & ~n699;
  assign n701 = n700 ^ x66;
  assign n702 = ~n627 & ~n689;
  assign n703 = n625 & ~n702;
  assign n704 = n293 & ~n605;
  assign n705 = n704 ^ x65;
  assign n706 = ~x53 & n705;
  assign n707 = x53 & x65;
  assign n708 = ~n605 & n707;
  assign n709 = ~n202 & ~n708;
  assign n710 = ~n706 & n709;
  assign n711 = ~n689 & ~n710;
  assign n712 = ~n703 & ~n711;
  assign n713 = n712 ^ x54;
  assign n714 = n713 ^ n700;
  assign n715 = ~n701 & n714;
  assign n716 = n715 ^ x66;
  assign n717 = n716 ^ x67;
  assign n718 = n632 ^ x66;
  assign n719 = ~n689 & ~n718;
  assign n720 = n719 ^ n618;
  assign n721 = n720 ^ n716;
  assign n722 = n717 & ~n721;
  assign n723 = n722 ^ x67;
  assign n724 = n723 ^ x68;
  assign n725 = n636 & ~n689;
  assign n726 = n725 ^ n639;
  assign n727 = n726 ^ n723;
  assign n728 = n724 & ~n727;
  assign n729 = n728 ^ x68;
  assign n730 = n729 ^ x69;
  assign n731 = n643 & ~n689;
  assign n732 = n731 ^ n645;
  assign n733 = n732 ^ n729;
  assign n734 = n730 & ~n733;
  assign n735 = n734 ^ x69;
  assign n736 = n735 ^ x70;
  assign n737 = n649 & ~n689;
  assign n738 = n737 ^ n651;
  assign n739 = n738 ^ n735;
  assign n740 = n736 & ~n739;
  assign n741 = n740 ^ x70;
  assign n742 = n741 ^ x71;
  assign n743 = n655 & ~n689;
  assign n744 = n743 ^ n657;
  assign n745 = n744 ^ n741;
  assign n746 = n742 & ~n745;
  assign n747 = n746 ^ x71;
  assign n748 = n747 ^ x72;
  assign n749 = n661 & ~n689;
  assign n750 = n749 ^ n664;
  assign n751 = n750 ^ n747;
  assign n752 = n748 & ~n751;
  assign n753 = n752 ^ x72;
  assign n754 = n753 ^ x73;
  assign n755 = n668 & ~n689;
  assign n756 = n755 ^ n672;
  assign n757 = n756 ^ n753;
  assign n758 = n754 & ~n757;
  assign n759 = n758 ^ x73;
  assign n760 = n759 ^ x74;
  assign n761 = n675 ^ x73;
  assign n762 = ~n689 & n761;
  assign n763 = n762 ^ n679;
  assign n764 = n763 ^ n759;
  assign n765 = n760 & n764;
  assign n766 = n765 ^ x74;
  assign n767 = x75 & n766;
  assign n768 = n180 & ~n767;
  assign n769 = ~x75 & ~n766;
  assign n770 = ~n242 & ~n689;
  assign n771 = ~n683 & ~n770;
  assign n772 = ~n769 & ~n771;
  assign n773 = n768 & ~n772;
  assign n774 = n760 & n773;
  assign n775 = n774 ^ n763;
  assign n776 = ~x75 & n775;
  assign n777 = ~n768 & n771;
  assign n778 = ~x76 & n777;
  assign n779 = ~n776 & ~n778;
  assign n780 = x64 & n773;
  assign n781 = x52 & n780;
  assign n782 = ~x52 & ~n773;
  assign n783 = x52 ^ x51;
  assign n784 = ~x64 & n783;
  assign n785 = n784 ^ x51;
  assign n786 = ~n782 & n785;
  assign n787 = ~n781 & n786;
  assign n788 = x65 & ~n787;
  assign n789 = ~x51 & x64;
  assign n790 = n773 ^ x52;
  assign n791 = n789 & ~n790;
  assign n792 = ~n788 & ~n791;
  assign n793 = n792 ^ x66;
  assign n794 = ~n695 & n773;
  assign n795 = n694 & ~n794;
  assign n796 = x52 & n694;
  assign n797 = n689 & n691;
  assign n798 = n797 ^ x65;
  assign n799 = ~n796 & n798;
  assign n800 = n773 & n799;
  assign n801 = ~n795 & ~n800;
  assign n802 = n801 ^ x53;
  assign n803 = n802 ^ n792;
  assign n804 = ~n793 & n803;
  assign n805 = n804 ^ x66;
  assign n806 = n805 ^ x67;
  assign n807 = ~n701 & n773;
  assign n808 = n807 ^ n713;
  assign n809 = n808 ^ n805;
  assign n810 = n806 & ~n809;
  assign n811 = n810 ^ x67;
  assign n812 = n811 ^ x68;
  assign n813 = n717 & n773;
  assign n814 = n813 ^ n720;
  assign n815 = n814 ^ n811;
  assign n816 = n812 & ~n815;
  assign n817 = n816 ^ x68;
  assign n818 = n817 ^ x69;
  assign n819 = n724 & n773;
  assign n820 = n819 ^ n726;
  assign n821 = n820 ^ n817;
  assign n822 = n818 & ~n821;
  assign n823 = n822 ^ x69;
  assign n824 = n823 ^ x70;
  assign n825 = n730 & n773;
  assign n826 = n825 ^ n732;
  assign n827 = n826 ^ n823;
  assign n828 = n824 & ~n827;
  assign n829 = n828 ^ x70;
  assign n830 = n829 ^ x71;
  assign n831 = n736 & n773;
  assign n832 = n831 ^ n738;
  assign n833 = n832 ^ n829;
  assign n834 = n830 & ~n833;
  assign n835 = n834 ^ x71;
  assign n836 = n835 ^ x72;
  assign n837 = n742 & n773;
  assign n838 = n837 ^ n744;
  assign n839 = n838 ^ n835;
  assign n840 = n836 & ~n839;
  assign n841 = n840 ^ x72;
  assign n842 = n841 ^ x73;
  assign n843 = n748 & n773;
  assign n844 = n843 ^ n750;
  assign n845 = n844 ^ n841;
  assign n846 = n842 & ~n845;
  assign n847 = n846 ^ x73;
  assign n848 = n847 ^ x74;
  assign n849 = n754 & n773;
  assign n850 = n849 ^ n756;
  assign n851 = n850 ^ n847;
  assign n852 = n848 & ~n851;
  assign n853 = n852 ^ x74;
  assign n854 = n779 & n853;
  assign n855 = x75 & ~n778;
  assign n856 = ~n775 & n855;
  assign n857 = x76 & ~n771;
  assign n858 = n179 & ~n857;
  assign n859 = ~n856 & n858;
  assign n860 = ~n854 & n859;
  assign n861 = n853 ^ x75;
  assign n862 = n860 & n861;
  assign n863 = n862 ^ n775;
  assign n864 = ~x76 & n863;
  assign n865 = x64 & n860;
  assign n866 = x50 & ~x65;
  assign n867 = x51 & ~n866;
  assign n868 = n865 & n867;
  assign n869 = ~x50 & n789;
  assign n870 = ~n860 & n869;
  assign n871 = ~x50 & x65;
  assign n872 = x64 & n871;
  assign n873 = ~n870 & ~n872;
  assign n874 = ~n868 & n873;
  assign n875 = ~x51 & x65;
  assign n876 = ~n865 & n875;
  assign n877 = n874 & ~n876;
  assign n878 = n877 ^ x66;
  assign n879 = x65 & n773;
  assign n880 = x51 & ~n879;
  assign n881 = n860 & ~n880;
  assign n882 = n780 & ~n881;
  assign n883 = n773 ^ x65;
  assign n884 = n789 & ~n883;
  assign n885 = ~n202 & ~n884;
  assign n886 = x65 & n880;
  assign n887 = n885 & ~n886;
  assign n888 = n860 & ~n887;
  assign n889 = ~n882 & ~n888;
  assign n890 = n889 ^ x52;
  assign n891 = n890 ^ n877;
  assign n892 = ~n878 & n891;
  assign n893 = n892 ^ x66;
  assign n894 = n893 ^ x67;
  assign n895 = ~n793 & n860;
  assign n896 = n895 ^ n802;
  assign n897 = n896 ^ n893;
  assign n898 = n894 & ~n897;
  assign n899 = n898 ^ x67;
  assign n900 = n899 ^ x68;
  assign n901 = n806 & n860;
  assign n902 = n901 ^ n808;
  assign n903 = n902 ^ n899;
  assign n904 = n900 & ~n903;
  assign n905 = n904 ^ x68;
  assign n906 = n905 ^ x69;
  assign n907 = n812 & n860;
  assign n908 = n907 ^ n814;
  assign n909 = n908 ^ n905;
  assign n910 = n906 & ~n909;
  assign n911 = n910 ^ x69;
  assign n912 = n911 ^ x70;
  assign n913 = n818 & n860;
  assign n914 = n913 ^ n820;
  assign n915 = n914 ^ n911;
  assign n916 = n912 & ~n915;
  assign n917 = n916 ^ x70;
  assign n918 = n917 ^ x71;
  assign n919 = n824 & n860;
  assign n920 = n919 ^ n826;
  assign n921 = n920 ^ n917;
  assign n922 = n918 & ~n921;
  assign n923 = n922 ^ x71;
  assign n924 = n923 ^ x72;
  assign n925 = n830 & n860;
  assign n926 = n925 ^ n832;
  assign n927 = n926 ^ n923;
  assign n928 = n924 & ~n927;
  assign n929 = n928 ^ x72;
  assign n930 = n929 ^ x73;
  assign n931 = n836 & n860;
  assign n932 = n931 ^ n838;
  assign n933 = n932 ^ n929;
  assign n934 = n930 & ~n933;
  assign n935 = n934 ^ x73;
  assign n936 = n935 ^ x74;
  assign n937 = n842 & n860;
  assign n938 = n937 ^ n844;
  assign n939 = n938 ^ n935;
  assign n940 = n936 & ~n939;
  assign n941 = n940 ^ x74;
  assign n942 = n941 ^ x75;
  assign n943 = n848 & n860;
  assign n944 = n943 ^ n850;
  assign n945 = n944 ^ n941;
  assign n946 = n942 & ~n945;
  assign n947 = n946 ^ x75;
  assign n948 = ~n864 & n947;
  assign n949 = n777 & ~n860;
  assign n950 = ~n242 & ~n949;
  assign n951 = x77 & n950;
  assign n952 = x76 & ~n863;
  assign n953 = ~n951 & ~n952;
  assign n954 = ~n948 & n953;
  assign n955 = ~x77 & ~n950;
  assign n956 = ~n954 & ~n955;
  assign n957 = n178 & ~n956;
  assign n958 = n957 ^ x50;
  assign n959 = n243 & ~n958;
  assign n960 = x64 & x65;
  assign n961 = x50 & n960;
  assign n962 = n961 ^ n871;
  assign n963 = n957 & n962;
  assign n964 = n963 ^ n871;
  assign n965 = ~n959 & ~n964;
  assign n966 = x65 & n243;
  assign n967 = ~x50 & n202;
  assign n968 = ~n966 & ~n967;
  assign n969 = n965 & n968;
  assign n970 = n969 ^ x66;
  assign n971 = x65 & n178;
  assign n972 = ~n860 & n971;
  assign n973 = ~n956 & n972;
  assign n974 = n219 & n860;
  assign n975 = ~n973 & ~n974;
  assign n976 = x50 & ~n975;
  assign n977 = n860 ^ x65;
  assign n978 = n341 & ~n977;
  assign n979 = x50 & n978;
  assign n980 = n979 ^ n340;
  assign n981 = n957 & n980;
  assign n982 = n981 ^ n865;
  assign n983 = ~n976 & ~n982;
  assign n984 = n983 ^ x51;
  assign n985 = n984 ^ n969;
  assign n986 = ~n970 & n985;
  assign n987 = n986 ^ x66;
  assign n988 = n987 ^ x67;
  assign n989 = ~n878 & n957;
  assign n990 = n989 ^ n890;
  assign n991 = n990 ^ n987;
  assign n992 = n988 & ~n991;
  assign n993 = n992 ^ x67;
  assign n994 = n993 ^ x68;
  assign n995 = n894 & n957;
  assign n996 = n995 ^ n896;
  assign n997 = n996 ^ n993;
  assign n998 = n994 & ~n997;
  assign n999 = n998 ^ x68;
  assign n1000 = n999 ^ x69;
  assign n1001 = n900 & n957;
  assign n1002 = n1001 ^ n902;
  assign n1003 = n1002 ^ n999;
  assign n1004 = n1000 & ~n1003;
  assign n1005 = n1004 ^ x69;
  assign n1006 = n1005 ^ x70;
  assign n1007 = n906 & n957;
  assign n1008 = n1007 ^ n908;
  assign n1009 = n1008 ^ n1005;
  assign n1010 = n1006 & ~n1009;
  assign n1011 = n1010 ^ x70;
  assign n1012 = n1011 ^ x71;
  assign n1013 = n912 & n957;
  assign n1014 = n1013 ^ n914;
  assign n1015 = n1014 ^ n1011;
  assign n1016 = n1012 & ~n1015;
  assign n1017 = n1016 ^ x71;
  assign n1018 = n1017 ^ x72;
  assign n1019 = n918 & n957;
  assign n1020 = n1019 ^ n920;
  assign n1021 = n1020 ^ n1017;
  assign n1022 = n1018 & ~n1021;
  assign n1023 = n1022 ^ x72;
  assign n1024 = n1023 ^ x73;
  assign n1025 = n924 & n957;
  assign n1026 = n1025 ^ n926;
  assign n1027 = n1026 ^ n1023;
  assign n1028 = n1024 & ~n1027;
  assign n1029 = n1028 ^ x73;
  assign n1030 = n1029 ^ x74;
  assign n1031 = n930 & n957;
  assign n1032 = n1031 ^ n932;
  assign n1033 = n1032 ^ n1029;
  assign n1034 = n1030 & ~n1033;
  assign n1035 = n1034 ^ x74;
  assign n1036 = n1035 ^ x75;
  assign n1037 = n936 & n957;
  assign n1038 = n1037 ^ n938;
  assign n1039 = n1038 ^ n1035;
  assign n1040 = n1036 & ~n1039;
  assign n1041 = n1040 ^ x75;
  assign n1042 = n1041 ^ x76;
  assign n1043 = n942 & n957;
  assign n1044 = n1043 ^ n944;
  assign n1045 = n1044 ^ n1041;
  assign n1046 = n1042 & ~n1045;
  assign n1047 = n1046 ^ x76;
  assign n1048 = ~x77 & ~n1047;
  assign n1049 = n947 ^ x76;
  assign n1050 = n957 & n1049;
  assign n1051 = n1050 ^ n863;
  assign n1052 = ~n1048 & ~n1051;
  assign n1053 = x77 & n1047;
  assign n1054 = n949 & ~n957;
  assign n1055 = ~n242 & ~n1054;
  assign n1056 = n1055 ^ x78;
  assign n1057 = n177 & n1056;
  assign n1058 = ~n1053 & n1057;
  assign n1059 = ~n1052 & n1058;
  assign n1060 = ~n178 & n949;
  assign n1061 = ~n1059 & n1060;
  assign n1062 = n178 & ~n1055;
  assign n1063 = ~n1059 & ~n1062;
  assign n1064 = n1047 ^ x77;
  assign n1065 = ~n1063 & n1064;
  assign n1066 = n1065 ^ n1051;
  assign n1067 = ~x78 & n1066;
  assign n1068 = ~n242 & ~n1061;
  assign n1069 = ~x79 & ~n1068;
  assign n1070 = ~n1067 & ~n1069;
  assign n1071 = ~x48 & x64;
  assign n1072 = x64 & ~n1063;
  assign n1073 = n1072 ^ x49;
  assign n1074 = ~n1071 & n1073;
  assign n1075 = x65 & n1074;
  assign n1076 = n1075 ^ x65;
  assign n1077 = n1063 ^ x49;
  assign n1078 = n1071 & n1077;
  assign n1079 = ~n1076 & ~n1078;
  assign n1080 = n1079 ^ x66;
  assign n1081 = ~x49 & ~n1063;
  assign n1082 = x64 & n957;
  assign n1083 = ~n1081 & n1082;
  assign n1084 = x65 & ~n1063;
  assign n1085 = n1083 & ~n1084;
  assign n1086 = n293 & ~n957;
  assign n1087 = n1086 ^ x65;
  assign n1088 = n1081 & n1087;
  assign n1089 = x65 & ~n243;
  assign n1090 = ~n1082 & n1089;
  assign n1091 = ~n1063 & n1090;
  assign n1092 = ~n1088 & ~n1091;
  assign n1093 = ~n1085 & n1092;
  assign n1094 = n1093 ^ x50;
  assign n1095 = n1094 ^ n1079;
  assign n1096 = ~n1080 & n1095;
  assign n1097 = n1096 ^ x66;
  assign n1098 = n1097 ^ x67;
  assign n1099 = ~n970 & ~n1063;
  assign n1100 = n1099 ^ n984;
  assign n1101 = n1100 ^ n1097;
  assign n1102 = n1098 & ~n1101;
  assign n1103 = n1102 ^ x67;
  assign n1104 = n1103 ^ x68;
  assign n1105 = n988 & ~n1063;
  assign n1106 = n1105 ^ n990;
  assign n1107 = n1106 ^ n1103;
  assign n1108 = n1104 & ~n1107;
  assign n1109 = n1108 ^ x68;
  assign n1110 = n1109 ^ x69;
  assign n1111 = n994 & ~n1063;
  assign n1112 = n1111 ^ n996;
  assign n1113 = n1112 ^ n1109;
  assign n1114 = n1110 & ~n1113;
  assign n1115 = n1114 ^ x69;
  assign n1116 = n1115 ^ x70;
  assign n1117 = n1000 & ~n1063;
  assign n1118 = n1117 ^ n1002;
  assign n1119 = n1118 ^ n1115;
  assign n1120 = n1116 & ~n1119;
  assign n1121 = n1120 ^ x70;
  assign n1122 = n1121 ^ x71;
  assign n1123 = n1006 & ~n1063;
  assign n1124 = n1123 ^ n1008;
  assign n1125 = n1124 ^ n1121;
  assign n1126 = n1122 & ~n1125;
  assign n1127 = n1126 ^ x71;
  assign n1128 = n1127 ^ x72;
  assign n1129 = n1012 & ~n1063;
  assign n1130 = n1129 ^ n1014;
  assign n1131 = n1130 ^ n1127;
  assign n1132 = n1128 & ~n1131;
  assign n1133 = n1132 ^ x72;
  assign n1134 = n1133 ^ x73;
  assign n1135 = n1018 & ~n1063;
  assign n1136 = n1135 ^ n1020;
  assign n1137 = n1136 ^ n1133;
  assign n1138 = n1134 & ~n1137;
  assign n1139 = n1138 ^ x73;
  assign n1140 = n1139 ^ x74;
  assign n1141 = n1024 & ~n1063;
  assign n1142 = n1141 ^ n1026;
  assign n1143 = n1142 ^ n1139;
  assign n1144 = n1140 & ~n1143;
  assign n1145 = n1144 ^ x74;
  assign n1146 = n1145 ^ x75;
  assign n1147 = n1030 & ~n1063;
  assign n1148 = n1147 ^ n1032;
  assign n1149 = n1148 ^ n1145;
  assign n1150 = n1146 & ~n1149;
  assign n1151 = n1150 ^ x75;
  assign n1152 = n1151 ^ x76;
  assign n1153 = n1036 & ~n1063;
  assign n1154 = n1153 ^ n1038;
  assign n1155 = n1154 ^ n1151;
  assign n1156 = n1152 & ~n1155;
  assign n1157 = n1156 ^ x76;
  assign n1158 = n1157 ^ x77;
  assign n1159 = n1042 & ~n1063;
  assign n1160 = n1159 ^ n1044;
  assign n1161 = n1160 ^ n1157;
  assign n1162 = n1158 & ~n1161;
  assign n1163 = n1162 ^ x77;
  assign n1164 = n1070 & n1163;
  assign n1165 = x78 & ~n1069;
  assign n1166 = ~n1066 & n1165;
  assign n1167 = n176 & ~n1068;
  assign n1168 = ~n177 & ~n1167;
  assign n1169 = ~n1166 & ~n1168;
  assign n1170 = ~n1164 & n1169;
  assign n1171 = n1061 & ~n1170;
  assign n1172 = ~n242 & ~n1171;
  assign n1173 = ~x80 & ~n1172;
  assign n1174 = n1163 ^ x78;
  assign n1175 = n1170 & n1174;
  assign n1176 = n1175 ^ n1066;
  assign n1177 = ~n1173 & ~n1176;
  assign n1178 = x79 & x80;
  assign n1179 = ~n1177 & ~n1178;
  assign n1180 = ~x47 & n1071;
  assign n1181 = ~n1170 & n1180;
  assign n1182 = ~x47 & x65;
  assign n1183 = x64 & n1182;
  assign n1184 = ~n1181 & ~n1183;
  assign n1185 = x64 & n1170;
  assign n1187 = x47 & ~x65;
  assign n1188 = x48 & ~n1187;
  assign n1186 = ~x48 & x65;
  assign n1189 = n1188 ^ n1186;
  assign n1190 = ~n1185 & n1189;
  assign n1191 = n1190 ^ n1188;
  assign n1192 = n1184 & ~n1191;
  assign n1193 = ~x66 & n1192;
  assign n1194 = x48 & ~n1084;
  assign n1195 = n1170 & ~n1194;
  assign n1196 = n1072 & ~n1195;
  assign n1197 = n1063 ^ x65;
  assign n1198 = n1071 & n1197;
  assign n1199 = ~n202 & ~n1198;
  assign n1200 = x65 & n1194;
  assign n1201 = n1199 & ~n1200;
  assign n1202 = n1170 & ~n1201;
  assign n1203 = ~n1196 & ~n1202;
  assign n1204 = n1203 ^ x49;
  assign n1205 = ~n1193 & n1204;
  assign n1206 = x66 & ~n1192;
  assign n1207 = ~n1080 & n1170;
  assign n1208 = n1207 ^ n1094;
  assign n1209 = x67 & n1208;
  assign n1210 = ~n1206 & ~n1209;
  assign n1211 = ~n1205 & n1210;
  assign n1212 = ~x67 & ~n1208;
  assign n1213 = ~n1211 & ~n1212;
  assign n1214 = n1213 ^ x68;
  assign n1215 = n1098 & n1170;
  assign n1216 = n1215 ^ n1100;
  assign n1217 = n1216 ^ n1213;
  assign n1218 = n1214 & ~n1217;
  assign n1219 = n1218 ^ x68;
  assign n1220 = n1219 ^ x69;
  assign n1221 = n1104 & n1170;
  assign n1222 = n1221 ^ n1106;
  assign n1223 = n1222 ^ n1219;
  assign n1224 = n1220 & ~n1223;
  assign n1225 = n1224 ^ x69;
  assign n1226 = n1225 ^ x70;
  assign n1227 = n1110 & n1170;
  assign n1228 = n1227 ^ n1112;
  assign n1229 = n1228 ^ n1225;
  assign n1230 = n1226 & ~n1229;
  assign n1231 = n1230 ^ x70;
  assign n1232 = n1231 ^ x71;
  assign n1233 = n1116 & n1170;
  assign n1234 = n1233 ^ n1118;
  assign n1235 = n1234 ^ n1231;
  assign n1236 = n1232 & ~n1235;
  assign n1237 = n1236 ^ x71;
  assign n1238 = n1237 ^ x72;
  assign n1239 = n1122 & n1170;
  assign n1240 = n1239 ^ n1124;
  assign n1241 = n1240 ^ n1237;
  assign n1242 = n1238 & ~n1241;
  assign n1243 = n1242 ^ x72;
  assign n1244 = n1243 ^ x73;
  assign n1245 = n1128 & n1170;
  assign n1246 = n1245 ^ n1130;
  assign n1247 = n1246 ^ n1243;
  assign n1248 = n1244 & ~n1247;
  assign n1249 = n1248 ^ x73;
  assign n1250 = n1249 ^ x74;
  assign n1251 = n1134 & n1170;
  assign n1252 = n1251 ^ n1136;
  assign n1253 = n1252 ^ n1249;
  assign n1254 = n1250 & ~n1253;
  assign n1255 = n1254 ^ x74;
  assign n1256 = n1255 ^ x75;
  assign n1257 = n1140 & n1170;
  assign n1258 = n1257 ^ n1142;
  assign n1259 = n1258 ^ n1255;
  assign n1260 = n1256 & ~n1259;
  assign n1261 = n1260 ^ x75;
  assign n1262 = n1261 ^ x76;
  assign n1263 = n1146 & n1170;
  assign n1264 = n1263 ^ n1148;
  assign n1265 = n1264 ^ n1261;
  assign n1266 = n1262 & ~n1265;
  assign n1267 = n1266 ^ x76;
  assign n1268 = n1267 ^ x77;
  assign n1269 = n1152 & n1170;
  assign n1270 = n1269 ^ n1154;
  assign n1271 = n1270 ^ n1267;
  assign n1272 = n1268 & ~n1271;
  assign n1273 = n1272 ^ x77;
  assign n1274 = n1273 ^ x78;
  assign n1275 = n1158 & n1170;
  assign n1276 = n1275 ^ n1160;
  assign n1277 = n1276 ^ n1273;
  assign n1278 = n1274 & ~n1277;
  assign n1279 = n1278 ^ x78;
  assign n1280 = ~n1179 & n1279;
  assign n1281 = x79 & n1177;
  assign n1282 = x80 & n1172;
  assign n1283 = ~n1281 & ~n1282;
  assign n1284 = ~n1280 & n1283;
  assign n1285 = x79 & n1172;
  assign n1286 = n1279 & n1285;
  assign n1287 = n1284 & ~n1286;
  assign n1288 = n175 & n1287;
  assign n1289 = ~n242 & n1288;
  assign n1290 = ~n1172 & ~n1289;
  assign n1291 = n1290 ^ x81;
  assign n1292 = n174 & ~n1291;
  assign n1293 = ~x46 & ~x47;
  assign n1294 = ~n1288 & n1293;
  assign n1295 = ~x46 & x65;
  assign n1296 = ~n1294 & ~n1295;
  assign n1297 = x64 & ~n1296;
  assign n1298 = x64 & n1288;
  assign n1299 = x46 & ~x65;
  assign n1300 = x47 & ~n1299;
  assign n1301 = n1300 ^ n1182;
  assign n1302 = n1298 & n1301;
  assign n1303 = n1302 ^ n1182;
  assign n1304 = ~n1297 & ~n1303;
  assign n1305 = n1304 ^ x66;
  assign n1306 = x65 & n175;
  assign n1307 = ~n1170 & n1306;
  assign n1308 = n1287 & n1307;
  assign n1309 = n219 & n1170;
  assign n1310 = ~n1308 & ~n1309;
  assign n1311 = x47 & ~n1310;
  assign n1312 = n1170 ^ x65;
  assign n1313 = n341 & ~n1312;
  assign n1314 = x47 & n1313;
  assign n1315 = n1314 ^ n340;
  assign n1316 = n1288 & n1315;
  assign n1317 = n1316 ^ n1185;
  assign n1318 = ~n1311 & ~n1317;
  assign n1319 = n1318 ^ x48;
  assign n1320 = n1319 ^ n1304;
  assign n1321 = ~n1305 & n1320;
  assign n1322 = n1321 ^ x66;
  assign n1323 = n1322 ^ x67;
  assign n1324 = n1192 ^ x66;
  assign n1325 = n1288 & ~n1324;
  assign n1326 = n1325 ^ n1204;
  assign n1327 = n1326 ^ n1322;
  assign n1328 = n1323 & ~n1327;
  assign n1329 = n1328 ^ x67;
  assign n1330 = n1329 ^ x68;
  assign n1331 = ~n1205 & ~n1206;
  assign n1332 = n1331 ^ x67;
  assign n1333 = n1288 & ~n1332;
  assign n1334 = n1333 ^ n1208;
  assign n1335 = n1334 ^ n1329;
  assign n1336 = n1330 & ~n1335;
  assign n1337 = n1336 ^ x68;
  assign n1338 = n1337 ^ x69;
  assign n1339 = n1214 & n1288;
  assign n1340 = n1339 ^ n1216;
  assign n1341 = n1340 ^ n1337;
  assign n1342 = n1338 & ~n1341;
  assign n1343 = n1342 ^ x69;
  assign n1344 = n1343 ^ x70;
  assign n1345 = n1220 & n1288;
  assign n1346 = n1345 ^ n1222;
  assign n1347 = n1346 ^ n1343;
  assign n1348 = n1344 & ~n1347;
  assign n1349 = n1348 ^ x70;
  assign n1350 = n1349 ^ x71;
  assign n1351 = n1226 & n1288;
  assign n1352 = n1351 ^ n1228;
  assign n1353 = n1352 ^ n1349;
  assign n1354 = n1350 & ~n1353;
  assign n1355 = n1354 ^ x71;
  assign n1356 = n1355 ^ x72;
  assign n1357 = n1232 & n1288;
  assign n1358 = n1357 ^ n1234;
  assign n1359 = n1358 ^ n1355;
  assign n1360 = n1356 & ~n1359;
  assign n1361 = n1360 ^ x72;
  assign n1362 = n1361 ^ x73;
  assign n1363 = n1238 & n1288;
  assign n1364 = n1363 ^ n1240;
  assign n1365 = n1364 ^ n1361;
  assign n1366 = n1362 & ~n1365;
  assign n1367 = n1366 ^ x73;
  assign n1368 = n1367 ^ x74;
  assign n1369 = n1244 & n1288;
  assign n1370 = n1369 ^ n1246;
  assign n1371 = n1370 ^ n1367;
  assign n1372 = n1368 & ~n1371;
  assign n1373 = n1372 ^ x74;
  assign n1374 = n1373 ^ x75;
  assign n1375 = n1250 & n1288;
  assign n1376 = n1375 ^ n1252;
  assign n1377 = n1376 ^ n1373;
  assign n1378 = n1374 & ~n1377;
  assign n1379 = n1378 ^ x75;
  assign n1380 = n1379 ^ x76;
  assign n1381 = n1256 & n1288;
  assign n1382 = n1381 ^ n1258;
  assign n1383 = n1382 ^ n1379;
  assign n1384 = n1380 & ~n1383;
  assign n1385 = n1384 ^ x76;
  assign n1386 = n1385 ^ x77;
  assign n1387 = n1262 & n1288;
  assign n1388 = n1387 ^ n1264;
  assign n1389 = n1388 ^ n1385;
  assign n1390 = n1386 & ~n1389;
  assign n1391 = n1390 ^ x77;
  assign n1392 = n1391 ^ x78;
  assign n1393 = n1268 & n1288;
  assign n1394 = n1393 ^ n1270;
  assign n1395 = n1394 ^ n1391;
  assign n1396 = n1392 & ~n1395;
  assign n1397 = n1396 ^ x78;
  assign n1398 = n1397 ^ x79;
  assign n1399 = n1274 & n1288;
  assign n1400 = n1399 ^ n1276;
  assign n1401 = n1400 ^ n1397;
  assign n1402 = n1398 & ~n1401;
  assign n1403 = n1402 ^ x79;
  assign n1404 = n1403 ^ x80;
  assign n1405 = n1279 ^ x79;
  assign n1406 = n1288 & n1405;
  assign n1407 = n1406 ^ n1176;
  assign n1408 = n1407 ^ n1403;
  assign n1409 = n1404 & n1408;
  assign n1410 = n1409 ^ x80;
  assign n1411 = n1292 & ~n1410;
  assign n1412 = ~n175 & n1171;
  assign n1413 = ~n1411 & n1412;
  assign n1414 = n175 & n1290;
  assign n1415 = ~n1411 & ~n1414;
  assign n1416 = n1404 & ~n1415;
  assign n1417 = n1416 ^ n1407;
  assign n1418 = x81 & ~n1417;
  assign n1419 = n1323 & ~n1415;
  assign n1420 = n1419 ^ n1326;
  assign n1421 = ~x68 & ~n1420;
  assign n1422 = n1330 & ~n1415;
  assign n1423 = n1422 ^ n1334;
  assign n1424 = ~x69 & ~n1423;
  assign n1425 = ~n1421 & ~n1424;
  assign n1426 = x64 & ~n1415;
  assign n1427 = x46 & n1426;
  assign n1428 = ~x46 & n1415;
  assign n1429 = ~x45 & x64;
  assign n1430 = ~x46 & ~x64;
  assign n1431 = ~n1429 & ~n1430;
  assign n1432 = ~n1428 & n1431;
  assign n1433 = ~n1427 & n1432;
  assign n1434 = x65 & ~n1433;
  assign n1435 = n1415 ^ x46;
  assign n1436 = n1429 & n1435;
  assign n1437 = ~n1434 & ~n1436;
  assign n1438 = n1437 ^ x66;
  assign n1439 = ~n1299 & ~n1415;
  assign n1440 = n1298 & ~n1439;
  assign n1441 = x65 ^ x46;
  assign n1442 = ~n1430 & ~n1441;
  assign n1443 = ~n1288 & n1442;
  assign n1444 = ~n202 & ~n1443;
  assign n1445 = n1288 & n1295;
  assign n1446 = n1444 & ~n1445;
  assign n1447 = ~n1415 & ~n1446;
  assign n1448 = ~n1440 & ~n1447;
  assign n1449 = n1448 ^ x47;
  assign n1450 = n1449 ^ n1437;
  assign n1451 = ~n1438 & n1450;
  assign n1452 = n1451 ^ x66;
  assign n1453 = n1452 ^ x67;
  assign n1454 = ~n1305 & ~n1415;
  assign n1455 = n1454 ^ n1319;
  assign n1456 = n1455 ^ n1452;
  assign n1457 = n1453 & ~n1456;
  assign n1458 = n1457 ^ x67;
  assign n1459 = n1425 & n1458;
  assign n1460 = n1423 ^ x69;
  assign n1461 = x68 & n1420;
  assign n1462 = n1461 ^ n1423;
  assign n1463 = n1460 & ~n1462;
  assign n1464 = n1463 ^ x69;
  assign n1465 = ~n1459 & ~n1464;
  assign n1466 = n1465 ^ x70;
  assign n1467 = n1338 & ~n1415;
  assign n1468 = n1467 ^ n1340;
  assign n1469 = n1468 ^ n1465;
  assign n1470 = ~n1466 & n1469;
  assign n1471 = n1470 ^ x70;
  assign n1472 = n1471 ^ x71;
  assign n1473 = n1344 & ~n1415;
  assign n1474 = n1473 ^ n1346;
  assign n1475 = n1474 ^ n1471;
  assign n1476 = n1472 & ~n1475;
  assign n1477 = n1476 ^ x71;
  assign n1478 = n1477 ^ x72;
  assign n1479 = n1350 & ~n1415;
  assign n1480 = n1479 ^ n1352;
  assign n1481 = n1480 ^ n1477;
  assign n1482 = n1478 & ~n1481;
  assign n1483 = n1482 ^ x72;
  assign n1484 = n1483 ^ x73;
  assign n1485 = n1356 & ~n1415;
  assign n1486 = n1485 ^ n1358;
  assign n1487 = n1486 ^ n1483;
  assign n1488 = n1484 & ~n1487;
  assign n1489 = n1488 ^ x73;
  assign n1490 = n1489 ^ x74;
  assign n1491 = n1362 & ~n1415;
  assign n1492 = n1491 ^ n1364;
  assign n1493 = n1492 ^ n1489;
  assign n1494 = n1490 & ~n1493;
  assign n1495 = n1494 ^ x74;
  assign n1496 = n1495 ^ x75;
  assign n1497 = n1368 & ~n1415;
  assign n1498 = n1497 ^ n1370;
  assign n1499 = n1498 ^ n1495;
  assign n1500 = n1496 & ~n1499;
  assign n1501 = n1500 ^ x75;
  assign n1502 = n1501 ^ x76;
  assign n1503 = n1374 & ~n1415;
  assign n1504 = n1503 ^ n1376;
  assign n1505 = n1504 ^ n1501;
  assign n1506 = n1502 & ~n1505;
  assign n1507 = n1506 ^ x76;
  assign n1508 = n1507 ^ x77;
  assign n1509 = n1380 & ~n1415;
  assign n1510 = n1509 ^ n1382;
  assign n1511 = n1510 ^ n1507;
  assign n1512 = n1508 & ~n1511;
  assign n1513 = n1512 ^ x77;
  assign n1514 = n1513 ^ x78;
  assign n1515 = n1386 & ~n1415;
  assign n1516 = n1515 ^ n1388;
  assign n1517 = n1516 ^ n1513;
  assign n1518 = n1514 & ~n1517;
  assign n1519 = n1518 ^ x78;
  assign n1520 = n1519 ^ x79;
  assign n1521 = n1392 & ~n1415;
  assign n1522 = n1521 ^ n1394;
  assign n1523 = n1522 ^ n1519;
  assign n1524 = n1520 & ~n1523;
  assign n1525 = n1524 ^ x79;
  assign n1526 = n1525 ^ x80;
  assign n1527 = n1398 & ~n1415;
  assign n1528 = n1527 ^ n1400;
  assign n1529 = n1528 ^ n1525;
  assign n1530 = n1526 & ~n1529;
  assign n1531 = n1530 ^ x80;
  assign n1532 = ~n1418 & ~n1531;
  assign n1533 = ~x81 & n1417;
  assign n1534 = ~n242 & ~n1413;
  assign n1535 = ~x82 & ~n1534;
  assign n1536 = ~n1533 & ~n1535;
  assign n1537 = ~n1532 & n1536;
  assign n1538 = x82 & n1534;
  assign n1539 = ~n1537 & ~n1538;
  assign n1540 = n173 & n1539;
  assign n1541 = n1413 & ~n1540;
  assign n1542 = ~n242 & ~n1541;
  assign n1543 = n1531 ^ x81;
  assign n1544 = n1540 & n1543;
  assign n1545 = n1544 ^ n1417;
  assign n1546 = ~x82 & n1545;
  assign n1547 = x65 & n1415;
  assign n1548 = n173 & n1547;
  assign n1549 = n1539 & n1548;
  assign n1550 = n219 & ~n1415;
  assign n1551 = ~n1549 & ~n1550;
  assign n1552 = x45 & ~n1551;
  assign n1553 = n1415 ^ x65;
  assign n1554 = n341 & n1553;
  assign n1555 = x45 & n1554;
  assign n1556 = n1555 ^ n340;
  assign n1557 = n1540 & n1556;
  assign n1558 = n1557 ^ n1426;
  assign n1559 = ~n1552 & ~n1558;
  assign n1560 = n1559 ^ x46;
  assign n1561 = n1560 ^ x66;
  assign n1562 = x64 & n1540;
  assign n1563 = x44 & ~x65;
  assign n1564 = x45 & ~n1563;
  assign n1565 = n1562 & n1564;
  assign n1566 = ~x44 & n1429;
  assign n1567 = ~x45 & x65;
  assign n1568 = ~n1566 & ~n1567;
  assign n1569 = ~n1540 & ~n1568;
  assign n1570 = ~x44 & x65;
  assign n1571 = n1570 ^ n1567;
  assign n1572 = x64 & n1571;
  assign n1573 = n1572 ^ n1567;
  assign n1574 = ~n1569 & ~n1573;
  assign n1575 = ~n1565 & n1574;
  assign n1576 = n1575 ^ n1560;
  assign n1577 = n1561 & n1576;
  assign n1578 = n1577 ^ x66;
  assign n1579 = n1578 ^ x67;
  assign n1580 = ~n1438 & n1540;
  assign n1581 = n1580 ^ n1449;
  assign n1582 = n1581 ^ n1578;
  assign n1583 = n1579 & ~n1582;
  assign n1584 = n1583 ^ x67;
  assign n1585 = n1584 ^ x68;
  assign n1586 = n1453 & n1540;
  assign n1587 = n1586 ^ n1455;
  assign n1588 = n1587 ^ n1584;
  assign n1589 = n1585 & ~n1588;
  assign n1590 = n1589 ^ x68;
  assign n1591 = n1590 ^ x69;
  assign n1592 = n1458 ^ x68;
  assign n1593 = n1540 & n1592;
  assign n1594 = n1593 ^ n1420;
  assign n1595 = n1594 ^ n1590;
  assign n1596 = n1591 & ~n1595;
  assign n1597 = n1596 ^ x69;
  assign n1598 = n1597 ^ x70;
  assign n1599 = n1458 ^ n1420;
  assign n1600 = n1592 & ~n1599;
  assign n1601 = n1600 ^ x68;
  assign n1602 = n1601 ^ x69;
  assign n1603 = n1540 & n1602;
  assign n1604 = n1603 ^ n1423;
  assign n1605 = n1604 ^ n1597;
  assign n1606 = n1598 & ~n1605;
  assign n1607 = n1606 ^ x70;
  assign n1608 = n1607 ^ x71;
  assign n1609 = ~n1466 & n1540;
  assign n1610 = n1609 ^ n1468;
  assign n1611 = n1610 ^ n1607;
  assign n1612 = n1608 & ~n1611;
  assign n1613 = n1612 ^ x71;
  assign n1614 = n1613 ^ x72;
  assign n1615 = n1472 & n1540;
  assign n1616 = n1615 ^ n1474;
  assign n1617 = n1616 ^ n1613;
  assign n1618 = n1614 & ~n1617;
  assign n1619 = n1618 ^ x72;
  assign n1620 = n1619 ^ x73;
  assign n1621 = n1478 & n1540;
  assign n1622 = n1621 ^ n1480;
  assign n1623 = n1622 ^ n1619;
  assign n1624 = n1620 & ~n1623;
  assign n1625 = n1624 ^ x73;
  assign n1626 = n1625 ^ x74;
  assign n1627 = n1484 & n1540;
  assign n1628 = n1627 ^ n1486;
  assign n1629 = n1628 ^ n1625;
  assign n1630 = n1626 & ~n1629;
  assign n1631 = n1630 ^ x74;
  assign n1632 = n1631 ^ x75;
  assign n1633 = n1490 & n1540;
  assign n1634 = n1633 ^ n1492;
  assign n1635 = n1634 ^ n1631;
  assign n1636 = n1632 & ~n1635;
  assign n1637 = n1636 ^ x75;
  assign n1638 = n1637 ^ x76;
  assign n1639 = n1496 & n1540;
  assign n1640 = n1639 ^ n1498;
  assign n1641 = n1640 ^ n1637;
  assign n1642 = n1638 & ~n1641;
  assign n1643 = n1642 ^ x76;
  assign n1644 = n1643 ^ x77;
  assign n1645 = n1502 & n1540;
  assign n1646 = n1645 ^ n1504;
  assign n1647 = n1646 ^ n1643;
  assign n1648 = n1644 & ~n1647;
  assign n1649 = n1648 ^ x77;
  assign n1650 = n1649 ^ x78;
  assign n1651 = n1508 & n1540;
  assign n1652 = n1651 ^ n1510;
  assign n1653 = n1652 ^ n1649;
  assign n1654 = n1650 & ~n1653;
  assign n1655 = n1654 ^ x78;
  assign n1656 = n1655 ^ x79;
  assign n1657 = n1514 & n1540;
  assign n1658 = n1657 ^ n1516;
  assign n1659 = n1658 ^ n1655;
  assign n1660 = n1656 & ~n1659;
  assign n1661 = n1660 ^ x79;
  assign n1662 = n1661 ^ x80;
  assign n1663 = n1520 & n1540;
  assign n1664 = n1663 ^ n1522;
  assign n1665 = n1664 ^ n1661;
  assign n1666 = n1662 & ~n1665;
  assign n1667 = n1666 ^ x80;
  assign n1668 = n1667 ^ x81;
  assign n1669 = n1526 & n1540;
  assign n1670 = n1669 ^ n1528;
  assign n1671 = n1670 ^ n1667;
  assign n1672 = n1668 & ~n1671;
  assign n1673 = n1672 ^ x81;
  assign n1674 = ~n1546 & n1673;
  assign n1675 = x83 & n1542;
  assign n1676 = x82 & ~n1545;
  assign n1677 = ~n1675 & ~n1676;
  assign n1678 = ~n1674 & n1677;
  assign n1679 = ~x83 & ~n1542;
  assign n1680 = ~n1678 & ~n1679;
  assign n1681 = n172 & ~n1680;
  assign n1682 = ~n242 & n1681;
  assign n1683 = ~n1542 & ~n1682;
  assign n1684 = x85 & ~n1683;
  assign n1685 = x65 & ~n1540;
  assign n1686 = n1681 & n1685;
  assign n1687 = ~x65 & n1540;
  assign n1688 = x64 & n1687;
  assign n1689 = ~n1686 & ~n1688;
  assign n1690 = x44 & ~n1689;
  assign n1691 = n1540 ^ x65;
  assign n1692 = n341 & ~n1691;
  assign n1693 = x44 & n1692;
  assign n1694 = n1693 ^ n340;
  assign n1695 = n1681 & n1694;
  assign n1696 = n1695 ^ n1562;
  assign n1697 = ~n1690 & ~n1696;
  assign n1698 = n1697 ^ x45;
  assign n1699 = ~x43 & ~x44;
  assign n1700 = ~n1681 & n1699;
  assign n1701 = ~x43 & x65;
  assign n1702 = ~n1700 & ~n1701;
  assign n1703 = x64 & ~n1702;
  assign n1704 = x64 & n1681;
  assign n1705 = x43 & n1563;
  assign n1706 = n1705 ^ x44;
  assign n1707 = n1706 ^ n1570;
  assign n1708 = n1704 & n1707;
  assign n1709 = n1708 ^ n1570;
  assign n1710 = ~n1703 & ~n1709;
  assign n1711 = ~x66 & n1710;
  assign n1712 = n1698 & ~n1711;
  assign n1713 = n1575 ^ x66;
  assign n1714 = n1681 & ~n1713;
  assign n1715 = n1714 ^ n1560;
  assign n1716 = n1712 & n1715;
  assign n1717 = x67 & ~n1710;
  assign n1718 = n1698 & n1717;
  assign n1719 = x66 & ~n1710;
  assign n1720 = ~x67 & ~n1715;
  assign n1721 = n1719 & ~n1720;
  assign n1722 = ~n1718 & ~n1721;
  assign n1723 = ~n1716 & n1722;
  assign n1724 = x66 & x67;
  assign n1725 = n1698 & n1724;
  assign n1726 = x67 & n1715;
  assign n1727 = ~n1725 & ~n1726;
  assign n1728 = n1723 & n1727;
  assign n1729 = n1728 ^ x68;
  assign n1730 = n1579 & n1681;
  assign n1731 = n1730 ^ n1581;
  assign n1732 = n1731 ^ n1728;
  assign n1733 = ~n1729 & n1732;
  assign n1734 = n1733 ^ x68;
  assign n1735 = n1734 ^ x69;
  assign n1736 = n1585 & n1681;
  assign n1737 = n1736 ^ n1587;
  assign n1738 = n1737 ^ n1734;
  assign n1739 = n1735 & ~n1738;
  assign n1740 = n1739 ^ x69;
  assign n1741 = n1740 ^ x70;
  assign n1742 = n1591 & n1681;
  assign n1743 = n1742 ^ n1594;
  assign n1744 = n1743 ^ n1740;
  assign n1745 = n1741 & ~n1744;
  assign n1746 = n1745 ^ x70;
  assign n1747 = n1746 ^ x71;
  assign n1748 = n1598 & n1681;
  assign n1749 = n1748 ^ n1604;
  assign n1750 = n1749 ^ n1746;
  assign n1751 = n1747 & ~n1750;
  assign n1752 = n1751 ^ x71;
  assign n1753 = n1752 ^ x72;
  assign n1754 = n1608 & n1681;
  assign n1755 = n1754 ^ n1610;
  assign n1756 = n1755 ^ n1752;
  assign n1757 = n1753 & ~n1756;
  assign n1758 = n1757 ^ x72;
  assign n1759 = n1758 ^ x73;
  assign n1760 = n1614 & n1681;
  assign n1761 = n1760 ^ n1616;
  assign n1762 = n1761 ^ n1758;
  assign n1763 = n1759 & ~n1762;
  assign n1764 = n1763 ^ x73;
  assign n1765 = n1764 ^ x74;
  assign n1766 = ~x87 & n168;
  assign n1767 = n169 & n1766;
  assign n1768 = n1620 & n1681;
  assign n1769 = n1768 ^ n1622;
  assign n1770 = n1769 ^ n1764;
  assign n1771 = n1765 & ~n1770;
  assign n1772 = n1771 ^ x74;
  assign n1773 = n1772 ^ x75;
  assign n1774 = n1626 & n1681;
  assign n1775 = n1774 ^ n1628;
  assign n1776 = n1775 ^ n1772;
  assign n1777 = n1773 & ~n1776;
  assign n1778 = n1777 ^ x75;
  assign n1779 = n1778 ^ x76;
  assign n1780 = n1632 & n1681;
  assign n1781 = n1780 ^ n1634;
  assign n1782 = n1781 ^ n1778;
  assign n1783 = n1779 & ~n1782;
  assign n1784 = n1783 ^ x76;
  assign n1785 = n1784 ^ x77;
  assign n1786 = n1638 & n1681;
  assign n1787 = n1786 ^ n1640;
  assign n1788 = n1787 ^ n1784;
  assign n1789 = n1785 & ~n1788;
  assign n1790 = n1789 ^ x77;
  assign n1791 = n1790 ^ x78;
  assign n1792 = n1644 & n1681;
  assign n1793 = n1792 ^ n1646;
  assign n1794 = n1793 ^ n1790;
  assign n1795 = n1791 & ~n1794;
  assign n1796 = n1795 ^ x78;
  assign n1797 = n1796 ^ x79;
  assign n1798 = n1650 & n1681;
  assign n1799 = n1798 ^ n1652;
  assign n1800 = n1799 ^ n1796;
  assign n1801 = n1797 & ~n1800;
  assign n1802 = n1801 ^ x79;
  assign n1803 = n1802 ^ x80;
  assign n1804 = n1656 & n1681;
  assign n1805 = n1804 ^ n1658;
  assign n1806 = n1805 ^ n1802;
  assign n1807 = n1803 & ~n1806;
  assign n1808 = n1807 ^ x80;
  assign n1809 = n1808 ^ x81;
  assign n1810 = n1662 & n1681;
  assign n1811 = n1810 ^ n1664;
  assign n1812 = n1811 ^ n1808;
  assign n1813 = n1809 & ~n1812;
  assign n1814 = n1813 ^ x81;
  assign n1815 = n1814 ^ x82;
  assign n1816 = n1668 & n1681;
  assign n1817 = n1816 ^ n1670;
  assign n1818 = n1817 ^ n1814;
  assign n1819 = n1815 & ~n1818;
  assign n1820 = n1819 ^ x82;
  assign n1821 = n1820 ^ x83;
  assign n1822 = n1673 ^ x82;
  assign n1823 = n1681 & n1822;
  assign n1824 = n1823 ^ n1545;
  assign n1825 = n1824 ^ n1820;
  assign n1826 = n1821 & n1825;
  assign n1827 = n1826 ^ x83;
  assign n1828 = n1827 ^ x84;
  assign n1829 = n1827 ^ n1683;
  assign n1830 = n1828 & n1829;
  assign n1831 = n1830 ^ x84;
  assign n1832 = n1767 & ~n1831;
  assign n1833 = n1765 & n1832;
  assign n1834 = n1833 ^ n1769;
  assign n1835 = ~x75 & ~n1834;
  assign n1836 = x65 & n1767;
  assign n1837 = ~n1681 & n1836;
  assign n1838 = ~n1831 & n1837;
  assign n1839 = n219 & n1681;
  assign n1840 = ~n1838 & ~n1839;
  assign n1841 = x43 & ~n1840;
  assign n1842 = n1681 ^ x65;
  assign n1843 = n341 & ~n1842;
  assign n1844 = x43 & n1843;
  assign n1845 = n1844 ^ n340;
  assign n1846 = n1832 & n1845;
  assign n1847 = n1846 ^ n1704;
  assign n1848 = ~n1841 & ~n1847;
  assign n1849 = n1848 ^ x44;
  assign n1850 = n1849 ^ x66;
  assign n1851 = x64 & n1832;
  assign n1852 = x42 & ~x65;
  assign n1853 = x43 & ~n1852;
  assign n1854 = n1851 & n1853;
  assign n1855 = ~x42 & x64;
  assign n1856 = ~x65 & ~n1855;
  assign n1857 = ~x43 & ~n1856;
  assign n1858 = ~n1832 & n1857;
  assign n1859 = x43 ^ x42;
  assign n1860 = ~x64 & n1859;
  assign n1861 = n1860 ^ x42;
  assign n1862 = x65 & ~n1861;
  assign n1863 = ~n1858 & ~n1862;
  assign n1864 = ~n1854 & n1863;
  assign n1865 = n1864 ^ n1849;
  assign n1866 = n1850 & n1865;
  assign n1867 = n1866 ^ x66;
  assign n1868 = n1867 ^ x67;
  assign n1869 = n1710 ^ x66;
  assign n1870 = n1832 & ~n1869;
  assign n1871 = n1870 ^ n1698;
  assign n1872 = n1871 ^ n1867;
  assign n1873 = n1868 & ~n1872;
  assign n1874 = n1873 ^ x67;
  assign n1875 = n1874 ^ x68;
  assign n1876 = ~n1712 & ~n1719;
  assign n1877 = n1876 ^ x67;
  assign n1878 = n1832 & ~n1877;
  assign n1879 = n1878 ^ n1715;
  assign n1880 = n1879 ^ n1874;
  assign n1881 = n1875 & ~n1880;
  assign n1882 = n1881 ^ x68;
  assign n1883 = n1882 ^ x69;
  assign n1884 = ~n1729 & n1832;
  assign n1885 = n1884 ^ n1731;
  assign n1886 = n1885 ^ n1882;
  assign n1887 = n1883 & ~n1886;
  assign n1888 = n1887 ^ x69;
  assign n1889 = n1888 ^ x70;
  assign n1890 = n1735 & n1832;
  assign n1891 = n1890 ^ n1737;
  assign n1892 = n1891 ^ n1888;
  assign n1893 = n1889 & ~n1892;
  assign n1894 = n1893 ^ x70;
  assign n1895 = n1894 ^ x71;
  assign n1896 = n1741 & n1832;
  assign n1897 = n1896 ^ n1743;
  assign n1898 = n1897 ^ n1894;
  assign n1899 = n1895 & ~n1898;
  assign n1900 = n1899 ^ x71;
  assign n1901 = n1900 ^ x72;
  assign n1902 = n1747 & n1832;
  assign n1903 = n1902 ^ n1749;
  assign n1904 = n1903 ^ n1900;
  assign n1905 = n1901 & ~n1904;
  assign n1906 = n1905 ^ x72;
  assign n1907 = n1906 ^ x73;
  assign n1908 = n1753 & n1832;
  assign n1909 = n1908 ^ n1755;
  assign n1910 = n1909 ^ n1906;
  assign n1911 = n1907 & ~n1910;
  assign n1912 = n1911 ^ x73;
  assign n1913 = n1912 ^ x74;
  assign n1914 = n1759 & n1832;
  assign n1915 = n1914 ^ n1761;
  assign n1916 = n1915 ^ n1912;
  assign n1917 = n1913 & ~n1916;
  assign n1918 = n1917 ^ x74;
  assign n1919 = ~n1835 & n1918;
  assign n1920 = x75 & n1834;
  assign n1921 = n1773 & n1832;
  assign n1922 = n1921 ^ n1775;
  assign n1923 = ~n1920 & ~n1922;
  assign n1924 = ~n1919 & n1923;
  assign n1925 = x76 & ~n1924;
  assign n1926 = ~n1919 & ~n1920;
  assign n1927 = n1922 & ~n1926;
  assign n1928 = ~n1925 & ~n1927;
  assign n1929 = n1928 ^ x77;
  assign n1930 = n1779 & n1832;
  assign n1931 = n1930 ^ n1781;
  assign n1932 = n1931 ^ n1928;
  assign n1933 = ~n1929 & n1932;
  assign n1934 = n1933 ^ x77;
  assign n1935 = n1934 ^ x78;
  assign n1936 = n1785 & n1832;
  assign n1937 = n1936 ^ n1787;
  assign n1938 = n1937 ^ n1934;
  assign n1939 = n1935 & ~n1938;
  assign n1940 = n1939 ^ x78;
  assign n1941 = n1940 ^ x79;
  assign n1942 = n1791 & n1832;
  assign n1943 = n1942 ^ n1793;
  assign n1944 = n1943 ^ n1940;
  assign n1945 = n1941 & ~n1944;
  assign n1946 = n1945 ^ x79;
  assign n1947 = n1946 ^ x80;
  assign n1948 = n1797 & n1832;
  assign n1949 = n1948 ^ n1799;
  assign n1950 = n1949 ^ n1946;
  assign n1951 = n1947 & ~n1950;
  assign n1952 = n1951 ^ x80;
  assign n1953 = n1952 ^ x81;
  assign n1954 = n1803 & n1832;
  assign n1955 = n1954 ^ n1805;
  assign n1956 = n1955 ^ n1952;
  assign n1957 = n1953 & ~n1956;
  assign n1958 = n1957 ^ x81;
  assign n1959 = n1958 ^ x82;
  assign n1960 = n1809 & n1832;
  assign n1961 = n1960 ^ n1811;
  assign n1962 = n1961 ^ n1958;
  assign n1963 = n1959 & ~n1962;
  assign n1964 = n1963 ^ x82;
  assign n1965 = n1964 ^ x83;
  assign n1966 = n1815 & n1832;
  assign n1967 = n1966 ^ n1817;
  assign n1968 = n1967 ^ n1964;
  assign n1969 = n1965 & ~n1968;
  assign n1970 = n1969 ^ x83;
  assign n1971 = n1970 ^ x84;
  assign n1972 = n1821 & n1832;
  assign n1973 = n1972 ^ n1824;
  assign n1974 = n1973 ^ n1970;
  assign n1975 = n1971 & n1974;
  assign n1976 = n1975 ^ x84;
  assign n1977 = ~n1684 & ~n1976;
  assign n1978 = x84 & n1827;
  assign n1979 = n1767 & ~n1978;
  assign n1980 = n1683 & ~n1979;
  assign n1981 = ~x85 & n1980;
  assign n1982 = ~n1977 & ~n1981;
  assign n1983 = ~x86 & n1766;
  assign n1984 = x42 & x65;
  assign n1985 = n1983 & n1984;
  assign n1986 = ~n1832 & n1985;
  assign n1987 = ~n1982 & n1986;
  assign n1988 = n1851 & n1852;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = ~n1982 & n1983;
  assign n1991 = n1832 ^ x65;
  assign n1992 = n1855 & ~n1991;
  assign n1993 = ~n202 & ~n1992;
  assign n1994 = n1993 ^ n1851;
  assign n1995 = n1990 & ~n1994;
  assign n1996 = n1995 ^ n1851;
  assign n1997 = n1989 & ~n1996;
  assign n1998 = n1997 ^ x43;
  assign n1999 = n1998 ^ x66;
  assign n2000 = x64 & n1990;
  assign n2001 = x41 & n1852;
  assign n2002 = n2001 ^ x42;
  assign n2003 = n2000 & n2002;
  assign n2004 = ~x41 & n1855;
  assign n2005 = ~x42 & x65;
  assign n2006 = ~n2004 & ~n2005;
  assign n2007 = ~n1990 & ~n2006;
  assign n2008 = ~x41 & x65;
  assign n2009 = n2008 ^ n2005;
  assign n2010 = x64 & n2009;
  assign n2011 = n2010 ^ n2005;
  assign n2012 = ~n2007 & ~n2011;
  assign n2013 = ~n2003 & n2012;
  assign n2014 = n2013 ^ n1998;
  assign n2015 = n1999 & n2014;
  assign n2016 = n2015 ^ x66;
  assign n2017 = n2016 ^ x67;
  assign n2018 = n1965 & n1990;
  assign n2019 = n2018 ^ n1967;
  assign n2020 = x84 & n2019;
  assign n2021 = n1941 & n1990;
  assign n2022 = n2021 ^ n1943;
  assign n2023 = x80 & n2022;
  assign n2024 = n1864 ^ x66;
  assign n2025 = n1990 & ~n2024;
  assign n2026 = n2025 ^ n1849;
  assign n2027 = n2026 ^ n2016;
  assign n2028 = n2017 & ~n2027;
  assign n2029 = n2028 ^ x67;
  assign n2030 = n2029 ^ x68;
  assign n2031 = n1868 & n1990;
  assign n2032 = n2031 ^ n1871;
  assign n2033 = n2032 ^ n2029;
  assign n2034 = n2030 & ~n2033;
  assign n2035 = n2034 ^ x68;
  assign n2036 = n2035 ^ x69;
  assign n2037 = n1875 & n1990;
  assign n2038 = n2037 ^ n1879;
  assign n2039 = n2038 ^ n2035;
  assign n2040 = n2036 & ~n2039;
  assign n2041 = n2040 ^ x69;
  assign n2042 = n2041 ^ x70;
  assign n2043 = n1883 & n1990;
  assign n2044 = n2043 ^ n1885;
  assign n2045 = n2044 ^ n2041;
  assign n2046 = n2042 & ~n2045;
  assign n2047 = n2046 ^ x70;
  assign n2048 = n2047 ^ x71;
  assign n2049 = n1889 & n1990;
  assign n2050 = n2049 ^ n1891;
  assign n2051 = n2050 ^ n2047;
  assign n2052 = n2048 & ~n2051;
  assign n2053 = n2052 ^ x71;
  assign n2054 = n2053 ^ x72;
  assign n2055 = n1895 & n1990;
  assign n2056 = n2055 ^ n1897;
  assign n2057 = n2056 ^ n2053;
  assign n2058 = n2054 & ~n2057;
  assign n2059 = n2058 ^ x72;
  assign n2060 = n2059 ^ x73;
  assign n2061 = n1901 & n1990;
  assign n2062 = n2061 ^ n1903;
  assign n2063 = n2062 ^ n2059;
  assign n2064 = n2060 & ~n2063;
  assign n2065 = n2064 ^ x73;
  assign n2066 = n2065 ^ x74;
  assign n2067 = n1907 & n1990;
  assign n2068 = n2067 ^ n1909;
  assign n2069 = n2068 ^ n2065;
  assign n2070 = n2066 & ~n2069;
  assign n2071 = n2070 ^ x74;
  assign n2072 = n2071 ^ x75;
  assign n2073 = n1913 & n1990;
  assign n2074 = n2073 ^ n1915;
  assign n2075 = n2074 ^ n2071;
  assign n2076 = n2072 & ~n2075;
  assign n2077 = n2076 ^ x75;
  assign n2078 = n2077 ^ x76;
  assign n2079 = n1918 ^ x75;
  assign n2080 = n1990 & n2079;
  assign n2081 = n2080 ^ n1834;
  assign n2082 = n2081 ^ n2077;
  assign n2083 = n2078 & ~n2082;
  assign n2084 = n2083 ^ x76;
  assign n2085 = n2084 ^ x77;
  assign n2086 = n1926 ^ x76;
  assign n2087 = n1990 & ~n2086;
  assign n2088 = n2087 ^ n1922;
  assign n2089 = n2088 ^ n2084;
  assign n2090 = n2085 & ~n2089;
  assign n2091 = n2090 ^ x77;
  assign n2092 = n2091 ^ x78;
  assign n2093 = ~n1929 & n1990;
  assign n2094 = n2093 ^ n1931;
  assign n2095 = n2094 ^ n2091;
  assign n2096 = n2092 & ~n2095;
  assign n2097 = n2096 ^ x78;
  assign n2098 = n2097 ^ x79;
  assign n2099 = n1935 & n1990;
  assign n2100 = n2099 ^ n1937;
  assign n2101 = n2100 ^ n2097;
  assign n2102 = n2098 & ~n2101;
  assign n2103 = n2102 ^ x79;
  assign n2104 = ~n2023 & ~n2103;
  assign n2105 = ~x80 & ~n2022;
  assign n2106 = n1947 & n1990;
  assign n2107 = n2106 ^ n1949;
  assign n2108 = ~x81 & ~n2107;
  assign n2109 = ~n2105 & ~n2108;
  assign n2110 = ~n2104 & n2109;
  assign n2111 = x81 & n2107;
  assign n2112 = ~n2110 & ~n2111;
  assign n2113 = n2112 ^ x82;
  assign n2114 = n1953 & n1990;
  assign n2115 = n2114 ^ n1955;
  assign n2116 = n2115 ^ n2112;
  assign n2117 = ~n2113 & n2116;
  assign n2118 = n2117 ^ x82;
  assign n2119 = n2118 ^ x83;
  assign n2120 = n1959 & n1990;
  assign n2121 = n2120 ^ n1961;
  assign n2122 = n2121 ^ n2118;
  assign n2123 = n2119 & ~n2122;
  assign n2124 = n2123 ^ x83;
  assign n2125 = ~n2020 & ~n2124;
  assign n2126 = ~x84 & ~n2019;
  assign n2127 = n1971 & n1990;
  assign n2128 = n2127 ^ n1973;
  assign n2129 = ~x85 & n2128;
  assign n2130 = ~n2126 & ~n2129;
  assign n2131 = ~n2125 & n2130;
  assign n2132 = n1980 & ~n1990;
  assign n2133 = ~n242 & ~n2132;
  assign n2134 = x86 & n2133;
  assign n2135 = n1766 & ~n2134;
  assign n2136 = x85 & ~n2128;
  assign n2137 = n2135 & ~n2136;
  assign n2138 = ~n2131 & n2137;
  assign n2139 = n1983 & ~n2133;
  assign n2140 = ~n2138 & ~n2139;
  assign n2141 = n2017 & ~n2140;
  assign n2142 = n2141 ^ n2026;
  assign n2143 = x68 & n2142;
  assign n2144 = x65 & ~n1990;
  assign n2145 = ~n2140 & n2144;
  assign n2146 = n219 & n1990;
  assign n2147 = ~n2145 & ~n2146;
  assign n2148 = x41 & ~n2147;
  assign n2149 = n1990 ^ x65;
  assign n2150 = n341 & ~n2149;
  assign n2151 = x41 & n2150;
  assign n2152 = n2151 ^ n340;
  assign n2153 = ~n2140 & n2152;
  assign n2154 = n2153 ^ n2000;
  assign n2155 = ~n2148 & ~n2154;
  assign n2156 = n2155 ^ x42;
  assign n2157 = n2156 ^ x66;
  assign n2158 = x64 & ~n2140;
  assign n2159 = x41 & ~x65;
  assign n2160 = x40 & n2159;
  assign n2161 = n2160 ^ x41;
  assign n2162 = n2158 & n2161;
  assign n2163 = ~x40 & x64;
  assign n2164 = ~x65 & ~n2163;
  assign n2165 = ~x41 & ~n2164;
  assign n2166 = n2140 & n2165;
  assign n2167 = ~x40 & x65;
  assign n2168 = x64 & n2167;
  assign n2169 = ~x41 & n202;
  assign n2170 = ~n2168 & ~n2169;
  assign n2171 = ~n2166 & n2170;
  assign n2172 = ~n2162 & n2171;
  assign n2173 = n2172 ^ n2156;
  assign n2174 = n2157 & n2173;
  assign n2175 = n2174 ^ x66;
  assign n2176 = n2175 ^ x67;
  assign n2177 = n2013 ^ x66;
  assign n2178 = ~n2140 & ~n2177;
  assign n2179 = n2178 ^ n1998;
  assign n2180 = n2179 ^ n2175;
  assign n2181 = n2176 & ~n2180;
  assign n2182 = n2181 ^ x67;
  assign n2183 = ~n2143 & ~n2182;
  assign n2184 = ~x68 & ~n2142;
  assign n2185 = n2030 & ~n2140;
  assign n2186 = n2185 ^ n2032;
  assign n2187 = ~x69 & ~n2186;
  assign n2188 = ~n2184 & ~n2187;
  assign n2189 = ~n2183 & n2188;
  assign n2190 = x69 & n2186;
  assign n2191 = ~n2189 & ~n2190;
  assign n2192 = n2191 ^ x70;
  assign n2193 = n2036 & ~n2140;
  assign n2194 = n2193 ^ n2038;
  assign n2195 = n2194 ^ n2191;
  assign n2196 = ~n2192 & n2195;
  assign n2197 = n2196 ^ x70;
  assign n2198 = n2197 ^ x71;
  assign n2199 = n2042 & ~n2140;
  assign n2200 = n2199 ^ n2044;
  assign n2201 = n2200 ^ n2197;
  assign n2202 = n2198 & ~n2201;
  assign n2203 = n2202 ^ x71;
  assign n2204 = n2203 ^ x72;
  assign n2205 = n2048 & ~n2140;
  assign n2206 = n2205 ^ n2050;
  assign n2207 = n2206 ^ n2203;
  assign n2208 = n2204 & ~n2207;
  assign n2209 = n2208 ^ x72;
  assign n2210 = n2209 ^ x73;
  assign n2211 = n2054 & ~n2140;
  assign n2212 = n2211 ^ n2056;
  assign n2213 = n2212 ^ n2209;
  assign n2214 = n2210 & ~n2213;
  assign n2215 = n2214 ^ x73;
  assign n2216 = n2215 ^ x74;
  assign n2217 = n2060 & ~n2140;
  assign n2218 = n2217 ^ n2062;
  assign n2219 = n2218 ^ n2215;
  assign n2220 = n2216 & ~n2219;
  assign n2221 = n2220 ^ x74;
  assign n2222 = n2221 ^ x75;
  assign n2223 = n2066 & ~n2140;
  assign n2224 = n2223 ^ n2068;
  assign n2225 = n2224 ^ n2221;
  assign n2226 = n2222 & ~n2225;
  assign n2227 = n2226 ^ x75;
  assign n2228 = n2227 ^ x76;
  assign n2229 = n2072 & ~n2140;
  assign n2230 = n2229 ^ n2074;
  assign n2231 = n2230 ^ n2227;
  assign n2232 = n2228 & ~n2231;
  assign n2233 = n2232 ^ x76;
  assign n2234 = n2233 ^ x77;
  assign n2235 = n2078 & ~n2140;
  assign n2236 = n2235 ^ n2081;
  assign n2237 = n2236 ^ n2233;
  assign n2238 = n2234 & ~n2237;
  assign n2239 = n2238 ^ x77;
  assign n2240 = n2239 ^ x78;
  assign n2241 = n2085 & ~n2140;
  assign n2242 = n2241 ^ n2088;
  assign n2243 = n2242 ^ n2239;
  assign n2244 = n2240 & ~n2243;
  assign n2245 = n2244 ^ x78;
  assign n2246 = n2245 ^ x79;
  assign n2247 = n2092 & ~n2140;
  assign n2248 = n2247 ^ n2094;
  assign n2249 = n2248 ^ n2245;
  assign n2250 = n2246 & ~n2249;
  assign n2251 = n2250 ^ x79;
  assign n2252 = n2251 ^ x80;
  assign n2253 = n2098 & ~n2140;
  assign n2254 = n2253 ^ n2100;
  assign n2255 = n2254 ^ n2251;
  assign n2256 = n2252 & ~n2255;
  assign n2257 = n2256 ^ x80;
  assign n2258 = n2257 ^ x81;
  assign n2259 = n2103 ^ x80;
  assign n2260 = ~n2140 & n2259;
  assign n2261 = n2260 ^ n2022;
  assign n2262 = n2261 ^ n2257;
  assign n2263 = n2258 & ~n2262;
  assign n2264 = n2263 ^ x81;
  assign n2265 = n2264 ^ x82;
  assign n2266 = ~n2104 & ~n2105;
  assign n2267 = n2266 ^ x81;
  assign n2268 = ~n2140 & n2267;
  assign n2269 = n2268 ^ n2107;
  assign n2270 = n2269 ^ n2264;
  assign n2271 = n2265 & ~n2270;
  assign n2272 = n2271 ^ x82;
  assign n2273 = n2272 ^ x83;
  assign n2274 = ~n2113 & ~n2140;
  assign n2275 = n2274 ^ n2115;
  assign n2276 = n2275 ^ n2272;
  assign n2277 = n2273 & ~n2276;
  assign n2278 = n2277 ^ x83;
  assign n2279 = n2278 ^ x84;
  assign n2280 = n2119 & ~n2140;
  assign n2281 = n2280 ^ n2121;
  assign n2282 = n2281 ^ n2278;
  assign n2283 = n2279 & ~n2282;
  assign n2284 = n2283 ^ x84;
  assign n2285 = n2284 ^ x85;
  assign n2286 = n2124 ^ x84;
  assign n2287 = ~n2140 & n2286;
  assign n2288 = n2287 ^ n2019;
  assign n2289 = n2288 ^ n2284;
  assign n2290 = n2285 & ~n2289;
  assign n2291 = n2290 ^ x85;
  assign n2292 = n2291 ^ x86;
  assign n2293 = ~n2125 & ~n2126;
  assign n2294 = n2293 ^ x85;
  assign n2295 = ~n2140 & n2294;
  assign n2296 = n2295 ^ n2128;
  assign n2297 = n2296 ^ n2291;
  assign n2298 = n2292 & n2297;
  assign n2299 = n2298 ^ x86;
  assign n2300 = n2299 ^ x87;
  assign n2301 = ~n242 & ~n2140;
  assign n2302 = ~n2133 & ~n2301;
  assign n2303 = n2302 ^ n2299;
  assign n2304 = n2300 & n2303;
  assign n2305 = n2304 ^ x87;
  assign n2306 = n168 & ~n2305;
  assign n2307 = n2292 & n2306;
  assign n2308 = n2307 ^ n2296;
  assign n2309 = x87 & ~n2308;
  assign n2310 = n2204 & n2306;
  assign n2311 = n2310 ^ n2206;
  assign n2312 = x73 & n2311;
  assign n2313 = x65 & n168;
  assign n2314 = n2140 & n2313;
  assign n2315 = ~n2305 & n2314;
  assign n2316 = n219 & ~n2140;
  assign n2317 = ~n2315 & ~n2316;
  assign n2318 = x40 & ~n2317;
  assign n2319 = n2140 ^ x65;
  assign n2320 = n341 & n2319;
  assign n2321 = x40 & n2320;
  assign n2322 = n2321 ^ n340;
  assign n2323 = n2306 & n2322;
  assign n2324 = n2323 ^ n2158;
  assign n2325 = ~n2318 & ~n2324;
  assign n2326 = n2325 ^ x41;
  assign n2327 = n2326 ^ x66;
  assign n2328 = x64 & n2306;
  assign n2329 = x39 & ~x65;
  assign n2330 = x40 & ~n2329;
  assign n2331 = n2328 & n2330;
  assign n2332 = ~x39 & n2163;
  assign n2333 = ~n2167 & ~n2332;
  assign n2334 = ~n2306 & ~n2333;
  assign n2335 = ~x39 & x65;
  assign n2336 = n2335 ^ n2167;
  assign n2337 = x64 & n2336;
  assign n2338 = n2337 ^ n2167;
  assign n2339 = ~n2334 & ~n2338;
  assign n2340 = ~n2331 & n2339;
  assign n2341 = n2340 ^ n2326;
  assign n2342 = n2327 & n2341;
  assign n2343 = n2342 ^ x66;
  assign n2344 = n2343 ^ x67;
  assign n2345 = n2172 ^ x66;
  assign n2346 = n2306 & ~n2345;
  assign n2347 = n2346 ^ n2156;
  assign n2348 = n2347 ^ n2343;
  assign n2349 = n2344 & ~n2348;
  assign n2350 = n2349 ^ x67;
  assign n2351 = n2350 ^ x68;
  assign n2352 = n2176 & n2306;
  assign n2353 = n2352 ^ n2179;
  assign n2354 = n2353 ^ n2350;
  assign n2355 = n2351 & ~n2354;
  assign n2356 = n2355 ^ x68;
  assign n2357 = n2356 ^ x69;
  assign n2358 = n2182 ^ x68;
  assign n2359 = n2306 & n2358;
  assign n2360 = n2359 ^ n2142;
  assign n2361 = n2360 ^ n2356;
  assign n2362 = n2357 & ~n2361;
  assign n2363 = n2362 ^ x69;
  assign n2364 = n2363 ^ x70;
  assign n2366 = ~n2183 & ~n2184;
  assign n2365 = n2186 ^ x69;
  assign n2367 = n2366 ^ n2365;
  assign n2368 = n2367 ^ n2186;
  assign n2369 = n2306 & n2368;
  assign n2370 = n2369 ^ n2186;
  assign n2371 = n2370 ^ n2363;
  assign n2372 = n2364 & ~n2371;
  assign n2373 = n2372 ^ x70;
  assign n2374 = n2373 ^ x71;
  assign n2375 = ~n2192 & n2306;
  assign n2376 = n2375 ^ n2194;
  assign n2377 = n2376 ^ n2373;
  assign n2378 = n2374 & ~n2377;
  assign n2379 = n2378 ^ x71;
  assign n2380 = n2379 ^ x72;
  assign n2381 = n2198 & n2306;
  assign n2382 = n2381 ^ n2200;
  assign n2383 = n2382 ^ n2379;
  assign n2384 = n2380 & ~n2383;
  assign n2385 = n2384 ^ x72;
  assign n2386 = ~n2312 & ~n2385;
  assign n2387 = ~x73 & ~n2311;
  assign n2388 = n2210 & n2306;
  assign n2389 = n2388 ^ n2212;
  assign n2390 = ~x74 & ~n2389;
  assign n2391 = ~n2387 & ~n2390;
  assign n2392 = ~n2386 & n2391;
  assign n2393 = x74 & n2389;
  assign n2394 = ~n2392 & ~n2393;
  assign n2395 = n2394 ^ x75;
  assign n2396 = n2216 & n2306;
  assign n2397 = n2396 ^ n2218;
  assign n2398 = n2397 ^ n2394;
  assign n2399 = ~n2395 & n2398;
  assign n2400 = n2399 ^ x75;
  assign n2401 = n2400 ^ x76;
  assign n2402 = n2222 & n2306;
  assign n2403 = n2402 ^ n2224;
  assign n2404 = n2403 ^ n2400;
  assign n2405 = n2401 & ~n2404;
  assign n2406 = n2405 ^ x76;
  assign n2407 = n2406 ^ x77;
  assign n2408 = n2228 & n2306;
  assign n2409 = n2408 ^ n2230;
  assign n2410 = n2409 ^ n2406;
  assign n2411 = n2407 & ~n2410;
  assign n2412 = n2411 ^ x77;
  assign n2413 = n2412 ^ x78;
  assign n2414 = n2234 & n2306;
  assign n2415 = n2414 ^ n2236;
  assign n2416 = n2415 ^ n2412;
  assign n2417 = n2413 & ~n2416;
  assign n2418 = n2417 ^ x78;
  assign n2419 = n2418 ^ x79;
  assign n2420 = n2240 & n2306;
  assign n2421 = n2420 ^ n2242;
  assign n2422 = n2421 ^ n2418;
  assign n2423 = n2419 & ~n2422;
  assign n2424 = n2423 ^ x79;
  assign n2425 = n2424 ^ x80;
  assign n2426 = n2246 & n2306;
  assign n2427 = n2426 ^ n2248;
  assign n2428 = n2427 ^ n2424;
  assign n2429 = n2425 & ~n2428;
  assign n2430 = n2429 ^ x80;
  assign n2431 = n2430 ^ x81;
  assign n2432 = n2252 & n2306;
  assign n2433 = n2432 ^ n2254;
  assign n2434 = n2433 ^ n2430;
  assign n2435 = n2431 & ~n2434;
  assign n2436 = n2435 ^ x81;
  assign n2437 = n2436 ^ x82;
  assign n2438 = n2258 & n2306;
  assign n2439 = n2438 ^ n2261;
  assign n2440 = n2439 ^ n2436;
  assign n2441 = n2437 & ~n2440;
  assign n2442 = n2441 ^ x82;
  assign n2443 = n2442 ^ x83;
  assign n2444 = n2265 & n2306;
  assign n2445 = n2444 ^ n2269;
  assign n2446 = n2445 ^ n2442;
  assign n2447 = n2443 & ~n2446;
  assign n2448 = n2447 ^ x83;
  assign n2449 = n2448 ^ x84;
  assign n2450 = n2273 & n2306;
  assign n2451 = n2450 ^ n2275;
  assign n2452 = n2451 ^ n2448;
  assign n2453 = n2449 & ~n2452;
  assign n2454 = n2453 ^ x84;
  assign n2455 = n2454 ^ x85;
  assign n2456 = n2279 & n2306;
  assign n2457 = n2456 ^ n2281;
  assign n2458 = n2457 ^ n2454;
  assign n2459 = n2455 & ~n2458;
  assign n2460 = n2459 ^ x85;
  assign n2461 = n2460 ^ x86;
  assign n2462 = n2285 & n2306;
  assign n2463 = n2462 ^ n2288;
  assign n2464 = n2463 ^ n2460;
  assign n2465 = n2461 & ~n2464;
  assign n2466 = n2465 ^ x86;
  assign n2467 = ~n2309 & ~n2466;
  assign n2468 = ~x87 & n2308;
  assign n2469 = n168 & ~n2299;
  assign n2470 = ~n1766 & n2302;
  assign n2471 = ~n2469 & n2470;
  assign n2472 = ~x88 & n2471;
  assign n2473 = ~n2468 & ~n2472;
  assign n2474 = ~n2467 & n2473;
  assign n2475 = x88 & ~n2302;
  assign n2476 = n167 & ~n2475;
  assign n2477 = ~n2474 & n2476;
  assign n2478 = x65 & ~n2306;
  assign n2479 = n2477 & n2478;
  assign n2480 = ~x65 & n2306;
  assign n2481 = x64 & n2480;
  assign n2482 = ~n2479 & ~n2481;
  assign n2483 = x39 & ~n2482;
  assign n2484 = n2306 ^ x65;
  assign n2485 = n341 & ~n2484;
  assign n2486 = x39 & n2485;
  assign n2487 = n2486 ^ n340;
  assign n2488 = n2477 & n2487;
  assign n2489 = n2488 ^ n2328;
  assign n2490 = ~n2483 & ~n2489;
  assign n2491 = n2490 ^ x40;
  assign n2492 = n2491 ^ x66;
  assign n2493 = ~x38 & ~n2477;
  assign n2494 = ~x38 & x65;
  assign n2495 = ~n2493 & ~n2494;
  assign n2496 = x64 & ~n2329;
  assign n2497 = ~n2495 & n2496;
  assign n2498 = x64 & n2477;
  assign n2499 = x38 & n2329;
  assign n2500 = n2499 ^ x39;
  assign n2501 = n2500 ^ n2335;
  assign n2502 = n2498 & n2501;
  assign n2503 = n2502 ^ n2335;
  assign n2504 = ~n2497 & ~n2503;
  assign n2505 = n2504 ^ n2491;
  assign n2506 = n2492 & n2505;
  assign n2507 = n2506 ^ x66;
  assign n2508 = n2507 ^ x67;
  assign n2509 = n2340 ^ x66;
  assign n2510 = n2477 & ~n2509;
  assign n2511 = n2510 ^ n2326;
  assign n2512 = n2511 ^ n2507;
  assign n2513 = n2508 & ~n2512;
  assign n2514 = n2513 ^ x67;
  assign n2515 = n2514 ^ x68;
  assign n2516 = n2344 & n2477;
  assign n2517 = n2516 ^ n2347;
  assign n2518 = n2517 ^ n2514;
  assign n2519 = n2515 & ~n2518;
  assign n2520 = n2519 ^ x68;
  assign n2521 = n2520 ^ x69;
  assign n2522 = n2351 & n2477;
  assign n2523 = n2522 ^ n2353;
  assign n2524 = n2523 ^ n2520;
  assign n2525 = n2521 & ~n2524;
  assign n2526 = n2525 ^ x69;
  assign n2527 = n2526 ^ x70;
  assign n2528 = n2461 & n2477;
  assign n2529 = n2528 ^ n2463;
  assign n2530 = x87 & n2529;
  assign n2531 = n2360 ^ x69;
  assign n2532 = n2531 ^ n2356;
  assign n2533 = n2532 ^ n2360;
  assign n2534 = n2477 & n2533;
  assign n2535 = n2534 ^ n2360;
  assign n2536 = n2535 ^ n2526;
  assign n2537 = n2527 & ~n2536;
  assign n2538 = n2537 ^ x70;
  assign n2539 = n2538 ^ x71;
  assign n2540 = n2364 & n2477;
  assign n2541 = n2540 ^ n2370;
  assign n2542 = n2541 ^ n2538;
  assign n2543 = n2539 & ~n2542;
  assign n2544 = n2543 ^ x71;
  assign n2545 = n2544 ^ x72;
  assign n2546 = n2374 & n2477;
  assign n2547 = n2546 ^ n2376;
  assign n2548 = n2547 ^ n2544;
  assign n2549 = n2545 & ~n2548;
  assign n2550 = n2549 ^ x72;
  assign n2551 = n2550 ^ x73;
  assign n2552 = n2380 & n2477;
  assign n2553 = n2552 ^ n2382;
  assign n2554 = n2553 ^ n2550;
  assign n2555 = n2551 & ~n2554;
  assign n2556 = n2555 ^ x73;
  assign n2557 = n2556 ^ x74;
  assign n2558 = n2385 ^ x73;
  assign n2559 = n2477 & n2558;
  assign n2560 = n2559 ^ n2311;
  assign n2561 = n2560 ^ n2556;
  assign n2562 = n2557 & ~n2561;
  assign n2563 = n2562 ^ x74;
  assign n2564 = n2563 ^ x75;
  assign n2565 = ~n2386 & ~n2387;
  assign n2566 = n2565 ^ x74;
  assign n2567 = n2477 & n2566;
  assign n2568 = n2567 ^ n2389;
  assign n2569 = n2568 ^ n2563;
  assign n2570 = n2564 & ~n2569;
  assign n2571 = n2570 ^ x75;
  assign n2572 = n2571 ^ x76;
  assign n2573 = ~n2395 & n2477;
  assign n2574 = n2573 ^ n2397;
  assign n2575 = n2574 ^ n2571;
  assign n2576 = n2572 & ~n2575;
  assign n2577 = n2576 ^ x76;
  assign n2578 = n2577 ^ x77;
  assign n2579 = n2401 & n2477;
  assign n2580 = n2579 ^ n2403;
  assign n2581 = n2580 ^ n2577;
  assign n2582 = n2578 & ~n2581;
  assign n2583 = n2582 ^ x77;
  assign n2584 = n2583 ^ x78;
  assign n2585 = n2407 & n2477;
  assign n2586 = n2585 ^ n2409;
  assign n2587 = n2586 ^ n2583;
  assign n2588 = n2584 & ~n2587;
  assign n2589 = n2588 ^ x78;
  assign n2590 = n2589 ^ x79;
  assign n2591 = n2413 & n2477;
  assign n2592 = n2591 ^ n2415;
  assign n2593 = n2592 ^ n2589;
  assign n2594 = n2590 & ~n2593;
  assign n2595 = n2594 ^ x79;
  assign n2596 = n2595 ^ x80;
  assign n2597 = n2419 & n2477;
  assign n2598 = n2597 ^ n2421;
  assign n2599 = n2598 ^ n2595;
  assign n2600 = n2596 & ~n2599;
  assign n2601 = n2600 ^ x80;
  assign n2602 = n2601 ^ x81;
  assign n2603 = n2425 & n2477;
  assign n2604 = n2603 ^ n2427;
  assign n2605 = n2604 ^ n2601;
  assign n2606 = n2602 & ~n2605;
  assign n2607 = n2606 ^ x81;
  assign n2608 = n2607 ^ x82;
  assign n2609 = n2431 & n2477;
  assign n2610 = n2609 ^ n2433;
  assign n2611 = n2610 ^ n2607;
  assign n2612 = n2608 & ~n2611;
  assign n2613 = n2612 ^ x82;
  assign n2614 = n2613 ^ x83;
  assign n2615 = n2437 & n2477;
  assign n2616 = n2615 ^ n2439;
  assign n2617 = n2616 ^ n2613;
  assign n2618 = n2614 & ~n2617;
  assign n2619 = n2618 ^ x83;
  assign n2620 = n2619 ^ x84;
  assign n2621 = n2443 & n2477;
  assign n2622 = n2621 ^ n2445;
  assign n2623 = n2622 ^ n2619;
  assign n2624 = n2620 & ~n2623;
  assign n2625 = n2624 ^ x84;
  assign n2626 = n2625 ^ x85;
  assign n2627 = n2449 & n2477;
  assign n2628 = n2627 ^ n2451;
  assign n2629 = n2628 ^ n2625;
  assign n2630 = n2626 & ~n2629;
  assign n2631 = n2630 ^ x85;
  assign n2632 = n2631 ^ x86;
  assign n2633 = n2455 & n2477;
  assign n2634 = n2633 ^ n2457;
  assign n2635 = n2634 ^ n2631;
  assign n2636 = n2632 & ~n2635;
  assign n2637 = n2636 ^ x86;
  assign n2638 = ~n2530 & ~n2637;
  assign n2639 = ~x87 & ~n2529;
  assign n2640 = n2466 ^ x87;
  assign n2641 = n2477 & n2640;
  assign n2642 = n2641 ^ n2308;
  assign n2643 = ~n2639 & ~n2642;
  assign n2644 = ~n2638 & n2643;
  assign n2645 = ~x88 & ~n2644;
  assign n2646 = ~n2638 & ~n2639;
  assign n2647 = n2642 & ~n2646;
  assign n2648 = ~n2645 & ~n2647;
  assign n2649 = n2648 ^ x89;
  assign n2650 = n2471 & ~n2477;
  assign n2651 = ~n242 & ~n2650;
  assign n2652 = n2651 ^ n2648;
  assign n2653 = n2649 & ~n2652;
  assign n2654 = n2653 ^ x89;
  assign n2655 = n166 & ~n2654;
  assign n2656 = n2527 & n2655;
  assign n2657 = n2656 ^ n2535;
  assign n2658 = ~x71 & ~n2657;
  assign n2659 = n2539 & n2655;
  assign n2660 = n2659 ^ n2541;
  assign n2661 = ~x72 & ~n2660;
  assign n2662 = ~n2658 & ~n2661;
  assign n2663 = x65 & n2655;
  assign n2664 = ~n2498 & ~n2663;
  assign n2665 = x65 & n2477;
  assign n2666 = x38 & ~n2665;
  assign n2667 = ~n2664 & n2666;
  assign n2668 = n2477 ^ x65;
  assign n2669 = n341 & ~n2668;
  assign n2670 = x38 & n2669;
  assign n2671 = n2670 ^ n340;
  assign n2672 = n2655 & n2671;
  assign n2673 = n2672 ^ n2498;
  assign n2674 = ~n2667 & ~n2673;
  assign n2675 = n2674 ^ x39;
  assign n2676 = n2675 ^ x66;
  assign n2677 = ~x38 & ~n2655;
  assign n2678 = ~x65 & ~n2677;
  assign n2679 = ~x37 & x64;
  assign n2680 = ~n2678 & n2679;
  assign n2681 = x64 & n2655;
  assign n2682 = x38 & ~x65;
  assign n2683 = x37 & n2682;
  assign n2684 = n2683 ^ x38;
  assign n2685 = n2684 ^ n2494;
  assign n2686 = n2681 & n2685;
  assign n2687 = n2686 ^ n2494;
  assign n2688 = ~n2680 & ~n2687;
  assign n2689 = n2688 ^ n2675;
  assign n2690 = n2676 & n2689;
  assign n2691 = n2690 ^ x66;
  assign n2692 = n2691 ^ x67;
  assign n2693 = n2504 ^ x66;
  assign n2694 = n2655 & ~n2693;
  assign n2695 = n2694 ^ n2491;
  assign n2696 = n2695 ^ n2691;
  assign n2697 = n2692 & ~n2696;
  assign n2698 = n2697 ^ x67;
  assign n2699 = n2698 ^ x68;
  assign n2700 = n2508 & n2655;
  assign n2701 = n2700 ^ n2511;
  assign n2702 = n2701 ^ n2698;
  assign n2703 = n2699 & ~n2702;
  assign n2704 = n2703 ^ x68;
  assign n2705 = n2704 ^ x69;
  assign n2706 = n2515 & n2655;
  assign n2707 = n2706 ^ n2517;
  assign n2708 = n2707 ^ n2704;
  assign n2709 = n2705 & ~n2708;
  assign n2710 = n2709 ^ x69;
  assign n2711 = n2710 ^ x70;
  assign n2712 = n2521 & n2655;
  assign n2713 = n2712 ^ n2523;
  assign n2714 = n2713 ^ n2710;
  assign n2715 = n2711 & ~n2714;
  assign n2716 = n2715 ^ x70;
  assign n2717 = n2662 & n2716;
  assign n2718 = n2660 ^ x72;
  assign n2719 = x71 & n2657;
  assign n2720 = n2719 ^ n2660;
  assign n2721 = n2718 & ~n2720;
  assign n2722 = n2721 ^ x72;
  assign n2723 = ~n2717 & ~n2722;
  assign n2724 = n2723 ^ x73;
  assign n2725 = n2545 & n2655;
  assign n2726 = n2725 ^ n2547;
  assign n2727 = n2726 ^ n2723;
  assign n2728 = ~n2724 & n2727;
  assign n2729 = n2728 ^ x73;
  assign n2730 = n2729 ^ x74;
  assign n2731 = n2551 & n2655;
  assign n2732 = n2731 ^ n2553;
  assign n2733 = n2732 ^ n2729;
  assign n2734 = n2730 & ~n2733;
  assign n2735 = n2734 ^ x74;
  assign n2736 = n2735 ^ x75;
  assign n2737 = n2557 & n2655;
  assign n2738 = n2737 ^ n2560;
  assign n2739 = n2738 ^ n2735;
  assign n2740 = n2736 & ~n2739;
  assign n2741 = n2740 ^ x75;
  assign n2742 = n2741 ^ x76;
  assign n2743 = n2564 & n2655;
  assign n2744 = n2743 ^ n2568;
  assign n2745 = n2744 ^ n2741;
  assign n2746 = n2742 & ~n2745;
  assign n2747 = n2746 ^ x76;
  assign n2748 = n2747 ^ x77;
  assign n2749 = n2572 & n2655;
  assign n2750 = n2749 ^ n2574;
  assign n2751 = n2750 ^ n2747;
  assign n2752 = n2748 & ~n2751;
  assign n2753 = n2752 ^ x77;
  assign n2754 = n2753 ^ x78;
  assign n2755 = n2578 & n2655;
  assign n2756 = n2755 ^ n2580;
  assign n2757 = n2756 ^ n2753;
  assign n2758 = n2754 & ~n2757;
  assign n2759 = n2758 ^ x78;
  assign n2760 = n2759 ^ x79;
  assign n2761 = n2584 & n2655;
  assign n2762 = n2761 ^ n2586;
  assign n2763 = n2762 ^ n2759;
  assign n2764 = n2760 & ~n2763;
  assign n2765 = n2764 ^ x79;
  assign n2766 = n2765 ^ x80;
  assign n2767 = n2590 & n2655;
  assign n2768 = n2767 ^ n2592;
  assign n2769 = n2768 ^ n2765;
  assign n2770 = n2766 & ~n2769;
  assign n2771 = n2770 ^ x80;
  assign n2772 = n2771 ^ x81;
  assign n2773 = n2596 & n2655;
  assign n2774 = n2773 ^ n2598;
  assign n2775 = n2774 ^ n2771;
  assign n2776 = n2772 & ~n2775;
  assign n2777 = n2776 ^ x81;
  assign n2778 = n2777 ^ x82;
  assign n2779 = n2602 & n2655;
  assign n2780 = n2779 ^ n2604;
  assign n2781 = n2780 ^ n2777;
  assign n2782 = n2778 & ~n2781;
  assign n2783 = n2782 ^ x82;
  assign n2784 = n2783 ^ x83;
  assign n2785 = n2608 & n2655;
  assign n2786 = n2785 ^ n2610;
  assign n2787 = n2786 ^ n2783;
  assign n2788 = n2784 & ~n2787;
  assign n2789 = n2788 ^ x83;
  assign n2790 = n2789 ^ x84;
  assign n2791 = n2614 & n2655;
  assign n2792 = n2791 ^ n2616;
  assign n2793 = n2792 ^ n2789;
  assign n2794 = n2790 & ~n2793;
  assign n2795 = n2794 ^ x84;
  assign n2796 = n2795 ^ x85;
  assign n2797 = n2620 & n2655;
  assign n2798 = n2797 ^ n2622;
  assign n2799 = n2798 ^ n2795;
  assign n2800 = n2796 & ~n2799;
  assign n2801 = n2800 ^ x85;
  assign n2802 = n2801 ^ x86;
  assign n2803 = n2626 & n2655;
  assign n2804 = n2803 ^ n2628;
  assign n2805 = n2804 ^ n2801;
  assign n2806 = n2802 & ~n2805;
  assign n2807 = n2806 ^ x86;
  assign n2808 = n2807 ^ x87;
  assign n2809 = n2632 & n2655;
  assign n2810 = n2809 ^ n2634;
  assign n2811 = n2810 ^ n2807;
  assign n2812 = n2808 & ~n2811;
  assign n2813 = n2812 ^ x87;
  assign n2814 = n2813 ^ x88;
  assign n2815 = n2637 ^ x87;
  assign n2816 = n2655 & n2815;
  assign n2817 = n2816 ^ n2529;
  assign n2818 = n2817 ^ n2813;
  assign n2819 = n2814 & ~n2818;
  assign n2820 = n2819 ^ x88;
  assign n2821 = n2820 ^ x89;
  assign n2822 = n2646 ^ x88;
  assign n2823 = n2655 & n2822;
  assign n2824 = n2823 ^ n2642;
  assign n2825 = n2824 ^ n2820;
  assign n2826 = n2821 & n2825;
  assign n2827 = n2826 ^ x89;
  assign n2828 = n2827 ^ x90;
  assign n2829 = ~x90 & ~n2654;
  assign n2830 = ~n2651 & ~n2829;
  assign n2831 = ~n242 & ~n2830;
  assign n2832 = n2831 ^ n2827;
  assign n2833 = n2828 & ~n2832;
  assign n2834 = n2833 ^ x90;
  assign n2835 = n165 & ~n2834;
  assign n2836 = n2760 & n2835;
  assign n2837 = n2836 ^ n2762;
  assign n2838 = x80 & n2837;
  assign n2839 = x37 & ~n2663;
  assign n2840 = n2835 & ~n2839;
  assign n2841 = n2681 & ~n2840;
  assign n2842 = n2655 ^ x65;
  assign n2843 = n2679 & ~n2842;
  assign n2844 = ~n202 & ~n2843;
  assign n2845 = x65 & n2839;
  assign n2846 = n2844 & ~n2845;
  assign n2847 = n2835 & ~n2846;
  assign n2848 = ~n2841 & ~n2847;
  assign n2849 = n2848 ^ x38;
  assign n2850 = n2849 ^ x66;
  assign n2851 = x64 & n2835;
  assign n2852 = x37 & ~x65;
  assign n2853 = x36 & n2852;
  assign n2854 = n2853 ^ x37;
  assign n2855 = n2851 & n2854;
  assign n2856 = ~x36 & x64;
  assign n2857 = ~x65 & ~n2856;
  assign n2858 = ~x37 & ~n2857;
  assign n2859 = ~n2835 & n2858;
  assign n2860 = x37 ^ x36;
  assign n2861 = ~x64 & n2860;
  assign n2862 = n2861 ^ x36;
  assign n2863 = x65 & ~n2862;
  assign n2864 = ~n2859 & ~n2863;
  assign n2865 = ~n2855 & n2864;
  assign n2866 = n2865 ^ n2849;
  assign n2867 = n2850 & n2866;
  assign n2868 = n2867 ^ x66;
  assign n2869 = n2868 ^ x67;
  assign n2870 = n2688 ^ x66;
  assign n2871 = n2835 & ~n2870;
  assign n2872 = n2871 ^ n2675;
  assign n2873 = n2872 ^ n2868;
  assign n2874 = n2869 & ~n2873;
  assign n2875 = n2874 ^ x67;
  assign n2876 = n2875 ^ x68;
  assign n2877 = n2692 & n2835;
  assign n2878 = n2877 ^ n2695;
  assign n2879 = n2878 ^ n2875;
  assign n2880 = n2876 & ~n2879;
  assign n2881 = n2880 ^ x68;
  assign n2882 = n2881 ^ x69;
  assign n2883 = n2699 & n2835;
  assign n2884 = n2883 ^ n2701;
  assign n2885 = n2884 ^ n2881;
  assign n2886 = n2882 & ~n2885;
  assign n2887 = n2886 ^ x69;
  assign n2888 = n2887 ^ x70;
  assign n2889 = n2705 & n2835;
  assign n2890 = n2889 ^ n2707;
  assign n2891 = n2890 ^ n2887;
  assign n2892 = n2888 & ~n2891;
  assign n2893 = n2892 ^ x70;
  assign n2894 = n2893 ^ x71;
  assign n2895 = n2711 & n2835;
  assign n2896 = n2895 ^ n2713;
  assign n2897 = n2896 ^ n2893;
  assign n2898 = n2894 & ~n2897;
  assign n2899 = n2898 ^ x71;
  assign n2900 = n2899 ^ x72;
  assign n2901 = n2716 ^ x71;
  assign n2902 = n2835 & n2901;
  assign n2903 = n2902 ^ n2657;
  assign n2904 = n2903 ^ n2899;
  assign n2905 = n2900 & ~n2904;
  assign n2906 = n2905 ^ x72;
  assign n2907 = n2906 ^ x73;
  assign n2908 = n2716 ^ n2657;
  assign n2909 = n2901 & ~n2908;
  assign n2910 = n2909 ^ x71;
  assign n2911 = n2910 ^ x72;
  assign n2912 = n2835 & n2911;
  assign n2913 = n2912 ^ n2660;
  assign n2914 = n2913 ^ n2906;
  assign n2915 = n2907 & ~n2914;
  assign n2916 = n2915 ^ x73;
  assign n2917 = n2916 ^ x74;
  assign n2918 = ~n2724 & n2835;
  assign n2919 = n2918 ^ n2726;
  assign n2920 = n2919 ^ n2916;
  assign n2921 = n2917 & ~n2920;
  assign n2922 = n2921 ^ x74;
  assign n2923 = n2922 ^ x75;
  assign n2924 = n2730 & n2835;
  assign n2925 = n2924 ^ n2732;
  assign n2926 = n2925 ^ n2922;
  assign n2927 = n2923 & ~n2926;
  assign n2928 = n2927 ^ x75;
  assign n2929 = n2928 ^ x76;
  assign n2930 = n2736 & n2835;
  assign n2931 = n2930 ^ n2738;
  assign n2932 = n2931 ^ n2928;
  assign n2933 = n2929 & ~n2932;
  assign n2934 = n2933 ^ x76;
  assign n2935 = n2934 ^ x77;
  assign n2936 = n2742 & n2835;
  assign n2937 = n2936 ^ n2744;
  assign n2938 = n2937 ^ n2934;
  assign n2939 = n2935 & ~n2938;
  assign n2940 = n2939 ^ x77;
  assign n2941 = n2940 ^ x78;
  assign n2942 = n2748 & n2835;
  assign n2943 = n2942 ^ n2750;
  assign n2944 = n2943 ^ n2940;
  assign n2945 = n2941 & ~n2944;
  assign n2946 = n2945 ^ x78;
  assign n2947 = n2946 ^ x79;
  assign n2948 = n2754 & n2835;
  assign n2949 = n2948 ^ n2756;
  assign n2950 = n2949 ^ n2946;
  assign n2951 = n2947 & ~n2950;
  assign n2952 = n2951 ^ x79;
  assign n2953 = ~n2838 & ~n2952;
  assign n2954 = ~x80 & ~n2837;
  assign n2955 = n2766 & n2835;
  assign n2956 = n2955 ^ n2768;
  assign n2957 = ~x81 & ~n2956;
  assign n2958 = ~n2954 & ~n2957;
  assign n2959 = ~n2953 & n2958;
  assign n2960 = x81 & n2956;
  assign n2961 = ~n2959 & ~n2960;
  assign n2962 = n2961 ^ x82;
  assign n2963 = n2772 & n2835;
  assign n2964 = n2963 ^ n2774;
  assign n2965 = n2964 ^ n2961;
  assign n2966 = ~n2962 & n2965;
  assign n2967 = n2966 ^ x82;
  assign n2968 = n2967 ^ x83;
  assign n2969 = n2778 & n2835;
  assign n2970 = n2969 ^ n2780;
  assign n2971 = n2970 ^ n2967;
  assign n2972 = n2968 & ~n2971;
  assign n2973 = n2972 ^ x83;
  assign n2974 = n2973 ^ x84;
  assign n2975 = n2784 & n2835;
  assign n2976 = n2975 ^ n2786;
  assign n2977 = n2976 ^ n2973;
  assign n2978 = n2974 & ~n2977;
  assign n2979 = n2978 ^ x84;
  assign n2980 = n2979 ^ x85;
  assign n2981 = n2790 & n2835;
  assign n2982 = n2981 ^ n2792;
  assign n2983 = n2982 ^ n2979;
  assign n2984 = n2980 & ~n2983;
  assign n2985 = n2984 ^ x85;
  assign n2986 = n2985 ^ x86;
  assign n2987 = n2814 & n2835;
  assign n2988 = n2987 ^ n2817;
  assign n2989 = x89 & n2988;
  assign n2990 = n2796 & n2835;
  assign n2991 = n2990 ^ n2798;
  assign n2992 = n2991 ^ n2985;
  assign n2993 = n2986 & ~n2992;
  assign n2994 = n2993 ^ x86;
  assign n2995 = n2994 ^ x87;
  assign n2996 = n2802 & n2835;
  assign n2997 = n2996 ^ n2804;
  assign n2998 = n2997 ^ n2994;
  assign n2999 = n2995 & ~n2998;
  assign n3000 = n2999 ^ x87;
  assign n3001 = n3000 ^ x88;
  assign n3002 = n2808 & n2835;
  assign n3003 = n3002 ^ n2810;
  assign n3004 = n3003 ^ n3000;
  assign n3005 = n3001 & ~n3004;
  assign n3006 = n3005 ^ x88;
  assign n3007 = ~n2989 & ~n3006;
  assign n3008 = ~x89 & ~n2988;
  assign n3009 = n2821 & n2835;
  assign n3010 = n3009 ^ n2824;
  assign n3011 = ~n3008 & ~n3010;
  assign n3012 = ~n3007 & n3011;
  assign n3013 = ~x90 & ~n3012;
  assign n3014 = ~n3007 & ~n3008;
  assign n3015 = n3010 & ~n3014;
  assign n3016 = ~n3013 & ~n3015;
  assign n3017 = n3016 ^ x91;
  assign n3018 = x90 & n2827;
  assign n3019 = n165 & ~n242;
  assign n3020 = ~n3018 & n3019;
  assign n3021 = ~n2651 & ~n3020;
  assign n3022 = n3021 ^ n3016;
  assign n3023 = n3017 & n3022;
  assign n3024 = n3023 ^ x91;
  assign n3025 = n164 & ~n3024;
  assign n3026 = n2986 & n3025;
  assign n3027 = n3026 ^ n2991;
  assign n3028 = ~x87 & ~n3027;
  assign n3029 = n2995 & n3025;
  assign n3030 = n3029 ^ n2997;
  assign n3031 = ~x88 & ~n3030;
  assign n3032 = ~n3028 & ~n3031;
  assign n3033 = n2869 & n3025;
  assign n3034 = n3033 ^ n2872;
  assign n3035 = ~x68 & ~n3034;
  assign n3036 = n2876 & n3025;
  assign n3037 = n3036 ^ n2878;
  assign n3038 = ~x69 & ~n3037;
  assign n3039 = ~n3035 & ~n3038;
  assign n3040 = ~x35 & n2856;
  assign n3041 = ~n3025 & n3040;
  assign n3042 = ~x35 & x65;
  assign n3043 = x64 & n3042;
  assign n3044 = ~n3041 & ~n3043;
  assign n3045 = x64 & n3025;
  assign n3049 = ~x36 & x65;
  assign n3046 = x36 & ~x65;
  assign n3047 = x35 & n3046;
  assign n3048 = n3047 ^ x36;
  assign n3050 = n3049 ^ n3048;
  assign n3051 = n3045 & n3050;
  assign n3052 = n3051 ^ n3049;
  assign n3053 = n3044 & ~n3052;
  assign n3054 = n3053 ^ x66;
  assign n3055 = x65 & n164;
  assign n3056 = ~n2835 & n3055;
  assign n3057 = ~n3024 & n3056;
  assign n3058 = n219 & n2835;
  assign n3059 = ~n3057 & ~n3058;
  assign n3060 = x36 & ~n3059;
  assign n3061 = n2835 ^ x65;
  assign n3062 = n2856 & ~n3061;
  assign n3063 = ~n202 & ~n3062;
  assign n3064 = n3063 ^ n2851;
  assign n3065 = n3025 & ~n3064;
  assign n3066 = n3065 ^ n2851;
  assign n3067 = ~n3060 & ~n3066;
  assign n3068 = n3067 ^ x37;
  assign n3069 = n3068 ^ n3053;
  assign n3070 = ~n3054 & n3069;
  assign n3071 = n3070 ^ x66;
  assign n3072 = n3071 ^ x67;
  assign n3073 = n2865 ^ x66;
  assign n3074 = n3025 & ~n3073;
  assign n3075 = n3074 ^ n2849;
  assign n3076 = n3075 ^ n3071;
  assign n3077 = n3072 & ~n3076;
  assign n3078 = n3077 ^ x67;
  assign n3079 = n3039 & n3078;
  assign n3080 = n3037 ^ x69;
  assign n3081 = x68 & n3034;
  assign n3082 = n3081 ^ n3037;
  assign n3083 = n3080 & ~n3082;
  assign n3084 = n3083 ^ x69;
  assign n3085 = ~n3079 & ~n3084;
  assign n3086 = n3085 ^ x70;
  assign n3087 = n2882 & n3025;
  assign n3088 = n3087 ^ n2884;
  assign n3089 = n3088 ^ n3085;
  assign n3090 = ~n3086 & n3089;
  assign n3091 = n3090 ^ x70;
  assign n3092 = n3091 ^ x71;
  assign n3093 = n2888 & n3025;
  assign n3094 = n3093 ^ n2890;
  assign n3095 = n3094 ^ n3091;
  assign n3096 = n3092 & ~n3095;
  assign n3097 = n3096 ^ x71;
  assign n3098 = n3097 ^ x72;
  assign n3099 = n2894 & n3025;
  assign n3100 = n3099 ^ n2896;
  assign n3101 = n3100 ^ n3097;
  assign n3102 = n3098 & ~n3101;
  assign n3103 = n3102 ^ x72;
  assign n3104 = n3103 ^ x73;
  assign n3105 = n2900 & n3025;
  assign n3106 = n3105 ^ n2903;
  assign n3107 = n3106 ^ n3103;
  assign n3108 = n3104 & ~n3107;
  assign n3109 = n3108 ^ x73;
  assign n3110 = n3109 ^ x74;
  assign n3111 = n2907 & n3025;
  assign n3112 = n3111 ^ n2913;
  assign n3113 = n3112 ^ n3109;
  assign n3114 = n3110 & ~n3113;
  assign n3115 = n3114 ^ x74;
  assign n3116 = n3115 ^ x75;
  assign n3117 = n2917 & n3025;
  assign n3118 = n3117 ^ n2919;
  assign n3119 = n3118 ^ n3115;
  assign n3120 = n3116 & ~n3119;
  assign n3121 = n3120 ^ x75;
  assign n3122 = n3121 ^ x76;
  assign n3123 = n2923 & n3025;
  assign n3124 = n3123 ^ n2925;
  assign n3125 = n3124 ^ n3121;
  assign n3126 = n3122 & ~n3125;
  assign n3127 = n3126 ^ x76;
  assign n3128 = n3127 ^ x77;
  assign n3129 = n2929 & n3025;
  assign n3130 = n3129 ^ n2931;
  assign n3131 = n3130 ^ n3127;
  assign n3132 = n3128 & ~n3131;
  assign n3133 = n3132 ^ x77;
  assign n3134 = n3133 ^ x78;
  assign n3135 = n2935 & n3025;
  assign n3136 = n3135 ^ n2937;
  assign n3137 = n3136 ^ n3133;
  assign n3138 = n3134 & ~n3137;
  assign n3139 = n3138 ^ x78;
  assign n3140 = n3139 ^ x79;
  assign n3141 = n2941 & n3025;
  assign n3142 = n3141 ^ n2943;
  assign n3143 = n3142 ^ n3139;
  assign n3144 = n3140 & ~n3143;
  assign n3145 = n3144 ^ x79;
  assign n3146 = n3145 ^ x80;
  assign n3147 = n2947 & n3025;
  assign n3148 = n3147 ^ n2949;
  assign n3149 = n3148 ^ n3145;
  assign n3150 = n3146 & ~n3149;
  assign n3151 = n3150 ^ x80;
  assign n3152 = n3151 ^ x81;
  assign n3153 = n2952 ^ x80;
  assign n3154 = n3025 & n3153;
  assign n3155 = n3154 ^ n2837;
  assign n3156 = n3155 ^ n3151;
  assign n3157 = n3152 & ~n3156;
  assign n3158 = n3157 ^ x81;
  assign n3159 = n3158 ^ x82;
  assign n3160 = ~n2953 & ~n2954;
  assign n3161 = n3160 ^ x81;
  assign n3162 = n3025 & n3161;
  assign n3163 = n3162 ^ n2956;
  assign n3164 = n3163 ^ n3158;
  assign n3165 = n3159 & ~n3164;
  assign n3166 = n3165 ^ x82;
  assign n3167 = n3166 ^ x83;
  assign n3168 = ~n2962 & n3025;
  assign n3169 = n3168 ^ n2964;
  assign n3170 = n3169 ^ n3166;
  assign n3171 = n3167 & ~n3170;
  assign n3172 = n3171 ^ x83;
  assign n3173 = n3172 ^ x84;
  assign n3174 = n2968 & n3025;
  assign n3175 = n3174 ^ n2970;
  assign n3176 = n3175 ^ n3172;
  assign n3177 = n3173 & ~n3176;
  assign n3178 = n3177 ^ x84;
  assign n3179 = n3178 ^ x85;
  assign n3180 = n2974 & n3025;
  assign n3181 = n3180 ^ n2976;
  assign n3182 = n3181 ^ n3178;
  assign n3183 = n3179 & ~n3182;
  assign n3184 = n3183 ^ x85;
  assign n3185 = n3184 ^ x86;
  assign n3186 = n2980 & n3025;
  assign n3187 = n3186 ^ n2982;
  assign n3188 = n3187 ^ n3184;
  assign n3189 = n3185 & ~n3188;
  assign n3190 = n3189 ^ x86;
  assign n3191 = n3032 & n3190;
  assign n3192 = n3030 ^ x88;
  assign n3193 = x87 & n3027;
  assign n3194 = n3193 ^ n3030;
  assign n3195 = n3192 & ~n3194;
  assign n3196 = n3195 ^ x88;
  assign n3197 = ~n3191 & ~n3196;
  assign n3198 = n3001 & n3025;
  assign n3199 = n3198 ^ n3003;
  assign n3200 = x89 & n3199;
  assign n3201 = n3197 & ~n3200;
  assign n3202 = n3006 ^ x89;
  assign n3203 = n3025 & n3202;
  assign n3204 = n3203 ^ n2988;
  assign n3205 = ~x90 & ~n3204;
  assign n3206 = ~x89 & ~n3199;
  assign n3207 = ~n3205 & ~n3206;
  assign n3208 = ~n3201 & n3207;
  assign n3209 = x90 & n3204;
  assign n3210 = ~n3208 & ~n3209;
  assign n3211 = n3014 ^ x90;
  assign n3212 = n3025 & n3211;
  assign n3213 = n3212 ^ n3010;
  assign n3214 = ~x91 & n3213;
  assign n3215 = n3021 & ~n3025;
  assign n3216 = ~n242 & ~n3215;
  assign n3217 = ~x92 & ~n3216;
  assign n3218 = ~n3214 & ~n3217;
  assign n3219 = ~n3210 & n3218;
  assign n3220 = x91 & ~n3213;
  assign n3221 = ~n3217 & n3220;
  assign n3222 = x92 & n3216;
  assign n3223 = n163 & ~n3222;
  assign n3224 = ~n3221 & n3223;
  assign n3225 = ~n3219 & n3224;
  assign n3226 = n3197 ^ x89;
  assign n3227 = n3225 & ~n3226;
  assign n3228 = n3227 ^ n3199;
  assign n3229 = ~x90 & ~n3228;
  assign n3230 = ~n3201 & ~n3206;
  assign n3231 = n3230 ^ x90;
  assign n3232 = n3225 & n3231;
  assign n3233 = n3232 ^ n3204;
  assign n3234 = ~x91 & ~n3233;
  assign n3235 = ~n3229 & ~n3234;
  assign n3236 = n3116 & n3225;
  assign n3237 = n3236 ^ n3118;
  assign n3238 = ~x76 & ~n3237;
  assign n3239 = n3122 & n3225;
  assign n3240 = n3239 ^ n3124;
  assign n3241 = ~x77 & ~n3240;
  assign n3242 = ~n3238 & ~n3241;
  assign n3243 = ~x34 & ~x35;
  assign n3244 = ~n3225 & n3243;
  assign n3245 = ~x34 & x65;
  assign n3246 = ~n3244 & ~n3245;
  assign n3247 = x64 & ~n3246;
  assign n3248 = x64 & n3225;
  assign n3249 = x34 & ~x65;
  assign n3250 = x35 & ~n3249;
  assign n3251 = n3250 ^ n3042;
  assign n3252 = n3248 & n3251;
  assign n3253 = n3252 ^ n3042;
  assign n3254 = ~n3247 & ~n3253;
  assign n3255 = n3254 ^ x66;
  assign n3256 = x65 & n3025;
  assign n3257 = x35 & ~n3256;
  assign n3258 = n3225 & ~n3257;
  assign n3259 = n3045 & ~n3258;
  assign n3260 = n293 & ~n3025;
  assign n3261 = n3260 ^ x65;
  assign n3262 = ~x35 & n3261;
  assign n3263 = ~n202 & ~n3262;
  assign n3264 = x65 & n3257;
  assign n3265 = n3263 & ~n3264;
  assign n3266 = n3225 & ~n3265;
  assign n3267 = ~n3259 & ~n3266;
  assign n3268 = n3267 ^ x36;
  assign n3269 = n3268 ^ n3254;
  assign n3270 = ~n3255 & n3269;
  assign n3271 = n3270 ^ x66;
  assign n3272 = n3271 ^ x67;
  assign n3273 = ~n3054 & n3225;
  assign n3274 = n3273 ^ n3068;
  assign n3275 = n3274 ^ n3271;
  assign n3276 = n3272 & ~n3275;
  assign n3277 = n3276 ^ x67;
  assign n3278 = n3277 ^ x68;
  assign n3279 = n3072 & n3225;
  assign n3280 = n3279 ^ n3075;
  assign n3281 = n3280 ^ n3277;
  assign n3282 = n3278 & ~n3281;
  assign n3283 = n3282 ^ x68;
  assign n3284 = n3283 ^ x69;
  assign n3285 = n3078 ^ x68;
  assign n3286 = n3225 & n3285;
  assign n3287 = n3286 ^ n3034;
  assign n3288 = n3287 ^ n3283;
  assign n3289 = n3284 & ~n3288;
  assign n3290 = n3289 ^ x69;
  assign n3291 = n3290 ^ x70;
  assign n3292 = n3078 ^ n3034;
  assign n3293 = n3285 & ~n3292;
  assign n3294 = n3293 ^ x68;
  assign n3295 = n3294 ^ x69;
  assign n3296 = n3225 & n3295;
  assign n3297 = n3296 ^ n3037;
  assign n3298 = n3297 ^ n3290;
  assign n3299 = n3291 & ~n3298;
  assign n3300 = n3299 ^ x70;
  assign n3301 = n3300 ^ x71;
  assign n3302 = ~n3086 & n3225;
  assign n3303 = n3302 ^ n3088;
  assign n3304 = n3303 ^ n3300;
  assign n3305 = n3301 & ~n3304;
  assign n3306 = n3305 ^ x71;
  assign n3307 = n3306 ^ x72;
  assign n3308 = n3092 & n3225;
  assign n3309 = n3308 ^ n3094;
  assign n3310 = n3309 ^ n3306;
  assign n3311 = n3307 & ~n3310;
  assign n3312 = n3311 ^ x72;
  assign n3313 = n3312 ^ x73;
  assign n3314 = n3098 & n3225;
  assign n3315 = n3314 ^ n3100;
  assign n3316 = n3315 ^ n3312;
  assign n3317 = n3313 & ~n3316;
  assign n3318 = n3317 ^ x73;
  assign n3319 = n3318 ^ x74;
  assign n3320 = n3104 & n3225;
  assign n3321 = n3320 ^ n3106;
  assign n3322 = n3321 ^ n3318;
  assign n3323 = n3319 & ~n3322;
  assign n3324 = n3323 ^ x74;
  assign n3325 = n3324 ^ x75;
  assign n3326 = n3110 & n3225;
  assign n3327 = n3326 ^ n3112;
  assign n3328 = n3327 ^ n3324;
  assign n3329 = n3325 & ~n3328;
  assign n3330 = n3329 ^ x75;
  assign n3331 = n3242 & n3330;
  assign n3332 = n3240 ^ x77;
  assign n3333 = x76 & n3237;
  assign n3334 = n3333 ^ n3240;
  assign n3335 = n3332 & ~n3334;
  assign n3336 = n3335 ^ x77;
  assign n3337 = ~n3331 & ~n3336;
  assign n3338 = n3337 ^ x78;
  assign n3339 = n3128 & n3225;
  assign n3340 = n3339 ^ n3130;
  assign n3341 = n3340 ^ n3337;
  assign n3342 = ~n3338 & n3341;
  assign n3343 = n3342 ^ x78;
  assign n3344 = n3343 ^ x79;
  assign n3345 = n3134 & n3225;
  assign n3346 = n3345 ^ n3136;
  assign n3347 = n3346 ^ n3343;
  assign n3348 = n3344 & ~n3347;
  assign n3349 = n3348 ^ x79;
  assign n3350 = n3349 ^ x80;
  assign n3351 = n3140 & n3225;
  assign n3352 = n3351 ^ n3142;
  assign n3353 = n3352 ^ n3349;
  assign n3354 = n3350 & ~n3353;
  assign n3355 = n3354 ^ x80;
  assign n3356 = n3355 ^ x81;
  assign n3357 = n3146 & n3225;
  assign n3358 = n3357 ^ n3148;
  assign n3359 = n3358 ^ n3355;
  assign n3360 = n3356 & ~n3359;
  assign n3361 = n3360 ^ x81;
  assign n3362 = n3361 ^ x82;
  assign n3363 = n3152 & n3225;
  assign n3364 = n3363 ^ n3155;
  assign n3365 = n3364 ^ n3361;
  assign n3366 = n3362 & ~n3365;
  assign n3367 = n3366 ^ x82;
  assign n3368 = n3367 ^ x83;
  assign n3369 = n3159 & n3225;
  assign n3370 = n3369 ^ n3163;
  assign n3371 = n3370 ^ n3367;
  assign n3372 = n3368 & ~n3371;
  assign n3373 = n3372 ^ x83;
  assign n3374 = n3373 ^ x84;
  assign n3375 = n3167 & n3225;
  assign n3376 = n3375 ^ n3169;
  assign n3377 = n3376 ^ n3373;
  assign n3378 = n3374 & ~n3377;
  assign n3379 = n3378 ^ x84;
  assign n3380 = n3379 ^ x85;
  assign n3381 = n3173 & n3225;
  assign n3382 = n3381 ^ n3175;
  assign n3383 = n3382 ^ n3379;
  assign n3384 = n3380 & ~n3383;
  assign n3385 = n3384 ^ x85;
  assign n3386 = n3385 ^ x86;
  assign n3387 = n3179 & n3225;
  assign n3388 = n3387 ^ n3181;
  assign n3389 = n3388 ^ n3385;
  assign n3390 = n3386 & ~n3389;
  assign n3391 = n3390 ^ x86;
  assign n3392 = n3391 ^ x87;
  assign n3393 = n3185 & n3225;
  assign n3394 = n3393 ^ n3187;
  assign n3395 = n3394 ^ n3391;
  assign n3396 = n3392 & ~n3395;
  assign n3397 = n3396 ^ x87;
  assign n3398 = n3397 ^ x88;
  assign n3399 = n3190 ^ x87;
  assign n3400 = n3225 & n3399;
  assign n3401 = n3400 ^ n3027;
  assign n3402 = n3401 ^ n3397;
  assign n3403 = n3398 & ~n3402;
  assign n3404 = n3403 ^ x88;
  assign n3405 = n3404 ^ x89;
  assign n3406 = n3190 ^ n3027;
  assign n3407 = n3399 & ~n3406;
  assign n3408 = n3407 ^ x87;
  assign n3409 = n3408 ^ x88;
  assign n3410 = n3225 & n3409;
  assign n3411 = n3410 ^ n3030;
  assign n3412 = n3411 ^ n3404;
  assign n3413 = n3405 & ~n3412;
  assign n3414 = n3413 ^ x89;
  assign n3415 = n3235 & n3414;
  assign n3416 = n3233 ^ x91;
  assign n3417 = x90 & n3228;
  assign n3418 = n3417 ^ n3233;
  assign n3419 = n3416 & ~n3418;
  assign n3420 = n3419 ^ x91;
  assign n3421 = ~n3415 & ~n3420;
  assign n3422 = n3421 ^ x92;
  assign n3423 = ~n3216 & ~n3225;
  assign n3424 = ~n242 & ~n3423;
  assign n3425 = ~x93 & ~n3424;
  assign n3426 = n3210 ^ x91;
  assign n3427 = n3225 & ~n3426;
  assign n3428 = n3427 ^ n3213;
  assign n3429 = n3428 ^ n3421;
  assign n3430 = ~n3422 & ~n3429;
  assign n3431 = n3430 ^ x92;
  assign n3432 = ~n3425 & n3431;
  assign n3433 = x93 & n3424;
  assign n3434 = n162 & ~n3433;
  assign n3435 = ~n3432 & n3434;
  assign n3436 = ~n3422 & n3435;
  assign n3437 = n3436 ^ n3428;
  assign n3438 = ~x93 & n3437;
  assign n3439 = n162 & ~n3431;
  assign n3440 = ~n163 & ~n3424;
  assign n3441 = ~n3439 & n3440;
  assign n3442 = ~x94 & n3441;
  assign n3443 = ~n3438 & ~n3442;
  assign n3444 = n3362 & n3435;
  assign n3445 = n3444 ^ n3364;
  assign n3446 = ~x83 & ~n3445;
  assign n3447 = n3368 & n3435;
  assign n3448 = n3447 ^ n3370;
  assign n3449 = ~x84 & ~n3448;
  assign n3450 = ~n3446 & ~n3449;
  assign n3451 = x64 & n3435;
  assign n3452 = ~n3245 & ~n3451;
  assign n3453 = x33 & ~x65;
  assign n3454 = ~n3452 & ~n3453;
  assign n3455 = ~x34 & n3451;
  assign n3456 = n3454 & ~n3455;
  assign n3457 = ~x65 & n3435;
  assign n3458 = ~x33 & x64;
  assign n3459 = ~n3249 & n3458;
  assign n3460 = ~n3457 & n3459;
  assign n3461 = ~n3456 & ~n3460;
  assign n3462 = n3461 ^ x66;
  assign n3463 = x65 & n3225;
  assign n3464 = x34 & ~n3463;
  assign n3465 = n3435 & ~n3464;
  assign n3466 = n3248 & ~n3465;
  assign n3467 = n293 & ~n3225;
  assign n3468 = n3467 ^ x65;
  assign n3469 = ~x34 & n3468;
  assign n3470 = ~n202 & ~n3469;
  assign n3471 = x65 & n3464;
  assign n3472 = n3470 & ~n3471;
  assign n3473 = n3435 & ~n3472;
  assign n3474 = ~n3466 & ~n3473;
  assign n3475 = n3474 ^ x35;
  assign n3476 = n3475 ^ n3461;
  assign n3477 = ~n3462 & n3476;
  assign n3478 = n3477 ^ x66;
  assign n3479 = n3478 ^ x67;
  assign n3480 = ~n3255 & n3435;
  assign n3481 = n3480 ^ n3268;
  assign n3482 = n3481 ^ n3478;
  assign n3483 = n3479 & ~n3482;
  assign n3484 = n3483 ^ x67;
  assign n3485 = n3484 ^ x68;
  assign n3486 = n3272 & n3435;
  assign n3487 = n3486 ^ n3274;
  assign n3488 = n3487 ^ n3484;
  assign n3489 = n3485 & ~n3488;
  assign n3490 = n3489 ^ x68;
  assign n3491 = n3490 ^ x69;
  assign n3492 = n3278 & n3435;
  assign n3493 = n3492 ^ n3280;
  assign n3494 = n3493 ^ n3490;
  assign n3495 = n3491 & ~n3494;
  assign n3496 = n3495 ^ x69;
  assign n3497 = n3496 ^ x70;
  assign n3498 = n3284 & n3435;
  assign n3499 = n3498 ^ n3287;
  assign n3500 = n3499 ^ n3496;
  assign n3501 = n3497 & ~n3500;
  assign n3502 = n3501 ^ x70;
  assign n3503 = n3502 ^ x71;
  assign n3504 = n3291 & n3435;
  assign n3505 = n3504 ^ n3297;
  assign n3506 = n3505 ^ n3502;
  assign n3507 = n3503 & ~n3506;
  assign n3508 = n3507 ^ x71;
  assign n3509 = n3508 ^ x72;
  assign n3510 = n3301 & n3435;
  assign n3511 = n3510 ^ n3303;
  assign n3512 = n3511 ^ n3508;
  assign n3513 = n3509 & ~n3512;
  assign n3514 = n3513 ^ x72;
  assign n3515 = n3514 ^ x73;
  assign n3516 = n3307 & n3435;
  assign n3517 = n3516 ^ n3309;
  assign n3518 = n3517 ^ n3514;
  assign n3519 = n3515 & ~n3518;
  assign n3520 = n3519 ^ x73;
  assign n3521 = n3520 ^ x74;
  assign n3522 = n3313 & n3435;
  assign n3523 = n3522 ^ n3315;
  assign n3524 = n3523 ^ n3520;
  assign n3525 = n3521 & ~n3524;
  assign n3526 = n3525 ^ x74;
  assign n3527 = n3526 ^ x75;
  assign n3528 = n3319 & n3435;
  assign n3529 = n3528 ^ n3321;
  assign n3530 = n3529 ^ n3526;
  assign n3531 = n3527 & ~n3530;
  assign n3532 = n3531 ^ x75;
  assign n3533 = n3532 ^ x76;
  assign n3534 = n3325 & n3435;
  assign n3535 = n3534 ^ n3327;
  assign n3536 = n3535 ^ n3532;
  assign n3537 = n3533 & ~n3536;
  assign n3538 = n3537 ^ x76;
  assign n3539 = n3538 ^ x77;
  assign n3540 = n3330 ^ x76;
  assign n3541 = n3435 & n3540;
  assign n3542 = n3541 ^ n3237;
  assign n3543 = n3542 ^ n3538;
  assign n3544 = n3539 & ~n3543;
  assign n3545 = n3544 ^ x77;
  assign n3546 = n3545 ^ x78;
  assign n3547 = n3330 ^ n3237;
  assign n3548 = n3540 & ~n3547;
  assign n3549 = n3548 ^ x76;
  assign n3550 = n3549 ^ x77;
  assign n3551 = n3435 & n3550;
  assign n3552 = n3551 ^ n3240;
  assign n3553 = n3552 ^ n3545;
  assign n3554 = n3546 & ~n3553;
  assign n3555 = n3554 ^ x78;
  assign n3556 = n3555 ^ x79;
  assign n3557 = ~n3338 & n3435;
  assign n3558 = n3557 ^ n3340;
  assign n3559 = n3558 ^ n3555;
  assign n3560 = n3556 & ~n3559;
  assign n3561 = n3560 ^ x79;
  assign n3562 = n3561 ^ x80;
  assign n3563 = n3344 & n3435;
  assign n3564 = n3563 ^ n3346;
  assign n3565 = n3564 ^ n3561;
  assign n3566 = n3562 & ~n3565;
  assign n3567 = n3566 ^ x80;
  assign n3568 = n3567 ^ x81;
  assign n3569 = n3350 & n3435;
  assign n3570 = n3569 ^ n3352;
  assign n3571 = n3570 ^ n3567;
  assign n3572 = n3568 & ~n3571;
  assign n3573 = n3572 ^ x81;
  assign n3574 = n3573 ^ x82;
  assign n3575 = n3356 & n3435;
  assign n3576 = n3575 ^ n3358;
  assign n3577 = n3576 ^ n3573;
  assign n3578 = n3574 & ~n3577;
  assign n3579 = n3578 ^ x82;
  assign n3580 = n3450 & n3579;
  assign n3581 = n3448 ^ x84;
  assign n3582 = x83 & n3445;
  assign n3583 = n3582 ^ n3448;
  assign n3584 = n3581 & ~n3583;
  assign n3585 = n3584 ^ x84;
  assign n3586 = ~n3580 & ~n3585;
  assign n3587 = n3586 ^ x85;
  assign n3588 = n3374 & n3435;
  assign n3589 = n3588 ^ n3376;
  assign n3590 = n3589 ^ n3586;
  assign n3591 = ~n3587 & n3590;
  assign n3592 = n3591 ^ x85;
  assign n3593 = n3592 ^ x86;
  assign n3594 = n3380 & n3435;
  assign n3595 = n3594 ^ n3382;
  assign n3596 = n3595 ^ n3592;
  assign n3597 = n3593 & ~n3596;
  assign n3598 = n3597 ^ x86;
  assign n3599 = n3598 ^ x87;
  assign n3600 = n3386 & n3435;
  assign n3601 = n3600 ^ n3388;
  assign n3602 = n3601 ^ n3598;
  assign n3603 = n3599 & ~n3602;
  assign n3604 = n3603 ^ x87;
  assign n3605 = n3604 ^ x88;
  assign n3606 = n3392 & n3435;
  assign n3607 = n3606 ^ n3394;
  assign n3608 = n3607 ^ n3604;
  assign n3609 = n3605 & ~n3608;
  assign n3610 = n3609 ^ x88;
  assign n3611 = n3610 ^ x89;
  assign n3612 = n3398 & n3435;
  assign n3613 = n3612 ^ n3401;
  assign n3614 = n3613 ^ n3610;
  assign n3615 = n3611 & ~n3614;
  assign n3616 = n3615 ^ x89;
  assign n3617 = n3616 ^ x90;
  assign n3618 = n3405 & n3435;
  assign n3619 = n3618 ^ n3411;
  assign n3620 = n3619 ^ n3616;
  assign n3621 = n3617 & ~n3620;
  assign n3622 = n3621 ^ x90;
  assign n3623 = n3622 ^ x91;
  assign n3624 = n3414 ^ x90;
  assign n3625 = n3435 & n3624;
  assign n3626 = n3625 ^ n3228;
  assign n3627 = n3626 ^ n3622;
  assign n3628 = n3623 & ~n3627;
  assign n3629 = n3628 ^ x91;
  assign n3630 = n3629 ^ x92;
  assign n3631 = n3414 ^ n3228;
  assign n3632 = n3624 & ~n3631;
  assign n3633 = n3632 ^ x90;
  assign n3634 = n3633 ^ x91;
  assign n3635 = n3435 & n3634;
  assign n3636 = n3635 ^ n3233;
  assign n3637 = n3636 ^ n3629;
  assign n3638 = n3630 & ~n3637;
  assign n3639 = n3638 ^ x92;
  assign n3640 = n3443 & n3639;
  assign n3641 = x93 & ~n3442;
  assign n3642 = ~n3437 & n3641;
  assign n3643 = n161 & ~n3424;
  assign n3644 = ~n162 & ~n3643;
  assign n3645 = ~n3642 & ~n3644;
  assign n3646 = ~n3640 & n3645;
  assign n3647 = n3639 ^ x93;
  assign n3648 = n3646 & n3647;
  assign n3649 = n3648 ^ n3437;
  assign n3650 = ~x94 & n3649;
  assign n3651 = n3579 ^ x83;
  assign n3652 = n3579 ^ n3445;
  assign n3653 = n3651 & ~n3652;
  assign n3654 = n3653 ^ x83;
  assign n3655 = n3654 ^ x84;
  assign n3656 = n3646 & n3655;
  assign n3657 = n3656 ^ n3448;
  assign n3658 = ~x85 & ~n3657;
  assign n3659 = ~n3587 & n3646;
  assign n3660 = n3659 ^ n3589;
  assign n3661 = ~x86 & ~n3660;
  assign n3662 = ~n3658 & ~n3661;
  assign n3663 = x65 & n3435;
  assign n3664 = x33 & ~n3663;
  assign n3665 = n3646 & ~n3664;
  assign n3666 = n3451 & ~n3665;
  assign n3667 = n3435 ^ x65;
  assign n3668 = n3458 & ~n3667;
  assign n3669 = ~n202 & ~n3668;
  assign n3670 = x65 & n3664;
  assign n3671 = n3669 & ~n3670;
  assign n3672 = n3646 & ~n3671;
  assign n3673 = ~n3666 & ~n3672;
  assign n3674 = n3673 ^ x34;
  assign n3675 = n3674 ^ x66;
  assign n3676 = x64 & n3646;
  assign n3677 = x32 & n3453;
  assign n3678 = n3677 ^ x33;
  assign n3679 = n3676 & n3678;
  assign n3680 = ~x32 & n219;
  assign n3681 = n3680 ^ x65;
  assign n3682 = ~x33 & n3681;
  assign n3683 = ~n3646 & n3682;
  assign n3684 = x32 & x64;
  assign n3685 = x65 & ~n3684;
  assign n3686 = x33 & ~x64;
  assign n3687 = n3685 & ~n3686;
  assign n3688 = ~n3683 & ~n3687;
  assign n3689 = ~n3679 & n3688;
  assign n3690 = n3689 ^ n3674;
  assign n3691 = n3675 & n3690;
  assign n3692 = n3691 ^ x66;
  assign n3693 = n3692 ^ x67;
  assign n3694 = ~n3462 & n3646;
  assign n3695 = n3694 ^ n3475;
  assign n3696 = n3695 ^ n3692;
  assign n3697 = n3693 & ~n3696;
  assign n3698 = n3697 ^ x67;
  assign n3699 = n3698 ^ x68;
  assign n3700 = n3479 & n3646;
  assign n3701 = n3700 ^ n3481;
  assign n3702 = n3701 ^ n3698;
  assign n3703 = n3699 & ~n3702;
  assign n3704 = n3703 ^ x68;
  assign n3705 = n3704 ^ x69;
  assign n3706 = n3485 & n3646;
  assign n3707 = n3706 ^ n3487;
  assign n3708 = n3707 ^ n3704;
  assign n3709 = n3705 & ~n3708;
  assign n3710 = n3709 ^ x69;
  assign n3711 = n3710 ^ x70;
  assign n3712 = n3491 & n3646;
  assign n3713 = n3712 ^ n3493;
  assign n3714 = n3713 ^ n3710;
  assign n3715 = n3711 & ~n3714;
  assign n3716 = n3715 ^ x70;
  assign n3717 = n3716 ^ x71;
  assign n3718 = n3497 & n3646;
  assign n3719 = n3718 ^ n3499;
  assign n3720 = n3719 ^ n3716;
  assign n3721 = n3717 & ~n3720;
  assign n3722 = n3721 ^ x71;
  assign n3723 = n3722 ^ x72;
  assign n3724 = n3505 ^ x71;
  assign n3725 = n3724 ^ n3502;
  assign n3726 = n3725 ^ n3505;
  assign n3727 = n3646 & n3726;
  assign n3728 = n3727 ^ n3505;
  assign n3729 = n3728 ^ n3722;
  assign n3730 = n3723 & ~n3729;
  assign n3731 = n3730 ^ x72;
  assign n3732 = n3731 ^ x73;
  assign n3733 = n3509 & n3646;
  assign n3734 = n3733 ^ n3511;
  assign n3735 = n3734 ^ n3731;
  assign n3736 = n3732 & ~n3735;
  assign n3737 = n3736 ^ x73;
  assign n3738 = n3737 ^ x74;
  assign n3739 = n3515 & n3646;
  assign n3740 = n3739 ^ n3517;
  assign n3741 = n3740 ^ n3737;
  assign n3742 = n3738 & ~n3741;
  assign n3743 = n3742 ^ x74;
  assign n3744 = n3743 ^ x75;
  assign n3745 = n3521 & n3646;
  assign n3746 = n3745 ^ n3523;
  assign n3747 = n3746 ^ n3743;
  assign n3748 = n3744 & ~n3747;
  assign n3749 = n3748 ^ x75;
  assign n3750 = n3749 ^ x76;
  assign n3751 = n3527 & n3646;
  assign n3752 = n3751 ^ n3529;
  assign n3753 = n3752 ^ n3749;
  assign n3754 = n3750 & ~n3753;
  assign n3755 = n3754 ^ x76;
  assign n3756 = n3755 ^ x77;
  assign n3757 = n3533 & n3646;
  assign n3758 = n3757 ^ n3535;
  assign n3759 = n3758 ^ n3755;
  assign n3760 = n3756 & ~n3759;
  assign n3761 = n3760 ^ x77;
  assign n3762 = n3761 ^ x78;
  assign n3763 = n3539 & n3646;
  assign n3764 = n3763 ^ n3542;
  assign n3765 = n3764 ^ n3761;
  assign n3766 = n3762 & ~n3765;
  assign n3767 = n3766 ^ x78;
  assign n3768 = n3767 ^ x79;
  assign n3769 = n3546 & n3646;
  assign n3770 = n3769 ^ n3552;
  assign n3771 = n3770 ^ n3767;
  assign n3772 = n3768 & ~n3771;
  assign n3773 = n3772 ^ x79;
  assign n3774 = n3773 ^ x80;
  assign n3775 = n3556 & n3646;
  assign n3776 = n3775 ^ n3558;
  assign n3777 = n3776 ^ n3773;
  assign n3778 = n3774 & ~n3777;
  assign n3779 = n3778 ^ x80;
  assign n3780 = n3779 ^ x81;
  assign n3781 = n3562 & n3646;
  assign n3782 = n3781 ^ n3564;
  assign n3783 = n3782 ^ n3779;
  assign n3784 = n3780 & ~n3783;
  assign n3785 = n3784 ^ x81;
  assign n3786 = n3785 ^ x82;
  assign n3787 = n3568 & n3646;
  assign n3788 = n3787 ^ n3570;
  assign n3789 = n3788 ^ n3785;
  assign n3790 = n3786 & ~n3789;
  assign n3791 = n3790 ^ x82;
  assign n3792 = n3791 ^ x83;
  assign n3793 = n3574 & n3646;
  assign n3794 = n3793 ^ n3576;
  assign n3795 = n3794 ^ n3791;
  assign n3796 = n3792 & ~n3795;
  assign n3797 = n3796 ^ x83;
  assign n3798 = n3797 ^ x84;
  assign n3799 = n3646 & n3651;
  assign n3800 = n3799 ^ n3445;
  assign n3801 = n3800 ^ n3797;
  assign n3802 = n3798 & ~n3801;
  assign n3803 = n3802 ^ x84;
  assign n3804 = n3662 & n3803;
  assign n3805 = n3660 ^ x86;
  assign n3806 = x85 & n3657;
  assign n3807 = n3806 ^ n3660;
  assign n3808 = n3805 & ~n3807;
  assign n3809 = n3808 ^ x86;
  assign n3810 = ~n3804 & ~n3809;
  assign n3811 = n3810 ^ x87;
  assign n3812 = n3593 & n3646;
  assign n3813 = n3812 ^ n3595;
  assign n3814 = n3813 ^ n3810;
  assign n3815 = ~n3811 & n3814;
  assign n3816 = n3815 ^ x87;
  assign n3817 = n3816 ^ x88;
  assign n3818 = n3599 & n3646;
  assign n3819 = n3818 ^ n3601;
  assign n3820 = n3819 ^ n3816;
  assign n3821 = n3817 & ~n3820;
  assign n3822 = n3821 ^ x88;
  assign n3823 = n3822 ^ x89;
  assign n3824 = n3605 & n3646;
  assign n3825 = n3824 ^ n3607;
  assign n3826 = n3825 ^ n3822;
  assign n3827 = n3823 & ~n3826;
  assign n3828 = n3827 ^ x89;
  assign n3829 = n3828 ^ x90;
  assign n3830 = n3611 & n3646;
  assign n3831 = n3830 ^ n3613;
  assign n3832 = n3831 ^ n3828;
  assign n3833 = n3829 & ~n3832;
  assign n3834 = n3833 ^ x90;
  assign n3835 = n3834 ^ x91;
  assign n3836 = n3617 & n3646;
  assign n3837 = n3836 ^ n3619;
  assign n3838 = n3837 ^ n3834;
  assign n3839 = n3835 & ~n3838;
  assign n3840 = n3839 ^ x91;
  assign n3841 = n3840 ^ x92;
  assign n3842 = n3623 & n3646;
  assign n3843 = n3842 ^ n3626;
  assign n3844 = n3843 ^ n3840;
  assign n3845 = n3841 & ~n3844;
  assign n3846 = n3845 ^ x92;
  assign n3847 = n3846 ^ x93;
  assign n3848 = n3630 & n3646;
  assign n3849 = n3848 ^ n3636;
  assign n3850 = n3849 ^ n3846;
  assign n3851 = n3847 & ~n3850;
  assign n3852 = n3851 ^ x93;
  assign n3853 = ~n3650 & n3852;
  assign n3854 = n3441 & ~n3646;
  assign n3855 = ~n242 & ~n3854;
  assign n3856 = x95 & n3855;
  assign n3857 = n160 & ~n3856;
  assign n3858 = x94 & ~n3649;
  assign n3859 = n3857 & ~n3858;
  assign n3860 = ~n3853 & n3859;
  assign n3861 = n161 & ~n3855;
  assign n3862 = ~n3860 & ~n3861;
  assign n3863 = n3852 ^ x94;
  assign n3864 = ~n3862 & n3863;
  assign n3865 = n3864 ^ n3649;
  assign n3866 = ~x95 & n3865;
  assign n3867 = ~n3855 & n3862;
  assign n3868 = ~n242 & ~n3867;
  assign n3869 = ~x96 & ~n3868;
  assign n3870 = ~n3866 & ~n3869;
  assign n3871 = n3762 & ~n3862;
  assign n3872 = n3871 ^ n3764;
  assign n3873 = ~x79 & ~n3872;
  assign n3874 = n3768 & ~n3862;
  assign n3875 = n3874 ^ n3770;
  assign n3876 = ~x80 & ~n3875;
  assign n3877 = ~n3873 & ~n3876;
  assign n3878 = x65 & ~n3646;
  assign n3879 = ~n3862 & n3878;
  assign n3880 = n219 & n3646;
  assign n3881 = ~n3879 & ~n3880;
  assign n3882 = x32 & ~n3881;
  assign n3883 = n3646 ^ x65;
  assign n3884 = n341 & ~n3883;
  assign n3885 = x32 & n3884;
  assign n3886 = n3885 ^ n340;
  assign n3887 = ~n3862 & n3886;
  assign n3888 = n3887 ^ n3676;
  assign n3889 = ~n3882 & ~n3888;
  assign n3890 = n3889 ^ x33;
  assign n3891 = n3890 ^ x66;
  assign n3892 = ~x65 & n3862;
  assign n3893 = ~x31 & x64;
  assign n3894 = n3892 & ~n3893;
  assign n3895 = x31 & ~x65;
  assign n3896 = n3684 & ~n3895;
  assign n3897 = n3896 ^ x32;
  assign n3898 = ~n3862 & ~n3897;
  assign n3899 = n3898 ^ x32;
  assign n3900 = ~n3894 & ~n3899;
  assign n3901 = x32 ^ x31;
  assign n3902 = ~x64 & n3901;
  assign n3903 = n3902 ^ x31;
  assign n3904 = x65 & ~n3903;
  assign n3905 = ~n3900 & ~n3904;
  assign n3906 = n3905 ^ n3890;
  assign n3907 = n3891 & n3906;
  assign n3908 = n3907 ^ x66;
  assign n3909 = n3908 ^ x67;
  assign n3910 = n3689 ^ x66;
  assign n3911 = ~n3862 & ~n3910;
  assign n3912 = n3911 ^ n3674;
  assign n3913 = n3912 ^ n3908;
  assign n3914 = n3909 & ~n3913;
  assign n3915 = n3914 ^ x67;
  assign n3916 = n3915 ^ x68;
  assign n3917 = n3693 & ~n3862;
  assign n3918 = n3917 ^ n3695;
  assign n3919 = n3918 ^ n3915;
  assign n3920 = n3916 & ~n3919;
  assign n3921 = n3920 ^ x68;
  assign n3922 = n3921 ^ x69;
  assign n3923 = n3699 & ~n3862;
  assign n3924 = n3923 ^ n3701;
  assign n3925 = n3924 ^ n3921;
  assign n3926 = n3922 & ~n3925;
  assign n3927 = n3926 ^ x69;
  assign n3928 = n3927 ^ x70;
  assign n3929 = n3705 & ~n3862;
  assign n3930 = n3929 ^ n3707;
  assign n3931 = n3930 ^ n3927;
  assign n3932 = n3928 & ~n3931;
  assign n3933 = n3932 ^ x70;
  assign n3934 = n3933 ^ x71;
  assign n3935 = n3711 & ~n3862;
  assign n3936 = n3935 ^ n3713;
  assign n3937 = n3936 ^ n3933;
  assign n3938 = n3934 & ~n3937;
  assign n3939 = n3938 ^ x71;
  assign n3940 = n3939 ^ x72;
  assign n3941 = n3717 & ~n3862;
  assign n3942 = n3941 ^ n3719;
  assign n3943 = n3942 ^ n3939;
  assign n3944 = n3940 & ~n3943;
  assign n3945 = n3944 ^ x72;
  assign n3946 = n3945 ^ x73;
  assign n3947 = n3723 & ~n3862;
  assign n3948 = n3947 ^ n3728;
  assign n3949 = n3948 ^ n3945;
  assign n3950 = n3946 & ~n3949;
  assign n3951 = n3950 ^ x73;
  assign n3952 = n3951 ^ x74;
  assign n3953 = n3732 & ~n3862;
  assign n3954 = n3953 ^ n3734;
  assign n3955 = n3954 ^ n3951;
  assign n3956 = n3952 & ~n3955;
  assign n3957 = n3956 ^ x74;
  assign n3958 = n3957 ^ x75;
  assign n3959 = n3738 & ~n3862;
  assign n3960 = n3959 ^ n3740;
  assign n3961 = n3960 ^ n3957;
  assign n3962 = n3958 & ~n3961;
  assign n3963 = n3962 ^ x75;
  assign n3964 = n3963 ^ x76;
  assign n3965 = n3744 & ~n3862;
  assign n3966 = n3965 ^ n3746;
  assign n3967 = n3966 ^ n3963;
  assign n3968 = n3964 & ~n3967;
  assign n3969 = n3968 ^ x76;
  assign n3970 = n3969 ^ x77;
  assign n3971 = n3750 & ~n3862;
  assign n3972 = n3971 ^ n3752;
  assign n3973 = n3972 ^ n3969;
  assign n3974 = n3970 & ~n3973;
  assign n3975 = n3974 ^ x77;
  assign n3976 = n3975 ^ x78;
  assign n3977 = n3756 & ~n3862;
  assign n3978 = n3977 ^ n3758;
  assign n3979 = n3978 ^ n3975;
  assign n3980 = n3976 & ~n3979;
  assign n3981 = n3980 ^ x78;
  assign n3982 = n3877 & n3981;
  assign n3983 = n3875 ^ x80;
  assign n3984 = x79 & n3872;
  assign n3985 = n3984 ^ n3875;
  assign n3986 = n3983 & ~n3985;
  assign n3987 = n3986 ^ x80;
  assign n3988 = ~n3982 & ~n3987;
  assign n3989 = n3988 ^ x81;
  assign n3990 = n3774 & ~n3862;
  assign n3991 = n3990 ^ n3776;
  assign n3992 = n3991 ^ n3988;
  assign n3993 = ~n3989 & n3992;
  assign n3994 = n3993 ^ x81;
  assign n3995 = n3994 ^ x82;
  assign n3996 = n3780 & ~n3862;
  assign n3997 = n3996 ^ n3782;
  assign n3998 = n3997 ^ n3994;
  assign n3999 = n3995 & ~n3998;
  assign n4000 = n3999 ^ x82;
  assign n4001 = n4000 ^ x83;
  assign n4002 = n3786 & ~n3862;
  assign n4003 = n4002 ^ n3788;
  assign n4004 = n4003 ^ n4000;
  assign n4005 = n4001 & ~n4004;
  assign n4006 = n4005 ^ x83;
  assign n4007 = n4006 ^ x84;
  assign n4008 = n3792 & ~n3862;
  assign n4009 = n4008 ^ n3794;
  assign n4010 = n4009 ^ n4006;
  assign n4011 = n4007 & ~n4010;
  assign n4012 = n4011 ^ x84;
  assign n4013 = n4012 ^ x85;
  assign n4014 = n3798 & ~n3862;
  assign n4015 = n4014 ^ n3800;
  assign n4016 = n4015 ^ n4012;
  assign n4017 = n4013 & ~n4016;
  assign n4018 = n4017 ^ x85;
  assign n4019 = n4018 ^ x86;
  assign n4020 = n3803 ^ x85;
  assign n4021 = ~n3862 & n4020;
  assign n4022 = n4021 ^ n3657;
  assign n4023 = n4022 ^ n4018;
  assign n4024 = n4019 & ~n4023;
  assign n4025 = n4024 ^ x86;
  assign n4026 = n4025 ^ x87;
  assign n4027 = n3803 ^ n3657;
  assign n4028 = n4020 & ~n4027;
  assign n4029 = n4028 ^ x85;
  assign n4030 = n4029 ^ x86;
  assign n4031 = ~n3862 & n4030;
  assign n4032 = n4031 ^ n3660;
  assign n4033 = n4032 ^ n4025;
  assign n4034 = n4026 & ~n4033;
  assign n4035 = n4034 ^ x87;
  assign n4036 = n4035 ^ x88;
  assign n4037 = ~n3811 & ~n3862;
  assign n4038 = n4037 ^ n3813;
  assign n4039 = n4038 ^ n4035;
  assign n4040 = n4036 & ~n4039;
  assign n4041 = n4040 ^ x88;
  assign n4042 = n4041 ^ x89;
  assign n4043 = n3817 & ~n3862;
  assign n4044 = n4043 ^ n3819;
  assign n4045 = n4044 ^ n4041;
  assign n4046 = n4042 & ~n4045;
  assign n4047 = n4046 ^ x89;
  assign n4048 = n4047 ^ x90;
  assign n4049 = n3823 & ~n3862;
  assign n4050 = n4049 ^ n3825;
  assign n4051 = n4050 ^ n4047;
  assign n4052 = n4048 & ~n4051;
  assign n4053 = n4052 ^ x90;
  assign n4054 = n4053 ^ x91;
  assign n4055 = n3829 & ~n3862;
  assign n4056 = n4055 ^ n3831;
  assign n4057 = n4056 ^ n4053;
  assign n4058 = n4054 & ~n4057;
  assign n4059 = n4058 ^ x91;
  assign n4060 = n4059 ^ x92;
  assign n4061 = n3835 & ~n3862;
  assign n4062 = n4061 ^ n3837;
  assign n4063 = n4062 ^ n4059;
  assign n4064 = n4060 & ~n4063;
  assign n4065 = n4064 ^ x92;
  assign n4066 = n4065 ^ x93;
  assign n4067 = n3841 & ~n3862;
  assign n4068 = n4067 ^ n3843;
  assign n4069 = n4068 ^ n4065;
  assign n4070 = n4066 & ~n4069;
  assign n4071 = n4070 ^ x93;
  assign n4072 = n4071 ^ x94;
  assign n4073 = n3847 & ~n3862;
  assign n4074 = n4073 ^ n3849;
  assign n4075 = n4074 ^ n4071;
  assign n4076 = n4072 & ~n4075;
  assign n4077 = n4076 ^ x94;
  assign n4078 = n3870 & n4077;
  assign n4079 = x95 & ~n3869;
  assign n4080 = ~n3865 & n4079;
  assign n4081 = x96 & n3868;
  assign n4082 = n155 & n157;
  assign n4083 = n156 & n4082;
  assign n4084 = ~n4081 & n4083;
  assign n4085 = ~n4080 & n4084;
  assign n4086 = ~n4078 & n4085;
  assign n4087 = n4077 ^ x95;
  assign n4088 = n4086 & n4087;
  assign n4089 = n4088 ^ n3865;
  assign n4090 = x96 & ~n4089;
  assign n4091 = x65 & ~n3862;
  assign n4092 = x31 & ~n4091;
  assign n4093 = n4086 & ~n4092;
  assign n4094 = x64 & ~n3862;
  assign n4095 = ~n4093 & n4094;
  assign n4096 = n3862 ^ x65;
  assign n4097 = n3893 & n4096;
  assign n4098 = ~n202 & ~n4097;
  assign n4099 = x65 & n4092;
  assign n4100 = n4098 & ~n4099;
  assign n4101 = n4086 & ~n4100;
  assign n4102 = ~n4095 & ~n4101;
  assign n4103 = n4102 ^ x32;
  assign n4104 = n4103 ^ x66;
  assign n4105 = x64 & n4086;
  assign n4106 = x30 & n3895;
  assign n4107 = n4106 ^ x31;
  assign n4108 = n4105 & n4107;
  assign n4109 = ~x30 & n3893;
  assign n4110 = ~x31 & x65;
  assign n4111 = ~n4109 & ~n4110;
  assign n4112 = ~n4086 & ~n4111;
  assign n4113 = ~x30 & x65;
  assign n4114 = n4113 ^ n4110;
  assign n4115 = x64 & n4114;
  assign n4116 = n4115 ^ n4110;
  assign n4117 = ~n4112 & ~n4116;
  assign n4118 = ~n4108 & n4117;
  assign n4119 = n4118 ^ n4103;
  assign n4120 = n4104 & n4119;
  assign n4121 = n4120 ^ x66;
  assign n4122 = n4121 ^ x67;
  assign n4123 = n3905 ^ x66;
  assign n4124 = n4086 & ~n4123;
  assign n4125 = n4124 ^ n3890;
  assign n4126 = n4125 ^ n4121;
  assign n4127 = n4122 & ~n4126;
  assign n4128 = n4127 ^ x67;
  assign n4129 = n4128 ^ x68;
  assign n4130 = n3909 & n4086;
  assign n4131 = n4130 ^ n3912;
  assign n4132 = n4131 ^ n4128;
  assign n4133 = n4129 & ~n4132;
  assign n4134 = n4133 ^ x68;
  assign n4135 = n4134 ^ x69;
  assign n4136 = n3916 & n4086;
  assign n4137 = n4136 ^ n3918;
  assign n4138 = n4137 ^ n4134;
  assign n4139 = n4135 & ~n4138;
  assign n4140 = n4139 ^ x69;
  assign n4141 = n4140 ^ x70;
  assign n4142 = n3922 & n4086;
  assign n4143 = n4142 ^ n3924;
  assign n4144 = n4143 ^ n4140;
  assign n4145 = n4141 & ~n4144;
  assign n4146 = n4145 ^ x70;
  assign n4147 = n4146 ^ x71;
  assign n4148 = n3928 & n4086;
  assign n4149 = n4148 ^ n3930;
  assign n4150 = n4149 ^ n4146;
  assign n4151 = n4147 & ~n4150;
  assign n4152 = n4151 ^ x71;
  assign n4153 = n4152 ^ x72;
  assign n4154 = n3934 & n4086;
  assign n4155 = n4154 ^ n3936;
  assign n4156 = n4155 ^ n4152;
  assign n4157 = n4153 & ~n4156;
  assign n4158 = n4157 ^ x72;
  assign n4159 = n4158 ^ x73;
  assign n4160 = n3940 & n4086;
  assign n4161 = n4160 ^ n3942;
  assign n4162 = n4161 ^ n4158;
  assign n4163 = n4159 & ~n4162;
  assign n4164 = n4163 ^ x73;
  assign n4165 = n4164 ^ x74;
  assign n4166 = n3946 & n4086;
  assign n4167 = n4166 ^ n3948;
  assign n4168 = n4167 ^ n4164;
  assign n4169 = n4165 & ~n4168;
  assign n4170 = n4169 ^ x74;
  assign n4171 = n4170 ^ x75;
  assign n4172 = n3952 & n4086;
  assign n4173 = n4172 ^ n3954;
  assign n4174 = n4173 ^ n4170;
  assign n4175 = n4171 & ~n4174;
  assign n4176 = n4175 ^ x75;
  assign n4177 = n4176 ^ x76;
  assign n4178 = n3958 & n4086;
  assign n4179 = n4178 ^ n3960;
  assign n4180 = n4179 ^ n4176;
  assign n4181 = n4177 & ~n4180;
  assign n4182 = n4181 ^ x76;
  assign n4183 = n4182 ^ x77;
  assign n4184 = n3964 & n4086;
  assign n4185 = n4184 ^ n3966;
  assign n4186 = n4185 ^ n4182;
  assign n4187 = n4183 & ~n4186;
  assign n4188 = n4187 ^ x77;
  assign n4189 = n4188 ^ x78;
  assign n4190 = n3970 & n4086;
  assign n4191 = n4190 ^ n3972;
  assign n4192 = n4191 ^ n4188;
  assign n4193 = n4189 & ~n4192;
  assign n4194 = n4193 ^ x78;
  assign n4195 = n4194 ^ x79;
  assign n4196 = n3976 & n4086;
  assign n4197 = n4196 ^ n3978;
  assign n4198 = n4197 ^ n4194;
  assign n4199 = n4195 & ~n4198;
  assign n4200 = n4199 ^ x79;
  assign n4201 = n4200 ^ x80;
  assign n4202 = n3981 ^ x79;
  assign n4203 = n4086 & n4202;
  assign n4204 = n4203 ^ n3872;
  assign n4205 = n4204 ^ n4200;
  assign n4206 = n4201 & ~n4205;
  assign n4207 = n4206 ^ x80;
  assign n4208 = n4207 ^ x81;
  assign n4209 = n3981 ^ n3872;
  assign n4210 = n4202 & ~n4209;
  assign n4211 = n4210 ^ x79;
  assign n4212 = n4211 ^ x80;
  assign n4213 = n4086 & n4212;
  assign n4214 = n4213 ^ n3875;
  assign n4215 = n4214 ^ n4207;
  assign n4216 = n4208 & ~n4215;
  assign n4217 = n4216 ^ x81;
  assign n4218 = n4217 ^ x82;
  assign n4219 = ~n3989 & n4086;
  assign n4220 = n4219 ^ n3991;
  assign n4221 = n4220 ^ n4217;
  assign n4222 = n4218 & ~n4221;
  assign n4223 = n4222 ^ x82;
  assign n4224 = n4223 ^ x83;
  assign n4225 = n3995 & n4086;
  assign n4226 = n4225 ^ n3997;
  assign n4227 = n4226 ^ n4223;
  assign n4228 = n4224 & ~n4227;
  assign n4229 = n4228 ^ x83;
  assign n4230 = n4229 ^ x84;
  assign n4231 = n4001 & n4086;
  assign n4232 = n4231 ^ n4003;
  assign n4233 = n4232 ^ n4229;
  assign n4234 = n4230 & ~n4233;
  assign n4235 = n4234 ^ x84;
  assign n4236 = n4235 ^ x85;
  assign n4237 = n4007 & n4086;
  assign n4238 = n4237 ^ n4009;
  assign n4239 = n4238 ^ n4235;
  assign n4240 = n4236 & ~n4239;
  assign n4241 = n4240 ^ x85;
  assign n4242 = n4241 ^ x86;
  assign n4243 = n4013 & n4086;
  assign n4244 = n4243 ^ n4015;
  assign n4245 = n4244 ^ n4241;
  assign n4246 = n4242 & ~n4245;
  assign n4247 = n4246 ^ x86;
  assign n4248 = n4247 ^ x87;
  assign n4249 = n4019 & n4086;
  assign n4250 = n4249 ^ n4022;
  assign n4251 = n4250 ^ n4247;
  assign n4252 = n4248 & ~n4251;
  assign n4253 = n4252 ^ x87;
  assign n4254 = n4253 ^ x88;
  assign n4255 = n4026 & n4086;
  assign n4256 = n4255 ^ n4032;
  assign n4257 = n4256 ^ n4253;
  assign n4258 = n4254 & ~n4257;
  assign n4259 = n4258 ^ x88;
  assign n4260 = n4259 ^ x89;
  assign n4261 = n4036 & n4086;
  assign n4262 = n4261 ^ n4038;
  assign n4263 = n4262 ^ n4259;
  assign n4264 = n4260 & ~n4263;
  assign n4265 = n4264 ^ x89;
  assign n4266 = n4265 ^ x90;
  assign n4267 = n4042 & n4086;
  assign n4268 = n4267 ^ n4044;
  assign n4269 = n4268 ^ n4265;
  assign n4270 = n4266 & ~n4269;
  assign n4271 = n4270 ^ x90;
  assign n4272 = n4271 ^ x91;
  assign n4273 = n4048 & n4086;
  assign n4274 = n4273 ^ n4050;
  assign n4275 = n4274 ^ n4271;
  assign n4276 = n4272 & ~n4275;
  assign n4277 = n4276 ^ x91;
  assign n4278 = n4277 ^ x92;
  assign n4279 = n4054 & n4086;
  assign n4280 = n4279 ^ n4056;
  assign n4281 = n4280 ^ n4277;
  assign n4282 = n4278 & ~n4281;
  assign n4283 = n4282 ^ x92;
  assign n4284 = n4283 ^ x93;
  assign n4285 = n4060 & n4086;
  assign n4286 = n4285 ^ n4062;
  assign n4287 = n4286 ^ n4283;
  assign n4288 = n4284 & ~n4287;
  assign n4289 = n4288 ^ x93;
  assign n4290 = n4289 ^ x94;
  assign n4291 = n4066 & n4086;
  assign n4292 = n4291 ^ n4068;
  assign n4293 = n4292 ^ n4289;
  assign n4294 = n4290 & ~n4293;
  assign n4295 = n4294 ^ x94;
  assign n4296 = n4295 ^ x95;
  assign n4297 = n4072 & n4086;
  assign n4298 = n4297 ^ n4074;
  assign n4299 = n4298 ^ n4295;
  assign n4300 = n4296 & ~n4299;
  assign n4301 = n4300 ^ x95;
  assign n4302 = ~n4090 & ~n4301;
  assign n4303 = x96 & ~n3866;
  assign n4304 = n4077 & n4303;
  assign n4305 = x95 & x96;
  assign n4306 = ~n3865 & n4305;
  assign n4307 = n4083 & ~n4306;
  assign n4308 = ~n4304 & n4307;
  assign n4309 = ~n3868 & ~n4308;
  assign n4310 = ~n242 & ~n4309;
  assign n4311 = ~x97 & ~n4310;
  assign n4312 = ~x96 & n4089;
  assign n4313 = ~n4311 & ~n4312;
  assign n4314 = ~n4302 & n4313;
  assign n4315 = x97 & n3868;
  assign n4316 = ~x98 & n4082;
  assign n4317 = ~n4315 & n4316;
  assign n4318 = ~n4314 & n4317;
  assign n4319 = ~x29 & ~x30;
  assign n4320 = ~n4318 & n4319;
  assign n4321 = ~x29 & x65;
  assign n4322 = ~n4320 & ~n4321;
  assign n4323 = x64 & ~n4322;
  assign n4324 = x64 & n4318;
  assign n4325 = x29 & ~x65;
  assign n4326 = x30 & ~n4325;
  assign n4327 = n4326 ^ n4113;
  assign n4328 = n4324 & n4327;
  assign n4329 = n4328 ^ n4113;
  assign n4330 = ~n4323 & ~n4329;
  assign n4331 = n4330 ^ x66;
  assign n4332 = x65 & n4086;
  assign n4333 = x30 & ~n4332;
  assign n4334 = n4318 & ~n4333;
  assign n4335 = n4105 & ~n4334;
  assign n4336 = n293 & ~n4086;
  assign n4337 = n4336 ^ x65;
  assign n4338 = ~x30 & n4337;
  assign n4339 = ~n202 & ~n4338;
  assign n4340 = x65 & n4333;
  assign n4341 = n4339 & ~n4340;
  assign n4342 = n4318 & ~n4341;
  assign n4343 = ~n4335 & ~n4342;
  assign n4344 = n4343 ^ x31;
  assign n4345 = n4344 ^ n4330;
  assign n4346 = ~n4331 & n4345;
  assign n4347 = n4346 ^ x66;
  assign n4348 = ~x67 & ~n4347;
  assign n4349 = x67 & ~n4330;
  assign n4350 = ~x66 & ~n4344;
  assign n4351 = n4349 & ~n4350;
  assign n4352 = n1724 & n4344;
  assign n4353 = n4118 ^ x66;
  assign n4354 = n4318 & ~n4353;
  assign n4355 = n4354 ^ n4103;
  assign n4356 = ~n4352 & ~n4355;
  assign n4357 = ~n4351 & n4356;
  assign n4358 = ~n4348 & ~n4357;
  assign n4359 = n4122 & n4318;
  assign n4360 = n4359 ^ n4125;
  assign n4361 = ~x68 & ~n4360;
  assign n4362 = n4358 & ~n4361;
  assign n4363 = n4129 & n4318;
  assign n4364 = n4363 ^ n4131;
  assign n4365 = x69 & n4364;
  assign n4366 = x68 & n4360;
  assign n4367 = ~n4365 & ~n4366;
  assign n4368 = ~n4362 & n4367;
  assign n4369 = ~x69 & ~n4364;
  assign n4370 = ~n4368 & ~n4369;
  assign n4371 = n4370 ^ x70;
  assign n4372 = n4135 & n4318;
  assign n4373 = n4372 ^ n4137;
  assign n4374 = n4373 ^ n4370;
  assign n4375 = n4371 & ~n4374;
  assign n4376 = n4375 ^ x70;
  assign n4377 = n4376 ^ x71;
  assign n4378 = n4141 & n4318;
  assign n4379 = n4378 ^ n4143;
  assign n4380 = n4379 ^ n4376;
  assign n4381 = n4377 & ~n4380;
  assign n4382 = n4381 ^ x71;
  assign n4383 = n4382 ^ x72;
  assign n4384 = n4147 & n4318;
  assign n4385 = n4384 ^ n4149;
  assign n4386 = n4385 ^ n4382;
  assign n4387 = n4383 & ~n4386;
  assign n4388 = n4387 ^ x72;
  assign n4389 = n4388 ^ x73;
  assign n4390 = n4153 & n4318;
  assign n4391 = n4390 ^ n4155;
  assign n4392 = n4391 ^ n4388;
  assign n4393 = n4389 & ~n4392;
  assign n4394 = n4393 ^ x73;
  assign n4395 = n4394 ^ x74;
  assign n4396 = n4159 & n4318;
  assign n4397 = n4396 ^ n4161;
  assign n4398 = n4397 ^ n4394;
  assign n4399 = n4395 & ~n4398;
  assign n4400 = n4399 ^ x74;
  assign n4401 = n4400 ^ x75;
  assign n4402 = n4165 & n4318;
  assign n4403 = n4402 ^ n4167;
  assign n4404 = n4403 ^ n4400;
  assign n4405 = n4401 & ~n4404;
  assign n4406 = n4405 ^ x75;
  assign n4407 = n4406 ^ x76;
  assign n4408 = n4171 & n4318;
  assign n4409 = n4408 ^ n4173;
  assign n4410 = n4409 ^ n4406;
  assign n4411 = n4407 & ~n4410;
  assign n4412 = n4411 ^ x76;
  assign n4413 = n4412 ^ x77;
  assign n4414 = n4177 & n4318;
  assign n4415 = n4414 ^ n4179;
  assign n4416 = n4415 ^ n4412;
  assign n4417 = n4413 & ~n4416;
  assign n4418 = n4417 ^ x77;
  assign n4419 = n4418 ^ x78;
  assign n4420 = n4183 & n4318;
  assign n4421 = n4420 ^ n4185;
  assign n4422 = n4421 ^ n4418;
  assign n4423 = n4419 & ~n4422;
  assign n4424 = n4423 ^ x78;
  assign n4425 = n4424 ^ x79;
  assign n4426 = n4189 & n4318;
  assign n4427 = n4426 ^ n4191;
  assign n4428 = n4427 ^ n4424;
  assign n4429 = n4425 & ~n4428;
  assign n4430 = n4429 ^ x79;
  assign n4431 = n4430 ^ x80;
  assign n4432 = n4195 & n4318;
  assign n4433 = n4432 ^ n4197;
  assign n4434 = n4433 ^ n4430;
  assign n4435 = n4431 & ~n4434;
  assign n4436 = n4435 ^ x80;
  assign n4437 = n4436 ^ x81;
  assign n4438 = n4201 & n4318;
  assign n4439 = n4438 ^ n4204;
  assign n4440 = n4439 ^ n4436;
  assign n4441 = n4437 & ~n4440;
  assign n4442 = n4441 ^ x81;
  assign n4443 = n4442 ^ x82;
  assign n4444 = n4208 & n4318;
  assign n4445 = n4444 ^ n4214;
  assign n4446 = n4445 ^ n4442;
  assign n4447 = n4443 & ~n4446;
  assign n4448 = n4447 ^ x82;
  assign n4449 = n4448 ^ x83;
  assign n4450 = n4218 & n4318;
  assign n4451 = n4450 ^ n4220;
  assign n4452 = n4451 ^ n4448;
  assign n4453 = n4449 & ~n4452;
  assign n4454 = n4453 ^ x83;
  assign n4455 = n4454 ^ x84;
  assign n4456 = n4224 & n4318;
  assign n4457 = n4456 ^ n4226;
  assign n4458 = n4457 ^ n4454;
  assign n4459 = n4455 & ~n4458;
  assign n4460 = n4459 ^ x84;
  assign n4461 = n4460 ^ x85;
  assign n4462 = n4230 & n4318;
  assign n4463 = n4462 ^ n4232;
  assign n4464 = n4463 ^ n4460;
  assign n4465 = n4461 & ~n4464;
  assign n4466 = n4465 ^ x85;
  assign n4467 = n4466 ^ x86;
  assign n4468 = n4236 & n4318;
  assign n4469 = n4468 ^ n4238;
  assign n4470 = n4469 ^ n4466;
  assign n4471 = n4467 & ~n4470;
  assign n4472 = n4471 ^ x86;
  assign n4473 = n4472 ^ x87;
  assign n4474 = n4242 & n4318;
  assign n4475 = n4474 ^ n4244;
  assign n4476 = n4475 ^ n4472;
  assign n4477 = n4473 & ~n4476;
  assign n4478 = n4477 ^ x87;
  assign n4479 = n4478 ^ x88;
  assign n4480 = n4248 & n4318;
  assign n4481 = n4480 ^ n4250;
  assign n4482 = n4481 ^ n4478;
  assign n4483 = n4479 & ~n4482;
  assign n4484 = n4483 ^ x88;
  assign n4485 = n4484 ^ x89;
  assign n4486 = n4254 & n4318;
  assign n4487 = n4486 ^ n4256;
  assign n4488 = n4487 ^ n4484;
  assign n4489 = n4485 & ~n4488;
  assign n4490 = n4489 ^ x89;
  assign n4491 = n4490 ^ x90;
  assign n4492 = n4260 & n4318;
  assign n4493 = n4492 ^ n4262;
  assign n4494 = n4493 ^ n4490;
  assign n4495 = n4491 & ~n4494;
  assign n4496 = n4495 ^ x90;
  assign n4497 = n4496 ^ x91;
  assign n4498 = n4266 & n4318;
  assign n4499 = n4498 ^ n4268;
  assign n4500 = n4499 ^ n4496;
  assign n4501 = n4497 & ~n4500;
  assign n4502 = n4501 ^ x91;
  assign n4503 = n4502 ^ x92;
  assign n4504 = n4272 & n4318;
  assign n4505 = n4504 ^ n4274;
  assign n4506 = n4505 ^ n4502;
  assign n4507 = n4503 & ~n4506;
  assign n4508 = n4507 ^ x92;
  assign n4509 = n4508 ^ x93;
  assign n4510 = n4278 & n4318;
  assign n4511 = n4510 ^ n4280;
  assign n4512 = n4511 ^ n4508;
  assign n4513 = n4509 & ~n4512;
  assign n4514 = n4513 ^ x93;
  assign n4515 = n4514 ^ x94;
  assign n4516 = n4284 & n4318;
  assign n4517 = n4516 ^ n4286;
  assign n4518 = n4517 ^ n4514;
  assign n4519 = n4515 & ~n4518;
  assign n4520 = n4519 ^ x94;
  assign n4521 = n4520 ^ x95;
  assign n4522 = n4290 & n4318;
  assign n4523 = n4522 ^ n4292;
  assign n4524 = n4523 ^ n4520;
  assign n4525 = n4521 & ~n4524;
  assign n4526 = n4525 ^ x95;
  assign n4527 = n4526 ^ x96;
  assign n4528 = n4296 & n4318;
  assign n4529 = n4528 ^ n4298;
  assign n4530 = n4529 ^ n4526;
  assign n4531 = n4527 & ~n4530;
  assign n4532 = n4531 ^ x96;
  assign n4533 = x97 & n4532;
  assign n4534 = n4301 ^ x96;
  assign n4535 = n4318 & n4534;
  assign n4536 = n4535 ^ n4089;
  assign n4537 = ~n4533 & n4536;
  assign n4538 = ~x97 & ~n4532;
  assign n4539 = ~n242 & ~n4314;
  assign n4540 = ~x98 & ~n4310;
  assign n4541 = ~n4539 & n4540;
  assign n4542 = ~n4538 & ~n4541;
  assign n4543 = ~n4537 & n4542;
  assign n4544 = x98 & n4310;
  assign n4545 = n4082 & ~n4544;
  assign n4546 = ~n4543 & n4545;
  assign n4547 = n4527 & n4546;
  assign n4548 = n4547 ^ n4529;
  assign n4549 = ~x97 & ~n4548;
  assign n4550 = n4532 ^ x97;
  assign n4551 = n4546 & n4550;
  assign n4552 = n4551 ^ n4536;
  assign n4553 = ~x98 & n4552;
  assign n4554 = ~n4549 & ~n4553;
  assign n4555 = n4503 & n4546;
  assign n4556 = n4555 ^ n4505;
  assign n4557 = ~x93 & ~n4556;
  assign n4558 = n4509 & n4546;
  assign n4559 = n4558 ^ n4511;
  assign n4560 = ~x94 & ~n4559;
  assign n4561 = ~n4557 & ~n4560;
  assign n4562 = n4358 ^ x68;
  assign n4563 = n4546 & n4562;
  assign n4564 = n4563 ^ n4360;
  assign n4565 = ~x69 & ~n4564;
  assign n4566 = ~n4362 & ~n4366;
  assign n4567 = n4566 ^ x69;
  assign n4568 = n4546 & ~n4567;
  assign n4569 = n4568 ^ n4364;
  assign n4570 = ~x70 & ~n4569;
  assign n4571 = ~n4565 & ~n4570;
  assign n4572 = ~x29 & n4546;
  assign n4573 = ~x28 & ~n4572;
  assign n4574 = ~x65 & ~n4573;
  assign n4575 = ~x28 & ~n4325;
  assign n4576 = ~n4546 & ~n4575;
  assign n4577 = x28 & ~x29;
  assign n4578 = x64 & ~n4577;
  assign n4579 = ~n4576 & n4578;
  assign n4580 = ~n4574 & n4579;
  assign n4581 = x64 & n4546;
  assign n4582 = n4321 & ~n4581;
  assign n4583 = ~n4580 & ~n4582;
  assign n4584 = n4583 ^ x66;
  assign n4585 = x65 & n4546;
  assign n4586 = ~n4324 & ~n4585;
  assign n4587 = x65 & n4318;
  assign n4588 = x29 & ~n4587;
  assign n4589 = n4581 & ~n4588;
  assign n4590 = ~n4586 & ~n4589;
  assign n4591 = n293 & ~n4318;
  assign n4592 = n4591 ^ x65;
  assign n4593 = n4572 & n4592;
  assign n4594 = ~n4590 & ~n4593;
  assign n4595 = n4594 ^ x30;
  assign n4596 = n4595 ^ n4583;
  assign n4597 = ~n4584 & n4596;
  assign n4598 = n4597 ^ x66;
  assign n4599 = n4598 ^ x67;
  assign n4600 = ~n4331 & n4546;
  assign n4601 = n4600 ^ n4344;
  assign n4602 = n4601 ^ n4598;
  assign n4603 = n4599 & ~n4602;
  assign n4604 = n4603 ^ x67;
  assign n4605 = n4604 ^ x68;
  assign n4606 = n4347 ^ x67;
  assign n4607 = n4546 & n4606;
  assign n4608 = n4607 ^ n4355;
  assign n4609 = n4608 ^ n4604;
  assign n4610 = n4605 & ~n4609;
  assign n4611 = n4610 ^ x68;
  assign n4612 = n4571 & n4611;
  assign n4613 = n4569 ^ x70;
  assign n4614 = x69 & n4564;
  assign n4615 = n4614 ^ n4569;
  assign n4616 = n4613 & ~n4615;
  assign n4617 = n4616 ^ x70;
  assign n4618 = ~n4612 & ~n4617;
  assign n4619 = n4618 ^ x71;
  assign n4620 = n4371 & n4546;
  assign n4621 = n4620 ^ n4373;
  assign n4622 = n4621 ^ n4618;
  assign n4623 = ~n4619 & n4622;
  assign n4624 = n4623 ^ x71;
  assign n4625 = n4624 ^ x72;
  assign n4626 = n4377 & n4546;
  assign n4627 = n4626 ^ n4379;
  assign n4628 = n4627 ^ n4624;
  assign n4629 = n4625 & ~n4628;
  assign n4630 = n4629 ^ x72;
  assign n4631 = n4630 ^ x73;
  assign n4632 = n4383 & n4546;
  assign n4633 = n4632 ^ n4385;
  assign n4634 = n4633 ^ n4630;
  assign n4635 = n4631 & ~n4634;
  assign n4636 = n4635 ^ x73;
  assign n4637 = n4636 ^ x74;
  assign n4638 = n4389 & n4546;
  assign n4639 = n4638 ^ n4391;
  assign n4640 = n4639 ^ n4636;
  assign n4641 = n4637 & ~n4640;
  assign n4642 = n4641 ^ x74;
  assign n4643 = n4642 ^ x75;
  assign n4644 = n4395 & n4546;
  assign n4645 = n4644 ^ n4397;
  assign n4646 = n4645 ^ n4642;
  assign n4647 = n4643 & ~n4646;
  assign n4648 = n4647 ^ x75;
  assign n4649 = n4648 ^ x76;
  assign n4650 = n4401 & n4546;
  assign n4651 = n4650 ^ n4403;
  assign n4652 = n4651 ^ n4648;
  assign n4653 = n4649 & ~n4652;
  assign n4654 = n4653 ^ x76;
  assign n4655 = n4654 ^ x77;
  assign n4656 = n4407 & n4546;
  assign n4657 = n4656 ^ n4409;
  assign n4658 = n4657 ^ n4654;
  assign n4659 = n4655 & ~n4658;
  assign n4660 = n4659 ^ x77;
  assign n4661 = n4660 ^ x78;
  assign n4662 = n4413 & n4546;
  assign n4663 = n4662 ^ n4415;
  assign n4664 = n4663 ^ n4660;
  assign n4665 = n4661 & ~n4664;
  assign n4666 = n4665 ^ x78;
  assign n4667 = n4666 ^ x79;
  assign n4668 = n4419 & n4546;
  assign n4669 = n4668 ^ n4421;
  assign n4670 = n4669 ^ n4666;
  assign n4671 = n4667 & ~n4670;
  assign n4672 = n4671 ^ x79;
  assign n4673 = n4672 ^ x80;
  assign n4674 = n4425 & n4546;
  assign n4675 = n4674 ^ n4427;
  assign n4676 = n4675 ^ n4672;
  assign n4677 = n4673 & ~n4676;
  assign n4678 = n4677 ^ x80;
  assign n4679 = n4678 ^ x81;
  assign n4680 = n4431 & n4546;
  assign n4681 = n4680 ^ n4433;
  assign n4682 = n4681 ^ n4678;
  assign n4683 = n4679 & ~n4682;
  assign n4684 = n4683 ^ x81;
  assign n4685 = n4684 ^ x82;
  assign n4686 = n4437 & n4546;
  assign n4687 = n4686 ^ n4439;
  assign n4688 = n4687 ^ n4684;
  assign n4689 = n4685 & ~n4688;
  assign n4690 = n4689 ^ x82;
  assign n4691 = n4690 ^ x83;
  assign n4692 = n4443 & n4546;
  assign n4693 = n4692 ^ n4445;
  assign n4694 = n4693 ^ n4690;
  assign n4695 = n4691 & ~n4694;
  assign n4696 = n4695 ^ x83;
  assign n4697 = n4696 ^ x84;
  assign n4698 = n4449 & n4546;
  assign n4699 = n4698 ^ n4451;
  assign n4700 = n4699 ^ n4696;
  assign n4701 = n4697 & ~n4700;
  assign n4702 = n4701 ^ x84;
  assign n4703 = n4702 ^ x85;
  assign n4704 = n4455 & n4546;
  assign n4705 = n4704 ^ n4457;
  assign n4706 = n4705 ^ n4702;
  assign n4707 = n4703 & ~n4706;
  assign n4708 = n4707 ^ x85;
  assign n4709 = n4708 ^ x86;
  assign n4710 = n4461 & n4546;
  assign n4711 = n4710 ^ n4463;
  assign n4712 = n4711 ^ n4708;
  assign n4713 = n4709 & ~n4712;
  assign n4714 = n4713 ^ x86;
  assign n4715 = n4714 ^ x87;
  assign n4716 = n4467 & n4546;
  assign n4717 = n4716 ^ n4469;
  assign n4718 = n4717 ^ n4714;
  assign n4719 = n4715 & ~n4718;
  assign n4720 = n4719 ^ x87;
  assign n4721 = n4720 ^ x88;
  assign n4722 = n4473 & n4546;
  assign n4723 = n4722 ^ n4475;
  assign n4724 = n4723 ^ n4720;
  assign n4725 = n4721 & ~n4724;
  assign n4726 = n4725 ^ x88;
  assign n4727 = n4726 ^ x89;
  assign n4728 = n4479 & n4546;
  assign n4729 = n4728 ^ n4481;
  assign n4730 = n4729 ^ n4726;
  assign n4731 = n4727 & ~n4730;
  assign n4732 = n4731 ^ x89;
  assign n4733 = n4732 ^ x90;
  assign n4734 = n4485 & n4546;
  assign n4735 = n4734 ^ n4487;
  assign n4736 = n4735 ^ n4732;
  assign n4737 = n4733 & ~n4736;
  assign n4738 = n4737 ^ x90;
  assign n4739 = n4738 ^ x91;
  assign n4740 = n4491 & n4546;
  assign n4741 = n4740 ^ n4493;
  assign n4742 = n4741 ^ n4738;
  assign n4743 = n4739 & ~n4742;
  assign n4744 = n4743 ^ x91;
  assign n4745 = n4744 ^ x92;
  assign n4746 = n4497 & n4546;
  assign n4747 = n4746 ^ n4499;
  assign n4748 = n4747 ^ n4744;
  assign n4749 = n4745 & ~n4748;
  assign n4750 = n4749 ^ x92;
  assign n4751 = n4561 & n4750;
  assign n4752 = n4559 ^ x94;
  assign n4753 = x93 & n4556;
  assign n4754 = n4753 ^ n4559;
  assign n4755 = n4752 & ~n4754;
  assign n4756 = n4755 ^ x94;
  assign n4757 = ~n4751 & ~n4756;
  assign n4758 = n4757 ^ x95;
  assign n4759 = n4515 & n4546;
  assign n4760 = n4759 ^ n4517;
  assign n4761 = n4760 ^ n4757;
  assign n4762 = ~n4758 & n4761;
  assign n4763 = n4762 ^ x95;
  assign n4764 = n4763 ^ x96;
  assign n4765 = n4521 & n4546;
  assign n4766 = n4765 ^ n4523;
  assign n4767 = n4766 ^ n4763;
  assign n4768 = n4764 & ~n4767;
  assign n4769 = n4768 ^ x96;
  assign n4770 = n4554 & n4769;
  assign n4771 = n4552 ^ x98;
  assign n4772 = x97 & n4548;
  assign n4773 = n4772 ^ n4552;
  assign n4774 = ~n4771 & n4773;
  assign n4775 = n4774 ^ x98;
  assign n4776 = ~n4770 & ~n4775;
  assign n4777 = x99 & ~n4776;
  assign n4778 = ~x100 & n155;
  assign n4779 = ~n4777 & n4778;
  assign n4780 = n4309 & ~n4318;
  assign n4781 = ~n4546 & n4780;
  assign n4782 = ~n242 & ~n4781;
  assign n4783 = ~n4779 & ~n4782;
  assign n4784 = ~x99 & n4776;
  assign n4785 = n4782 & ~n4784;
  assign n4786 = n4779 & ~n4785;
  assign n4787 = n4769 ^ x97;
  assign n4788 = n4769 ^ n4548;
  assign n4789 = n4787 & ~n4788;
  assign n4790 = n4789 ^ x97;
  assign n4791 = n4790 ^ x98;
  assign n4792 = n4786 & n4791;
  assign n4793 = n4792 ^ n4552;
  assign n4794 = ~x99 & n4793;
  assign n4795 = n4739 & n4786;
  assign n4796 = n4795 ^ n4741;
  assign n4797 = ~x92 & ~n4796;
  assign n4798 = n4745 & n4786;
  assign n4799 = n4798 ^ n4747;
  assign n4800 = ~x93 & ~n4799;
  assign n4801 = ~n4797 & ~n4800;
  assign n4802 = n4709 & n4786;
  assign n4803 = n4802 ^ n4711;
  assign n4804 = ~x87 & ~n4803;
  assign n4805 = n4715 & n4786;
  assign n4806 = n4805 ^ n4717;
  assign n4807 = ~x88 & ~n4806;
  assign n4808 = ~n4804 & ~n4807;
  assign n4809 = n4679 & n4786;
  assign n4810 = n4809 ^ n4681;
  assign n4811 = ~x82 & ~n4810;
  assign n4812 = n4673 & n4786;
  assign n4813 = n4812 ^ n4675;
  assign n4814 = ~x81 & ~n4813;
  assign n4815 = ~n4811 & ~n4814;
  assign n4816 = n4649 & n4786;
  assign n4817 = n4816 ^ n4651;
  assign n4818 = ~x77 & ~n4817;
  assign n4819 = x28 & ~n4585;
  assign n4820 = n4786 & ~n4819;
  assign n4821 = n4581 & ~n4820;
  assign n4822 = n293 & ~n4546;
  assign n4823 = n4822 ^ x65;
  assign n4824 = ~x28 & n4823;
  assign n4825 = ~n202 & ~n4824;
  assign n4826 = x65 & n4819;
  assign n4827 = n4825 & ~n4826;
  assign n4828 = n4786 & ~n4827;
  assign n4829 = ~n4821 & ~n4828;
  assign n4830 = n4829 ^ x29;
  assign n4831 = n4830 ^ x66;
  assign n4832 = x64 & n4786;
  assign n4833 = x27 & ~x65;
  assign n4834 = x28 & ~n4833;
  assign n4835 = n4832 & n4834;
  assign n4836 = ~x27 & x64;
  assign n4837 = ~x65 & ~n4836;
  assign n4838 = ~x28 & ~n4837;
  assign n4839 = ~n4786 & n4838;
  assign n4840 = x28 ^ x27;
  assign n4841 = ~x64 & n4840;
  assign n4842 = n4841 ^ x27;
  assign n4843 = x65 & ~n4842;
  assign n4844 = ~n4839 & ~n4843;
  assign n4845 = ~n4835 & n4844;
  assign n4846 = n4845 ^ n4830;
  assign n4847 = n4831 & n4846;
  assign n4848 = n4847 ^ x66;
  assign n4849 = n4848 ^ x67;
  assign n4850 = ~n4584 & n4786;
  assign n4851 = n4850 ^ n4595;
  assign n4852 = n4851 ^ n4848;
  assign n4853 = n4849 & ~n4852;
  assign n4854 = n4853 ^ x67;
  assign n4855 = n4854 ^ x68;
  assign n4856 = n4599 & n4786;
  assign n4857 = n4856 ^ n4601;
  assign n4858 = n4857 ^ n4854;
  assign n4859 = n4855 & ~n4858;
  assign n4860 = n4859 ^ x68;
  assign n4861 = n4860 ^ x69;
  assign n4862 = n4605 & n4786;
  assign n4863 = n4862 ^ n4608;
  assign n4864 = n4863 ^ n4860;
  assign n4865 = n4861 & ~n4864;
  assign n4866 = n4865 ^ x69;
  assign n4867 = n4866 ^ x70;
  assign n4868 = n4611 ^ x69;
  assign n4869 = n4786 & n4868;
  assign n4870 = n4869 ^ n4564;
  assign n4871 = n4870 ^ n4866;
  assign n4872 = n4867 & ~n4871;
  assign n4873 = n4872 ^ x70;
  assign n4874 = n4873 ^ x71;
  assign n4875 = n4611 ^ n4564;
  assign n4876 = n4868 & ~n4875;
  assign n4877 = n4876 ^ x69;
  assign n4878 = n4877 ^ x70;
  assign n4879 = n4786 & n4878;
  assign n4880 = n4879 ^ n4569;
  assign n4881 = n4880 ^ n4873;
  assign n4882 = n4874 & ~n4881;
  assign n4883 = n4882 ^ x71;
  assign n4884 = n4883 ^ x72;
  assign n4885 = ~n4619 & n4786;
  assign n4886 = n4885 ^ n4621;
  assign n4887 = n4886 ^ n4883;
  assign n4888 = n4884 & ~n4887;
  assign n4889 = n4888 ^ x72;
  assign n4890 = n4889 ^ x73;
  assign n4891 = n4625 & n4786;
  assign n4892 = n4891 ^ n4627;
  assign n4893 = n4892 ^ n4889;
  assign n4894 = n4890 & ~n4893;
  assign n4895 = n4894 ^ x73;
  assign n4896 = n4895 ^ x74;
  assign n4897 = n4631 & n4786;
  assign n4898 = n4897 ^ n4633;
  assign n4899 = n4898 ^ n4895;
  assign n4900 = n4896 & ~n4899;
  assign n4901 = n4900 ^ x74;
  assign n4902 = n4901 ^ x75;
  assign n4903 = n4637 & n4786;
  assign n4904 = n4903 ^ n4639;
  assign n4905 = n4904 ^ n4901;
  assign n4906 = n4902 & ~n4905;
  assign n4907 = n4906 ^ x75;
  assign n4908 = n4907 ^ x76;
  assign n4909 = n4643 & n4786;
  assign n4910 = n4909 ^ n4645;
  assign n4911 = n4910 ^ n4907;
  assign n4912 = n4908 & ~n4911;
  assign n4913 = n4912 ^ x76;
  assign n4914 = ~n4818 & n4913;
  assign n4915 = n4655 & n4786;
  assign n4916 = n4915 ^ n4657;
  assign n4917 = x78 & n4916;
  assign n4918 = x77 & n4817;
  assign n4919 = ~n4917 & ~n4918;
  assign n4920 = ~n4914 & n4919;
  assign n4921 = ~x78 & ~n4916;
  assign n4922 = ~n4920 & ~n4921;
  assign n4923 = n4922 ^ x79;
  assign n4924 = n4663 ^ x78;
  assign n4925 = n4924 ^ n4660;
  assign n4926 = n4925 ^ n4663;
  assign n4927 = n4786 & n4926;
  assign n4928 = n4927 ^ n4663;
  assign n4929 = n4928 ^ n4922;
  assign n4930 = n4923 & ~n4929;
  assign n4931 = n4930 ^ x79;
  assign n4932 = n4931 ^ x80;
  assign n4933 = n4667 & n4786;
  assign n4934 = n4933 ^ n4669;
  assign n4935 = n4934 ^ n4931;
  assign n4936 = n4932 & ~n4935;
  assign n4937 = n4936 ^ x80;
  assign n4938 = n4815 & n4937;
  assign n4939 = n4810 ^ x82;
  assign n4940 = x81 & n4813;
  assign n4941 = n4940 ^ n4810;
  assign n4942 = n4939 & ~n4941;
  assign n4943 = n4942 ^ x82;
  assign n4944 = ~n4938 & ~n4943;
  assign n4945 = n4685 & n4786;
  assign n4946 = n4945 ^ n4687;
  assign n4947 = ~x83 & ~n4946;
  assign n4948 = n4691 & n4786;
  assign n4949 = n4948 ^ n4693;
  assign n4950 = ~x84 & ~n4949;
  assign n4951 = ~n4947 & ~n4950;
  assign n4952 = ~n4944 & n4951;
  assign n4953 = n4949 ^ x84;
  assign n4954 = x83 & n4946;
  assign n4955 = n4954 ^ n4949;
  assign n4956 = n4953 & ~n4955;
  assign n4957 = n4956 ^ x84;
  assign n4958 = ~n4952 & ~n4957;
  assign n4959 = n4958 ^ x85;
  assign n4960 = n4697 & n4786;
  assign n4961 = n4960 ^ n4699;
  assign n4962 = n4961 ^ n4958;
  assign n4963 = ~n4959 & n4962;
  assign n4964 = n4963 ^ x85;
  assign n4965 = n4964 ^ x86;
  assign n4966 = n4703 & n4786;
  assign n4967 = n4966 ^ n4705;
  assign n4968 = n4967 ^ n4964;
  assign n4969 = n4965 & ~n4968;
  assign n4970 = n4969 ^ x86;
  assign n4971 = n4808 & n4970;
  assign n4972 = n4806 ^ x88;
  assign n4973 = x87 & n4803;
  assign n4974 = n4973 ^ n4806;
  assign n4975 = n4972 & ~n4974;
  assign n4976 = n4975 ^ x88;
  assign n4977 = ~n4971 & ~n4976;
  assign n4978 = n4977 ^ x89;
  assign n4979 = n4721 & n4786;
  assign n4980 = n4979 ^ n4723;
  assign n4981 = n4980 ^ n4977;
  assign n4982 = ~n4978 & n4981;
  assign n4983 = n4982 ^ x89;
  assign n4984 = n4983 ^ x90;
  assign n4985 = n4727 & n4786;
  assign n4986 = n4985 ^ n4729;
  assign n4987 = n4986 ^ n4983;
  assign n4988 = n4984 & ~n4987;
  assign n4989 = n4988 ^ x90;
  assign n4990 = n4989 ^ x91;
  assign n4991 = n4733 & n4786;
  assign n4992 = n4991 ^ n4735;
  assign n4993 = n4992 ^ n4989;
  assign n4994 = n4990 & ~n4993;
  assign n4995 = n4994 ^ x91;
  assign n4996 = n4801 & n4995;
  assign n4997 = n4799 ^ x93;
  assign n4998 = x92 & n4796;
  assign n4999 = n4998 ^ n4799;
  assign n5000 = n4997 & ~n4999;
  assign n5001 = n5000 ^ x93;
  assign n5002 = ~n4996 & ~n5001;
  assign n5003 = n5002 ^ x94;
  assign n5004 = n4750 ^ x93;
  assign n5005 = n4786 & n5004;
  assign n5006 = n5005 ^ n4556;
  assign n5007 = n5006 ^ n5002;
  assign n5008 = ~n5003 & n5007;
  assign n5009 = n5008 ^ x94;
  assign n5010 = n5009 ^ x95;
  assign n5011 = n4750 ^ n4556;
  assign n5012 = n5004 & ~n5011;
  assign n5013 = n5012 ^ x93;
  assign n5014 = n5013 ^ x94;
  assign n5015 = n4786 & n5014;
  assign n5016 = n5015 ^ n4559;
  assign n5017 = n5016 ^ n5009;
  assign n5018 = n5010 & ~n5017;
  assign n5019 = n5018 ^ x95;
  assign n5020 = n5019 ^ x96;
  assign n5021 = ~n4758 & n4786;
  assign n5022 = n5021 ^ n4760;
  assign n5023 = n5022 ^ n5019;
  assign n5024 = n5020 & ~n5023;
  assign n5025 = n5024 ^ x96;
  assign n5026 = n5025 ^ x97;
  assign n5027 = n4764 & n4786;
  assign n5028 = n5027 ^ n4766;
  assign n5029 = n5028 ^ n5025;
  assign n5030 = n5026 & ~n5029;
  assign n5031 = n5030 ^ x97;
  assign n5032 = n5031 ^ x98;
  assign n5033 = n4786 & n4787;
  assign n5034 = n5033 ^ n4548;
  assign n5035 = n5034 ^ n5031;
  assign n5036 = n5032 & ~n5035;
  assign n5037 = n5036 ^ x98;
  assign n5038 = ~n4794 & n5037;
  assign n5039 = x99 & ~n4793;
  assign n5040 = ~n242 & ~n4783;
  assign n5041 = x100 & n5040;
  assign n5042 = n155 & ~n5041;
  assign n5043 = ~n5039 & n5042;
  assign n5044 = ~n5038 & n5043;
  assign n5045 = n4778 & ~n5040;
  assign n5046 = ~n5044 & ~n5045;
  assign n5047 = n4783 & n5046;
  assign n5048 = ~n242 & ~n5047;
  assign n5049 = ~x101 & ~n5048;
  assign n5050 = n5037 ^ x99;
  assign n5051 = ~n5046 & n5050;
  assign n5052 = n5051 ^ n4793;
  assign n5053 = ~n5049 & ~n5052;
  assign n5054 = x100 & x101;
  assign n5055 = ~n5053 & ~n5054;
  assign n5056 = n5020 & ~n5046;
  assign n5057 = n5056 ^ n5022;
  assign n5058 = ~x97 & ~n5057;
  assign n5059 = n5010 & ~n5046;
  assign n5060 = n5059 ^ n5016;
  assign n5061 = ~x96 & ~n5060;
  assign n5062 = ~n5058 & ~n5061;
  assign n5063 = n4995 ^ x92;
  assign n5064 = ~n5046 & n5063;
  assign n5065 = n5064 ^ n4796;
  assign n5066 = x93 & n5065;
  assign n5067 = n4970 ^ x87;
  assign n5068 = n4970 ^ n4803;
  assign n5069 = n5067 & ~n5068;
  assign n5070 = n5069 ^ x87;
  assign n5071 = n5070 ^ x88;
  assign n5072 = ~n5046 & n5071;
  assign n5073 = n5072 ^ n4806;
  assign n5074 = ~x89 & ~n5073;
  assign n5075 = ~n4978 & ~n5046;
  assign n5076 = n5075 ^ n4980;
  assign n5077 = ~x90 & ~n5076;
  assign n5078 = ~n5074 & ~n5077;
  assign n5079 = n4908 & ~n5046;
  assign n5080 = n5079 ^ n4910;
  assign n5081 = ~x77 & ~n5080;
  assign n5082 = n4913 ^ x77;
  assign n5083 = ~n5046 & n5082;
  assign n5084 = n5083 ^ n4817;
  assign n5085 = ~x78 & ~n5084;
  assign n5086 = ~n5081 & ~n5085;
  assign n5087 = x65 & n4786;
  assign n5088 = x27 & ~n5087;
  assign n5089 = ~n5046 & ~n5088;
  assign n5090 = n4832 & ~n5089;
  assign n5091 = n4786 ^ x65;
  assign n5092 = n4836 & ~n5091;
  assign n5093 = ~n202 & ~n5092;
  assign n5094 = x65 & n5088;
  assign n5095 = n5093 & ~n5094;
  assign n5096 = ~n5046 & ~n5095;
  assign n5097 = ~n5090 & ~n5096;
  assign n5098 = n5097 ^ x28;
  assign n5099 = n5098 ^ x66;
  assign n5100 = x64 & ~n5046;
  assign n5101 = x26 & n4833;
  assign n5102 = n5101 ^ x27;
  assign n5103 = n5100 & n5102;
  assign n5104 = ~x26 & n4836;
  assign n5105 = ~x27 & x65;
  assign n5106 = ~n5104 & ~n5105;
  assign n5107 = n5046 & ~n5106;
  assign n5108 = ~x26 & x65;
  assign n5109 = n5108 ^ n5105;
  assign n5110 = x64 & n5109;
  assign n5111 = n5110 ^ n5105;
  assign n5112 = ~n5107 & ~n5111;
  assign n5113 = ~n5103 & n5112;
  assign n5114 = n5113 ^ n5098;
  assign n5115 = n5099 & n5114;
  assign n5116 = n5115 ^ x66;
  assign n5117 = n5116 ^ x67;
  assign n5118 = n4845 ^ x66;
  assign n5119 = ~n5046 & ~n5118;
  assign n5120 = n5119 ^ n4830;
  assign n5121 = n5120 ^ n5116;
  assign n5122 = n5117 & ~n5121;
  assign n5123 = n5122 ^ x67;
  assign n5124 = n5123 ^ x68;
  assign n5125 = n4849 & ~n5046;
  assign n5126 = n5125 ^ n4851;
  assign n5127 = n5126 ^ n5123;
  assign n5128 = n5124 & ~n5127;
  assign n5129 = n5128 ^ x68;
  assign n5130 = n5129 ^ x69;
  assign n5131 = n4855 & ~n5046;
  assign n5132 = n5131 ^ n4857;
  assign n5133 = n5132 ^ n5129;
  assign n5134 = n5130 & ~n5133;
  assign n5135 = n5134 ^ x69;
  assign n5136 = n5135 ^ x70;
  assign n5137 = n4861 & ~n5046;
  assign n5138 = n5137 ^ n4863;
  assign n5139 = n5138 ^ n5135;
  assign n5140 = n5136 & ~n5139;
  assign n5141 = n5140 ^ x70;
  assign n5142 = n5141 ^ x71;
  assign n5143 = n4867 & ~n5046;
  assign n5144 = n5143 ^ n4870;
  assign n5145 = n5144 ^ n5141;
  assign n5146 = n5142 & ~n5145;
  assign n5147 = n5146 ^ x71;
  assign n5148 = n5147 ^ x72;
  assign n5149 = n4874 & ~n5046;
  assign n5150 = n5149 ^ n4880;
  assign n5151 = n5150 ^ n5147;
  assign n5152 = n5148 & ~n5151;
  assign n5153 = n5152 ^ x72;
  assign n5154 = n5153 ^ x73;
  assign n5155 = n4884 & ~n5046;
  assign n5156 = n5155 ^ n4886;
  assign n5157 = n5156 ^ n5153;
  assign n5158 = n5154 & ~n5157;
  assign n5159 = n5158 ^ x73;
  assign n5160 = n5159 ^ x74;
  assign n5161 = n4890 & ~n5046;
  assign n5162 = n5161 ^ n4892;
  assign n5163 = n5162 ^ n5159;
  assign n5164 = n5160 & ~n5163;
  assign n5165 = n5164 ^ x74;
  assign n5166 = n5165 ^ x75;
  assign n5167 = n4896 & ~n5046;
  assign n5168 = n5167 ^ n4898;
  assign n5169 = n5168 ^ n5165;
  assign n5170 = n5166 & ~n5169;
  assign n5171 = n5170 ^ x75;
  assign n5172 = n5171 ^ x76;
  assign n5173 = n4902 & ~n5046;
  assign n5174 = n5173 ^ n4904;
  assign n5175 = n5174 ^ n5171;
  assign n5176 = n5172 & ~n5175;
  assign n5177 = n5176 ^ x76;
  assign n5178 = n5086 & n5177;
  assign n5179 = n5084 ^ x78;
  assign n5180 = x77 & n5080;
  assign n5181 = n5180 ^ n5084;
  assign n5182 = n5179 & ~n5181;
  assign n5183 = n5182 ^ x78;
  assign n5184 = ~n5178 & ~n5183;
  assign n5185 = n5184 ^ x79;
  assign n5186 = ~n4914 & ~n4918;
  assign n5187 = n5186 ^ x78;
  assign n5188 = ~n5046 & ~n5187;
  assign n5189 = n5188 ^ n4916;
  assign n5190 = n5189 ^ n5184;
  assign n5191 = ~n5185 & n5190;
  assign n5192 = n5191 ^ x79;
  assign n5193 = n5192 ^ x80;
  assign n5194 = n4923 & ~n5046;
  assign n5195 = n5194 ^ n4928;
  assign n5196 = n5195 ^ n5192;
  assign n5197 = n5193 & ~n5196;
  assign n5198 = n5197 ^ x80;
  assign n5199 = n5198 ^ x81;
  assign n5200 = n4932 & ~n5046;
  assign n5201 = n5200 ^ n4934;
  assign n5202 = n5201 ^ n5198;
  assign n5203 = n5199 & ~n5202;
  assign n5204 = n5203 ^ x81;
  assign n5205 = n5204 ^ x82;
  assign n5206 = n4937 ^ x81;
  assign n5207 = ~n5046 & n5206;
  assign n5208 = n5207 ^ n4813;
  assign n5209 = n5208 ^ n5204;
  assign n5210 = n5205 & ~n5209;
  assign n5211 = n5210 ^ x82;
  assign n5212 = n5211 ^ x83;
  assign n5213 = n4937 ^ n4813;
  assign n5214 = n5206 & ~n5213;
  assign n5215 = n5214 ^ x81;
  assign n5216 = n5215 ^ x82;
  assign n5217 = ~n5046 & n5216;
  assign n5218 = n5217 ^ n4810;
  assign n5219 = n5218 ^ n5211;
  assign n5220 = n5212 & ~n5219;
  assign n5221 = n5220 ^ x83;
  assign n5222 = n5221 ^ x84;
  assign n5223 = n4944 ^ x83;
  assign n5224 = ~n5046 & ~n5223;
  assign n5225 = n5224 ^ n4946;
  assign n5226 = n5225 ^ n5221;
  assign n5227 = n5222 & ~n5226;
  assign n5228 = n5227 ^ x84;
  assign n5229 = n5228 ^ x85;
  assign n5230 = n4946 ^ n4944;
  assign n5231 = ~n5223 & n5230;
  assign n5232 = n5231 ^ x83;
  assign n5233 = n5232 ^ x84;
  assign n5234 = ~n5046 & n5233;
  assign n5235 = n5234 ^ n4949;
  assign n5236 = n5235 ^ n5228;
  assign n5237 = n5229 & ~n5236;
  assign n5238 = n5237 ^ x85;
  assign n5239 = n5238 ^ x86;
  assign n5240 = ~n4959 & ~n5046;
  assign n5241 = n5240 ^ n4961;
  assign n5242 = n5241 ^ n5238;
  assign n5243 = n5239 & ~n5242;
  assign n5244 = n5243 ^ x86;
  assign n5245 = n5244 ^ x87;
  assign n5246 = n4965 & ~n5046;
  assign n5247 = n5246 ^ n4967;
  assign n5248 = n5247 ^ n5244;
  assign n5249 = n5245 & ~n5248;
  assign n5250 = n5249 ^ x87;
  assign n5251 = n5250 ^ x88;
  assign n5252 = ~n5046 & n5067;
  assign n5253 = n5252 ^ n4803;
  assign n5254 = n5253 ^ n5250;
  assign n5255 = n5251 & ~n5254;
  assign n5256 = n5255 ^ x88;
  assign n5257 = n5078 & n5256;
  assign n5258 = n5076 ^ x90;
  assign n5259 = x89 & n5073;
  assign n5260 = n5259 ^ n5076;
  assign n5261 = n5258 & ~n5260;
  assign n5262 = n5261 ^ x90;
  assign n5263 = ~n5257 & ~n5262;
  assign n5264 = n5263 ^ x91;
  assign n5265 = n4984 & ~n5046;
  assign n5266 = n5265 ^ n4986;
  assign n5267 = n5266 ^ n5263;
  assign n5268 = ~n5264 & n5267;
  assign n5269 = n5268 ^ x91;
  assign n5270 = n5269 ^ x92;
  assign n5271 = n4990 & ~n5046;
  assign n5272 = n5271 ^ n4992;
  assign n5273 = n5272 ^ n5269;
  assign n5274 = n5270 & ~n5273;
  assign n5275 = n5274 ^ x92;
  assign n5276 = ~n5066 & ~n5275;
  assign n5277 = n4995 ^ n4796;
  assign n5278 = n5063 & ~n5277;
  assign n5279 = n5278 ^ x92;
  assign n5280 = n5279 ^ x93;
  assign n5281 = ~n5046 & n5280;
  assign n5282 = n5281 ^ n4799;
  assign n5283 = ~x94 & ~n5282;
  assign n5284 = ~x93 & ~n5065;
  assign n5285 = ~n5283 & ~n5284;
  assign n5286 = ~n5276 & n5285;
  assign n5287 = x94 & n5282;
  assign n5288 = ~n5286 & ~n5287;
  assign n5289 = n5288 ^ x95;
  assign n5290 = ~n5003 & ~n5046;
  assign n5291 = n5290 ^ n5006;
  assign n5292 = n5291 ^ n5288;
  assign n5293 = ~n5289 & n5292;
  assign n5294 = n5293 ^ x95;
  assign n5295 = n5062 & n5294;
  assign n5296 = n5057 ^ x97;
  assign n5297 = x96 & n5060;
  assign n5298 = n5297 ^ n5057;
  assign n5299 = n5296 & ~n5298;
  assign n5300 = n5299 ^ x97;
  assign n5301 = ~n5295 & ~n5300;
  assign n5302 = n5301 ^ x98;
  assign n5303 = n5026 & ~n5046;
  assign n5304 = n5303 ^ n5028;
  assign n5305 = n5304 ^ n5301;
  assign n5306 = ~n5302 & n5305;
  assign n5307 = n5306 ^ x98;
  assign n5308 = n5307 ^ x99;
  assign n5309 = n5032 & ~n5046;
  assign n5310 = n5309 ^ n5034;
  assign n5311 = n5310 ^ n5307;
  assign n5312 = n5308 & ~n5311;
  assign n5313 = n5312 ^ x99;
  assign n5314 = ~n5055 & n5313;
  assign n5315 = x100 & n5053;
  assign n5316 = x101 & n5048;
  assign n5317 = n154 & ~n5316;
  assign n5318 = ~n5315 & n5317;
  assign n5319 = ~n5314 & n5318;
  assign n5320 = x100 & n5048;
  assign n5321 = n5313 & n5320;
  assign n5322 = n5319 & ~n5321;
  assign n5323 = n5256 ^ x89;
  assign n5324 = n5322 & n5323;
  assign n5325 = n5324 ^ n5073;
  assign n5326 = ~x90 & ~n5325;
  assign n5327 = n5256 ^ n5073;
  assign n5328 = n5323 & ~n5327;
  assign n5329 = n5328 ^ x89;
  assign n5330 = n5329 ^ x90;
  assign n5331 = n5322 & n5330;
  assign n5332 = n5331 ^ n5076;
  assign n5333 = ~x91 & ~n5332;
  assign n5334 = ~n5326 & ~n5333;
  assign n5335 = x65 & n5046;
  assign n5336 = n5322 & n5335;
  assign n5337 = n219 & ~n5046;
  assign n5338 = ~n5336 & ~n5337;
  assign n5339 = x26 & ~n5338;
  assign n5340 = n5046 ^ x65;
  assign n5341 = n341 & n5340;
  assign n5342 = x26 & n5341;
  assign n5343 = n5342 ^ n340;
  assign n5344 = n5322 & n5343;
  assign n5345 = n5344 ^ n5100;
  assign n5346 = ~n5339 & ~n5345;
  assign n5347 = n5346 ^ x27;
  assign n5348 = n5347 ^ x66;
  assign n5349 = x64 & n5322;
  assign n5350 = x25 & ~x65;
  assign n5351 = x26 & ~n5350;
  assign n5352 = n5349 & n5351;
  assign n5353 = ~x25 & x64;
  assign n5354 = ~x26 & n5353;
  assign n5355 = ~n5108 & ~n5354;
  assign n5356 = ~n5322 & ~n5355;
  assign n5357 = ~x25 & x65;
  assign n5358 = x64 & n5357;
  assign n5359 = ~x26 & n202;
  assign n5360 = ~n5358 & ~n5359;
  assign n5361 = ~n5356 & n5360;
  assign n5362 = ~n5352 & n5361;
  assign n5363 = n5362 ^ n5347;
  assign n5364 = n5348 & n5363;
  assign n5365 = n5364 ^ x66;
  assign n5366 = n5365 ^ x67;
  assign n5367 = n5113 ^ x66;
  assign n5368 = n5322 & ~n5367;
  assign n5369 = n5368 ^ n5098;
  assign n5370 = n5369 ^ n5365;
  assign n5371 = n5366 & ~n5370;
  assign n5372 = n5371 ^ x67;
  assign n5373 = n5372 ^ x68;
  assign n5374 = n5117 & n5322;
  assign n5375 = n5374 ^ n5120;
  assign n5376 = n5375 ^ n5372;
  assign n5377 = n5373 & ~n5376;
  assign n5378 = n5377 ^ x68;
  assign n5379 = n5378 ^ x69;
  assign n5380 = n5124 & n5322;
  assign n5381 = n5380 ^ n5126;
  assign n5382 = n5381 ^ n5378;
  assign n5383 = n5379 & ~n5382;
  assign n5384 = n5383 ^ x69;
  assign n5385 = n5384 ^ x70;
  assign n5386 = n5130 & n5322;
  assign n5387 = n5386 ^ n5132;
  assign n5388 = n5387 ^ n5384;
  assign n5389 = n5385 & ~n5388;
  assign n5390 = n5389 ^ x70;
  assign n5391 = n5390 ^ x71;
  assign n5392 = n5136 & n5322;
  assign n5393 = n5392 ^ n5138;
  assign n5394 = n5393 ^ n5390;
  assign n5395 = n5391 & ~n5394;
  assign n5396 = n5395 ^ x71;
  assign n5397 = n5396 ^ x72;
  assign n5398 = n5142 & n5322;
  assign n5399 = n5398 ^ n5144;
  assign n5400 = n5399 ^ n5396;
  assign n5401 = n5397 & ~n5400;
  assign n5402 = n5401 ^ x72;
  assign n5403 = n5402 ^ x73;
  assign n5404 = n5148 & n5322;
  assign n5405 = n5404 ^ n5150;
  assign n5406 = n5405 ^ n5402;
  assign n5407 = n5403 & ~n5406;
  assign n5408 = n5407 ^ x73;
  assign n5409 = n5408 ^ x74;
  assign n5410 = n5154 & n5322;
  assign n5411 = n5410 ^ n5156;
  assign n5412 = n5411 ^ n5408;
  assign n5413 = n5409 & ~n5412;
  assign n5414 = n5413 ^ x74;
  assign n5415 = n5414 ^ x75;
  assign n5416 = n5160 & n5322;
  assign n5417 = n5416 ^ n5162;
  assign n5418 = n5417 ^ n5414;
  assign n5419 = n5415 & ~n5418;
  assign n5420 = n5419 ^ x75;
  assign n5421 = n5420 ^ x76;
  assign n5422 = n5166 & n5322;
  assign n5423 = n5422 ^ n5168;
  assign n5424 = n5423 ^ n5420;
  assign n5425 = n5421 & ~n5424;
  assign n5426 = n5425 ^ x76;
  assign n5427 = n5426 ^ x77;
  assign n5428 = n5172 & n5322;
  assign n5429 = n5428 ^ n5174;
  assign n5430 = n5429 ^ n5426;
  assign n5431 = n5427 & ~n5430;
  assign n5432 = n5431 ^ x77;
  assign n5433 = n5432 ^ x78;
  assign n5434 = n5177 ^ x77;
  assign n5435 = n5322 & n5434;
  assign n5436 = n5435 ^ n5080;
  assign n5437 = n5436 ^ n5432;
  assign n5438 = n5433 & ~n5437;
  assign n5439 = n5438 ^ x78;
  assign n5440 = n5439 ^ x79;
  assign n5441 = n5177 ^ n5080;
  assign n5442 = n5434 & ~n5441;
  assign n5443 = n5442 ^ x77;
  assign n5444 = n5443 ^ x78;
  assign n5445 = n5322 & n5444;
  assign n5446 = n5445 ^ n5084;
  assign n5447 = n5446 ^ n5439;
  assign n5448 = n5440 & ~n5447;
  assign n5449 = n5448 ^ x79;
  assign n5450 = n5449 ^ x80;
  assign n5451 = ~n5185 & n5322;
  assign n5452 = n5451 ^ n5189;
  assign n5453 = n5452 ^ n5449;
  assign n5454 = n5450 & ~n5453;
  assign n5455 = n5454 ^ x80;
  assign n5456 = n5455 ^ x81;
  assign n5457 = n5193 & n5322;
  assign n5458 = n5457 ^ n5195;
  assign n5459 = n5458 ^ n5455;
  assign n5460 = n5456 & ~n5459;
  assign n5461 = n5460 ^ x81;
  assign n5462 = n5461 ^ x82;
  assign n5463 = n5199 & n5322;
  assign n5464 = n5463 ^ n5201;
  assign n5465 = n5464 ^ n5461;
  assign n5466 = n5462 & ~n5465;
  assign n5467 = n5466 ^ x82;
  assign n5468 = n5467 ^ x83;
  assign n5469 = n5205 & n5322;
  assign n5470 = n5469 ^ n5208;
  assign n5471 = n5470 ^ n5467;
  assign n5472 = n5468 & ~n5471;
  assign n5473 = n5472 ^ x83;
  assign n5474 = n5473 ^ x84;
  assign n5475 = n5212 & n5322;
  assign n5476 = n5475 ^ n5218;
  assign n5477 = n5476 ^ n5473;
  assign n5478 = n5474 & ~n5477;
  assign n5479 = n5478 ^ x84;
  assign n5480 = n5479 ^ x85;
  assign n5481 = n5222 & n5322;
  assign n5482 = n5481 ^ n5225;
  assign n5483 = n5482 ^ n5479;
  assign n5484 = n5480 & ~n5483;
  assign n5485 = n5484 ^ x85;
  assign n5486 = n5485 ^ x86;
  assign n5487 = n5229 & n5322;
  assign n5488 = n5487 ^ n5235;
  assign n5489 = n5488 ^ n5485;
  assign n5490 = n5486 & ~n5489;
  assign n5491 = n5490 ^ x86;
  assign n5492 = n5491 ^ x87;
  assign n5493 = n5239 & n5322;
  assign n5494 = n5493 ^ n5241;
  assign n5495 = n5494 ^ n5491;
  assign n5496 = n5492 & ~n5495;
  assign n5497 = n5496 ^ x87;
  assign n5498 = n5497 ^ x88;
  assign n5499 = n5245 & n5322;
  assign n5500 = n5499 ^ n5247;
  assign n5501 = n5500 ^ n5497;
  assign n5502 = n5498 & ~n5501;
  assign n5503 = n5502 ^ x88;
  assign n5504 = n5503 ^ x89;
  assign n5505 = n5251 & n5322;
  assign n5506 = n5505 ^ n5253;
  assign n5507 = n5506 ^ n5503;
  assign n5508 = n5504 & ~n5507;
  assign n5509 = n5508 ^ x89;
  assign n5510 = n5334 & n5509;
  assign n5511 = n5332 ^ x91;
  assign n5512 = x90 & n5325;
  assign n5513 = n5512 ^ n5332;
  assign n5514 = n5511 & ~n5513;
  assign n5515 = n5514 ^ x91;
  assign n5516 = ~n5510 & ~n5515;
  assign n5517 = ~n5264 & n5322;
  assign n5518 = n5517 ^ n5266;
  assign n5519 = ~x92 & ~n5518;
  assign n5520 = n5270 & n5322;
  assign n5521 = n5520 ^ n5272;
  assign n5522 = ~x93 & ~n5521;
  assign n5523 = ~n5519 & ~n5522;
  assign n5524 = ~n5516 & n5523;
  assign n5525 = n5521 ^ x93;
  assign n5526 = x92 & n5518;
  assign n5527 = n5526 ^ n5521;
  assign n5528 = n5525 & ~n5527;
  assign n5529 = n5528 ^ x93;
  assign n5530 = ~n5524 & ~n5529;
  assign n5531 = n5530 ^ x94;
  assign n5532 = n5275 ^ x93;
  assign n5533 = n5322 & n5532;
  assign n5534 = n5533 ^ n5065;
  assign n5535 = n5534 ^ n5530;
  assign n5536 = ~n5531 & n5535;
  assign n5537 = n5536 ^ x94;
  assign n5538 = n5537 ^ x95;
  assign n5539 = ~n5276 & ~n5284;
  assign n5540 = n5539 ^ x94;
  assign n5541 = n5322 & n5540;
  assign n5542 = n5541 ^ n5282;
  assign n5543 = n5542 ^ n5537;
  assign n5544 = n5538 & ~n5543;
  assign n5545 = n5544 ^ x95;
  assign n5546 = n5545 ^ x96;
  assign n5547 = ~n5289 & n5322;
  assign n5548 = n5547 ^ n5291;
  assign n5549 = n5548 ^ n5545;
  assign n5550 = n5546 & ~n5549;
  assign n5551 = n5550 ^ x96;
  assign n5552 = n5551 ^ x97;
  assign n5553 = n5294 ^ x96;
  assign n5554 = n5322 & n5553;
  assign n5555 = n5554 ^ n5060;
  assign n5556 = n5555 ^ n5551;
  assign n5557 = n5552 & ~n5556;
  assign n5558 = n5557 ^ x97;
  assign n5559 = n5558 ^ x98;
  assign n5560 = n5294 ^ n5060;
  assign n5561 = n5553 & ~n5560;
  assign n5562 = n5561 ^ x96;
  assign n5563 = n5562 ^ x97;
  assign n5564 = n5322 & n5563;
  assign n5565 = n5564 ^ n5057;
  assign n5566 = n5565 ^ n5558;
  assign n5567 = n5559 & ~n5566;
  assign n5568 = n5567 ^ x98;
  assign n5569 = n5568 ^ x99;
  assign n5570 = ~n5302 & n5322;
  assign n5571 = n5570 ^ n5304;
  assign n5572 = n5571 ^ n5568;
  assign n5573 = n5569 & ~n5572;
  assign n5574 = n5573 ^ x99;
  assign n5575 = n5574 ^ x100;
  assign n5576 = n5308 & n5322;
  assign n5577 = n5576 ^ n5310;
  assign n5578 = n5577 ^ n5574;
  assign n5579 = n5575 & ~n5578;
  assign n5580 = n5579 ^ x100;
  assign n5581 = n5580 ^ x101;
  assign n5582 = n5313 ^ x100;
  assign n5583 = n5319 & n5582;
  assign n5584 = n5583 ^ n5052;
  assign n5585 = n5584 ^ n5580;
  assign n5586 = n5581 & n5585;
  assign n5587 = n5586 ^ x101;
  assign n5588 = n153 & ~n5587;
  assign n5589 = ~n154 & n5047;
  assign n5590 = ~n5588 & n5589;
  assign n5591 = ~n242 & n5319;
  assign n5592 = ~n5048 & ~n5591;
  assign n5593 = ~x102 & n5592;
  assign n5594 = n5587 & ~n5593;
  assign n5595 = x102 & ~n5592;
  assign n5596 = n153 & ~n5595;
  assign n5597 = ~n5594 & n5596;
  assign n5598 = n5581 & n5597;
  assign n5599 = n5598 ^ n5584;
  assign n5600 = ~x102 & n5599;
  assign n5601 = ~n242 & ~n5590;
  assign n5602 = ~x103 & ~n5601;
  assign n5603 = ~n5600 & ~n5602;
  assign n5604 = n5546 & n5597;
  assign n5605 = n5604 ^ n5548;
  assign n5606 = ~x97 & ~n5605;
  assign n5607 = n5385 & n5597;
  assign n5608 = n5607 ^ n5387;
  assign n5609 = ~x71 & ~n5608;
  assign n5610 = n5391 & n5597;
  assign n5611 = n5610 ^ n5393;
  assign n5612 = ~x72 & ~n5611;
  assign n5613 = ~n5609 & ~n5612;
  assign n5614 = x65 & ~n5322;
  assign n5615 = x25 & n5614;
  assign n5616 = n5597 & n5615;
  assign n5617 = n5349 & n5350;
  assign n5618 = ~n5616 & ~n5617;
  assign n5619 = n5322 ^ x65;
  assign n5620 = n341 & ~n5619;
  assign n5621 = x25 & n5620;
  assign n5622 = n5621 ^ n340;
  assign n5623 = n5597 & n5622;
  assign n5624 = n5623 ^ n5349;
  assign n5625 = n5618 & ~n5624;
  assign n5626 = n5625 ^ x26;
  assign n5627 = n5626 ^ x66;
  assign n5628 = x64 & n5597;
  assign n5629 = x24 & n5350;
  assign n5630 = n5629 ^ x25;
  assign n5631 = n5628 & n5630;
  assign n5632 = ~x24 & n5353;
  assign n5633 = ~n5357 & ~n5632;
  assign n5634 = ~n5597 & ~n5633;
  assign n5635 = ~x24 & x65;
  assign n5636 = n5635 ^ n5357;
  assign n5637 = x64 & n5636;
  assign n5638 = n5637 ^ n5357;
  assign n5639 = ~n5634 & ~n5638;
  assign n5640 = ~n5631 & n5639;
  assign n5641 = n5640 ^ n5626;
  assign n5642 = n5627 & n5641;
  assign n5643 = n5642 ^ x66;
  assign n5644 = n5643 ^ x67;
  assign n5645 = n5362 ^ x66;
  assign n5646 = n5597 & ~n5645;
  assign n5647 = n5646 ^ n5347;
  assign n5648 = n5647 ^ n5643;
  assign n5649 = n5644 & ~n5648;
  assign n5650 = n5649 ^ x67;
  assign n5651 = n5650 ^ x68;
  assign n5652 = n5366 & n5597;
  assign n5653 = n5652 ^ n5369;
  assign n5654 = n5653 ^ n5650;
  assign n5655 = n5651 & ~n5654;
  assign n5656 = n5655 ^ x68;
  assign n5657 = n5656 ^ x69;
  assign n5658 = n5373 & n5597;
  assign n5659 = n5658 ^ n5375;
  assign n5660 = n5659 ^ n5656;
  assign n5661 = n5657 & ~n5660;
  assign n5662 = n5661 ^ x69;
  assign n5663 = n5662 ^ x70;
  assign n5664 = n5379 & n5597;
  assign n5665 = n5664 ^ n5381;
  assign n5666 = n5665 ^ n5662;
  assign n5667 = n5663 & ~n5666;
  assign n5668 = n5667 ^ x70;
  assign n5669 = n5613 & n5668;
  assign n5670 = n5611 ^ x72;
  assign n5671 = x71 & n5608;
  assign n5672 = n5671 ^ n5611;
  assign n5673 = n5670 & ~n5672;
  assign n5674 = n5673 ^ x72;
  assign n5675 = ~n5669 & ~n5674;
  assign n5676 = n5675 ^ x73;
  assign n5677 = n5397 & n5597;
  assign n5678 = n5677 ^ n5399;
  assign n5679 = n5678 ^ n5675;
  assign n5680 = ~n5676 & n5679;
  assign n5681 = n5680 ^ x73;
  assign n5682 = n5681 ^ x74;
  assign n5683 = n5403 & n5597;
  assign n5684 = n5683 ^ n5405;
  assign n5685 = n5684 ^ n5681;
  assign n5686 = n5682 & ~n5685;
  assign n5687 = n5686 ^ x74;
  assign n5688 = n5687 ^ x75;
  assign n5689 = n5409 & n5597;
  assign n5690 = n5689 ^ n5411;
  assign n5691 = n5690 ^ n5687;
  assign n5692 = n5688 & ~n5691;
  assign n5693 = n5692 ^ x75;
  assign n5694 = n5693 ^ x76;
  assign n5695 = n5415 & n5597;
  assign n5696 = n5695 ^ n5417;
  assign n5697 = n5696 ^ n5693;
  assign n5698 = n5694 & ~n5697;
  assign n5699 = n5698 ^ x76;
  assign n5700 = n5699 ^ x77;
  assign n5701 = n5421 & n5597;
  assign n5702 = n5701 ^ n5423;
  assign n5703 = n5702 ^ n5699;
  assign n5704 = n5700 & ~n5703;
  assign n5705 = n5704 ^ x77;
  assign n5706 = n5705 ^ x78;
  assign n5707 = n5427 & n5597;
  assign n5708 = n5707 ^ n5429;
  assign n5709 = n5708 ^ n5705;
  assign n5710 = n5706 & ~n5709;
  assign n5711 = n5710 ^ x78;
  assign n5712 = n5711 ^ x79;
  assign n5713 = n5433 & n5597;
  assign n5714 = n5713 ^ n5436;
  assign n5715 = n5714 ^ n5711;
  assign n5716 = n5712 & ~n5715;
  assign n5717 = n5716 ^ x79;
  assign n5718 = n5717 ^ x80;
  assign n5719 = n5440 & n5597;
  assign n5720 = n5719 ^ n5446;
  assign n5721 = n5720 ^ n5717;
  assign n5722 = n5718 & ~n5721;
  assign n5723 = n5722 ^ x80;
  assign n5724 = n5723 ^ x81;
  assign n5725 = n5450 & n5597;
  assign n5726 = n5725 ^ n5452;
  assign n5727 = n5726 ^ n5723;
  assign n5728 = n5724 & ~n5727;
  assign n5729 = n5728 ^ x81;
  assign n5730 = n5729 ^ x82;
  assign n5731 = n5456 & n5597;
  assign n5732 = n5731 ^ n5458;
  assign n5733 = n5732 ^ n5729;
  assign n5734 = n5730 & ~n5733;
  assign n5735 = n5734 ^ x82;
  assign n5736 = n5735 ^ x83;
  assign n5737 = n5462 & n5597;
  assign n5738 = n5737 ^ n5464;
  assign n5739 = n5738 ^ n5735;
  assign n5740 = n5736 & ~n5739;
  assign n5741 = n5740 ^ x83;
  assign n5742 = n5741 ^ x84;
  assign n5743 = n5468 & n5597;
  assign n5744 = n5743 ^ n5470;
  assign n5745 = n5744 ^ n5741;
  assign n5746 = n5742 & ~n5745;
  assign n5747 = n5746 ^ x84;
  assign n5748 = n5747 ^ x85;
  assign n5749 = n5474 & n5597;
  assign n5750 = n5749 ^ n5476;
  assign n5751 = n5750 ^ n5747;
  assign n5752 = n5748 & ~n5751;
  assign n5753 = n5752 ^ x85;
  assign n5754 = n5753 ^ x86;
  assign n5755 = n5480 & n5597;
  assign n5756 = n5755 ^ n5482;
  assign n5757 = n5756 ^ n5753;
  assign n5758 = n5754 & ~n5757;
  assign n5759 = n5758 ^ x86;
  assign n5760 = n5759 ^ x87;
  assign n5761 = n5486 & n5597;
  assign n5762 = n5761 ^ n5488;
  assign n5763 = n5762 ^ n5759;
  assign n5764 = n5760 & ~n5763;
  assign n5765 = n5764 ^ x87;
  assign n5766 = n5765 ^ x88;
  assign n5767 = n5492 & n5597;
  assign n5768 = n5767 ^ n5494;
  assign n5769 = n5768 ^ n5765;
  assign n5770 = n5766 & ~n5769;
  assign n5771 = n5770 ^ x88;
  assign n5772 = n5771 ^ x89;
  assign n5773 = n5498 & n5597;
  assign n5774 = n5773 ^ n5500;
  assign n5775 = n5774 ^ n5771;
  assign n5776 = n5772 & ~n5775;
  assign n5777 = n5776 ^ x89;
  assign n5778 = n5777 ^ x90;
  assign n5779 = n5504 & n5597;
  assign n5780 = n5779 ^ n5506;
  assign n5781 = n5780 ^ n5777;
  assign n5782 = n5778 & ~n5781;
  assign n5783 = n5782 ^ x90;
  assign n5784 = n5783 ^ x91;
  assign n5785 = n5509 ^ x90;
  assign n5786 = n5597 & n5785;
  assign n5787 = n5786 ^ n5325;
  assign n5788 = n5787 ^ n5783;
  assign n5789 = n5784 & ~n5788;
  assign n5790 = n5789 ^ x91;
  assign n5791 = n5790 ^ x92;
  assign n5792 = n5509 ^ n5325;
  assign n5793 = n5785 & ~n5792;
  assign n5794 = n5793 ^ x90;
  assign n5795 = n5794 ^ x91;
  assign n5796 = n5597 & n5795;
  assign n5797 = n5796 ^ n5332;
  assign n5798 = n5797 ^ n5790;
  assign n5799 = n5791 & ~n5798;
  assign n5800 = n5799 ^ x92;
  assign n5801 = n5800 ^ x93;
  assign n5802 = n5516 ^ x92;
  assign n5803 = n5597 & ~n5802;
  assign n5804 = n5803 ^ n5518;
  assign n5805 = n5804 ^ n5800;
  assign n5806 = n5801 & ~n5805;
  assign n5807 = n5806 ^ x93;
  assign n5808 = n5807 ^ x94;
  assign n5809 = n5518 ^ n5516;
  assign n5810 = ~n5802 & n5809;
  assign n5811 = n5810 ^ x92;
  assign n5812 = n5811 ^ x93;
  assign n5813 = n5597 & n5812;
  assign n5814 = n5813 ^ n5521;
  assign n5815 = n5814 ^ n5807;
  assign n5816 = n5808 & ~n5815;
  assign n5817 = n5816 ^ x94;
  assign n5818 = n5817 ^ x95;
  assign n5819 = ~n5531 & n5597;
  assign n5820 = n5819 ^ n5534;
  assign n5821 = n5820 ^ n5817;
  assign n5822 = n5818 & ~n5821;
  assign n5823 = n5822 ^ x95;
  assign n5824 = n5823 ^ x96;
  assign n5825 = n5538 & n5597;
  assign n5826 = n5825 ^ n5542;
  assign n5827 = n5826 ^ n5823;
  assign n5828 = n5824 & ~n5827;
  assign n5829 = n5828 ^ x96;
  assign n5830 = ~n5606 & n5829;
  assign n5831 = x97 & n5605;
  assign n5832 = n5552 & n5597;
  assign n5833 = n5832 ^ n5555;
  assign n5834 = x98 & n5833;
  assign n5835 = ~n5831 & ~n5834;
  assign n5836 = ~n5830 & n5835;
  assign n5837 = ~x98 & ~n5833;
  assign n5838 = ~n5836 & ~n5837;
  assign n5839 = n5838 ^ x99;
  assign n5840 = n5559 & n5597;
  assign n5841 = n5840 ^ n5565;
  assign n5842 = n5841 ^ n5838;
  assign n5843 = n5839 & ~n5842;
  assign n5844 = n5843 ^ x99;
  assign n5845 = n5844 ^ x100;
  assign n5846 = n5569 & n5597;
  assign n5847 = n5846 ^ n5571;
  assign n5848 = n5847 ^ n5844;
  assign n5849 = n5845 & ~n5848;
  assign n5850 = n5849 ^ x100;
  assign n5851 = n5850 ^ x101;
  assign n5852 = n5575 & n5597;
  assign n5853 = n5852 ^ n5577;
  assign n5854 = n5853 ^ n5850;
  assign n5855 = n5851 & ~n5854;
  assign n5856 = n5855 ^ x101;
  assign n5857 = n5603 & n5856;
  assign n5858 = x102 & ~n5602;
  assign n5859 = ~n5599 & n5858;
  assign n5860 = n152 & ~n5048;
  assign n5861 = ~n153 & ~n5860;
  assign n5862 = ~n5859 & ~n5861;
  assign n5863 = ~n5857 & n5862;
  assign n5864 = n5590 & ~n5863;
  assign n5865 = n5851 & n5863;
  assign n5866 = n5865 ^ n5853;
  assign n5867 = x102 & n5866;
  assign n5868 = n5818 & n5863;
  assign n5869 = n5868 ^ n5820;
  assign n5870 = ~x96 & ~n5869;
  assign n5871 = n5784 & n5863;
  assign n5872 = n5871 ^ n5787;
  assign n5873 = ~x92 & ~n5872;
  assign n5874 = n5791 & n5863;
  assign n5875 = n5874 ^ n5797;
  assign n5876 = ~x93 & ~n5875;
  assign n5877 = ~n5873 & ~n5876;
  assign n5878 = n5748 & n5863;
  assign n5879 = n5878 ^ n5750;
  assign n5880 = ~x86 & ~n5879;
  assign n5881 = n5754 & n5863;
  assign n5882 = n5881 ^ n5756;
  assign n5883 = ~x87 & ~n5882;
  assign n5884 = ~n5880 & ~n5883;
  assign n5885 = n293 & ~n5597;
  assign n5886 = n5885 ^ x65;
  assign n5887 = ~x24 & n5886;
  assign n5888 = ~x65 & ~n5887;
  assign n5889 = n5863 & ~n5888;
  assign n5890 = ~n5628 & ~n5889;
  assign n5891 = x65 & n5597;
  assign n5892 = x24 & ~n5891;
  assign n5893 = ~n202 & ~n5892;
  assign n5894 = ~n5887 & n5893;
  assign n5895 = n5863 & n5894;
  assign n5896 = ~n5890 & ~n5895;
  assign n5897 = n5896 ^ x25;
  assign n5898 = n5897 ^ x66;
  assign n5899 = x64 & n5863;
  assign n5900 = x24 & ~x65;
  assign n5901 = x23 & n5900;
  assign n5902 = n5901 ^ x24;
  assign n5903 = n5899 & n5902;
  assign n5904 = ~x23 & x64;
  assign n5905 = ~x24 & n5904;
  assign n5906 = ~n5635 & ~n5905;
  assign n5907 = ~n5863 & ~n5906;
  assign n5908 = x24 ^ x23;
  assign n5909 = ~x64 & n5908;
  assign n5910 = n5909 ^ x23;
  assign n5911 = x65 & ~n5910;
  assign n5912 = ~n5907 & ~n5911;
  assign n5913 = ~n5903 & n5912;
  assign n5914 = n5913 ^ n5897;
  assign n5915 = ~n5898 & ~n5914;
  assign n5916 = n5915 ^ x66;
  assign n5917 = n5916 ^ x67;
  assign n5918 = n5640 ^ x66;
  assign n5919 = n5863 & ~n5918;
  assign n5920 = n5919 ^ n5626;
  assign n5921 = n5920 ^ n5916;
  assign n5922 = n5917 & ~n5921;
  assign n5923 = n5922 ^ x67;
  assign n5924 = n5923 ^ x68;
  assign n5925 = n5644 & n5863;
  assign n5926 = n5925 ^ n5647;
  assign n5927 = n5926 ^ n5923;
  assign n5928 = n5924 & ~n5927;
  assign n5929 = n5928 ^ x68;
  assign n5930 = n5929 ^ x69;
  assign n5931 = n5651 & n5863;
  assign n5932 = n5931 ^ n5653;
  assign n5933 = n5932 ^ n5929;
  assign n5934 = n5930 & ~n5933;
  assign n5935 = n5934 ^ x69;
  assign n5936 = n5935 ^ x70;
  assign n5937 = n5657 & n5863;
  assign n5938 = n5937 ^ n5659;
  assign n5939 = n5938 ^ n5935;
  assign n5940 = n5936 & ~n5939;
  assign n5941 = n5940 ^ x70;
  assign n5942 = n5941 ^ x71;
  assign n5943 = n5663 & n5863;
  assign n5944 = n5943 ^ n5665;
  assign n5945 = n5944 ^ n5941;
  assign n5946 = n5942 & ~n5945;
  assign n5947 = n5946 ^ x71;
  assign n5948 = n5947 ^ x72;
  assign n5949 = n5668 ^ x71;
  assign n5950 = n5863 & n5949;
  assign n5951 = n5950 ^ n5608;
  assign n5952 = n5951 ^ n5947;
  assign n5953 = n5948 & ~n5952;
  assign n5954 = n5953 ^ x72;
  assign n5955 = n5954 ^ x73;
  assign n5956 = n5668 ^ n5608;
  assign n5957 = n5949 & ~n5956;
  assign n5958 = n5957 ^ x71;
  assign n5959 = n5958 ^ x72;
  assign n5960 = n5863 & n5959;
  assign n5961 = n5960 ^ n5611;
  assign n5962 = n5961 ^ n5954;
  assign n5963 = n5955 & ~n5962;
  assign n5964 = n5963 ^ x73;
  assign n5965 = n5964 ^ x74;
  assign n5966 = ~n5676 & n5863;
  assign n5967 = n5966 ^ n5678;
  assign n5968 = n5967 ^ n5964;
  assign n5969 = n5965 & ~n5968;
  assign n5970 = n5969 ^ x74;
  assign n5971 = n5970 ^ x75;
  assign n5972 = n5682 & n5863;
  assign n5973 = n5972 ^ n5684;
  assign n5974 = n5973 ^ n5970;
  assign n5975 = n5971 & ~n5974;
  assign n5976 = n5975 ^ x75;
  assign n5977 = n5976 ^ x76;
  assign n5978 = n5688 & n5863;
  assign n5979 = n5978 ^ n5690;
  assign n5980 = n5979 ^ n5976;
  assign n5981 = n5977 & ~n5980;
  assign n5982 = n5981 ^ x76;
  assign n5983 = n5982 ^ x77;
  assign n5984 = n5694 & n5863;
  assign n5985 = n5984 ^ n5696;
  assign n5986 = n5985 ^ n5982;
  assign n5987 = n5983 & ~n5986;
  assign n5988 = n5987 ^ x77;
  assign n5989 = n5988 ^ x78;
  assign n5990 = n5700 & n5863;
  assign n5991 = n5990 ^ n5702;
  assign n5992 = n5991 ^ n5988;
  assign n5993 = n5989 & ~n5992;
  assign n5994 = n5993 ^ x78;
  assign n5995 = n5994 ^ x79;
  assign n5996 = n5706 & n5863;
  assign n5997 = n5996 ^ n5708;
  assign n5998 = n5997 ^ n5994;
  assign n5999 = n5995 & ~n5998;
  assign n6000 = n5999 ^ x79;
  assign n6001 = n6000 ^ x80;
  assign n6002 = n5712 & n5863;
  assign n6003 = n6002 ^ n5714;
  assign n6004 = n6003 ^ n6000;
  assign n6005 = n6001 & ~n6004;
  assign n6006 = n6005 ^ x80;
  assign n6007 = n6006 ^ x81;
  assign n6008 = n5718 & n5863;
  assign n6009 = n6008 ^ n5720;
  assign n6010 = n6009 ^ n6006;
  assign n6011 = n6007 & ~n6010;
  assign n6012 = n6011 ^ x81;
  assign n6013 = n6012 ^ x82;
  assign n6014 = n5724 & n5863;
  assign n6015 = n6014 ^ n5726;
  assign n6016 = n6015 ^ n6012;
  assign n6017 = n6013 & ~n6016;
  assign n6018 = n6017 ^ x82;
  assign n6019 = n6018 ^ x83;
  assign n6020 = n5730 & n5863;
  assign n6021 = n6020 ^ n5732;
  assign n6022 = n6021 ^ n6018;
  assign n6023 = n6019 & ~n6022;
  assign n6024 = n6023 ^ x83;
  assign n6025 = n6024 ^ x84;
  assign n6026 = n5736 & n5863;
  assign n6027 = n6026 ^ n5738;
  assign n6028 = n6027 ^ n6024;
  assign n6029 = n6025 & ~n6028;
  assign n6030 = n6029 ^ x84;
  assign n6031 = n6030 ^ x85;
  assign n6032 = n5742 & n5863;
  assign n6033 = n6032 ^ n5744;
  assign n6034 = n6033 ^ n6030;
  assign n6035 = n6031 & ~n6034;
  assign n6036 = n6035 ^ x85;
  assign n6037 = n5884 & n6036;
  assign n6038 = n5882 ^ x87;
  assign n6039 = x86 & n5879;
  assign n6040 = n6039 ^ n5882;
  assign n6041 = n6038 & ~n6040;
  assign n6042 = n6041 ^ x87;
  assign n6043 = ~n6037 & ~n6042;
  assign n6044 = n5760 & n5863;
  assign n6045 = n6044 ^ n5762;
  assign n6046 = ~x88 & ~n6045;
  assign n6047 = n5766 & n5863;
  assign n6048 = n6047 ^ n5768;
  assign n6049 = ~x89 & ~n6048;
  assign n6050 = ~n6046 & ~n6049;
  assign n6051 = ~n6043 & n6050;
  assign n6052 = n6048 ^ x89;
  assign n6053 = x88 & n6045;
  assign n6054 = n6053 ^ n6048;
  assign n6055 = n6052 & ~n6054;
  assign n6056 = n6055 ^ x89;
  assign n6057 = ~n6051 & ~n6056;
  assign n6058 = n6057 ^ x90;
  assign n6059 = n5772 & n5863;
  assign n6060 = n6059 ^ n5774;
  assign n6061 = n6060 ^ n6057;
  assign n6062 = ~n6058 & n6061;
  assign n6063 = n6062 ^ x90;
  assign n6064 = n6063 ^ x91;
  assign n6065 = n5778 & n5863;
  assign n6066 = n6065 ^ n5780;
  assign n6067 = n6066 ^ n6063;
  assign n6068 = n6064 & ~n6067;
  assign n6069 = n6068 ^ x91;
  assign n6070 = n5877 & n6069;
  assign n6071 = n5875 ^ x93;
  assign n6072 = x92 & n5872;
  assign n6073 = n6072 ^ n5875;
  assign n6074 = n6071 & ~n6073;
  assign n6075 = n6074 ^ x93;
  assign n6076 = ~n6070 & ~n6075;
  assign n6077 = n6076 ^ x94;
  assign n6078 = n5801 & n5863;
  assign n6079 = n6078 ^ n5804;
  assign n6080 = n6079 ^ n6076;
  assign n6081 = ~n6077 & n6080;
  assign n6082 = n6081 ^ x94;
  assign n6083 = n6082 ^ x95;
  assign n6084 = n5808 & n5863;
  assign n6085 = n6084 ^ n5814;
  assign n6086 = n6085 ^ n6082;
  assign n6087 = n6083 & ~n6086;
  assign n6088 = n6087 ^ x95;
  assign n6089 = ~n5870 & n6088;
  assign n6090 = n5824 & n5863;
  assign n6091 = n6090 ^ n5826;
  assign n6092 = x97 & n6091;
  assign n6093 = x96 & n5869;
  assign n6094 = ~n6092 & ~n6093;
  assign n6095 = ~n6089 & n6094;
  assign n6096 = ~x97 & ~n6091;
  assign n6097 = ~n6095 & ~n6096;
  assign n6098 = n6097 ^ x98;
  assign n6099 = n5829 ^ x97;
  assign n6100 = n5863 & n6099;
  assign n6101 = n6100 ^ n5605;
  assign n6102 = n6101 ^ n6097;
  assign n6103 = n6098 & ~n6102;
  assign n6104 = n6103 ^ x98;
  assign n6105 = n6104 ^ x99;
  assign n6106 = ~n5830 & ~n5831;
  assign n6107 = n6106 ^ x98;
  assign n6108 = n5863 & ~n6107;
  assign n6109 = n6108 ^ n5833;
  assign n6110 = n6109 ^ n6104;
  assign n6111 = n6105 & ~n6110;
  assign n6112 = n6111 ^ x99;
  assign n6113 = n6112 ^ x100;
  assign n6114 = n5839 & n5863;
  assign n6115 = n6114 ^ n5841;
  assign n6116 = n6115 ^ n6112;
  assign n6117 = n6113 & ~n6116;
  assign n6118 = n6117 ^ x100;
  assign n6119 = n6118 ^ x101;
  assign n6120 = n5845 & n5863;
  assign n6121 = n6120 ^ n5847;
  assign n6122 = n6121 ^ n6118;
  assign n6123 = n6119 & ~n6122;
  assign n6124 = n6123 ^ x101;
  assign n6125 = ~n5867 & ~n6124;
  assign n6126 = ~x102 & ~n5866;
  assign n6127 = n5856 ^ x102;
  assign n6128 = n5863 & n6127;
  assign n6129 = n6128 ^ n5599;
  assign n6130 = ~x103 & n6129;
  assign n6131 = ~n6126 & ~n6130;
  assign n6132 = ~n6125 & n6131;
  assign n6133 = ~n242 & ~n5864;
  assign n6134 = x104 & n6133;
  assign n6135 = x103 & ~n6129;
  assign n6136 = ~n6134 & ~n6135;
  assign n6137 = ~n6132 & n6136;
  assign n6138 = ~x104 & ~n6133;
  assign n6139 = ~n6137 & ~n6138;
  assign n6140 = ~x108 & n147;
  assign n6141 = n150 & n6140;
  assign n6142 = ~x105 & n6141;
  assign n6143 = ~n6139 & n6142;
  assign n6144 = n5864 & ~n6143;
  assign n6145 = ~n242 & ~n6144;
  assign n6146 = ~x107 & n6140;
  assign n6147 = x105 & n6145;
  assign n6148 = n6141 & ~n6147;
  assign n6149 = n5936 & n6143;
  assign n6150 = n6149 ^ n5938;
  assign n6151 = ~x71 & ~n6150;
  assign n6152 = n5942 & n6143;
  assign n6153 = n6152 ^ n5944;
  assign n6154 = ~x72 & ~n6153;
  assign n6155 = ~n6151 & ~n6154;
  assign n6156 = x65 & ~n5863;
  assign n6157 = n6143 & n6156;
  assign n6158 = ~x65 & n5863;
  assign n6159 = x64 & n6158;
  assign n6160 = ~n6157 & ~n6159;
  assign n6161 = x23 & ~n6160;
  assign n6162 = n5863 ^ x65;
  assign n6163 = n341 & ~n6162;
  assign n6164 = x23 & n6163;
  assign n6165 = n6164 ^ n340;
  assign n6166 = n6143 & n6165;
  assign n6167 = n6166 ^ n5899;
  assign n6168 = ~n6161 & ~n6167;
  assign n6169 = n6168 ^ x24;
  assign n6170 = n6169 ^ x66;
  assign n6171 = x64 & n6143;
  assign n6172 = n6171 ^ x23;
  assign n6173 = n6172 ^ x65;
  assign n6174 = ~x22 & x64;
  assign n6175 = n6174 ^ n6172;
  assign n6176 = ~n6173 & n6175;
  assign n6177 = n6176 ^ x65;
  assign n6178 = n6177 ^ n6169;
  assign n6179 = n6170 & ~n6178;
  assign n6180 = n6179 ^ x66;
  assign n6181 = n6180 ^ x67;
  assign n6182 = n5913 ^ x66;
  assign n6183 = n6143 & ~n6182;
  assign n6184 = n6183 ^ n5897;
  assign n6185 = n6184 ^ n6180;
  assign n6186 = n6181 & n6185;
  assign n6187 = n6186 ^ x67;
  assign n6188 = n6187 ^ x68;
  assign n6189 = n5917 & n6143;
  assign n6190 = n6189 ^ n5920;
  assign n6191 = n6190 ^ n6187;
  assign n6192 = n6188 & ~n6191;
  assign n6193 = n6192 ^ x68;
  assign n6194 = n6193 ^ x69;
  assign n6195 = n5924 & n6143;
  assign n6196 = n6195 ^ n5926;
  assign n6197 = n6196 ^ n6193;
  assign n6198 = n6194 & ~n6197;
  assign n6199 = n6198 ^ x69;
  assign n6200 = n6199 ^ x70;
  assign n6201 = n5930 & n6143;
  assign n6202 = n6201 ^ n5932;
  assign n6203 = n6202 ^ n6199;
  assign n6204 = n6200 & ~n6203;
  assign n6205 = n6204 ^ x70;
  assign n6206 = n6155 & n6205;
  assign n6207 = n6153 ^ x72;
  assign n6208 = x71 & n6150;
  assign n6209 = n6208 ^ n6153;
  assign n6210 = n6207 & ~n6209;
  assign n6211 = n6210 ^ x72;
  assign n6212 = ~n6206 & ~n6211;
  assign n6213 = n6212 ^ x73;
  assign n6214 = n5948 & n6143;
  assign n6215 = n6214 ^ n5951;
  assign n6216 = n6215 ^ n6212;
  assign n6217 = ~n6213 & n6216;
  assign n6218 = n6217 ^ x73;
  assign n6219 = n6218 ^ x74;
  assign n6220 = n5955 & n6143;
  assign n6221 = n6220 ^ n5961;
  assign n6222 = n6221 ^ n6218;
  assign n6223 = n6219 & ~n6222;
  assign n6224 = n6223 ^ x74;
  assign n6225 = n6224 ^ x75;
  assign n6226 = n5965 & n6143;
  assign n6227 = n6226 ^ n5967;
  assign n6228 = n6227 ^ n6224;
  assign n6229 = n6225 & ~n6228;
  assign n6230 = n6229 ^ x75;
  assign n6231 = n6230 ^ x76;
  assign n6232 = n5971 & n6143;
  assign n6233 = n6232 ^ n5973;
  assign n6234 = n6233 ^ n6230;
  assign n6235 = n6231 & ~n6234;
  assign n6236 = n6235 ^ x76;
  assign n6237 = n6236 ^ x77;
  assign n6238 = n5977 & n6143;
  assign n6239 = n6238 ^ n5979;
  assign n6240 = n6239 ^ n6236;
  assign n6241 = n6237 & ~n6240;
  assign n6242 = n6241 ^ x77;
  assign n6243 = n6242 ^ x78;
  assign n6244 = n5983 & n6143;
  assign n6245 = n6244 ^ n5985;
  assign n6246 = n6245 ^ n6242;
  assign n6247 = n6243 & ~n6246;
  assign n6248 = n6247 ^ x78;
  assign n6249 = n6248 ^ x79;
  assign n6250 = n5989 & n6143;
  assign n6251 = n6250 ^ n5991;
  assign n6252 = n6251 ^ n6248;
  assign n6253 = n6249 & ~n6252;
  assign n6254 = n6253 ^ x79;
  assign n6255 = n6254 ^ x80;
  assign n6256 = n5995 & n6143;
  assign n6257 = n6256 ^ n5997;
  assign n6258 = n6257 ^ n6254;
  assign n6259 = n6255 & ~n6258;
  assign n6260 = n6259 ^ x80;
  assign n6261 = n6260 ^ x81;
  assign n6262 = n6001 & n6143;
  assign n6263 = n6262 ^ n6003;
  assign n6264 = n6263 ^ n6260;
  assign n6265 = n6261 & ~n6264;
  assign n6266 = n6265 ^ x81;
  assign n6267 = n6266 ^ x82;
  assign n6268 = n6007 & n6143;
  assign n6269 = n6268 ^ n6009;
  assign n6270 = n6269 ^ n6266;
  assign n6271 = n6267 & ~n6270;
  assign n6272 = n6271 ^ x82;
  assign n6273 = n6272 ^ x83;
  assign n6274 = n6013 & n6143;
  assign n6275 = n6274 ^ n6015;
  assign n6276 = n6275 ^ n6272;
  assign n6277 = n6273 & ~n6276;
  assign n6278 = n6277 ^ x83;
  assign n6279 = n6278 ^ x84;
  assign n6280 = n6019 & n6143;
  assign n6281 = n6280 ^ n6021;
  assign n6282 = n6281 ^ n6278;
  assign n6283 = n6279 & ~n6282;
  assign n6284 = n6283 ^ x84;
  assign n6285 = n6284 ^ x85;
  assign n6286 = n6025 & n6143;
  assign n6287 = n6286 ^ n6027;
  assign n6288 = n6287 ^ n6284;
  assign n6289 = n6285 & ~n6288;
  assign n6290 = n6289 ^ x85;
  assign n6291 = n6290 ^ x86;
  assign n6292 = n6031 & n6143;
  assign n6293 = n6292 ^ n6033;
  assign n6294 = n6293 ^ n6290;
  assign n6295 = n6291 & ~n6294;
  assign n6296 = n6295 ^ x86;
  assign n6297 = n6296 ^ x87;
  assign n6298 = n6036 ^ x86;
  assign n6299 = n6143 & n6298;
  assign n6300 = n6299 ^ n5879;
  assign n6301 = n6300 ^ n6296;
  assign n6302 = n6297 & ~n6301;
  assign n6303 = n6302 ^ x87;
  assign n6304 = n6303 ^ x88;
  assign n6305 = n6036 ^ n5879;
  assign n6306 = n6298 & ~n6305;
  assign n6307 = n6306 ^ x86;
  assign n6308 = n6307 ^ x87;
  assign n6309 = n6143 & n6308;
  assign n6310 = n6309 ^ n5882;
  assign n6311 = n6310 ^ n6303;
  assign n6312 = n6304 & ~n6311;
  assign n6313 = n6312 ^ x88;
  assign n6314 = n6313 ^ x89;
  assign n6315 = n6043 ^ x88;
  assign n6316 = n6143 & ~n6315;
  assign n6317 = n6316 ^ n6045;
  assign n6318 = n6317 ^ n6313;
  assign n6319 = n6314 & ~n6318;
  assign n6320 = n6319 ^ x89;
  assign n6321 = n6320 ^ x90;
  assign n6322 = n6045 ^ n6043;
  assign n6323 = ~n6315 & n6322;
  assign n6324 = n6323 ^ x88;
  assign n6325 = n6324 ^ x89;
  assign n6326 = n6143 & n6325;
  assign n6327 = n6326 ^ n6048;
  assign n6328 = n6327 ^ n6320;
  assign n6329 = n6321 & ~n6328;
  assign n6330 = n6329 ^ x90;
  assign n6331 = n6330 ^ x91;
  assign n6332 = ~n6058 & n6143;
  assign n6333 = n6332 ^ n6060;
  assign n6334 = n6333 ^ n6330;
  assign n6335 = n6331 & ~n6334;
  assign n6336 = n6335 ^ x91;
  assign n6337 = n6336 ^ x92;
  assign n6338 = n6064 & n6143;
  assign n6339 = n6338 ^ n6066;
  assign n6340 = n6339 ^ n6336;
  assign n6341 = n6337 & ~n6340;
  assign n6342 = n6341 ^ x92;
  assign n6343 = n6342 ^ x93;
  assign n6344 = n6069 ^ x92;
  assign n6345 = n6143 & n6344;
  assign n6346 = n6345 ^ n5872;
  assign n6347 = n6346 ^ n6342;
  assign n6348 = n6343 & ~n6347;
  assign n6349 = n6348 ^ x93;
  assign n6350 = n6349 ^ x94;
  assign n6351 = n6069 ^ n5872;
  assign n6352 = n6344 & ~n6351;
  assign n6353 = n6352 ^ x92;
  assign n6354 = n6353 ^ x93;
  assign n6355 = n6143 & n6354;
  assign n6356 = n6355 ^ n5875;
  assign n6357 = n6356 ^ n6349;
  assign n6358 = n6350 & ~n6357;
  assign n6359 = n6358 ^ x94;
  assign n6360 = n6359 ^ x95;
  assign n6361 = ~n6077 & n6143;
  assign n6362 = n6361 ^ n6079;
  assign n6363 = n6362 ^ n6359;
  assign n6364 = n6360 & ~n6363;
  assign n6365 = n6364 ^ x95;
  assign n6366 = n6365 ^ x96;
  assign n6367 = n6083 & n6143;
  assign n6368 = n6367 ^ n6085;
  assign n6369 = n6368 ^ n6365;
  assign n6370 = n6366 & ~n6369;
  assign n6371 = n6370 ^ x96;
  assign n6372 = n6371 ^ x97;
  assign n6373 = n6088 ^ x96;
  assign n6374 = n6143 & n6373;
  assign n6375 = n6374 ^ n5869;
  assign n6376 = n6375 ^ n6371;
  assign n6377 = n6372 & ~n6376;
  assign n6378 = n6377 ^ x97;
  assign n6379 = x98 & n6378;
  assign n6380 = ~n6089 & ~n6093;
  assign n6381 = n6380 ^ x97;
  assign n6382 = n6143 & ~n6381;
  assign n6383 = n6382 ^ n6091;
  assign n6384 = x98 & n6383;
  assign n6385 = ~x99 & ~n6384;
  assign n6386 = ~n6379 & n6385;
  assign n6387 = n6098 & n6143;
  assign n6388 = n6387 ^ n6101;
  assign n6389 = ~n6386 & n6388;
  assign n6390 = ~n6378 & ~n6383;
  assign n6391 = x98 & x99;
  assign n6392 = ~n6390 & n6391;
  assign n6393 = ~x99 & ~n6388;
  assign n6394 = n6383 & ~n6393;
  assign n6395 = n6378 & n6394;
  assign n6396 = ~n6392 & ~n6395;
  assign n6397 = ~n6389 & n6396;
  assign n6398 = n6397 ^ x100;
  assign n6399 = n6105 & n6143;
  assign n6400 = n6399 ^ n6109;
  assign n6401 = n6400 ^ n6397;
  assign n6402 = ~n6398 & n6401;
  assign n6403 = n6402 ^ x100;
  assign n6404 = n6403 ^ x101;
  assign n6405 = n6113 & n6143;
  assign n6406 = n6405 ^ n6115;
  assign n6407 = n6406 ^ n6403;
  assign n6408 = n6404 & ~n6407;
  assign n6409 = n6408 ^ x101;
  assign n6410 = n6409 ^ x102;
  assign n6411 = n6119 & n6143;
  assign n6412 = n6411 ^ n6121;
  assign n6413 = n6412 ^ n6409;
  assign n6414 = n6410 & ~n6413;
  assign n6415 = n6414 ^ x102;
  assign n6416 = n6415 ^ x103;
  assign n6417 = n6124 ^ x102;
  assign n6418 = n6143 & n6417;
  assign n6419 = n6418 ^ n5866;
  assign n6420 = n6419 ^ n6415;
  assign n6421 = n6416 & ~n6420;
  assign n6422 = n6421 ^ x103;
  assign n6423 = n6422 ^ x104;
  assign n6424 = ~n6125 & ~n6126;
  assign n6425 = n6424 ^ x103;
  assign n6426 = n6143 & n6425;
  assign n6427 = n6426 ^ n6129;
  assign n6428 = n6427 ^ n6422;
  assign n6429 = n6423 & n6428;
  assign n6430 = n6429 ^ x104;
  assign n6431 = n6148 & ~n6430;
  assign n6432 = n6142 & ~n6145;
  assign n6433 = ~n6431 & ~n6432;
  assign n6434 = n6378 ^ x98;
  assign n6435 = ~n6433 & n6434;
  assign n6436 = n6435 ^ n6383;
  assign n6437 = x99 & n6436;
  assign n6438 = n6383 ^ n6378;
  assign n6439 = n6434 & ~n6438;
  assign n6440 = n6439 ^ x98;
  assign n6441 = n6440 ^ x99;
  assign n6442 = ~n6433 & n6441;
  assign n6443 = n6442 ^ n6388;
  assign n6444 = x100 & n6443;
  assign n6445 = ~n6437 & ~n6444;
  assign n6446 = n6331 & ~n6433;
  assign n6447 = n6446 ^ n6333;
  assign n6448 = ~x92 & ~n6447;
  assign n6449 = n6337 & ~n6433;
  assign n6450 = n6449 ^ n6339;
  assign n6451 = ~x93 & ~n6450;
  assign n6452 = ~n6448 & ~n6451;
  assign n6453 = x64 & ~n6433;
  assign n6454 = x21 & ~x65;
  assign n6455 = x22 & ~n6454;
  assign n6456 = ~n6173 & n6455;
  assign n6457 = n6453 & n6456;
  assign n6458 = ~x66 & ~n6457;
  assign n6459 = ~x21 & x65;
  assign n6460 = ~x22 & n6459;
  assign n6461 = ~n6172 & n6460;
  assign n6462 = ~n6433 & ~n6461;
  assign n6463 = ~x21 & ~x22;
  assign n6464 = ~n6459 & ~n6463;
  assign n6465 = x64 & ~n6464;
  assign n6466 = ~n6172 & n6465;
  assign n6467 = ~n6462 & n6466;
  assign n6468 = n6458 & ~n6467;
  assign n6469 = ~x22 & x65;
  assign n6470 = ~n6453 & n6469;
  assign n6471 = n6433 ^ n6172;
  assign n6472 = n6470 & n6471;
  assign n6473 = n6468 & ~n6472;
  assign n6474 = ~x21 & x64;
  assign n6475 = ~n6433 & n6474;
  assign n6476 = ~n6465 & ~n6469;
  assign n6477 = ~n6475 & n6476;
  assign n6478 = ~x65 & ~n6174;
  assign n6479 = ~n6433 & ~n6478;
  assign n6480 = n6172 & ~n6479;
  assign n6481 = n6477 & n6480;
  assign n6482 = n6174 & ~n6459;
  assign n6483 = ~n6173 & n6482;
  assign n6484 = x22 & n202;
  assign n6485 = ~n6172 & n6484;
  assign n6486 = ~n6483 & ~n6485;
  assign n6487 = ~n6433 & ~n6486;
  assign n6488 = ~n6481 & ~n6487;
  assign n6489 = ~n6473 & n6488;
  assign n6490 = n6489 ^ x67;
  assign n6491 = n6177 ^ x66;
  assign n6492 = ~n6433 & n6491;
  assign n6493 = n6492 ^ n6169;
  assign n6494 = n6493 ^ n6489;
  assign n6495 = n6490 & ~n6494;
  assign n6496 = n6495 ^ x67;
  assign n6497 = n6496 ^ x68;
  assign n6498 = n6181 & ~n6433;
  assign n6499 = n6498 ^ n6184;
  assign n6500 = n6499 ^ n6496;
  assign n6501 = n6497 & n6500;
  assign n6502 = n6501 ^ x68;
  assign n6503 = n6502 ^ x69;
  assign n6504 = n6188 & ~n6433;
  assign n6505 = n6504 ^ n6190;
  assign n6506 = n6505 ^ n6502;
  assign n6507 = n6503 & ~n6506;
  assign n6508 = n6507 ^ x69;
  assign n6509 = n6508 ^ x70;
  assign n6510 = n6194 & ~n6433;
  assign n6511 = n6510 ^ n6196;
  assign n6512 = n6511 ^ n6508;
  assign n6513 = n6509 & ~n6512;
  assign n6514 = n6513 ^ x70;
  assign n6515 = n6514 ^ x71;
  assign n6516 = n6200 & ~n6433;
  assign n6517 = n6516 ^ n6202;
  assign n6518 = n6517 ^ n6514;
  assign n6519 = n6515 & ~n6518;
  assign n6520 = n6519 ^ x71;
  assign n6521 = n6520 ^ x72;
  assign n6522 = n6205 ^ x71;
  assign n6523 = ~n6433 & n6522;
  assign n6524 = n6523 ^ n6150;
  assign n6525 = n6524 ^ n6520;
  assign n6526 = n6521 & ~n6525;
  assign n6527 = n6526 ^ x72;
  assign n6528 = n6527 ^ x73;
  assign n6529 = n6205 ^ n6150;
  assign n6530 = n6522 & ~n6529;
  assign n6531 = n6530 ^ x71;
  assign n6532 = n6531 ^ x72;
  assign n6533 = ~n6433 & n6532;
  assign n6534 = n6533 ^ n6153;
  assign n6535 = n6534 ^ n6527;
  assign n6536 = n6528 & ~n6535;
  assign n6537 = n6536 ^ x73;
  assign n6538 = n6537 ^ x74;
  assign n6539 = ~n6213 & ~n6433;
  assign n6540 = n6539 ^ n6215;
  assign n6541 = n6540 ^ n6537;
  assign n6542 = n6538 & ~n6541;
  assign n6543 = n6542 ^ x74;
  assign n6544 = n6543 ^ x75;
  assign n6545 = n6219 & ~n6433;
  assign n6546 = n6545 ^ n6221;
  assign n6547 = n6546 ^ n6543;
  assign n6548 = n6544 & ~n6547;
  assign n6549 = n6548 ^ x75;
  assign n6550 = n6549 ^ x76;
  assign n6551 = n6225 & ~n6433;
  assign n6552 = n6551 ^ n6227;
  assign n6553 = n6552 ^ n6549;
  assign n6554 = n6550 & ~n6553;
  assign n6555 = n6554 ^ x76;
  assign n6556 = n6555 ^ x77;
  assign n6557 = n6231 & ~n6433;
  assign n6558 = n6557 ^ n6233;
  assign n6559 = n6558 ^ n6555;
  assign n6560 = n6556 & ~n6559;
  assign n6561 = n6560 ^ x77;
  assign n6562 = n6561 ^ x78;
  assign n6563 = n6237 & ~n6433;
  assign n6564 = n6563 ^ n6239;
  assign n6565 = n6564 ^ n6561;
  assign n6566 = n6562 & ~n6565;
  assign n6567 = n6566 ^ x78;
  assign n6568 = n6567 ^ x79;
  assign n6569 = n6243 & ~n6433;
  assign n6570 = n6569 ^ n6245;
  assign n6571 = n6570 ^ n6567;
  assign n6572 = n6568 & ~n6571;
  assign n6573 = n6572 ^ x79;
  assign n6574 = n6573 ^ x80;
  assign n6575 = n6249 & ~n6433;
  assign n6576 = n6575 ^ n6251;
  assign n6577 = n6576 ^ n6573;
  assign n6578 = n6574 & ~n6577;
  assign n6579 = n6578 ^ x80;
  assign n6580 = n6579 ^ x81;
  assign n6581 = n6255 & ~n6433;
  assign n6582 = n6581 ^ n6257;
  assign n6583 = n6582 ^ n6579;
  assign n6584 = n6580 & ~n6583;
  assign n6585 = n6584 ^ x81;
  assign n6586 = n6585 ^ x82;
  assign n6587 = n6261 & ~n6433;
  assign n6588 = n6587 ^ n6263;
  assign n6589 = n6588 ^ n6585;
  assign n6590 = n6586 & ~n6589;
  assign n6591 = n6590 ^ x82;
  assign n6592 = n6591 ^ x83;
  assign n6593 = n6267 & ~n6433;
  assign n6594 = n6593 ^ n6269;
  assign n6595 = n6594 ^ n6591;
  assign n6596 = n6592 & ~n6595;
  assign n6597 = n6596 ^ x83;
  assign n6598 = n6597 ^ x84;
  assign n6599 = n6273 & ~n6433;
  assign n6600 = n6599 ^ n6275;
  assign n6601 = n6600 ^ n6597;
  assign n6602 = n6598 & ~n6601;
  assign n6603 = n6602 ^ x84;
  assign n6604 = n6603 ^ x85;
  assign n6605 = n6279 & ~n6433;
  assign n6606 = n6605 ^ n6281;
  assign n6607 = n6606 ^ n6603;
  assign n6608 = n6604 & ~n6607;
  assign n6609 = n6608 ^ x85;
  assign n6610 = n6609 ^ x86;
  assign n6611 = n6285 & ~n6433;
  assign n6612 = n6611 ^ n6287;
  assign n6613 = n6612 ^ n6609;
  assign n6614 = n6610 & ~n6613;
  assign n6615 = n6614 ^ x86;
  assign n6616 = n6615 ^ x87;
  assign n6617 = n6291 & ~n6433;
  assign n6618 = n6617 ^ n6293;
  assign n6619 = n6618 ^ n6615;
  assign n6620 = n6616 & ~n6619;
  assign n6621 = n6620 ^ x87;
  assign n6622 = n6621 ^ x88;
  assign n6623 = n6297 & ~n6433;
  assign n6624 = n6623 ^ n6300;
  assign n6625 = n6624 ^ n6621;
  assign n6626 = n6622 & ~n6625;
  assign n6627 = n6626 ^ x88;
  assign n6628 = n6627 ^ x89;
  assign n6629 = n6304 & ~n6433;
  assign n6630 = n6629 ^ n6310;
  assign n6631 = n6630 ^ n6627;
  assign n6632 = n6628 & ~n6631;
  assign n6633 = n6632 ^ x89;
  assign n6634 = n6633 ^ x90;
  assign n6635 = n6314 & ~n6433;
  assign n6636 = n6635 ^ n6317;
  assign n6637 = n6636 ^ n6633;
  assign n6638 = n6634 & ~n6637;
  assign n6639 = n6638 ^ x90;
  assign n6640 = n6639 ^ x91;
  assign n6641 = n6321 & ~n6433;
  assign n6642 = n6641 ^ n6327;
  assign n6643 = n6642 ^ n6639;
  assign n6644 = n6640 & ~n6643;
  assign n6645 = n6644 ^ x91;
  assign n6646 = n6452 & n6645;
  assign n6647 = n6450 ^ x93;
  assign n6648 = x92 & n6447;
  assign n6649 = n6648 ^ n6450;
  assign n6650 = n6647 & ~n6649;
  assign n6651 = n6650 ^ x93;
  assign n6652 = ~n6646 & ~n6651;
  assign n6653 = n6343 & ~n6433;
  assign n6654 = n6653 ^ n6346;
  assign n6655 = ~x94 & ~n6654;
  assign n6656 = n6350 & ~n6433;
  assign n6657 = n6656 ^ n6356;
  assign n6658 = ~x95 & ~n6657;
  assign n6659 = ~n6655 & ~n6658;
  assign n6660 = ~n6652 & n6659;
  assign n6661 = n6657 ^ x95;
  assign n6662 = x94 & n6654;
  assign n6663 = n6662 ^ n6657;
  assign n6664 = n6661 & ~n6663;
  assign n6665 = n6664 ^ x95;
  assign n6666 = ~n6660 & ~n6665;
  assign n6667 = n6666 ^ x96;
  assign n6668 = n6360 & ~n6433;
  assign n6669 = n6668 ^ n6362;
  assign n6670 = n6669 ^ n6666;
  assign n6671 = ~n6667 & n6670;
  assign n6672 = n6671 ^ x96;
  assign n6673 = n6672 ^ x97;
  assign n6674 = n6366 & ~n6433;
  assign n6675 = n6674 ^ n6368;
  assign n6676 = n6675 ^ n6672;
  assign n6677 = n6673 & ~n6676;
  assign n6678 = n6677 ^ x97;
  assign n6679 = n6678 ^ x98;
  assign n6680 = n6372 & ~n6433;
  assign n6681 = n6680 ^ n6375;
  assign n6682 = n6681 ^ n6678;
  assign n6683 = n6679 & ~n6682;
  assign n6684 = n6683 ^ x98;
  assign n6685 = n6445 & ~n6684;
  assign n6686 = n6443 ^ x100;
  assign n6687 = ~x99 & ~n6436;
  assign n6688 = n6687 ^ n6443;
  assign n6689 = n6686 & n6688;
  assign n6690 = n6689 ^ x100;
  assign n6691 = ~n6685 & n6690;
  assign n6692 = ~n6398 & ~n6433;
  assign n6693 = n6692 ^ n6400;
  assign n6694 = ~x101 & ~n6693;
  assign n6695 = n6404 & ~n6433;
  assign n6696 = n6695 ^ n6406;
  assign n6697 = ~x102 & ~n6696;
  assign n6698 = ~n6694 & ~n6697;
  assign n6699 = n6691 & n6698;
  assign n6700 = n6696 ^ x102;
  assign n6701 = x101 & n6693;
  assign n6702 = n6701 ^ n6696;
  assign n6703 = n6700 & ~n6702;
  assign n6704 = n6703 ^ x102;
  assign n6705 = ~n6699 & ~n6704;
  assign n6706 = n6705 ^ x103;
  assign n6707 = n6410 & ~n6433;
  assign n6708 = n6707 ^ n6412;
  assign n6709 = n6708 ^ n6705;
  assign n6710 = ~n6706 & n6709;
  assign n6711 = n6710 ^ x103;
  assign n6712 = n6711 ^ x104;
  assign n6713 = n6416 & ~n6433;
  assign n6714 = n6713 ^ n6419;
  assign n6715 = n6714 ^ n6711;
  assign n6716 = n6712 & ~n6715;
  assign n6717 = n6716 ^ x104;
  assign n6718 = ~x105 & ~n6717;
  assign n6719 = n6423 & ~n6433;
  assign n6720 = n6719 ^ n6427;
  assign n6721 = ~x105 & n6720;
  assign n6722 = ~n6430 & ~n6721;
  assign n6723 = ~n6718 & n6722;
  assign n6724 = ~x105 & n6430;
  assign n6725 = ~x106 & ~n6724;
  assign n6726 = ~n6723 & n6725;
  assign n6727 = n6717 ^ x105;
  assign n6728 = n6720 ^ n6717;
  assign n6729 = n6727 & n6728;
  assign n6730 = n6729 ^ x105;
  assign n6731 = n6726 & ~n6730;
  assign n6732 = n6146 & ~n6731;
  assign n6733 = x106 & n6730;
  assign n6734 = n6732 & ~n6733;
  assign n6735 = ~n6145 & ~n6734;
  assign n6736 = x106 & n6145;
  assign n6737 = ~n6730 & ~n6736;
  assign n6738 = n6430 ^ x105;
  assign n6739 = ~x106 & ~n6145;
  assign n6740 = ~n6738 & n6739;
  assign n6741 = ~n6737 & ~n6740;
  assign n6742 = n6146 & ~n6741;
  assign n6743 = n6691 ^ x101;
  assign n6744 = n6742 & n6743;
  assign n6745 = n6744 ^ n6693;
  assign n6746 = x102 & n6745;
  assign n6747 = n6673 & n6742;
  assign n6748 = n6747 ^ n6675;
  assign n6749 = ~x98 & ~n6748;
  assign n6750 = n6679 & n6742;
  assign n6751 = n6750 ^ n6681;
  assign n6752 = ~x99 & ~n6751;
  assign n6753 = ~n6749 & ~n6752;
  assign n6754 = n6574 & n6742;
  assign n6755 = n6754 ^ n6576;
  assign n6756 = ~x81 & ~n6755;
  assign n6757 = n6580 & n6742;
  assign n6758 = n6757 ^ n6582;
  assign n6759 = ~x82 & ~n6758;
  assign n6760 = ~n6756 & ~n6759;
  assign n6761 = n6503 & n6742;
  assign n6762 = n6761 ^ n6505;
  assign n6763 = ~x70 & ~n6762;
  assign n6764 = x64 & n6742;
  assign n6765 = n6764 ^ x21;
  assign n6766 = n6765 ^ x65;
  assign n6767 = ~x20 & x64;
  assign n6768 = n6767 ^ n6765;
  assign n6769 = ~n6766 & n6768;
  assign n6770 = n6769 ^ x65;
  assign n6771 = n6770 ^ x66;
  assign n6772 = ~n6454 & n6742;
  assign n6773 = n6453 & ~n6772;
  assign n6774 = x65 & n6433;
  assign n6775 = x21 & n6774;
  assign n6776 = ~n202 & ~n6775;
  assign n6777 = n6433 ^ x65;
  assign n6778 = n6474 & n6777;
  assign n6779 = n6776 & ~n6778;
  assign n6780 = n6742 & ~n6779;
  assign n6781 = ~n6773 & ~n6780;
  assign n6782 = n6781 ^ x22;
  assign n6783 = n6782 ^ n6770;
  assign n6784 = n6771 & ~n6783;
  assign n6785 = n6784 ^ x66;
  assign n6786 = n6785 ^ x67;
  assign n6790 = ~n6433 & n6455;
  assign n6791 = ~n6459 & ~n6790;
  assign n6792 = n6433 & n6463;
  assign n6793 = n6791 & ~n6792;
  assign n6794 = x64 & ~n6793;
  assign n6795 = ~n6470 & ~n6794;
  assign n6796 = n6795 ^ x66;
  assign n6797 = n6742 & ~n6796;
  assign n6787 = n6174 ^ x65;
  assign n6788 = ~n6433 & n6787;
  assign n6789 = n6788 ^ n6172;
  assign n6798 = n6797 ^ n6789;
  assign n6799 = n6798 ^ n6785;
  assign n6800 = n6786 & n6799;
  assign n6801 = n6800 ^ x67;
  assign n6802 = n6801 ^ x68;
  assign n6803 = n6490 & n6742;
  assign n6804 = n6803 ^ n6493;
  assign n6805 = n6804 ^ n6801;
  assign n6806 = n6802 & ~n6805;
  assign n6807 = n6806 ^ x68;
  assign n6808 = n6807 ^ x69;
  assign n6809 = n6497 & n6742;
  assign n6810 = n6809 ^ n6499;
  assign n6811 = n6810 ^ n6807;
  assign n6812 = n6808 & n6811;
  assign n6813 = n6812 ^ x69;
  assign n6814 = ~n6763 & n6813;
  assign n6815 = n6509 & n6742;
  assign n6816 = n6815 ^ n6511;
  assign n6817 = x71 & n6816;
  assign n6818 = x70 & n6762;
  assign n6819 = ~n6817 & ~n6818;
  assign n6820 = ~n6814 & n6819;
  assign n6821 = ~x71 & ~n6816;
  assign n6822 = ~n6820 & ~n6821;
  assign n6823 = n6822 ^ x72;
  assign n6824 = n6515 & n6742;
  assign n6825 = n6824 ^ n6517;
  assign n6826 = n6825 ^ n6822;
  assign n6827 = n6823 & ~n6826;
  assign n6828 = n6827 ^ x72;
  assign n6829 = n6828 ^ x73;
  assign n6830 = n6521 & n6742;
  assign n6831 = n6830 ^ n6524;
  assign n6832 = n6831 ^ n6828;
  assign n6833 = n6829 & ~n6832;
  assign n6834 = n6833 ^ x73;
  assign n6835 = n6834 ^ x74;
  assign n6836 = n6528 & n6742;
  assign n6837 = n6836 ^ n6534;
  assign n6838 = n6837 ^ n6834;
  assign n6839 = n6835 & ~n6838;
  assign n6840 = n6839 ^ x74;
  assign n6841 = n6840 ^ x75;
  assign n6842 = n6538 & n6742;
  assign n6843 = n6842 ^ n6540;
  assign n6844 = n6843 ^ n6840;
  assign n6845 = n6841 & ~n6844;
  assign n6846 = n6845 ^ x75;
  assign n6847 = n6846 ^ x76;
  assign n6848 = n6544 & n6742;
  assign n6849 = n6848 ^ n6546;
  assign n6850 = n6849 ^ n6846;
  assign n6851 = n6847 & ~n6850;
  assign n6852 = n6851 ^ x76;
  assign n6853 = n6852 ^ x77;
  assign n6854 = n6550 & n6742;
  assign n6855 = n6854 ^ n6552;
  assign n6856 = n6855 ^ n6852;
  assign n6857 = n6853 & ~n6856;
  assign n6858 = n6857 ^ x77;
  assign n6859 = n6858 ^ x78;
  assign n6860 = n6556 & n6742;
  assign n6861 = n6860 ^ n6558;
  assign n6862 = n6861 ^ n6858;
  assign n6863 = n6859 & ~n6862;
  assign n6864 = n6863 ^ x78;
  assign n6865 = n6864 ^ x79;
  assign n6866 = n6562 & n6742;
  assign n6867 = n6866 ^ n6564;
  assign n6868 = n6867 ^ n6864;
  assign n6869 = n6865 & ~n6868;
  assign n6870 = n6869 ^ x79;
  assign n6871 = n6870 ^ x80;
  assign n6872 = n6568 & n6742;
  assign n6873 = n6872 ^ n6570;
  assign n6874 = n6873 ^ n6870;
  assign n6875 = n6871 & ~n6874;
  assign n6876 = n6875 ^ x80;
  assign n6877 = n6760 & n6876;
  assign n6878 = n6758 ^ x82;
  assign n6879 = x81 & n6755;
  assign n6880 = n6879 ^ n6758;
  assign n6881 = n6878 & ~n6880;
  assign n6882 = n6881 ^ x82;
  assign n6883 = ~n6877 & ~n6882;
  assign n6884 = n6883 ^ x83;
  assign n6885 = n6586 & n6742;
  assign n6886 = n6885 ^ n6588;
  assign n6887 = n6886 ^ n6883;
  assign n6888 = ~n6884 & n6887;
  assign n6889 = n6888 ^ x83;
  assign n6890 = n6889 ^ x84;
  assign n6891 = n6592 & n6742;
  assign n6892 = n6891 ^ n6594;
  assign n6893 = n6892 ^ n6889;
  assign n6894 = n6890 & ~n6893;
  assign n6895 = n6894 ^ x84;
  assign n6896 = n6895 ^ x85;
  assign n6897 = n6598 & n6742;
  assign n6898 = n6897 ^ n6600;
  assign n6899 = n6898 ^ n6895;
  assign n6900 = n6896 & ~n6899;
  assign n6901 = n6900 ^ x85;
  assign n6902 = n6901 ^ x86;
  assign n6903 = n6604 & n6742;
  assign n6904 = n6903 ^ n6606;
  assign n6905 = n6904 ^ n6901;
  assign n6906 = n6902 & ~n6905;
  assign n6907 = n6906 ^ x86;
  assign n6908 = n6907 ^ x87;
  assign n6909 = n6610 & n6742;
  assign n6910 = n6909 ^ n6612;
  assign n6911 = n6910 ^ n6907;
  assign n6912 = n6908 & ~n6911;
  assign n6913 = n6912 ^ x87;
  assign n6914 = n6913 ^ x88;
  assign n6915 = n6616 & n6742;
  assign n6916 = n6915 ^ n6618;
  assign n6917 = n6916 ^ n6913;
  assign n6918 = n6914 & ~n6917;
  assign n6919 = n6918 ^ x88;
  assign n6920 = n6919 ^ x89;
  assign n6921 = n6622 & n6742;
  assign n6922 = n6921 ^ n6624;
  assign n6923 = n6922 ^ n6919;
  assign n6924 = n6920 & ~n6923;
  assign n6925 = n6924 ^ x89;
  assign n6926 = n6925 ^ x90;
  assign n6927 = n6628 & n6742;
  assign n6928 = n6927 ^ n6630;
  assign n6929 = n6928 ^ n6925;
  assign n6930 = n6926 & ~n6929;
  assign n6931 = n6930 ^ x90;
  assign n6932 = n6931 ^ x91;
  assign n6933 = n6634 & n6742;
  assign n6934 = n6933 ^ n6636;
  assign n6935 = n6934 ^ n6931;
  assign n6936 = n6932 & ~n6935;
  assign n6937 = n6936 ^ x91;
  assign n6938 = n6937 ^ x92;
  assign n6939 = n6640 & n6742;
  assign n6940 = n6939 ^ n6642;
  assign n6941 = n6940 ^ n6937;
  assign n6942 = n6938 & ~n6941;
  assign n6943 = n6942 ^ x92;
  assign n6944 = n6943 ^ x93;
  assign n6945 = n6645 ^ x92;
  assign n6946 = n6742 & n6945;
  assign n6947 = n6946 ^ n6447;
  assign n6948 = n6947 ^ n6943;
  assign n6949 = n6944 & ~n6948;
  assign n6950 = n6949 ^ x93;
  assign n6951 = n6950 ^ x94;
  assign n6952 = n6645 ^ n6447;
  assign n6953 = n6945 & ~n6952;
  assign n6954 = n6953 ^ x92;
  assign n6955 = n6954 ^ x93;
  assign n6956 = n6742 & n6955;
  assign n6957 = n6956 ^ n6450;
  assign n6958 = n6957 ^ n6950;
  assign n6959 = n6951 & ~n6958;
  assign n6960 = n6959 ^ x94;
  assign n6961 = n6960 ^ x95;
  assign n6962 = n6652 ^ x94;
  assign n6963 = n6742 & ~n6962;
  assign n6964 = n6963 ^ n6654;
  assign n6965 = n6964 ^ n6960;
  assign n6966 = n6961 & ~n6965;
  assign n6967 = n6966 ^ x95;
  assign n6968 = n6967 ^ x96;
  assign n6969 = n6654 ^ n6652;
  assign n6970 = ~n6962 & n6969;
  assign n6971 = n6970 ^ x94;
  assign n6972 = n6971 ^ x95;
  assign n6973 = n6742 & n6972;
  assign n6974 = n6973 ^ n6657;
  assign n6975 = n6974 ^ n6967;
  assign n6976 = n6968 & ~n6975;
  assign n6977 = n6976 ^ x96;
  assign n6978 = n6977 ^ x97;
  assign n6979 = ~n6667 & n6742;
  assign n6980 = n6979 ^ n6669;
  assign n6981 = n6980 ^ n6977;
  assign n6982 = n6978 & ~n6981;
  assign n6983 = n6982 ^ x97;
  assign n6984 = n6753 & n6983;
  assign n6985 = n6751 ^ x99;
  assign n6986 = x98 & n6748;
  assign n6987 = n6986 ^ n6751;
  assign n6988 = n6985 & ~n6987;
  assign n6989 = n6988 ^ x99;
  assign n6990 = ~n6984 & ~n6989;
  assign n6991 = n6990 ^ x100;
  assign n6992 = n6684 ^ x99;
  assign n6993 = n6742 & n6992;
  assign n6994 = n6993 ^ n6436;
  assign n6995 = n6994 ^ n6990;
  assign n6996 = ~n6991 & n6995;
  assign n6997 = n6996 ^ x100;
  assign n6998 = n6997 ^ x101;
  assign n6999 = n6684 ^ n6436;
  assign n7000 = n6992 & ~n6999;
  assign n7001 = n7000 ^ x99;
  assign n7002 = n7001 ^ x100;
  assign n7003 = n6742 & n7002;
  assign n7004 = n7003 ^ n6443;
  assign n7005 = n7004 ^ n6997;
  assign n7006 = n6998 & ~n7005;
  assign n7007 = n7006 ^ x101;
  assign n7008 = ~n6746 & ~n7007;
  assign n7009 = n6693 ^ n6691;
  assign n7010 = n6743 & ~n7009;
  assign n7011 = n7010 ^ x101;
  assign n7012 = n7011 ^ x102;
  assign n7013 = n6742 & n7012;
  assign n7014 = n7013 ^ n6696;
  assign n7015 = ~x103 & ~n7014;
  assign n7016 = ~x102 & ~n6745;
  assign n7017 = ~n7015 & ~n7016;
  assign n7018 = ~n7008 & n7017;
  assign n7019 = x103 & n7014;
  assign n7020 = ~n7018 & ~n7019;
  assign n7021 = ~n6706 & n6742;
  assign n7022 = n7021 ^ n6708;
  assign n7023 = ~x104 & ~n7022;
  assign n7024 = ~n7020 & ~n7023;
  assign n7025 = n6712 & n6742;
  assign n7026 = n7025 ^ n6714;
  assign n7027 = x104 & x105;
  assign n7028 = ~n7026 & ~n7027;
  assign n7029 = n7024 & ~n7028;
  assign n7030 = x105 & n7022;
  assign n7031 = ~n7020 & n7030;
  assign n7032 = n7026 ^ x105;
  assign n7033 = x104 & n7022;
  assign n7034 = n7033 ^ n7026;
  assign n7035 = n7032 & ~n7034;
  assign n7036 = n7035 ^ x105;
  assign n7037 = ~n7031 & ~n7036;
  assign n7038 = ~n7029 & n7037;
  assign n7039 = n7038 ^ x106;
  assign n7040 = ~x107 & n6735;
  assign n7041 = n6727 & n6742;
  assign n7042 = n7041 ^ n6720;
  assign n7043 = n7042 ^ n7038;
  assign n7044 = ~n7039 & ~n7043;
  assign n7045 = n7044 ^ x106;
  assign n7046 = ~n7040 & n7045;
  assign n7047 = x107 & n6145;
  assign n7048 = n6140 & ~n7047;
  assign n7049 = ~n7046 & n7048;
  assign n7050 = ~n7039 & n7049;
  assign n7051 = n7050 ^ n7042;
  assign n7052 = x107 & ~n7051;
  assign n7053 = ~x65 & n7049;
  assign n7054 = x20 & ~x65;
  assign n7055 = ~x19 & ~n7054;
  assign n7056 = ~n7053 & n7055;
  assign n7057 = ~n6765 & n7056;
  assign n7058 = x20 & n7049;
  assign n7059 = ~n7057 & ~n7058;
  assign n7060 = x19 & ~x65;
  assign n7061 = n7058 & ~n7060;
  assign n7062 = ~n6766 & n7061;
  assign n7063 = n7062 ^ n7058;
  assign n7064 = x64 & ~n7063;
  assign n7065 = ~n7059 & n7064;
  assign n7066 = x64 & n7049;
  assign n7067 = ~x20 & x65;
  assign n7068 = ~n7066 & n7067;
  assign n7069 = n7049 ^ n6765;
  assign n7070 = n7068 & ~n7069;
  assign n7071 = ~x66 & ~n7070;
  assign n7072 = ~n7065 & n7071;
  assign n7073 = ~x19 & x64;
  assign n7074 = ~n7054 & n7073;
  assign n7075 = ~n7049 & ~n7074;
  assign n7076 = ~x65 & ~n6767;
  assign n7077 = ~n7073 & n7076;
  assign n7078 = ~n7075 & ~n7077;
  assign n7079 = n6765 & ~n7067;
  assign n7080 = ~n7078 & n7079;
  assign n7081 = ~x21 & n202;
  assign n7082 = n7058 & n7081;
  assign n7083 = ~x19 & x65;
  assign n7084 = n6767 & ~n7083;
  assign n7085 = ~n6766 & n7084;
  assign n7086 = n7049 & n7085;
  assign n7087 = ~n7082 & ~n7086;
  assign n7088 = ~n7080 & n7087;
  assign n7089 = ~n7072 & n7088;
  assign n7090 = n7089 ^ x67;
  assign n7091 = n6771 & n7049;
  assign n7092 = n7091 ^ n6782;
  assign n7093 = n7092 ^ n7089;
  assign n7094 = n7090 & ~n7093;
  assign n7095 = n7094 ^ x67;
  assign n7096 = n7095 ^ x68;
  assign n7097 = n6786 & n7049;
  assign n7098 = n7097 ^ n6798;
  assign n7099 = n7098 ^ n7095;
  assign n7100 = n7096 & n7099;
  assign n7101 = n7100 ^ x68;
  assign n7102 = n7101 ^ x69;
  assign n7103 = n6802 & n7049;
  assign n7104 = n7103 ^ n6804;
  assign n7105 = n7104 ^ n7101;
  assign n7106 = n7102 & ~n7105;
  assign n7107 = n7106 ^ x69;
  assign n7108 = n7107 ^ x70;
  assign n7109 = n6808 & n7049;
  assign n7110 = n7109 ^ n6810;
  assign n7111 = n7110 ^ n7107;
  assign n7112 = n7108 & n7111;
  assign n7113 = n7112 ^ x70;
  assign n7114 = n7113 ^ x71;
  assign n7115 = n6813 ^ x70;
  assign n7116 = n7049 & n7115;
  assign n7117 = n7116 ^ n6762;
  assign n7118 = n7117 ^ n7113;
  assign n7119 = n7114 & ~n7118;
  assign n7120 = n7119 ^ x71;
  assign n7121 = n7120 ^ x72;
  assign n7122 = ~n6814 & ~n6818;
  assign n7123 = n7122 ^ x71;
  assign n7124 = n7049 & ~n7123;
  assign n7125 = n7124 ^ n6816;
  assign n7126 = n7125 ^ n7120;
  assign n7127 = n7121 & ~n7126;
  assign n7128 = n7127 ^ x72;
  assign n7129 = n7128 ^ x73;
  assign n7130 = n6823 & n7049;
  assign n7131 = n7130 ^ n6825;
  assign n7132 = n7131 ^ n7128;
  assign n7133 = n7129 & ~n7132;
  assign n7134 = n7133 ^ x73;
  assign n7135 = n7134 ^ x74;
  assign n7136 = n6829 & n7049;
  assign n7137 = n7136 ^ n6831;
  assign n7138 = n7137 ^ n7134;
  assign n7139 = n7135 & ~n7138;
  assign n7140 = n7139 ^ x74;
  assign n7141 = n7140 ^ x75;
  assign n7142 = n6835 & n7049;
  assign n7143 = n7142 ^ n6837;
  assign n7144 = n7143 ^ n7140;
  assign n7145 = n7141 & ~n7144;
  assign n7146 = n7145 ^ x75;
  assign n7147 = n7146 ^ x76;
  assign n7148 = n6841 & n7049;
  assign n7149 = n7148 ^ n6843;
  assign n7150 = n7149 ^ n7146;
  assign n7151 = n7147 & ~n7150;
  assign n7152 = n7151 ^ x76;
  assign n7153 = n7152 ^ x77;
  assign n7154 = n6847 & n7049;
  assign n7155 = n7154 ^ n6849;
  assign n7156 = n7155 ^ n7152;
  assign n7157 = n7153 & ~n7156;
  assign n7158 = n7157 ^ x77;
  assign n7159 = n7158 ^ x78;
  assign n7160 = n6853 & n7049;
  assign n7161 = n7160 ^ n6855;
  assign n7162 = n7161 ^ n7158;
  assign n7163 = n7159 & ~n7162;
  assign n7164 = n7163 ^ x78;
  assign n7165 = n7164 ^ x79;
  assign n7166 = n6859 & n7049;
  assign n7167 = n7166 ^ n6861;
  assign n7168 = n7167 ^ n7164;
  assign n7169 = n7165 & ~n7168;
  assign n7170 = n7169 ^ x79;
  assign n7171 = n7170 ^ x80;
  assign n7172 = n6865 & n7049;
  assign n7173 = n7172 ^ n6867;
  assign n7174 = n7173 ^ n7170;
  assign n7175 = n7171 & ~n7174;
  assign n7176 = n7175 ^ x80;
  assign n7177 = n7176 ^ x81;
  assign n7178 = n6871 & n7049;
  assign n7179 = n7178 ^ n6873;
  assign n7180 = n7179 ^ n7176;
  assign n7181 = n7177 & ~n7180;
  assign n7182 = n7181 ^ x81;
  assign n7183 = n7182 ^ x82;
  assign n7184 = n6876 ^ x81;
  assign n7185 = n7049 & n7184;
  assign n7186 = n7185 ^ n6755;
  assign n7187 = n7186 ^ n7182;
  assign n7188 = n7183 & ~n7187;
  assign n7189 = n7188 ^ x82;
  assign n7190 = n7189 ^ x83;
  assign n7191 = n6876 ^ n6755;
  assign n7192 = n7184 & ~n7191;
  assign n7193 = n7192 ^ x81;
  assign n7194 = n7193 ^ x82;
  assign n7195 = n7049 & n7194;
  assign n7196 = n7195 ^ n6758;
  assign n7197 = n7196 ^ n7189;
  assign n7198 = n7190 & ~n7197;
  assign n7199 = n7198 ^ x83;
  assign n7200 = n7199 ^ x84;
  assign n7201 = ~n6884 & n7049;
  assign n7202 = n7201 ^ n6886;
  assign n7203 = n7202 ^ n7199;
  assign n7204 = n7200 & ~n7203;
  assign n7205 = n7204 ^ x84;
  assign n7206 = n7205 ^ x85;
  assign n7207 = n6890 & n7049;
  assign n7208 = n7207 ^ n6892;
  assign n7209 = n7208 ^ n7205;
  assign n7210 = n7206 & ~n7209;
  assign n7211 = n7210 ^ x85;
  assign n7212 = n7211 ^ x86;
  assign n7213 = n6896 & n7049;
  assign n7214 = n7213 ^ n6898;
  assign n7215 = n7214 ^ n7211;
  assign n7216 = n7212 & ~n7215;
  assign n7217 = n7216 ^ x86;
  assign n7218 = n7217 ^ x87;
  assign n7219 = n6902 & n7049;
  assign n7220 = n7219 ^ n6904;
  assign n7221 = n7220 ^ n7217;
  assign n7222 = n7218 & ~n7221;
  assign n7223 = n7222 ^ x87;
  assign n7224 = n7223 ^ x88;
  assign n7225 = n6908 & n7049;
  assign n7226 = n7225 ^ n6910;
  assign n7227 = n7226 ^ n7223;
  assign n7228 = n7224 & ~n7227;
  assign n7229 = n7228 ^ x88;
  assign n7230 = n7229 ^ x89;
  assign n7231 = n6914 & n7049;
  assign n7232 = n7231 ^ n6916;
  assign n7233 = n7232 ^ n7229;
  assign n7234 = n7230 & ~n7233;
  assign n7235 = n7234 ^ x89;
  assign n7236 = n7235 ^ x90;
  assign n7237 = n6920 & n7049;
  assign n7238 = n7237 ^ n6922;
  assign n7239 = n7238 ^ n7235;
  assign n7240 = n7236 & ~n7239;
  assign n7241 = n7240 ^ x90;
  assign n7242 = n7241 ^ x91;
  assign n7243 = n6926 & n7049;
  assign n7244 = n7243 ^ n6928;
  assign n7245 = n7244 ^ n7241;
  assign n7246 = n7242 & ~n7245;
  assign n7247 = n7246 ^ x91;
  assign n7248 = n7247 ^ x92;
  assign n7249 = n6932 & n7049;
  assign n7250 = n7249 ^ n6934;
  assign n7251 = n7250 ^ n7247;
  assign n7252 = n7248 & ~n7251;
  assign n7253 = n7252 ^ x92;
  assign n7254 = n7253 ^ x93;
  assign n7255 = n6938 & n7049;
  assign n7256 = n7255 ^ n6940;
  assign n7257 = n7256 ^ n7253;
  assign n7258 = n7254 & ~n7257;
  assign n7259 = n7258 ^ x93;
  assign n7260 = n7259 ^ x94;
  assign n7261 = n6944 & n7049;
  assign n7262 = n7261 ^ n6947;
  assign n7263 = n7262 ^ n7259;
  assign n7264 = n7260 & ~n7263;
  assign n7265 = n7264 ^ x94;
  assign n7266 = n7265 ^ x95;
  assign n7267 = n6951 & n7049;
  assign n7268 = n7267 ^ n6957;
  assign n7269 = n7268 ^ n7265;
  assign n7270 = n7266 & ~n7269;
  assign n7271 = n7270 ^ x95;
  assign n7272 = n7271 ^ x96;
  assign n7273 = n6961 & n7049;
  assign n7274 = n7273 ^ n6964;
  assign n7275 = n7274 ^ n7271;
  assign n7276 = n7272 & ~n7275;
  assign n7277 = n7276 ^ x96;
  assign n7278 = n7277 ^ x97;
  assign n7279 = n6968 & n7049;
  assign n7280 = n7279 ^ n6974;
  assign n7281 = n7280 ^ n7277;
  assign n7282 = n7278 & ~n7281;
  assign n7283 = n7282 ^ x97;
  assign n7284 = n7283 ^ x98;
  assign n7285 = n6978 & n7049;
  assign n7286 = n7285 ^ n6980;
  assign n7287 = n7286 ^ n7283;
  assign n7288 = n7284 & ~n7287;
  assign n7289 = n7288 ^ x98;
  assign n7290 = n7289 ^ x99;
  assign n7291 = n6983 ^ x98;
  assign n7292 = n7049 & n7291;
  assign n7293 = n7292 ^ n6748;
  assign n7294 = n7293 ^ n7289;
  assign n7295 = n7290 & ~n7294;
  assign n7296 = n7295 ^ x99;
  assign n7297 = n7296 ^ x100;
  assign n7298 = n6983 ^ n6748;
  assign n7299 = n7291 & ~n7298;
  assign n7300 = n7299 ^ x98;
  assign n7301 = n7300 ^ x99;
  assign n7302 = n7049 & n7301;
  assign n7303 = n7302 ^ n6751;
  assign n7304 = n7303 ^ n7296;
  assign n7305 = n7297 & ~n7304;
  assign n7306 = n7305 ^ x100;
  assign n7307 = n7306 ^ x101;
  assign n7308 = ~n6991 & n7049;
  assign n7309 = n7308 ^ n6994;
  assign n7310 = n7309 ^ n7306;
  assign n7311 = n7307 & ~n7310;
  assign n7312 = n7311 ^ x101;
  assign n7313 = n7312 ^ x102;
  assign n7314 = n6998 & n7049;
  assign n7315 = n7314 ^ n7004;
  assign n7316 = n7315 ^ n7312;
  assign n7317 = n7313 & ~n7316;
  assign n7318 = n7317 ^ x102;
  assign n7319 = n7318 ^ x103;
  assign n7320 = n7007 ^ x102;
  assign n7321 = n7049 & n7320;
  assign n7322 = n7321 ^ n6745;
  assign n7323 = n7322 ^ n7318;
  assign n7324 = n7319 & ~n7323;
  assign n7325 = n7324 ^ x103;
  assign n7326 = n7325 ^ x104;
  assign n7327 = ~n7008 & ~n7016;
  assign n7328 = n7327 ^ x103;
  assign n7329 = n7049 & n7328;
  assign n7330 = n7329 ^ n7014;
  assign n7331 = n7330 ^ n7325;
  assign n7332 = n7326 & ~n7331;
  assign n7333 = n7332 ^ x104;
  assign n7334 = n7333 ^ x105;
  assign n7335 = n7020 ^ x104;
  assign n7336 = n7049 & ~n7335;
  assign n7337 = n7336 ^ n7022;
  assign n7338 = n7337 ^ n7333;
  assign n7339 = n7334 & ~n7338;
  assign n7340 = n7339 ^ x105;
  assign n7341 = n7340 ^ x106;
  assign n7342 = ~n7024 & ~n7033;
  assign n7343 = n7342 ^ x105;
  assign n7344 = n7049 & ~n7343;
  assign n7345 = n7344 ^ n7026;
  assign n7346 = n7345 ^ n7340;
  assign n7347 = n7341 & ~n7346;
  assign n7348 = n7347 ^ x106;
  assign n7349 = ~n7052 & ~n7348;
  assign n7350 = ~x107 & n7051;
  assign n7351 = ~n7349 & ~n7350;
  assign n7352 = n7045 ^ x107;
  assign n7353 = ~x108 & ~n7352;
  assign n7354 = n7353 ^ x108;
  assign n7355 = ~n7351 & n7354;
  assign n7356 = n7355 ^ x108;
  assign n7357 = n147 & ~n7356;
  assign n7358 = n6735 & ~n7357;
  assign n7359 = ~n6734 & n7353;
  assign n7360 = ~n7350 & ~n7359;
  assign n7361 = ~n7349 & n7360;
  assign n7362 = n147 & ~n6145;
  assign n7363 = ~n7361 & n7362;
  assign n7364 = n6140 & ~n7351;
  assign n7365 = ~n7363 & ~n7364;
  assign n7366 = n7334 & ~n7365;
  assign n7367 = n7366 ^ n7337;
  assign n7368 = ~x106 & ~n7367;
  assign n7369 = n7341 & ~n7365;
  assign n7370 = n7369 ^ n7345;
  assign n7371 = ~x107 & ~n7370;
  assign n7372 = ~n7368 & ~n7371;
  assign n7373 = n7272 & ~n7365;
  assign n7374 = n7373 ^ n7274;
  assign n7375 = x97 & n7374;
  assign n7376 = n7278 & ~n7365;
  assign n7377 = n7376 ^ n7280;
  assign n7378 = x98 & n7377;
  assign n7379 = ~n7375 & ~n7378;
  assign n7380 = n7165 & ~n7365;
  assign n7381 = n7380 ^ n7167;
  assign n7382 = x80 & n7381;
  assign n7383 = n7171 & ~n7365;
  assign n7384 = n7383 ^ n7173;
  assign n7385 = x81 & n7384;
  assign n7386 = ~n7382 & ~n7385;
  assign n7387 = x65 & ~n7049;
  assign n7388 = ~n7365 & n7387;
  assign n7389 = ~x65 & n7066;
  assign n7390 = ~n7388 & ~n7389;
  assign n7391 = x19 & ~n7390;
  assign n7392 = n7049 ^ x65;
  assign n7393 = n341 & ~n7392;
  assign n7394 = x19 & n7393;
  assign n7395 = n7394 ^ n340;
  assign n7396 = ~n7365 & n7395;
  assign n7397 = n7396 ^ n7066;
  assign n7398 = ~n7391 & ~n7397;
  assign n7399 = n7398 ^ x20;
  assign n7400 = n7399 ^ x66;
  assign n7401 = x64 & ~n7365;
  assign n7402 = x18 & n7060;
  assign n7403 = n7402 ^ x19;
  assign n7404 = n7401 & n7403;
  assign n7405 = ~x18 & n7073;
  assign n7406 = ~n7083 & ~n7405;
  assign n7407 = n7365 & ~n7406;
  assign n7408 = ~x18 & x65;
  assign n7409 = n7408 ^ n7083;
  assign n7410 = x64 & n7409;
  assign n7411 = n7410 ^ n7083;
  assign n7412 = ~n7407 & ~n7411;
  assign n7413 = ~n7404 & n7412;
  assign n7414 = n7413 ^ n7399;
  assign n7415 = n7400 & n7414;
  assign n7416 = n7415 ^ x66;
  assign n7417 = n7416 ^ x67;
  assign n7421 = ~n7056 & ~n7061;
  assign n7422 = x64 & ~n7421;
  assign n7423 = ~n7068 & ~n7422;
  assign n7424 = n7423 ^ x66;
  assign n7425 = ~n7365 & ~n7424;
  assign n7418 = n6767 ^ x65;
  assign n7419 = n7049 & n7418;
  assign n7420 = n7419 ^ n6765;
  assign n7426 = n7425 ^ n7420;
  assign n7427 = n7426 ^ n7416;
  assign n7428 = n7417 & n7427;
  assign n7429 = n7428 ^ x67;
  assign n7430 = n7429 ^ x68;
  assign n7431 = n7090 & ~n7365;
  assign n7432 = n7431 ^ n7092;
  assign n7433 = n7432 ^ n7429;
  assign n7434 = n7430 & ~n7433;
  assign n7435 = n7434 ^ x68;
  assign n7436 = n7435 ^ x69;
  assign n7437 = n7096 & ~n7365;
  assign n7438 = n7437 ^ n7098;
  assign n7439 = n7438 ^ n7435;
  assign n7440 = n7436 & n7439;
  assign n7441 = n7440 ^ x69;
  assign n7442 = n7441 ^ x70;
  assign n7443 = n7102 & ~n7365;
  assign n7444 = n7443 ^ n7104;
  assign n7445 = n7444 ^ n7441;
  assign n7446 = n7442 & ~n7445;
  assign n7447 = n7446 ^ x70;
  assign n7448 = n7447 ^ x71;
  assign n7449 = n7108 & ~n7365;
  assign n7450 = n7449 ^ n7110;
  assign n7451 = n7450 ^ n7447;
  assign n7452 = n7448 & n7451;
  assign n7453 = n7452 ^ x71;
  assign n7454 = n7453 ^ x72;
  assign n7455 = n7114 & ~n7365;
  assign n7456 = n7455 ^ n7117;
  assign n7457 = n7456 ^ n7453;
  assign n7458 = n7454 & ~n7457;
  assign n7459 = n7458 ^ x72;
  assign n7460 = n7459 ^ x73;
  assign n7461 = n7121 & ~n7365;
  assign n7462 = n7461 ^ n7125;
  assign n7463 = n7462 ^ n7459;
  assign n7464 = n7460 & ~n7463;
  assign n7465 = n7464 ^ x73;
  assign n7466 = n7465 ^ x74;
  assign n7467 = n7129 & ~n7365;
  assign n7468 = n7467 ^ n7131;
  assign n7469 = n7468 ^ n7465;
  assign n7470 = n7466 & ~n7469;
  assign n7471 = n7470 ^ x74;
  assign n7472 = n7471 ^ x75;
  assign n7473 = n7135 & ~n7365;
  assign n7474 = n7473 ^ n7137;
  assign n7475 = n7474 ^ n7471;
  assign n7476 = n7472 & ~n7475;
  assign n7477 = n7476 ^ x75;
  assign n7478 = n7477 ^ x76;
  assign n7479 = n7141 & ~n7365;
  assign n7480 = n7479 ^ n7143;
  assign n7481 = n7480 ^ n7477;
  assign n7482 = n7478 & ~n7481;
  assign n7483 = n7482 ^ x76;
  assign n7484 = n7483 ^ x77;
  assign n7485 = n7147 & ~n7365;
  assign n7486 = n7485 ^ n7149;
  assign n7487 = n7486 ^ n7483;
  assign n7488 = n7484 & ~n7487;
  assign n7489 = n7488 ^ x77;
  assign n7490 = n7489 ^ x78;
  assign n7491 = n7153 & ~n7365;
  assign n7492 = n7491 ^ n7155;
  assign n7493 = n7492 ^ n7489;
  assign n7494 = n7490 & ~n7493;
  assign n7495 = n7494 ^ x78;
  assign n7496 = n7495 ^ x79;
  assign n7497 = n7159 & ~n7365;
  assign n7498 = n7497 ^ n7161;
  assign n7499 = n7498 ^ n7495;
  assign n7500 = n7496 & ~n7499;
  assign n7501 = n7500 ^ x79;
  assign n7502 = n7386 & ~n7501;
  assign n7503 = n7384 ^ x81;
  assign n7504 = ~x80 & ~n7381;
  assign n7505 = n7504 ^ n7384;
  assign n7506 = n7503 & n7505;
  assign n7507 = n7506 ^ x81;
  assign n7508 = ~n7502 & n7507;
  assign n7509 = n7508 ^ x82;
  assign n7510 = n7177 & ~n7365;
  assign n7511 = n7510 ^ n7179;
  assign n7512 = n7511 ^ n7508;
  assign n7513 = n7509 & ~n7512;
  assign n7514 = n7513 ^ x82;
  assign n7515 = n7514 ^ x83;
  assign n7516 = n7183 & ~n7365;
  assign n7517 = n7516 ^ n7186;
  assign n7518 = n7517 ^ n7514;
  assign n7519 = n7515 & ~n7518;
  assign n7520 = n7519 ^ x83;
  assign n7521 = n7520 ^ x84;
  assign n7522 = n7190 & ~n7365;
  assign n7523 = n7522 ^ n7196;
  assign n7524 = n7523 ^ n7520;
  assign n7525 = n7521 & ~n7524;
  assign n7526 = n7525 ^ x84;
  assign n7527 = n7526 ^ x85;
  assign n7528 = n7200 & ~n7365;
  assign n7529 = n7528 ^ n7202;
  assign n7530 = n7529 ^ n7526;
  assign n7531 = n7527 & ~n7530;
  assign n7532 = n7531 ^ x85;
  assign n7533 = n7532 ^ x86;
  assign n7534 = n7206 & ~n7365;
  assign n7535 = n7534 ^ n7208;
  assign n7536 = n7535 ^ n7532;
  assign n7537 = n7533 & ~n7536;
  assign n7538 = n7537 ^ x86;
  assign n7539 = n7538 ^ x87;
  assign n7540 = n7212 & ~n7365;
  assign n7541 = n7540 ^ n7214;
  assign n7542 = n7541 ^ n7538;
  assign n7543 = n7539 & ~n7542;
  assign n7544 = n7543 ^ x87;
  assign n7545 = n7544 ^ x88;
  assign n7546 = n7218 & ~n7365;
  assign n7547 = n7546 ^ n7220;
  assign n7548 = n7547 ^ n7544;
  assign n7549 = n7545 & ~n7548;
  assign n7550 = n7549 ^ x88;
  assign n7551 = n7550 ^ x89;
  assign n7552 = n7224 & ~n7365;
  assign n7553 = n7552 ^ n7226;
  assign n7554 = n7553 ^ n7550;
  assign n7555 = n7551 & ~n7554;
  assign n7556 = n7555 ^ x89;
  assign n7557 = n7556 ^ x90;
  assign n7558 = n7230 & ~n7365;
  assign n7559 = n7558 ^ n7232;
  assign n7560 = n7559 ^ n7556;
  assign n7561 = n7557 & ~n7560;
  assign n7562 = n7561 ^ x90;
  assign n7563 = n7562 ^ x91;
  assign n7564 = n7236 & ~n7365;
  assign n7565 = n7564 ^ n7238;
  assign n7566 = n7565 ^ n7562;
  assign n7567 = n7563 & ~n7566;
  assign n7568 = n7567 ^ x91;
  assign n7569 = n7568 ^ x92;
  assign n7570 = n7242 & ~n7365;
  assign n7571 = n7570 ^ n7244;
  assign n7572 = n7571 ^ n7568;
  assign n7573 = n7569 & ~n7572;
  assign n7574 = n7573 ^ x92;
  assign n7575 = n7574 ^ x93;
  assign n7576 = n7248 & ~n7365;
  assign n7577 = n7576 ^ n7250;
  assign n7578 = n7577 ^ n7574;
  assign n7579 = n7575 & ~n7578;
  assign n7580 = n7579 ^ x93;
  assign n7581 = n7580 ^ x94;
  assign n7582 = n7254 & ~n7365;
  assign n7583 = n7582 ^ n7256;
  assign n7584 = n7583 ^ n7580;
  assign n7585 = n7581 & ~n7584;
  assign n7586 = n7585 ^ x94;
  assign n7587 = n7586 ^ x95;
  assign n7588 = n7260 & ~n7365;
  assign n7589 = n7588 ^ n7262;
  assign n7590 = n7589 ^ n7586;
  assign n7591 = n7587 & ~n7590;
  assign n7592 = n7591 ^ x95;
  assign n7593 = n7592 ^ x96;
  assign n7594 = n7266 & ~n7365;
  assign n7595 = n7594 ^ n7268;
  assign n7596 = n7595 ^ n7592;
  assign n7597 = n7593 & ~n7596;
  assign n7598 = n7597 ^ x96;
  assign n7599 = n7379 & ~n7598;
  assign n7600 = n7377 ^ x98;
  assign n7601 = ~x97 & ~n7374;
  assign n7602 = n7601 ^ n7377;
  assign n7603 = n7600 & n7602;
  assign n7604 = n7603 ^ x98;
  assign n7605 = ~n7599 & n7604;
  assign n7606 = n7284 & ~n7365;
  assign n7607 = n7606 ^ n7286;
  assign n7608 = ~x99 & ~n7607;
  assign n7609 = n7290 & ~n7365;
  assign n7610 = n7609 ^ n7293;
  assign n7611 = ~x100 & ~n7610;
  assign n7612 = ~n7608 & ~n7611;
  assign n7613 = n7605 & n7612;
  assign n7614 = n7610 ^ x100;
  assign n7615 = x99 & n7607;
  assign n7616 = n7615 ^ n7610;
  assign n7617 = n7614 & ~n7616;
  assign n7618 = n7617 ^ x100;
  assign n7619 = ~n7613 & ~n7618;
  assign n7620 = n7619 ^ x101;
  assign n7621 = n7297 & ~n7365;
  assign n7622 = n7621 ^ n7303;
  assign n7623 = n7622 ^ n7619;
  assign n7624 = ~n7620 & n7623;
  assign n7625 = n7624 ^ x101;
  assign n7626 = n7625 ^ x102;
  assign n7627 = n7307 & ~n7365;
  assign n7628 = n7627 ^ n7309;
  assign n7629 = n7628 ^ n7625;
  assign n7630 = n7626 & ~n7629;
  assign n7631 = n7630 ^ x102;
  assign n7632 = n7631 ^ x103;
  assign n7633 = n7313 & ~n7365;
  assign n7634 = n7633 ^ n7315;
  assign n7635 = n7634 ^ n7631;
  assign n7636 = n7632 & ~n7635;
  assign n7637 = n7636 ^ x103;
  assign n7638 = n7637 ^ x104;
  assign n7639 = n7319 & ~n7365;
  assign n7640 = n7639 ^ n7322;
  assign n7641 = n7640 ^ n7637;
  assign n7642 = n7638 & ~n7641;
  assign n7643 = n7642 ^ x104;
  assign n7644 = n7643 ^ x105;
  assign n7645 = n7326 & ~n7365;
  assign n7646 = n7645 ^ n7330;
  assign n7647 = n7646 ^ n7643;
  assign n7648 = n7644 & ~n7647;
  assign n7649 = n7648 ^ x105;
  assign n7650 = n7372 & n7649;
  assign n7651 = n7370 ^ x107;
  assign n7652 = x106 & n7367;
  assign n7653 = n7652 ^ n7370;
  assign n7654 = n7651 & ~n7653;
  assign n7655 = n7654 ^ x107;
  assign n7656 = ~n7650 & ~n7655;
  assign n7657 = n7656 ^ x108;
  assign n7658 = n7348 ^ x107;
  assign n7659 = ~n7365 & n7658;
  assign n7660 = n7659 ^ n7051;
  assign n7661 = n7660 ^ n7656;
  assign n7662 = ~n7657 & ~n7661;
  assign n7663 = n7662 ^ x108;
  assign n7664 = n7663 ^ x109;
  assign n7665 = n146 & n7664;
  assign n7666 = n7358 & ~n7665;
  assign n7667 = ~x109 & n7358;
  assign n7668 = n7663 & ~n7667;
  assign n7669 = x109 & n6145;
  assign n7670 = n146 & ~n7669;
  assign n7671 = ~n7668 & n7670;
  assign n7672 = n7521 & n7671;
  assign n7673 = n7672 ^ n7523;
  assign n7674 = ~x85 & ~n7673;
  assign n7675 = n7527 & n7671;
  assign n7676 = n7675 ^ n7529;
  assign n7677 = ~x86 & ~n7676;
  assign n7678 = ~n7674 & ~n7677;
  assign n7679 = x65 & n7365;
  assign n7680 = n7671 & n7679;
  assign n7681 = ~x65 & n7401;
  assign n7682 = ~n7680 & ~n7681;
  assign n7683 = x18 & ~n7682;
  assign n7684 = n7365 ^ x65;
  assign n7685 = n341 & n7684;
  assign n7686 = x18 & n7685;
  assign n7687 = n7686 ^ n340;
  assign n7688 = n7671 & n7687;
  assign n7689 = n7688 ^ n7401;
  assign n7690 = ~n7683 & ~n7689;
  assign n7691 = n7690 ^ x19;
  assign n7692 = n7691 ^ x66;
  assign n7693 = x64 & n7671;
  assign n7694 = n7693 ^ x18;
  assign n7695 = n7694 ^ x65;
  assign n7696 = ~x17 & x64;
  assign n7697 = n7696 ^ n7694;
  assign n7698 = ~n7695 & n7697;
  assign n7699 = n7698 ^ x65;
  assign n7700 = n7699 ^ n7691;
  assign n7701 = n7692 & ~n7700;
  assign n7702 = n7701 ^ x66;
  assign n7703 = n7702 ^ x67;
  assign n7704 = n7413 ^ x66;
  assign n7705 = n7671 & ~n7704;
  assign n7706 = n7705 ^ n7399;
  assign n7707 = n7706 ^ n7702;
  assign n7708 = n7703 & ~n7707;
  assign n7709 = n7708 ^ x67;
  assign n7710 = n7709 ^ x68;
  assign n7711 = n7417 & n7671;
  assign n7712 = n7711 ^ n7426;
  assign n7713 = n7712 ^ n7709;
  assign n7714 = n7710 & n7713;
  assign n7715 = n7714 ^ x68;
  assign n7716 = n7715 ^ x69;
  assign n7717 = n7430 & n7671;
  assign n7718 = n7717 ^ n7432;
  assign n7719 = n7718 ^ n7715;
  assign n7720 = n7716 & ~n7719;
  assign n7721 = n7720 ^ x69;
  assign n7722 = n7721 ^ x70;
  assign n7723 = n7436 & n7671;
  assign n7724 = n7723 ^ n7438;
  assign n7725 = n7724 ^ n7721;
  assign n7726 = n7722 & n7725;
  assign n7727 = n7726 ^ x70;
  assign n7728 = n7727 ^ x71;
  assign n7729 = n7442 & n7671;
  assign n7730 = n7729 ^ n7444;
  assign n7731 = n7730 ^ n7727;
  assign n7732 = n7728 & ~n7731;
  assign n7733 = n7732 ^ x71;
  assign n7734 = n7733 ^ x72;
  assign n7735 = n7448 & n7671;
  assign n7736 = n7735 ^ n7450;
  assign n7737 = n7736 ^ n7733;
  assign n7738 = n7734 & n7737;
  assign n7739 = n7738 ^ x72;
  assign n7740 = n7739 ^ x73;
  assign n7741 = n7454 & n7671;
  assign n7742 = n7741 ^ n7456;
  assign n7743 = n7742 ^ n7739;
  assign n7744 = n7740 & ~n7743;
  assign n7745 = n7744 ^ x73;
  assign n7746 = n7745 ^ x74;
  assign n7747 = n7462 ^ x73;
  assign n7748 = n7747 ^ n7459;
  assign n7749 = n7748 ^ n7462;
  assign n7750 = n7671 & n7749;
  assign n7751 = n7750 ^ n7462;
  assign n7752 = n7751 ^ n7745;
  assign n7753 = n7746 & ~n7752;
  assign n7754 = n7753 ^ x74;
  assign n7755 = n7754 ^ x75;
  assign n7756 = n7466 & n7671;
  assign n7757 = n7756 ^ n7468;
  assign n7758 = n7757 ^ n7754;
  assign n7759 = n7755 & ~n7758;
  assign n7760 = n7759 ^ x75;
  assign n7761 = n7760 ^ x76;
  assign n7762 = n7472 & n7671;
  assign n7763 = n7762 ^ n7474;
  assign n7764 = n7763 ^ n7760;
  assign n7765 = n7761 & ~n7764;
  assign n7766 = n7765 ^ x76;
  assign n7767 = n7766 ^ x77;
  assign n7768 = n7478 & n7671;
  assign n7769 = n7768 ^ n7480;
  assign n7770 = n7769 ^ n7766;
  assign n7771 = n7767 & ~n7770;
  assign n7772 = n7771 ^ x77;
  assign n7773 = n7772 ^ x78;
  assign n7774 = n7484 & n7671;
  assign n7775 = n7774 ^ n7486;
  assign n7776 = n7775 ^ n7772;
  assign n7777 = n7773 & ~n7776;
  assign n7778 = n7777 ^ x78;
  assign n7779 = n7778 ^ x79;
  assign n7780 = n7490 & n7671;
  assign n7781 = n7780 ^ n7492;
  assign n7782 = n7781 ^ n7778;
  assign n7783 = n7779 & ~n7782;
  assign n7784 = n7783 ^ x79;
  assign n7785 = n7784 ^ x80;
  assign n7786 = n7496 & n7671;
  assign n7787 = n7786 ^ n7498;
  assign n7788 = n7787 ^ n7784;
  assign n7789 = n7785 & ~n7788;
  assign n7790 = n7789 ^ x80;
  assign n7791 = n7790 ^ x81;
  assign n7792 = n7501 ^ x80;
  assign n7793 = n7671 & n7792;
  assign n7794 = n7793 ^ n7381;
  assign n7795 = n7794 ^ n7790;
  assign n7796 = n7791 & ~n7795;
  assign n7797 = n7796 ^ x81;
  assign n7798 = n7797 ^ x82;
  assign n7799 = n7501 ^ n7381;
  assign n7800 = n7792 & ~n7799;
  assign n7801 = n7800 ^ x80;
  assign n7802 = n7801 ^ x81;
  assign n7803 = n7671 & n7802;
  assign n7804 = n7803 ^ n7384;
  assign n7805 = n7804 ^ n7797;
  assign n7806 = n7798 & ~n7805;
  assign n7807 = n7806 ^ x82;
  assign n7808 = n7807 ^ x83;
  assign n7809 = n7509 & n7671;
  assign n7810 = n7809 ^ n7511;
  assign n7811 = n7810 ^ n7807;
  assign n7812 = n7808 & ~n7811;
  assign n7813 = n7812 ^ x83;
  assign n7814 = n7813 ^ x84;
  assign n7815 = n7515 & n7671;
  assign n7816 = n7815 ^ n7517;
  assign n7817 = n7816 ^ n7813;
  assign n7818 = n7814 & ~n7817;
  assign n7819 = n7818 ^ x84;
  assign n7820 = n7678 & n7819;
  assign n7821 = n7676 ^ x86;
  assign n7822 = x85 & n7673;
  assign n7823 = n7822 ^ n7676;
  assign n7824 = n7821 & ~n7823;
  assign n7825 = n7824 ^ x86;
  assign n7826 = ~n7820 & ~n7825;
  assign n7827 = n7826 ^ x87;
  assign n7828 = n7533 & n7671;
  assign n7829 = n7828 ^ n7535;
  assign n7830 = n7829 ^ n7826;
  assign n7831 = ~n7827 & n7830;
  assign n7832 = n7831 ^ x87;
  assign n7833 = n7832 ^ x88;
  assign n7834 = n7539 & n7671;
  assign n7835 = n7834 ^ n7541;
  assign n7836 = n7835 ^ n7832;
  assign n7837 = n7833 & ~n7836;
  assign n7838 = n7837 ^ x88;
  assign n7839 = n7838 ^ x89;
  assign n7840 = n7545 & n7671;
  assign n7841 = n7840 ^ n7547;
  assign n7842 = n7841 ^ n7838;
  assign n7843 = n7839 & ~n7842;
  assign n7844 = n7843 ^ x89;
  assign n7845 = n7844 ^ x90;
  assign n7846 = n7551 & n7671;
  assign n7847 = n7846 ^ n7553;
  assign n7848 = n7847 ^ n7844;
  assign n7849 = n7845 & ~n7848;
  assign n7850 = n7849 ^ x90;
  assign n7851 = n7850 ^ x91;
  assign n7852 = n7557 & n7671;
  assign n7853 = n7852 ^ n7559;
  assign n7854 = n7853 ^ n7850;
  assign n7855 = n7851 & ~n7854;
  assign n7856 = n7855 ^ x91;
  assign n7857 = n7856 ^ x92;
  assign n7858 = n7563 & n7671;
  assign n7859 = n7858 ^ n7565;
  assign n7860 = n7859 ^ n7856;
  assign n7861 = n7857 & ~n7860;
  assign n7862 = n7861 ^ x92;
  assign n7863 = n7862 ^ x93;
  assign n7864 = n7569 & n7671;
  assign n7865 = n7864 ^ n7571;
  assign n7866 = n7865 ^ n7862;
  assign n7867 = n7863 & ~n7866;
  assign n7868 = n7867 ^ x93;
  assign n7869 = n7868 ^ x94;
  assign n7870 = n7575 & n7671;
  assign n7871 = n7870 ^ n7577;
  assign n7872 = n7871 ^ n7868;
  assign n7873 = n7869 & ~n7872;
  assign n7874 = n7873 ^ x94;
  assign n7875 = n7874 ^ x95;
  assign n7876 = n7581 & n7671;
  assign n7877 = n7876 ^ n7583;
  assign n7878 = n7877 ^ n7874;
  assign n7879 = n7875 & ~n7878;
  assign n7880 = n7879 ^ x95;
  assign n7881 = n7880 ^ x96;
  assign n7882 = n7587 & n7671;
  assign n7883 = n7882 ^ n7589;
  assign n7884 = n7883 ^ n7880;
  assign n7885 = n7881 & ~n7884;
  assign n7886 = n7885 ^ x96;
  assign n7887 = n7886 ^ x97;
  assign n7888 = n7593 & n7671;
  assign n7889 = n7888 ^ n7595;
  assign n7890 = n7889 ^ n7886;
  assign n7891 = n7887 & ~n7890;
  assign n7892 = n7891 ^ x97;
  assign n7893 = n7892 ^ x98;
  assign n7894 = n7598 ^ x97;
  assign n7895 = n7671 & n7894;
  assign n7896 = n7895 ^ n7374;
  assign n7897 = n7896 ^ n7892;
  assign n7898 = n7893 & ~n7897;
  assign n7899 = n7898 ^ x98;
  assign n7900 = n7899 ^ x99;
  assign n7901 = n7598 ^ n7374;
  assign n7902 = n7894 & ~n7901;
  assign n7903 = n7902 ^ x97;
  assign n7904 = n7903 ^ x98;
  assign n7905 = n7671 & n7904;
  assign n7906 = n7905 ^ n7377;
  assign n7907 = n7906 ^ n7899;
  assign n7908 = n7900 & ~n7907;
  assign n7909 = n7908 ^ x99;
  assign n7910 = n7909 ^ x100;
  assign n7911 = n7605 ^ x99;
  assign n7912 = n7671 & n7911;
  assign n7913 = n7912 ^ n7607;
  assign n7914 = n7913 ^ n7909;
  assign n7915 = n7910 & ~n7914;
  assign n7916 = n7915 ^ x100;
  assign n7917 = n7916 ^ x101;
  assign n7918 = n7607 ^ n7605;
  assign n7919 = n7911 & ~n7918;
  assign n7920 = n7919 ^ x99;
  assign n7921 = n7920 ^ x100;
  assign n7922 = n7671 & n7921;
  assign n7923 = n7922 ^ n7610;
  assign n7924 = n7923 ^ n7916;
  assign n7925 = n7917 & ~n7924;
  assign n7926 = n7925 ^ x101;
  assign n7927 = n7926 ^ x102;
  assign n7928 = ~n7620 & n7671;
  assign n7929 = n7928 ^ n7622;
  assign n7930 = n7929 ^ n7926;
  assign n7931 = n7927 & ~n7930;
  assign n7932 = n7931 ^ x102;
  assign n7933 = n7932 ^ x103;
  assign n7934 = n7626 & n7671;
  assign n7935 = n7934 ^ n7628;
  assign n7936 = n7935 ^ n7932;
  assign n7937 = n7933 & ~n7936;
  assign n7938 = n7937 ^ x103;
  assign n7939 = n7938 ^ x104;
  assign n7940 = n7632 & n7671;
  assign n7941 = n7940 ^ n7634;
  assign n7942 = n7941 ^ n7938;
  assign n7943 = n7939 & ~n7942;
  assign n7944 = n7943 ^ x104;
  assign n7945 = n7944 ^ x105;
  assign n7946 = n7638 & n7671;
  assign n7947 = n7946 ^ n7640;
  assign n7948 = n7947 ^ n7944;
  assign n7949 = n7945 & ~n7948;
  assign n7950 = n7949 ^ x105;
  assign n7951 = n7950 ^ x106;
  assign n7952 = n7644 & n7671;
  assign n7953 = n7952 ^ n7646;
  assign n7954 = n7953 ^ n7950;
  assign n7955 = n7951 & ~n7954;
  assign n7956 = n7955 ^ x106;
  assign n7957 = n7956 ^ x107;
  assign n7958 = n7649 ^ x106;
  assign n7959 = n7671 & n7958;
  assign n7960 = n7959 ^ n7367;
  assign n7961 = n7960 ^ n7956;
  assign n7962 = n7957 & ~n7961;
  assign n7963 = n7962 ^ x107;
  assign n7964 = n7963 ^ x108;
  assign n7965 = n7649 ^ n7367;
  assign n7966 = n7958 & ~n7965;
  assign n7967 = n7966 ^ x106;
  assign n7968 = n7967 ^ x107;
  assign n7969 = n7671 & n7968;
  assign n7970 = n7969 ^ n7370;
  assign n7971 = n7970 ^ n7963;
  assign n7972 = n7964 & ~n7971;
  assign n7973 = n7972 ^ x108;
  assign n7974 = n7973 ^ x109;
  assign n7975 = ~n7657 & n7671;
  assign n7976 = n7975 ^ n7660;
  assign n7977 = n7976 ^ n7973;
  assign n7978 = n7974 & n7977;
  assign n7979 = n7978 ^ x109;
  assign n7980 = n7979 ^ x110;
  assign n7981 = n145 & n7980;
  assign n7982 = n7666 & ~n7981;
  assign n7983 = n141 & n143;
  assign n7986 = ~n7666 & n7981;
  assign n7984 = n145 & ~n7979;
  assign n7985 = ~n146 & ~n7984;
  assign n7987 = n7986 ^ n7985;
  assign n7991 = n7945 & ~n7987;
  assign n7992 = n7991 ^ n7947;
  assign n7993 = x106 & n7992;
  assign n7994 = n7900 & ~n7987;
  assign n7995 = n7994 ^ n7906;
  assign n7996 = ~x100 & ~n7995;
  assign n7997 = n7863 & ~n7987;
  assign n7998 = n7997 ^ n7865;
  assign n7999 = x94 & n7998;
  assign n8000 = n7710 & ~n7987;
  assign n8001 = n8000 ^ n7712;
  assign n8002 = ~x69 & n8001;
  assign n8003 = ~n7694 & n7987;
  assign n8004 = ~x16 & x65;
  assign n8005 = n8003 & n8004;
  assign n8006 = x17 & ~n7987;
  assign n8007 = x16 & ~x65;
  assign n8008 = n8006 & ~n8007;
  assign n8009 = ~n7695 & n8008;
  assign n8010 = ~n8005 & ~n8009;
  assign n8011 = x64 & ~n8010;
  assign n8012 = x64 & ~n7987;
  assign n8013 = ~x17 & x65;
  assign n8014 = ~n8012 & n8013;
  assign n8015 = n7987 ^ n7694;
  assign n8016 = n8014 & n8015;
  assign n8017 = ~x65 & ~n7987;
  assign n8018 = ~x16 & x64;
  assign n8019 = ~x17 & n8018;
  assign n8020 = ~n7694 & n8019;
  assign n8021 = ~n8017 & n8020;
  assign n8022 = ~x66 & ~n8021;
  assign n8023 = ~n8016 & n8022;
  assign n8024 = ~n8011 & n8023;
  assign n8025 = x17 & ~x65;
  assign n8026 = n7987 & n8025;
  assign n8027 = n8018 & ~n8026;
  assign n8028 = ~x65 & ~n7696;
  assign n8029 = ~n7987 & ~n8028;
  assign n8030 = n7694 & ~n8013;
  assign n8031 = ~n8029 & n8030;
  assign n8032 = ~n8027 & n8031;
  assign n8033 = n7696 & ~n8004;
  assign n8034 = ~n7695 & n8033;
  assign n8035 = ~x18 & n202;
  assign n8036 = x17 & n8035;
  assign n8037 = ~n8034 & ~n8036;
  assign n8038 = ~n7987 & ~n8037;
  assign n8039 = ~n8032 & ~n8038;
  assign n8040 = ~n8024 & n8039;
  assign n8041 = n8040 ^ x67;
  assign n8042 = n7699 ^ x66;
  assign n8043 = ~n7987 & n8042;
  assign n8044 = n8043 ^ n7691;
  assign n8045 = n8044 ^ n8040;
  assign n8046 = n8041 & ~n8045;
  assign n8047 = n8046 ^ x67;
  assign n8048 = n8047 ^ x68;
  assign n8049 = n7703 & ~n7987;
  assign n8050 = n8049 ^ n7706;
  assign n8051 = n8050 ^ n8047;
  assign n8052 = n8048 & ~n8051;
  assign n8053 = n8052 ^ x68;
  assign n8054 = ~n8002 & n8053;
  assign n8055 = n7716 & ~n7987;
  assign n8056 = n8055 ^ n7718;
  assign n8057 = x70 & n8056;
  assign n8058 = x69 & ~n8001;
  assign n8059 = ~n8057 & ~n8058;
  assign n8060 = ~n8054 & n8059;
  assign n8061 = ~x70 & ~n8056;
  assign n8062 = ~n8060 & ~n8061;
  assign n8063 = n8062 ^ x71;
  assign n8064 = n7722 & ~n7987;
  assign n8065 = n8064 ^ n7724;
  assign n8066 = n8065 ^ n8062;
  assign n8067 = n8063 & n8066;
  assign n8068 = n8067 ^ x71;
  assign n8069 = n8068 ^ x72;
  assign n8070 = n7728 & ~n7987;
  assign n8071 = n8070 ^ n7730;
  assign n8072 = n8071 ^ n8068;
  assign n8073 = n8069 & ~n8072;
  assign n8074 = n8073 ^ x72;
  assign n8075 = n8074 ^ x73;
  assign n8076 = n7734 & ~n7987;
  assign n8077 = n8076 ^ n7736;
  assign n8078 = n8077 ^ n8074;
  assign n8079 = n8075 & n8078;
  assign n8080 = n8079 ^ x73;
  assign n8081 = n8080 ^ x74;
  assign n8082 = n7740 & ~n7987;
  assign n8083 = n8082 ^ n7742;
  assign n8084 = n8083 ^ n8080;
  assign n8085 = n8081 & ~n8084;
  assign n8086 = n8085 ^ x74;
  assign n8087 = n8086 ^ x75;
  assign n8088 = n7746 & ~n7987;
  assign n8089 = n8088 ^ n7751;
  assign n8090 = n8089 ^ n8086;
  assign n8091 = n8087 & ~n8090;
  assign n8092 = n8091 ^ x75;
  assign n8093 = n8092 ^ x76;
  assign n8094 = n7755 & ~n7987;
  assign n8095 = n8094 ^ n7757;
  assign n8096 = n8095 ^ n8092;
  assign n8097 = n8093 & ~n8096;
  assign n8098 = n8097 ^ x76;
  assign n8099 = n8098 ^ x77;
  assign n8100 = n7761 & ~n7987;
  assign n8101 = n8100 ^ n7763;
  assign n8102 = n8101 ^ n8098;
  assign n8103 = n8099 & ~n8102;
  assign n8104 = n8103 ^ x77;
  assign n8105 = n8104 ^ x78;
  assign n8106 = n7767 & ~n7987;
  assign n8107 = n8106 ^ n7769;
  assign n8108 = n8107 ^ n8104;
  assign n8109 = n8105 & ~n8108;
  assign n8110 = n8109 ^ x78;
  assign n8111 = n8110 ^ x79;
  assign n8112 = n7773 & ~n7987;
  assign n8113 = n8112 ^ n7775;
  assign n8114 = n8113 ^ n8110;
  assign n8115 = n8111 & ~n8114;
  assign n8116 = n8115 ^ x79;
  assign n8117 = n8116 ^ x80;
  assign n8118 = n7779 & ~n7987;
  assign n8119 = n8118 ^ n7781;
  assign n8120 = n8119 ^ n8116;
  assign n8121 = n8117 & ~n8120;
  assign n8122 = n8121 ^ x80;
  assign n8123 = n8122 ^ x81;
  assign n8124 = n7785 & ~n7987;
  assign n8125 = n8124 ^ n7787;
  assign n8126 = n8125 ^ n8122;
  assign n8127 = n8123 & ~n8126;
  assign n8128 = n8127 ^ x81;
  assign n8129 = n8128 ^ x82;
  assign n8130 = n7791 & ~n7987;
  assign n8131 = n8130 ^ n7794;
  assign n8132 = n8131 ^ n8128;
  assign n8133 = n8129 & ~n8132;
  assign n8134 = n8133 ^ x82;
  assign n8135 = n8134 ^ x83;
  assign n8136 = n7798 & ~n7987;
  assign n8137 = n8136 ^ n7804;
  assign n8138 = n8137 ^ n8134;
  assign n8139 = n8135 & ~n8138;
  assign n8140 = n8139 ^ x83;
  assign n8141 = n8140 ^ x84;
  assign n8142 = n7808 & ~n7987;
  assign n8143 = n8142 ^ n7810;
  assign n8144 = n8143 ^ n8140;
  assign n8145 = n8141 & ~n8144;
  assign n8146 = n8145 ^ x84;
  assign n8147 = n8146 ^ x85;
  assign n8148 = n7814 & ~n7987;
  assign n8149 = n8148 ^ n7816;
  assign n8150 = n8149 ^ n8146;
  assign n8151 = n8147 & ~n8150;
  assign n8152 = n8151 ^ x85;
  assign n8153 = n8152 ^ x86;
  assign n8154 = n7819 ^ x85;
  assign n8155 = ~n7987 & n8154;
  assign n8156 = n8155 ^ n7673;
  assign n8157 = n8156 ^ n8152;
  assign n8158 = n8153 & ~n8157;
  assign n8159 = n8158 ^ x86;
  assign n8160 = n8159 ^ x87;
  assign n8161 = n7819 ^ n7673;
  assign n8162 = n8154 & ~n8161;
  assign n8163 = n8162 ^ x85;
  assign n8164 = n8163 ^ x86;
  assign n8165 = ~n7987 & n8164;
  assign n8166 = n8165 ^ n7676;
  assign n8167 = n8166 ^ n8159;
  assign n8168 = n8160 & ~n8167;
  assign n8169 = n8168 ^ x87;
  assign n8170 = n8169 ^ x88;
  assign n8171 = ~n7827 & ~n7987;
  assign n8172 = n8171 ^ n7829;
  assign n8173 = n8172 ^ n8169;
  assign n8174 = n8170 & ~n8173;
  assign n8175 = n8174 ^ x88;
  assign n8176 = n8175 ^ x89;
  assign n8177 = n7833 & ~n7987;
  assign n8178 = n8177 ^ n7835;
  assign n8179 = n8178 ^ n8175;
  assign n8180 = n8176 & ~n8179;
  assign n8181 = n8180 ^ x89;
  assign n8182 = n8181 ^ x90;
  assign n8183 = n7839 & ~n7987;
  assign n8184 = n8183 ^ n7841;
  assign n8185 = n8184 ^ n8181;
  assign n8186 = n8182 & ~n8185;
  assign n8187 = n8186 ^ x90;
  assign n8188 = n8187 ^ x91;
  assign n8189 = n7845 & ~n7987;
  assign n8190 = n8189 ^ n7847;
  assign n8191 = n8190 ^ n8187;
  assign n8192 = n8188 & ~n8191;
  assign n8193 = n8192 ^ x91;
  assign n8194 = n8193 ^ x92;
  assign n8195 = n7851 & ~n7987;
  assign n8196 = n8195 ^ n7853;
  assign n8197 = n8196 ^ n8193;
  assign n8198 = n8194 & ~n8197;
  assign n8199 = n8198 ^ x92;
  assign n8200 = n8199 ^ x93;
  assign n8201 = n7857 & ~n7987;
  assign n8202 = n8201 ^ n7859;
  assign n8203 = n8202 ^ n8199;
  assign n8204 = n8200 & ~n8203;
  assign n8205 = n8204 ^ x93;
  assign n8206 = ~n7999 & ~n8205;
  assign n8207 = ~x94 & ~n7998;
  assign n8208 = n7869 & ~n7987;
  assign n8209 = n8208 ^ n7871;
  assign n8210 = ~x95 & ~n8209;
  assign n8211 = ~n8207 & ~n8210;
  assign n8212 = ~n8206 & n8211;
  assign n8213 = x95 & n8209;
  assign n8214 = ~n8212 & ~n8213;
  assign n8215 = n8214 ^ x96;
  assign n8216 = n7875 & ~n7987;
  assign n8217 = n8216 ^ n7877;
  assign n8218 = n8217 ^ n8214;
  assign n8219 = ~n8215 & n8218;
  assign n8220 = n8219 ^ x96;
  assign n8221 = n8220 ^ x97;
  assign n8222 = n7881 & ~n7987;
  assign n8223 = n8222 ^ n7883;
  assign n8224 = n8223 ^ n8220;
  assign n8225 = n8221 & ~n8224;
  assign n8226 = n8225 ^ x97;
  assign n8227 = n8226 ^ x98;
  assign n8228 = n7887 & ~n7987;
  assign n8229 = n8228 ^ n7889;
  assign n8230 = n8229 ^ n8226;
  assign n8231 = n8227 & ~n8230;
  assign n8232 = n8231 ^ x98;
  assign n8233 = n8232 ^ x99;
  assign n8234 = n7893 & ~n7987;
  assign n8235 = n8234 ^ n7896;
  assign n8236 = n8235 ^ n8232;
  assign n8237 = n8233 & ~n8236;
  assign n8238 = n8237 ^ x99;
  assign n8239 = ~n7996 & n8238;
  assign n8240 = n7910 & ~n7987;
  assign n8241 = n8240 ^ n7913;
  assign n8242 = x101 & n8241;
  assign n8243 = x100 & n7995;
  assign n8244 = ~n8242 & ~n8243;
  assign n8245 = ~n8239 & n8244;
  assign n8246 = ~x101 & ~n8241;
  assign n8247 = ~n8245 & ~n8246;
  assign n8248 = n8247 ^ x102;
  assign n8249 = n7917 & ~n7987;
  assign n8250 = n8249 ^ n7923;
  assign n8251 = n8250 ^ n8247;
  assign n8252 = n8248 & ~n8251;
  assign n8253 = n8252 ^ x102;
  assign n8254 = n8253 ^ x103;
  assign n8255 = n7927 & ~n7987;
  assign n8256 = n8255 ^ n7929;
  assign n8257 = n8256 ^ n8253;
  assign n8258 = n8254 & ~n8257;
  assign n8259 = n8258 ^ x103;
  assign n8260 = n8259 ^ x104;
  assign n8261 = n7933 & ~n7987;
  assign n8262 = n8261 ^ n7935;
  assign n8263 = n8262 ^ n8259;
  assign n8264 = n8260 & ~n8263;
  assign n8265 = n8264 ^ x104;
  assign n8266 = n8265 ^ x105;
  assign n8267 = n7939 & ~n7987;
  assign n8268 = n8267 ^ n7941;
  assign n8269 = n8268 ^ n8265;
  assign n8270 = n8266 & ~n8269;
  assign n8271 = n8270 ^ x105;
  assign n8272 = ~n7993 & ~n8271;
  assign n8273 = ~x106 & ~n7992;
  assign n8274 = n7951 & ~n7987;
  assign n8275 = n8274 ^ n7953;
  assign n8276 = ~x107 & ~n8275;
  assign n8277 = ~n8273 & ~n8276;
  assign n8278 = ~n8272 & n8277;
  assign n8279 = x107 & n8275;
  assign n8280 = ~n8278 & ~n8279;
  assign n8281 = n8280 ^ x108;
  assign n7988 = n7974 & ~n7987;
  assign n7989 = n7988 ^ n7976;
  assign n7990 = n7989 ^ x110;
  assign n8282 = n7957 & ~n7987;
  assign n8283 = n8282 ^ n7960;
  assign n8284 = n8283 ^ n8280;
  assign n8285 = ~n8281 & n8284;
  assign n8286 = n8285 ^ x108;
  assign n8287 = n8286 ^ x109;
  assign n8288 = n7964 & ~n7987;
  assign n8289 = n8288 ^ n7970;
  assign n8290 = n8289 ^ n8286;
  assign n8291 = n8287 & ~n8290;
  assign n8292 = n8291 ^ x109;
  assign n8293 = n8292 ^ n7989;
  assign n8294 = ~n7990 & n8293;
  assign n8295 = n8294 ^ x110;
  assign n8296 = n7666 & ~n8295;
  assign n8297 = ~n7982 & n8295;
  assign n8298 = ~x111 & ~n8297;
  assign n8299 = ~n8296 & ~n8298;
  assign n8300 = ~x112 & n7983;
  assign n8301 = ~n8299 & n8300;
  assign n8302 = ~n8281 & n8301;
  assign n8303 = n8302 ^ n8283;
  assign n8304 = ~x109 & ~n8303;
  assign n8305 = n8254 & n8301;
  assign n8306 = n8305 ^ n8256;
  assign n8307 = ~x104 & ~n8306;
  assign n8308 = n8260 & n8301;
  assign n8309 = n8308 ^ n8262;
  assign n8310 = ~x105 & ~n8309;
  assign n8311 = ~n8307 & ~n8310;
  assign n8312 = n8117 & n8301;
  assign n8313 = n8312 ^ n8119;
  assign n8314 = ~x81 & ~n8313;
  assign n8315 = n8123 & n8301;
  assign n8316 = n8315 ^ n8125;
  assign n8317 = ~x82 & ~n8316;
  assign n8318 = ~n8314 & ~n8317;
  assign n8319 = n8012 & ~n8301;
  assign n8320 = x65 & n8300;
  assign n8321 = x16 & n8320;
  assign n8322 = n7987 & n8321;
  assign n8323 = ~n8299 & n8322;
  assign n8324 = n8007 & n8012;
  assign n8325 = ~n8323 & ~n8324;
  assign n8326 = ~n8319 & n8325;
  assign n8327 = ~x16 & ~n8017;
  assign n8328 = ~n219 & n7987;
  assign n8329 = n8327 & ~n8328;
  assign n8330 = ~n202 & ~n8329;
  assign n8331 = n8301 & ~n8330;
  assign n8332 = n8326 & ~n8331;
  assign n8333 = n8332 ^ x17;
  assign n8334 = n8333 ^ x66;
  assign n8335 = x64 & n8301;
  assign n8336 = x15 & n8007;
  assign n8337 = n8336 ^ x16;
  assign n8338 = n8335 & n8337;
  assign n8339 = ~x15 & n8018;
  assign n8340 = ~n8004 & ~n8339;
  assign n8341 = ~n8301 & ~n8340;
  assign n8342 = ~x15 & x65;
  assign n8343 = n8342 ^ n8004;
  assign n8344 = x64 & n8343;
  assign n8345 = n8344 ^ n8004;
  assign n8346 = ~n8341 & ~n8345;
  assign n8347 = ~n8338 & n8346;
  assign n8348 = n8347 ^ n8333;
  assign n8349 = n8334 & n8348;
  assign n8350 = n8349 ^ x66;
  assign n8351 = n8350 ^ x67;
  assign n8355 = ~n8025 & n8327;
  assign n8356 = ~n8008 & ~n8355;
  assign n8357 = x64 & ~n8356;
  assign n8358 = ~n8014 & ~n8357;
  assign n8359 = n8358 ^ x66;
  assign n8360 = n8301 & ~n8359;
  assign n8352 = n7696 ^ x65;
  assign n8353 = ~n7987 & n8352;
  assign n8354 = n8353 ^ n7694;
  assign n8361 = n8360 ^ n8354;
  assign n8362 = n8361 ^ n8350;
  assign n8363 = n8351 & n8362;
  assign n8364 = n8363 ^ x67;
  assign n8365 = n8364 ^ x68;
  assign n8366 = n8041 & n8301;
  assign n8367 = n8366 ^ n8044;
  assign n8368 = n8367 ^ n8364;
  assign n8369 = n8365 & ~n8368;
  assign n8370 = n8369 ^ x68;
  assign n8371 = n8370 ^ x69;
  assign n8372 = n8048 & n8301;
  assign n8373 = n8372 ^ n8050;
  assign n8374 = n8373 ^ n8370;
  assign n8375 = n8371 & ~n8374;
  assign n8376 = n8375 ^ x69;
  assign n8377 = n8376 ^ x70;
  assign n8378 = n8053 ^ x69;
  assign n8379 = n8301 & n8378;
  assign n8380 = n8379 ^ n8001;
  assign n8381 = n8380 ^ n8376;
  assign n8382 = n8377 & n8381;
  assign n8383 = n8382 ^ x70;
  assign n8384 = n8383 ^ x71;
  assign n8385 = ~n8054 & ~n8058;
  assign n8386 = n8385 ^ x70;
  assign n8387 = n8301 & ~n8386;
  assign n8388 = n8387 ^ n8056;
  assign n8389 = n8388 ^ n8383;
  assign n8390 = n8384 & ~n8389;
  assign n8391 = n8390 ^ x71;
  assign n8392 = n8391 ^ x72;
  assign n8393 = n8063 & n8301;
  assign n8394 = n8393 ^ n8065;
  assign n8395 = n8394 ^ n8391;
  assign n8396 = n8392 & n8395;
  assign n8397 = n8396 ^ x72;
  assign n8398 = n8397 ^ x73;
  assign n8399 = n8069 & n8301;
  assign n8400 = n8399 ^ n8071;
  assign n8401 = n8400 ^ n8397;
  assign n8402 = n8398 & ~n8401;
  assign n8403 = n8402 ^ x73;
  assign n8404 = n8403 ^ x74;
  assign n8405 = n8075 & n8301;
  assign n8406 = n8405 ^ n8077;
  assign n8407 = n8406 ^ n8403;
  assign n8408 = n8404 & n8407;
  assign n8409 = n8408 ^ x74;
  assign n8410 = n8409 ^ x75;
  assign n8411 = n8081 & n8301;
  assign n8412 = n8411 ^ n8083;
  assign n8413 = n8412 ^ n8409;
  assign n8414 = n8410 & ~n8413;
  assign n8415 = n8414 ^ x75;
  assign n8416 = n8415 ^ x76;
  assign n8417 = n8087 & n8301;
  assign n8418 = n8417 ^ n8089;
  assign n8419 = n8418 ^ n8415;
  assign n8420 = n8416 & ~n8419;
  assign n8421 = n8420 ^ x76;
  assign n8422 = n8421 ^ x77;
  assign n8423 = n8093 & n8301;
  assign n8424 = n8423 ^ n8095;
  assign n8425 = n8424 ^ n8421;
  assign n8426 = n8422 & ~n8425;
  assign n8427 = n8426 ^ x77;
  assign n8428 = n8427 ^ x78;
  assign n8429 = n8099 & n8301;
  assign n8430 = n8429 ^ n8101;
  assign n8431 = n8430 ^ n8427;
  assign n8432 = n8428 & ~n8431;
  assign n8433 = n8432 ^ x78;
  assign n8434 = n8433 ^ x79;
  assign n8435 = n8105 & n8301;
  assign n8436 = n8435 ^ n8107;
  assign n8437 = n8436 ^ n8433;
  assign n8438 = n8434 & ~n8437;
  assign n8439 = n8438 ^ x79;
  assign n8440 = n8439 ^ x80;
  assign n8441 = n8111 & n8301;
  assign n8442 = n8441 ^ n8113;
  assign n8443 = n8442 ^ n8439;
  assign n8444 = n8440 & ~n8443;
  assign n8445 = n8444 ^ x80;
  assign n8446 = n8318 & n8445;
  assign n8447 = n8316 ^ x82;
  assign n8448 = x81 & n8313;
  assign n8449 = n8448 ^ n8316;
  assign n8450 = n8447 & ~n8449;
  assign n8451 = n8450 ^ x82;
  assign n8452 = ~n8446 & ~n8451;
  assign n8453 = n8452 ^ x83;
  assign n8454 = n8129 & n8301;
  assign n8455 = n8454 ^ n8131;
  assign n8456 = n8455 ^ n8452;
  assign n8457 = ~n8453 & n8456;
  assign n8458 = n8457 ^ x83;
  assign n8459 = n8458 ^ x84;
  assign n8460 = n8135 & n8301;
  assign n8461 = n8460 ^ n8137;
  assign n8462 = n8461 ^ n8458;
  assign n8463 = n8459 & ~n8462;
  assign n8464 = n8463 ^ x84;
  assign n8465 = n8464 ^ x85;
  assign n8466 = n8141 & n8301;
  assign n8467 = n8466 ^ n8143;
  assign n8468 = n8467 ^ n8464;
  assign n8469 = n8465 & ~n8468;
  assign n8470 = n8469 ^ x85;
  assign n8471 = n8470 ^ x86;
  assign n8472 = n8147 & n8301;
  assign n8473 = n8472 ^ n8149;
  assign n8474 = n8473 ^ n8470;
  assign n8475 = n8471 & ~n8474;
  assign n8476 = n8475 ^ x86;
  assign n8477 = n8476 ^ x87;
  assign n8478 = n8153 & n8301;
  assign n8479 = n8478 ^ n8156;
  assign n8480 = n8479 ^ n8476;
  assign n8481 = n8477 & ~n8480;
  assign n8482 = n8481 ^ x87;
  assign n8483 = n8482 ^ x88;
  assign n8484 = n8160 & n8301;
  assign n8485 = n8484 ^ n8166;
  assign n8486 = n8485 ^ n8482;
  assign n8487 = n8483 & ~n8486;
  assign n8488 = n8487 ^ x88;
  assign n8489 = n8488 ^ x89;
  assign n8490 = n8170 & n8301;
  assign n8491 = n8490 ^ n8172;
  assign n8492 = n8491 ^ n8488;
  assign n8493 = n8489 & ~n8492;
  assign n8494 = n8493 ^ x89;
  assign n8495 = n8494 ^ x90;
  assign n8496 = n8176 & n8301;
  assign n8497 = n8496 ^ n8178;
  assign n8498 = n8497 ^ n8494;
  assign n8499 = n8495 & ~n8498;
  assign n8500 = n8499 ^ x90;
  assign n8501 = n8500 ^ x91;
  assign n8502 = n8182 & n8301;
  assign n8503 = n8502 ^ n8184;
  assign n8504 = n8503 ^ n8500;
  assign n8505 = n8501 & ~n8504;
  assign n8506 = n8505 ^ x91;
  assign n8507 = n8506 ^ x92;
  assign n8508 = n8188 & n8301;
  assign n8509 = n8508 ^ n8190;
  assign n8510 = n8509 ^ n8506;
  assign n8511 = n8507 & ~n8510;
  assign n8512 = n8511 ^ x92;
  assign n8513 = n8512 ^ x93;
  assign n8514 = n8194 & n8301;
  assign n8515 = n8514 ^ n8196;
  assign n8516 = n8515 ^ n8512;
  assign n8517 = n8513 & ~n8516;
  assign n8518 = n8517 ^ x93;
  assign n8519 = n8518 ^ x94;
  assign n8520 = n8200 & n8301;
  assign n8521 = n8520 ^ n8202;
  assign n8522 = n8521 ^ n8518;
  assign n8523 = n8519 & ~n8522;
  assign n8524 = n8523 ^ x94;
  assign n8525 = n8524 ^ x95;
  assign n8526 = n8205 ^ x94;
  assign n8527 = n8301 & n8526;
  assign n8528 = n8527 ^ n7998;
  assign n8529 = n8528 ^ n8524;
  assign n8530 = n8525 & ~n8529;
  assign n8531 = n8530 ^ x95;
  assign n8532 = n8531 ^ x96;
  assign n8533 = ~n8206 & ~n8207;
  assign n8534 = n8533 ^ x95;
  assign n8535 = n8301 & n8534;
  assign n8536 = n8535 ^ n8209;
  assign n8537 = n8536 ^ n8531;
  assign n8538 = n8532 & ~n8537;
  assign n8539 = n8538 ^ x96;
  assign n8540 = n8539 ^ x97;
  assign n8541 = ~n8215 & n8301;
  assign n8542 = n8541 ^ n8217;
  assign n8543 = n8542 ^ n8539;
  assign n8544 = n8540 & ~n8543;
  assign n8545 = n8544 ^ x97;
  assign n8546 = n8545 ^ x98;
  assign n8547 = n8221 & n8301;
  assign n8548 = n8547 ^ n8223;
  assign n8549 = n8548 ^ n8545;
  assign n8550 = n8546 & ~n8549;
  assign n8551 = n8550 ^ x98;
  assign n8552 = n8551 ^ x99;
  assign n8553 = n8227 & n8301;
  assign n8554 = n8553 ^ n8229;
  assign n8555 = n8554 ^ n8551;
  assign n8556 = n8552 & ~n8555;
  assign n8557 = n8556 ^ x99;
  assign n8558 = n8557 ^ x100;
  assign n8559 = n8233 & n8301;
  assign n8560 = n8559 ^ n8235;
  assign n8561 = n8560 ^ n8557;
  assign n8562 = n8558 & ~n8561;
  assign n8563 = n8562 ^ x100;
  assign n8564 = n8563 ^ x101;
  assign n8565 = n8238 ^ x100;
  assign n8566 = n8301 & n8565;
  assign n8567 = n8566 ^ n7995;
  assign n8568 = n8567 ^ n8563;
  assign n8569 = n8564 & ~n8568;
  assign n8570 = n8569 ^ x101;
  assign n8571 = n8570 ^ x102;
  assign n8572 = ~n8239 & ~n8243;
  assign n8573 = n8572 ^ x101;
  assign n8574 = n8301 & ~n8573;
  assign n8575 = n8574 ^ n8241;
  assign n8576 = n8575 ^ n8570;
  assign n8577 = n8571 & ~n8576;
  assign n8578 = n8577 ^ x102;
  assign n8579 = n8578 ^ x103;
  assign n8580 = n8248 & n8301;
  assign n8581 = n8580 ^ n8250;
  assign n8582 = n8581 ^ n8578;
  assign n8583 = n8579 & ~n8582;
  assign n8584 = n8583 ^ x103;
  assign n8585 = n8311 & n8584;
  assign n8586 = n8309 ^ x105;
  assign n8587 = x104 & n8306;
  assign n8588 = n8587 ^ n8309;
  assign n8589 = n8586 & ~n8588;
  assign n8590 = n8589 ^ x105;
  assign n8591 = ~n8585 & ~n8590;
  assign n8592 = n8591 ^ x106;
  assign n8593 = n8266 & n8301;
  assign n8594 = n8593 ^ n8268;
  assign n8595 = n8594 ^ n8591;
  assign n8596 = ~n8592 & n8595;
  assign n8597 = n8596 ^ x106;
  assign n8598 = n8597 ^ x107;
  assign n8599 = n8271 ^ x106;
  assign n8600 = n8301 & n8599;
  assign n8601 = n8600 ^ n7992;
  assign n8602 = n8601 ^ n8597;
  assign n8603 = n8598 & ~n8602;
  assign n8604 = n8603 ^ x107;
  assign n8605 = n8604 ^ x108;
  assign n8606 = ~n8272 & ~n8273;
  assign n8607 = n8606 ^ x107;
  assign n8608 = n8301 & n8607;
  assign n8609 = n8608 ^ n8275;
  assign n8610 = n8609 ^ n8604;
  assign n8611 = n8605 & ~n8610;
  assign n8612 = n8611 ^ x108;
  assign n8613 = ~n8304 & n8612;
  assign n8614 = n8287 & n8301;
  assign n8615 = n8614 ^ n8289;
  assign n8616 = x110 & n8615;
  assign n8617 = x109 & n8303;
  assign n8618 = ~n8616 & ~n8617;
  assign n8619 = ~n8613 & n8618;
  assign n8620 = ~x110 & ~n8615;
  assign n8621 = ~n8619 & ~n8620;
  assign n8622 = n8292 ^ x110;
  assign n8623 = n8301 & n8622;
  assign n8624 = n8623 ^ n7989;
  assign n8625 = n8621 & ~n8624;
  assign n8626 = ~x111 & ~n8625;
  assign n8628 = ~n8621 & n8624;
  assign n8629 = ~n8626 & ~n8628;
  assign n8627 = ~n8295 & n8626;
  assign n8630 = n8629 ^ n8627;
  assign n8631 = ~x112 & n8630;
  assign n8632 = n8631 ^ n8629;
  assign n8633 = n7983 & ~n8632;
  assign n8634 = n7982 & ~n8633;
  assign n8635 = ~x114 & n141;
  assign n8636 = n7358 & n7983;
  assign n8637 = ~n8629 & n8636;
  assign n8638 = ~x111 & n8295;
  assign n8639 = n8301 & n8638;
  assign n8640 = n7982 & ~n8639;
  assign n8641 = n8625 & ~n8640;
  assign n8642 = n8300 & ~n8641;
  assign n8643 = ~n8295 & n8301;
  assign n8644 = n7982 & ~n8643;
  assign n8645 = x111 & ~n8644;
  assign n8646 = ~n8628 & n8645;
  assign n8647 = n8642 & ~n8646;
  assign n8648 = ~n8637 & ~n8647;
  assign n8649 = n8477 & ~n8648;
  assign n8650 = n8649 ^ n8479;
  assign n8651 = ~x88 & ~n8650;
  assign n8652 = n8483 & ~n8648;
  assign n8653 = n8652 ^ n8485;
  assign n8654 = ~x89 & ~n8653;
  assign n8655 = ~n8651 & ~n8654;
  assign n8656 = n8459 & ~n8648;
  assign n8657 = n8656 ^ n8461;
  assign n8658 = x85 & n8657;
  assign n8659 = n8410 & ~n8648;
  assign n8660 = n8659 ^ n8412;
  assign n8661 = ~x76 & ~n8660;
  assign n8662 = n8416 & ~n8648;
  assign n8663 = n8662 ^ n8418;
  assign n8664 = ~x77 & ~n8663;
  assign n8665 = ~n8661 & ~n8664;
  assign n8666 = x64 & ~n8648;
  assign n8667 = n8666 ^ x15;
  assign n8668 = n8667 ^ x65;
  assign n8669 = ~x14 & x64;
  assign n8670 = n8669 ^ n8667;
  assign n8671 = ~n8668 & n8670;
  assign n8672 = n8671 ^ x65;
  assign n8673 = n8672 ^ x66;
  assign n8674 = n219 & ~n8301;
  assign n8675 = ~n8299 & n8320;
  assign n8676 = ~n8674 & ~n8675;
  assign n8677 = ~x15 & ~n8676;
  assign n8678 = ~x65 & ~n8677;
  assign n8679 = ~n8648 & ~n8678;
  assign n8680 = ~n8335 & ~n8679;
  assign n8681 = x15 & ~n8675;
  assign n8682 = ~n202 & ~n8681;
  assign n8683 = ~n8677 & n8682;
  assign n8684 = ~n8648 & n8683;
  assign n8685 = ~n8680 & ~n8684;
  assign n8686 = n8685 ^ x16;
  assign n8687 = n8686 ^ n8672;
  assign n8688 = n8673 & n8687;
  assign n8689 = n8688 ^ x66;
  assign n8690 = n8689 ^ x67;
  assign n8691 = n8347 ^ x66;
  assign n8692 = ~n8648 & ~n8691;
  assign n8693 = n8692 ^ n8333;
  assign n8694 = n8693 ^ n8689;
  assign n8695 = n8690 & ~n8694;
  assign n8696 = n8695 ^ x67;
  assign n8697 = n8696 ^ x68;
  assign n8698 = n8351 & ~n8648;
  assign n8699 = n8698 ^ n8361;
  assign n8700 = n8699 ^ n8696;
  assign n8701 = n8697 & n8700;
  assign n8702 = n8701 ^ x68;
  assign n8703 = n8702 ^ x69;
  assign n8704 = n8365 & ~n8648;
  assign n8705 = n8704 ^ n8367;
  assign n8706 = n8705 ^ n8702;
  assign n8707 = n8703 & ~n8706;
  assign n8708 = n8707 ^ x69;
  assign n8709 = n8708 ^ x70;
  assign n8710 = n8371 & ~n8648;
  assign n8711 = n8710 ^ n8373;
  assign n8712 = n8711 ^ n8708;
  assign n8713 = n8709 & ~n8712;
  assign n8714 = n8713 ^ x70;
  assign n8715 = n8714 ^ x71;
  assign n8716 = n8377 & ~n8648;
  assign n8717 = n8716 ^ n8380;
  assign n8718 = n8717 ^ n8714;
  assign n8719 = n8715 & n8718;
  assign n8720 = n8719 ^ x71;
  assign n8721 = n8720 ^ x72;
  assign n8722 = n8384 & ~n8648;
  assign n8723 = n8722 ^ n8388;
  assign n8724 = n8723 ^ n8720;
  assign n8725 = n8721 & ~n8724;
  assign n8726 = n8725 ^ x72;
  assign n8727 = n8726 ^ x73;
  assign n8728 = n8392 & ~n8648;
  assign n8729 = n8728 ^ n8394;
  assign n8730 = n8729 ^ n8726;
  assign n8731 = n8727 & n8730;
  assign n8732 = n8731 ^ x73;
  assign n8733 = n8732 ^ x74;
  assign n8734 = n8398 & ~n8648;
  assign n8735 = n8734 ^ n8400;
  assign n8736 = n8735 ^ n8732;
  assign n8737 = n8733 & ~n8736;
  assign n8738 = n8737 ^ x74;
  assign n8739 = n8738 ^ x75;
  assign n8740 = n8404 & ~n8648;
  assign n8741 = n8740 ^ n8406;
  assign n8742 = n8741 ^ n8738;
  assign n8743 = n8739 & n8742;
  assign n8744 = n8743 ^ x75;
  assign n8745 = n8665 & n8744;
  assign n8746 = n8663 ^ x77;
  assign n8747 = x76 & n8660;
  assign n8748 = n8747 ^ n8663;
  assign n8749 = n8746 & ~n8748;
  assign n8750 = n8749 ^ x77;
  assign n8751 = ~n8745 & ~n8750;
  assign n8752 = n8751 ^ x78;
  assign n8753 = n8422 & ~n8648;
  assign n8754 = n8753 ^ n8424;
  assign n8755 = n8754 ^ n8751;
  assign n8756 = ~n8752 & n8755;
  assign n8757 = n8756 ^ x78;
  assign n8758 = n8757 ^ x79;
  assign n8759 = n8428 & ~n8648;
  assign n8760 = n8759 ^ n8430;
  assign n8761 = n8760 ^ n8757;
  assign n8762 = n8758 & ~n8761;
  assign n8763 = n8762 ^ x79;
  assign n8764 = n8763 ^ x80;
  assign n8765 = n8434 & ~n8648;
  assign n8766 = n8765 ^ n8436;
  assign n8767 = n8766 ^ n8763;
  assign n8768 = n8764 & ~n8767;
  assign n8769 = n8768 ^ x80;
  assign n8770 = n8769 ^ x81;
  assign n8771 = n8440 & ~n8648;
  assign n8772 = n8771 ^ n8442;
  assign n8773 = n8772 ^ n8769;
  assign n8774 = n8770 & ~n8773;
  assign n8775 = n8774 ^ x81;
  assign n8776 = n8775 ^ x82;
  assign n8777 = n8445 ^ x81;
  assign n8778 = ~n8648 & n8777;
  assign n8779 = n8778 ^ n8313;
  assign n8780 = n8779 ^ n8775;
  assign n8781 = n8776 & ~n8780;
  assign n8782 = n8781 ^ x82;
  assign n8783 = n8782 ^ x83;
  assign n8784 = n8445 ^ n8313;
  assign n8785 = n8777 & ~n8784;
  assign n8786 = n8785 ^ x81;
  assign n8787 = n8786 ^ x82;
  assign n8788 = ~n8648 & n8787;
  assign n8789 = n8788 ^ n8316;
  assign n8790 = n8789 ^ n8782;
  assign n8791 = n8783 & ~n8790;
  assign n8792 = n8791 ^ x83;
  assign n8793 = n8792 ^ x84;
  assign n8794 = ~n8453 & ~n8648;
  assign n8795 = n8794 ^ n8455;
  assign n8796 = n8795 ^ n8792;
  assign n8797 = n8793 & ~n8796;
  assign n8798 = n8797 ^ x84;
  assign n8799 = ~n8658 & ~n8798;
  assign n8800 = ~x85 & ~n8657;
  assign n8801 = n8465 & ~n8648;
  assign n8802 = n8801 ^ n8467;
  assign n8803 = ~x86 & ~n8802;
  assign n8804 = ~n8800 & ~n8803;
  assign n8805 = ~n8799 & n8804;
  assign n8806 = x86 & n8802;
  assign n8807 = ~n8805 & ~n8806;
  assign n8808 = n8807 ^ x87;
  assign n8809 = n8471 & ~n8648;
  assign n8810 = n8809 ^ n8473;
  assign n8811 = n8810 ^ n8807;
  assign n8812 = ~n8808 & n8811;
  assign n8813 = n8812 ^ x87;
  assign n8814 = n8655 & n8813;
  assign n8815 = n8653 ^ x89;
  assign n8816 = x88 & n8650;
  assign n8817 = n8816 ^ n8653;
  assign n8818 = n8815 & ~n8817;
  assign n8819 = n8818 ^ x89;
  assign n8820 = ~n8814 & ~n8819;
  assign n8821 = n8489 & ~n8648;
  assign n8822 = n8821 ^ n8491;
  assign n8823 = ~x90 & ~n8822;
  assign n8824 = n8495 & ~n8648;
  assign n8825 = n8824 ^ n8497;
  assign n8826 = ~x91 & ~n8825;
  assign n8827 = ~n8823 & ~n8826;
  assign n8828 = ~n8820 & n8827;
  assign n8829 = n8825 ^ x91;
  assign n8830 = x90 & n8822;
  assign n8831 = n8830 ^ n8825;
  assign n8832 = n8829 & ~n8831;
  assign n8833 = n8832 ^ x91;
  assign n8834 = ~n8828 & ~n8833;
  assign n8835 = n8834 ^ x92;
  assign n8836 = n8501 & ~n8648;
  assign n8837 = n8836 ^ n8503;
  assign n8838 = n8837 ^ n8834;
  assign n8839 = ~n8835 & n8838;
  assign n8840 = n8839 ^ x92;
  assign n8841 = n8840 ^ x93;
  assign n8842 = n8507 & ~n8648;
  assign n8843 = n8842 ^ n8509;
  assign n8844 = n8843 ^ n8840;
  assign n8845 = n8841 & ~n8844;
  assign n8846 = n8845 ^ x93;
  assign n8847 = n8846 ^ x94;
  assign n8848 = n8513 & ~n8648;
  assign n8849 = n8848 ^ n8515;
  assign n8850 = n8849 ^ n8846;
  assign n8851 = n8847 & ~n8850;
  assign n8852 = n8851 ^ x94;
  assign n8853 = n8852 ^ x95;
  assign n8854 = n8519 & ~n8648;
  assign n8855 = n8854 ^ n8521;
  assign n8856 = n8855 ^ n8852;
  assign n8857 = n8853 & ~n8856;
  assign n8858 = n8857 ^ x95;
  assign n8859 = n8858 ^ x96;
  assign n8860 = n8525 & ~n8648;
  assign n8861 = n8860 ^ n8528;
  assign n8862 = n8861 ^ n8858;
  assign n8863 = n8859 & ~n8862;
  assign n8864 = n8863 ^ x96;
  assign n8865 = n8864 ^ x97;
  assign n8866 = n8532 & ~n8648;
  assign n8867 = n8866 ^ n8536;
  assign n8868 = n8867 ^ n8864;
  assign n8869 = n8865 & ~n8868;
  assign n8870 = n8869 ^ x97;
  assign n8871 = n8870 ^ x98;
  assign n8872 = n8540 & ~n8648;
  assign n8873 = n8872 ^ n8542;
  assign n8874 = n8873 ^ n8870;
  assign n8875 = n8871 & ~n8874;
  assign n8876 = n8875 ^ x98;
  assign n8877 = n8876 ^ x99;
  assign n8878 = n8546 & ~n8648;
  assign n8879 = n8878 ^ n8548;
  assign n8880 = n8879 ^ n8876;
  assign n8881 = n8877 & ~n8880;
  assign n8882 = n8881 ^ x99;
  assign n8883 = n8882 ^ x100;
  assign n8884 = n8552 & ~n8648;
  assign n8885 = n8884 ^ n8554;
  assign n8886 = n8885 ^ n8882;
  assign n8887 = n8883 & ~n8886;
  assign n8888 = n8887 ^ x100;
  assign n8889 = n8888 ^ x101;
  assign n8890 = n8558 & ~n8648;
  assign n8891 = n8890 ^ n8560;
  assign n8892 = n8891 ^ n8888;
  assign n8893 = n8889 & ~n8892;
  assign n8894 = n8893 ^ x101;
  assign n8895 = n8894 ^ x102;
  assign n8896 = n8564 & ~n8648;
  assign n8897 = n8896 ^ n8567;
  assign n8898 = n8897 ^ n8894;
  assign n8899 = n8895 & ~n8898;
  assign n8900 = n8899 ^ x102;
  assign n8901 = n8900 ^ x103;
  assign n8902 = n8571 & ~n8648;
  assign n8903 = n8902 ^ n8575;
  assign n8904 = n8903 ^ n8900;
  assign n8905 = n8901 & ~n8904;
  assign n8906 = n8905 ^ x103;
  assign n8907 = n8906 ^ x104;
  assign n8908 = n8579 & ~n8648;
  assign n8909 = n8908 ^ n8581;
  assign n8910 = n8909 ^ n8906;
  assign n8911 = n8907 & ~n8910;
  assign n8912 = n8911 ^ x104;
  assign n8913 = n8912 ^ x105;
  assign n8914 = n8584 ^ x104;
  assign n8915 = ~n8648 & n8914;
  assign n8916 = n8915 ^ n8306;
  assign n8917 = n8916 ^ n8912;
  assign n8918 = n8913 & ~n8917;
  assign n8919 = n8918 ^ x105;
  assign n8920 = n8919 ^ x106;
  assign n8921 = n8584 ^ n8306;
  assign n8922 = n8914 & ~n8921;
  assign n8923 = n8922 ^ x104;
  assign n8924 = n8923 ^ x105;
  assign n8925 = ~n8648 & n8924;
  assign n8926 = n8925 ^ n8309;
  assign n8927 = n8926 ^ n8919;
  assign n8928 = n8920 & ~n8927;
  assign n8929 = n8928 ^ x106;
  assign n8930 = n8929 ^ x107;
  assign n8931 = ~n8592 & ~n8648;
  assign n8932 = n8931 ^ n8594;
  assign n8933 = n8932 ^ n8929;
  assign n8934 = n8930 & ~n8933;
  assign n8935 = n8934 ^ x107;
  assign n8936 = n8935 ^ x108;
  assign n8937 = n8598 & ~n8648;
  assign n8938 = n8937 ^ n8601;
  assign n8939 = n8938 ^ n8935;
  assign n8940 = n8936 & ~n8939;
  assign n8941 = n8940 ^ x108;
  assign n8942 = n8941 ^ x109;
  assign n8943 = n8605 & ~n8648;
  assign n8944 = n8943 ^ n8609;
  assign n8945 = n8944 ^ n8941;
  assign n8946 = n8942 & ~n8945;
  assign n8947 = n8946 ^ x109;
  assign n8948 = n8947 ^ x110;
  assign n8949 = n8612 ^ x109;
  assign n8950 = ~n8648 & n8949;
  assign n8951 = n8950 ^ n8303;
  assign n8952 = n8951 ^ n8947;
  assign n8953 = n8948 & ~n8952;
  assign n8954 = n8953 ^ x110;
  assign n8955 = n8954 ^ x111;
  assign n8956 = ~n8613 & ~n8617;
  assign n8957 = n8956 ^ x110;
  assign n8958 = ~n8648 & ~n8957;
  assign n8959 = n8958 ^ n8615;
  assign n8960 = n8959 ^ n8954;
  assign n8961 = n8955 & ~n8960;
  assign n8962 = n8961 ^ x111;
  assign n8963 = n8962 ^ x112;
  assign n8964 = n8621 ^ x111;
  assign n8965 = ~n8648 & n8964;
  assign n8966 = n8965 ^ n8624;
  assign n8967 = n8966 ^ n8962;
  assign n8968 = n8963 & n8967;
  assign n8969 = n8968 ^ x112;
  assign n8970 = n8969 ^ x113;
  assign n8971 = n8635 & n8970;
  assign n8972 = n8634 & ~n8971;
  assign n8973 = ~n8634 & n8969;
  assign n8974 = ~x113 & ~n8973;
  assign n8975 = n7666 & ~n8969;
  assign n8976 = ~n8974 & ~n8975;
  assign n8977 = n8635 & ~n8976;
  assign n8978 = n8913 & n8977;
  assign n8979 = n8978 ^ n8916;
  assign n8980 = ~x106 & ~n8979;
  assign n8981 = n8920 & n8977;
  assign n8982 = n8981 ^ n8926;
  assign n8983 = ~x107 & ~n8982;
  assign n8984 = ~n8980 & ~n8983;
  assign n8985 = n8853 & n8977;
  assign n8986 = n8985 ^ n8855;
  assign n8987 = ~x96 & ~n8986;
  assign n8988 = n8783 & n8977;
  assign n8989 = n8988 ^ n8789;
  assign n8990 = ~x84 & ~n8989;
  assign n8991 = n8793 & n8977;
  assign n8992 = n8991 ^ n8795;
  assign n8993 = ~x85 & ~n8992;
  assign n8994 = ~n8990 & ~n8993;
  assign n8995 = x64 & n8977;
  assign n8996 = ~x14 & x65;
  assign n8997 = ~n8995 & n8996;
  assign n8998 = n8977 ^ n8667;
  assign n8999 = n8997 & ~n8998;
  assign n9000 = ~n8667 & ~n8977;
  assign n9001 = x14 & ~x65;
  assign n9002 = ~x13 & x64;
  assign n9003 = ~n9001 & n9002;
  assign n9004 = n9000 & n9003;
  assign n9005 = ~x66 & ~n9004;
  assign n9006 = ~n8999 & n9005;
  assign n9007 = x13 & n9001;
  assign n9008 = n9007 ^ x14;
  assign n9009 = ~n8668 & n9008;
  assign n9010 = n8977 & n9009;
  assign n9011 = ~x13 & n8996;
  assign n9012 = ~n8667 & n9011;
  assign n9013 = ~n9010 & ~n9012;
  assign n9014 = x64 & ~n9013;
  assign n9015 = n9006 & ~n9014;
  assign n9016 = ~x65 & ~n8669;
  assign n9017 = ~n9002 & n9016;
  assign n9018 = n8977 & ~n9017;
  assign n9019 = ~n8996 & ~n9003;
  assign n9020 = n8667 & n9019;
  assign n9021 = ~n9018 & n9020;
  assign n9022 = ~x13 & x65;
  assign n9023 = n8669 & ~n9022;
  assign n9024 = ~n8668 & n9023;
  assign n9025 = x14 & n202;
  assign n9026 = ~n8667 & n9025;
  assign n9027 = ~n9024 & ~n9026;
  assign n9028 = n8977 & ~n9027;
  assign n9029 = ~n9021 & ~n9028;
  assign n9030 = ~n9015 & n9029;
  assign n9031 = n9030 ^ x67;
  assign n9032 = n8673 & n8977;
  assign n9033 = n9032 ^ n8686;
  assign n9034 = n9033 ^ n9030;
  assign n9035 = n9031 & n9034;
  assign n9036 = n9035 ^ x67;
  assign n9037 = n9036 ^ x68;
  assign n9038 = n8690 & n8977;
  assign n9039 = n9038 ^ n8693;
  assign n9040 = n9039 ^ n9036;
  assign n9041 = n9037 & ~n9040;
  assign n9042 = n9041 ^ x68;
  assign n9043 = n9042 ^ x69;
  assign n9044 = n8697 & n8977;
  assign n9045 = n9044 ^ n8699;
  assign n9046 = n9045 ^ n9042;
  assign n9047 = n9043 & n9046;
  assign n9048 = n9047 ^ x69;
  assign n9049 = n9048 ^ x70;
  assign n9050 = n8703 & n8977;
  assign n9051 = n9050 ^ n8705;
  assign n9052 = n9051 ^ n9048;
  assign n9053 = n9049 & ~n9052;
  assign n9054 = n9053 ^ x70;
  assign n9055 = n9054 ^ x71;
  assign n9056 = n8709 & n8977;
  assign n9057 = n9056 ^ n8711;
  assign n9058 = n9057 ^ n9054;
  assign n9059 = n9055 & ~n9058;
  assign n9060 = n9059 ^ x71;
  assign n9061 = n9060 ^ x72;
  assign n9062 = n8715 & n8977;
  assign n9063 = n9062 ^ n8717;
  assign n9064 = n9063 ^ n9060;
  assign n9065 = n9061 & n9064;
  assign n9066 = n9065 ^ x72;
  assign n9067 = n9066 ^ x73;
  assign n9068 = n8721 & n8977;
  assign n9069 = n9068 ^ n8723;
  assign n9070 = n9069 ^ n9066;
  assign n9071 = n9067 & ~n9070;
  assign n9072 = n9071 ^ x73;
  assign n9073 = n9072 ^ x74;
  assign n9074 = n8727 & n8977;
  assign n9075 = n9074 ^ n8729;
  assign n9076 = n9075 ^ n9072;
  assign n9077 = n9073 & n9076;
  assign n9078 = n9077 ^ x74;
  assign n9079 = n9078 ^ x75;
  assign n9080 = n8733 & n8977;
  assign n9081 = n9080 ^ n8735;
  assign n9082 = n9081 ^ n9078;
  assign n9083 = n9079 & ~n9082;
  assign n9084 = n9083 ^ x75;
  assign n9085 = n9084 ^ x76;
  assign n9086 = n8739 & n8977;
  assign n9087 = n9086 ^ n8741;
  assign n9088 = n9087 ^ n9084;
  assign n9089 = n9085 & n9088;
  assign n9090 = n9089 ^ x76;
  assign n9091 = n9090 ^ x77;
  assign n9092 = n8744 ^ x76;
  assign n9093 = n8977 & n9092;
  assign n9094 = n9093 ^ n8660;
  assign n9095 = n9094 ^ n9090;
  assign n9096 = n9091 & ~n9095;
  assign n9097 = n9096 ^ x77;
  assign n9098 = n9097 ^ x78;
  assign n9099 = n8744 ^ n8660;
  assign n9100 = n9092 & ~n9099;
  assign n9101 = n9100 ^ x76;
  assign n9102 = n9101 ^ x77;
  assign n9103 = n8977 & n9102;
  assign n9104 = n9103 ^ n8663;
  assign n9105 = n9104 ^ n9097;
  assign n9106 = n9098 & ~n9105;
  assign n9107 = n9106 ^ x78;
  assign n9108 = n9107 ^ x79;
  assign n9109 = ~n8752 & n8977;
  assign n9110 = n9109 ^ n8754;
  assign n9111 = n9110 ^ n9107;
  assign n9112 = n9108 & ~n9111;
  assign n9113 = n9112 ^ x79;
  assign n9114 = n9113 ^ x80;
  assign n9115 = n8758 & n8977;
  assign n9116 = n9115 ^ n8760;
  assign n9117 = n9116 ^ n9113;
  assign n9118 = n9114 & ~n9117;
  assign n9119 = n9118 ^ x80;
  assign n9120 = n9119 ^ x81;
  assign n9121 = n8764 & n8977;
  assign n9122 = n9121 ^ n8766;
  assign n9123 = n9122 ^ n9119;
  assign n9124 = n9120 & ~n9123;
  assign n9125 = n9124 ^ x81;
  assign n9126 = n9125 ^ x82;
  assign n9127 = n8770 & n8977;
  assign n9128 = n9127 ^ n8772;
  assign n9129 = n9128 ^ n9125;
  assign n9130 = n9126 & ~n9129;
  assign n9131 = n9130 ^ x82;
  assign n9132 = n9131 ^ x83;
  assign n9133 = n8776 & n8977;
  assign n9134 = n9133 ^ n8779;
  assign n9135 = n9134 ^ n9131;
  assign n9136 = n9132 & ~n9135;
  assign n9137 = n9136 ^ x83;
  assign n9138 = n8994 & n9137;
  assign n9139 = n8992 ^ x85;
  assign n9140 = x84 & n8989;
  assign n9141 = n9140 ^ n8992;
  assign n9142 = n9139 & ~n9141;
  assign n9143 = n9142 ^ x85;
  assign n9144 = ~n9138 & ~n9143;
  assign n9145 = n9144 ^ x86;
  assign n9146 = n8798 ^ x85;
  assign n9147 = n8977 & n9146;
  assign n9148 = n9147 ^ n8657;
  assign n9149 = n9148 ^ n9144;
  assign n9150 = ~n9145 & n9149;
  assign n9151 = n9150 ^ x86;
  assign n9152 = n9151 ^ x87;
  assign n9153 = ~n8799 & ~n8800;
  assign n9154 = n9153 ^ x86;
  assign n9155 = n8977 & n9154;
  assign n9156 = n9155 ^ n8802;
  assign n9157 = n9156 ^ n9151;
  assign n9158 = n9152 & ~n9157;
  assign n9159 = n9158 ^ x87;
  assign n9160 = n9159 ^ x88;
  assign n9161 = ~n8808 & n8977;
  assign n9162 = n9161 ^ n8810;
  assign n9163 = n9162 ^ n9159;
  assign n9164 = n9160 & ~n9163;
  assign n9165 = n9164 ^ x88;
  assign n9166 = n9165 ^ x89;
  assign n9167 = n8813 ^ x88;
  assign n9168 = n8977 & n9167;
  assign n9169 = n9168 ^ n8650;
  assign n9170 = n9169 ^ n9165;
  assign n9171 = n9166 & ~n9170;
  assign n9172 = n9171 ^ x89;
  assign n9173 = n9172 ^ x90;
  assign n9174 = n8813 ^ n8650;
  assign n9175 = n9167 & ~n9174;
  assign n9176 = n9175 ^ x88;
  assign n9177 = n9176 ^ x89;
  assign n9178 = n8977 & n9177;
  assign n9179 = n9178 ^ n8653;
  assign n9180 = n9179 ^ n9172;
  assign n9181 = n9173 & ~n9180;
  assign n9182 = n9181 ^ x90;
  assign n9183 = n9182 ^ x91;
  assign n9184 = n8820 ^ x90;
  assign n9185 = n8977 & ~n9184;
  assign n9186 = n9185 ^ n8822;
  assign n9187 = n9186 ^ n9182;
  assign n9188 = n9183 & ~n9187;
  assign n9189 = n9188 ^ x91;
  assign n9190 = n9189 ^ x92;
  assign n9191 = n8822 ^ n8820;
  assign n9192 = ~n9184 & n9191;
  assign n9193 = n9192 ^ x90;
  assign n9194 = n9193 ^ x91;
  assign n9195 = n8977 & n9194;
  assign n9196 = n9195 ^ n8825;
  assign n9197 = n9196 ^ n9189;
  assign n9198 = n9190 & ~n9197;
  assign n9199 = n9198 ^ x92;
  assign n9200 = n9199 ^ x93;
  assign n9201 = ~n8835 & n8977;
  assign n9202 = n9201 ^ n8837;
  assign n9203 = n9202 ^ n9199;
  assign n9204 = n9200 & ~n9203;
  assign n9205 = n9204 ^ x93;
  assign n9206 = n9205 ^ x94;
  assign n9207 = n8841 & n8977;
  assign n9208 = n9207 ^ n8843;
  assign n9209 = n9208 ^ n9205;
  assign n9210 = n9206 & ~n9209;
  assign n9211 = n9210 ^ x94;
  assign n9212 = n9211 ^ x95;
  assign n9213 = n8847 & n8977;
  assign n9214 = n9213 ^ n8849;
  assign n9215 = n9214 ^ n9211;
  assign n9216 = n9212 & ~n9215;
  assign n9217 = n9216 ^ x95;
  assign n9218 = ~n8987 & n9217;
  assign n9219 = n8859 & n8977;
  assign n9220 = n9219 ^ n8861;
  assign n9221 = x97 & n9220;
  assign n9222 = x96 & n8986;
  assign n9223 = ~n9221 & ~n9222;
  assign n9224 = ~n9218 & n9223;
  assign n9225 = ~x97 & ~n9220;
  assign n9226 = ~n9224 & ~n9225;
  assign n9227 = n9226 ^ x98;
  assign n9228 = n8865 & n8977;
  assign n9229 = n9228 ^ n8867;
  assign n9230 = n9229 ^ n9226;
  assign n9231 = n9227 & ~n9230;
  assign n9232 = n9231 ^ x98;
  assign n9233 = n9232 ^ x99;
  assign n9234 = n8871 & n8977;
  assign n9235 = n9234 ^ n8873;
  assign n9236 = n9235 ^ n9232;
  assign n9237 = n9233 & ~n9236;
  assign n9238 = n9237 ^ x99;
  assign n9239 = n9238 ^ x100;
  assign n9240 = n8877 & n8977;
  assign n9241 = n9240 ^ n8879;
  assign n9242 = n9241 ^ n9238;
  assign n9243 = n9239 & ~n9242;
  assign n9244 = n9243 ^ x100;
  assign n9245 = n9244 ^ x101;
  assign n9246 = n8883 & n8977;
  assign n9247 = n9246 ^ n8885;
  assign n9248 = n9247 ^ n9244;
  assign n9249 = n9245 & ~n9248;
  assign n9250 = n9249 ^ x101;
  assign n9251 = n9250 ^ x102;
  assign n9252 = n8889 & n8977;
  assign n9253 = n9252 ^ n8891;
  assign n9254 = n9253 ^ n9250;
  assign n9255 = n9251 & ~n9254;
  assign n9256 = n9255 ^ x102;
  assign n9257 = n9256 ^ x103;
  assign n9258 = n8895 & n8977;
  assign n9259 = n9258 ^ n8897;
  assign n9260 = n9259 ^ n9256;
  assign n9261 = n9257 & ~n9260;
  assign n9262 = n9261 ^ x103;
  assign n9263 = n9262 ^ x104;
  assign n9264 = n8901 & n8977;
  assign n9265 = n9264 ^ n8903;
  assign n9266 = n9265 ^ n9262;
  assign n9267 = n9263 & ~n9266;
  assign n9268 = n9267 ^ x104;
  assign n9269 = n9268 ^ x105;
  assign n9270 = n8907 & n8977;
  assign n9271 = n9270 ^ n8909;
  assign n9272 = n9271 ^ n9268;
  assign n9273 = n9269 & ~n9272;
  assign n9274 = n9273 ^ x105;
  assign n9275 = n8984 & n9274;
  assign n9276 = n8982 ^ x107;
  assign n9277 = x106 & n8979;
  assign n9278 = n9277 ^ n8982;
  assign n9279 = n9276 & ~n9278;
  assign n9280 = n9279 ^ x107;
  assign n9281 = ~n9275 & ~n9280;
  assign n9282 = n9281 ^ x108;
  assign n9283 = n8930 & n8977;
  assign n9284 = n9283 ^ n8932;
  assign n9285 = n9284 ^ n9281;
  assign n9286 = ~n9282 & n9285;
  assign n9287 = n9286 ^ x108;
  assign n9288 = n9287 ^ x109;
  assign n9289 = n8936 & n8977;
  assign n9290 = n9289 ^ n8938;
  assign n9291 = n9290 ^ n9287;
  assign n9292 = n9288 & ~n9291;
  assign n9293 = n9292 ^ x109;
  assign n9294 = n9293 ^ x110;
  assign n9295 = n8942 & n8977;
  assign n9296 = n9295 ^ n8944;
  assign n9297 = n9296 ^ n9293;
  assign n9298 = n9294 & ~n9297;
  assign n9299 = n9298 ^ x110;
  assign n9300 = n9299 ^ x111;
  assign n9301 = n8948 & n8977;
  assign n9302 = n9301 ^ n8951;
  assign n9303 = n9302 ^ n9299;
  assign n9304 = n9300 & ~n9303;
  assign n9305 = n9304 ^ x111;
  assign n9306 = n9305 ^ x112;
  assign n9307 = n8955 & n8977;
  assign n9308 = n9307 ^ n8959;
  assign n9309 = n9308 ^ n9305;
  assign n9310 = n9306 & ~n9309;
  assign n9311 = n9310 ^ x112;
  assign n9312 = n9311 ^ x113;
  assign n9313 = n8963 & n8977;
  assign n9314 = n9313 ^ n8966;
  assign n9315 = n9314 ^ n9311;
  assign n9316 = n9312 & n9315;
  assign n9317 = n9316 ^ x113;
  assign n9318 = n9317 ^ x114;
  assign n9319 = n141 & n9318;
  assign n9320 = n8972 & ~n9319;
  assign n9321 = ~x120 & n135;
  assign n9322 = ~x119 & n9321;
  assign n9323 = ~x118 & n9322;
  assign n9324 = ~x117 & n9323;
  assign n9325 = n9317 ^ n8972;
  assign n9326 = n9318 & n9325;
  assign n9327 = n9326 ^ x114;
  assign n9328 = n141 & ~n9327;
  assign n9329 = n9312 & n9328;
  assign n9330 = n9329 ^ n9314;
  assign n9331 = ~x114 & n9330;
  assign n9332 = ~x115 & n9320;
  assign n9333 = ~n9331 & ~n9332;
  assign n9334 = n9233 & n9328;
  assign n9335 = n9334 ^ n9235;
  assign n9336 = ~x100 & ~n9335;
  assign n9337 = n9239 & n9328;
  assign n9338 = n9337 ^ n9241;
  assign n9339 = ~x101 & ~n9338;
  assign n9340 = ~n9336 & ~n9339;
  assign n9341 = n9073 & n9328;
  assign n9342 = n9341 ^ n9075;
  assign n9343 = ~x75 & n9342;
  assign n9344 = n9079 & n9328;
  assign n9345 = n9344 ^ n9081;
  assign n9346 = ~x76 & ~n9345;
  assign n9347 = ~n9343 & ~n9346;
  assign n9348 = x65 & n141;
  assign n9349 = ~n8977 & n9348;
  assign n9350 = ~n9327 & n9349;
  assign n9351 = ~x65 & n8977;
  assign n9352 = x64 & n9351;
  assign n9353 = ~n9350 & ~n9352;
  assign n9354 = x13 & ~n9353;
  assign n9355 = n8977 ^ x65;
  assign n9356 = n341 & ~n9355;
  assign n9357 = x13 & n9356;
  assign n9358 = n9357 ^ n340;
  assign n9359 = n9328 & n9358;
  assign n9360 = n9359 ^ n8995;
  assign n9361 = ~n9354 & ~n9360;
  assign n9362 = n9361 ^ x14;
  assign n9363 = n9362 ^ x66;
  assign n9364 = x64 & n9328;
  assign n9365 = x13 & ~x65;
  assign n9366 = x12 & n9365;
  assign n9367 = n9366 ^ x13;
  assign n9368 = n9364 & n9367;
  assign n9369 = ~x12 & n9002;
  assign n9370 = ~n9022 & ~n9369;
  assign n9371 = ~n9328 & ~n9370;
  assign n9372 = x12 & x64;
  assign n9373 = x65 & ~n9372;
  assign n9374 = x13 & ~x64;
  assign n9375 = n9373 & ~n9374;
  assign n9376 = ~n9371 & ~n9375;
  assign n9377 = ~n9368 & n9376;
  assign n9378 = n9377 ^ n9362;
  assign n9379 = n9363 & n9378;
  assign n9380 = n9379 ^ x66;
  assign n9381 = n9380 ^ x67;
  assign n9385 = n9003 & ~n9351;
  assign n9386 = n9008 ^ n8996;
  assign n9387 = n8995 & n9386;
  assign n9388 = n9387 ^ n8996;
  assign n9389 = ~n9385 & ~n9388;
  assign n9390 = n9389 ^ x66;
  assign n9391 = n9328 & ~n9390;
  assign n9382 = n8669 ^ x65;
  assign n9383 = n8977 & n9382;
  assign n9384 = n9383 ^ n8667;
  assign n9392 = n9391 ^ n9384;
  assign n9393 = n9392 ^ n9380;
  assign n9394 = n9381 & n9393;
  assign n9395 = n9394 ^ x67;
  assign n9396 = n9395 ^ x68;
  assign n9397 = n9031 & n9328;
  assign n9398 = n9397 ^ n9033;
  assign n9399 = n9398 ^ n9395;
  assign n9400 = n9396 & n9399;
  assign n9401 = n9400 ^ x68;
  assign n9402 = n9401 ^ x69;
  assign n9403 = n9037 & n9328;
  assign n9404 = n9403 ^ n9039;
  assign n9405 = n9404 ^ n9401;
  assign n9406 = n9402 & ~n9405;
  assign n9407 = n9406 ^ x69;
  assign n9408 = n9407 ^ x70;
  assign n9409 = n9043 & n9328;
  assign n9410 = n9409 ^ n9045;
  assign n9411 = n9410 ^ n9407;
  assign n9412 = n9408 & n9411;
  assign n9413 = n9412 ^ x70;
  assign n9414 = n9413 ^ x71;
  assign n9415 = n9049 & n9328;
  assign n9416 = n9415 ^ n9051;
  assign n9417 = n9416 ^ n9413;
  assign n9418 = n9414 & ~n9417;
  assign n9419 = n9418 ^ x71;
  assign n9420 = n9419 ^ x72;
  assign n9421 = n9055 & n9328;
  assign n9422 = n9421 ^ n9057;
  assign n9423 = n9422 ^ n9419;
  assign n9424 = n9420 & ~n9423;
  assign n9425 = n9424 ^ x72;
  assign n9426 = n9425 ^ x73;
  assign n9427 = n9061 & n9328;
  assign n9428 = n9427 ^ n9063;
  assign n9429 = n9428 ^ n9425;
  assign n9430 = n9426 & n9429;
  assign n9431 = n9430 ^ x73;
  assign n9432 = n9431 ^ x74;
  assign n9433 = n9067 & n9328;
  assign n9434 = n9433 ^ n9069;
  assign n9435 = n9434 ^ n9431;
  assign n9436 = n9432 & ~n9435;
  assign n9437 = n9436 ^ x74;
  assign n9438 = n9347 & n9437;
  assign n9439 = n9345 ^ x76;
  assign n9440 = x75 & ~n9342;
  assign n9441 = n9440 ^ n9345;
  assign n9442 = n9439 & ~n9441;
  assign n9443 = n9442 ^ x76;
  assign n9444 = ~n9438 & ~n9443;
  assign n9445 = n9444 ^ x77;
  assign n9446 = n9085 & n9328;
  assign n9447 = n9446 ^ n9087;
  assign n9448 = n9447 ^ n9444;
  assign n9449 = ~n9445 & ~n9448;
  assign n9450 = n9449 ^ x77;
  assign n9451 = n9450 ^ x78;
  assign n9452 = n9091 & n9328;
  assign n9453 = n9452 ^ n9094;
  assign n9454 = n9453 ^ n9450;
  assign n9455 = n9451 & ~n9454;
  assign n9456 = n9455 ^ x78;
  assign n9457 = n9456 ^ x79;
  assign n9458 = n9098 & n9328;
  assign n9459 = n9458 ^ n9104;
  assign n9460 = n9459 ^ n9456;
  assign n9461 = n9457 & ~n9460;
  assign n9462 = n9461 ^ x79;
  assign n9463 = n9462 ^ x80;
  assign n9464 = n9108 & n9328;
  assign n9465 = n9464 ^ n9110;
  assign n9466 = n9465 ^ n9462;
  assign n9467 = n9463 & ~n9466;
  assign n9468 = n9467 ^ x80;
  assign n9469 = n9468 ^ x81;
  assign n9470 = n9114 & n9328;
  assign n9471 = n9470 ^ n9116;
  assign n9472 = n9471 ^ n9468;
  assign n9473 = n9469 & ~n9472;
  assign n9474 = n9473 ^ x81;
  assign n9475 = n9474 ^ x82;
  assign n9476 = n9120 & n9328;
  assign n9477 = n9476 ^ n9122;
  assign n9478 = n9477 ^ n9474;
  assign n9479 = n9475 & ~n9478;
  assign n9480 = n9479 ^ x82;
  assign n9481 = n9480 ^ x83;
  assign n9482 = n9126 & n9328;
  assign n9483 = n9482 ^ n9128;
  assign n9484 = n9483 ^ n9480;
  assign n9485 = n9481 & ~n9484;
  assign n9486 = n9485 ^ x83;
  assign n9487 = n9486 ^ x84;
  assign n9488 = n9132 & n9328;
  assign n9489 = n9488 ^ n9134;
  assign n9490 = n9489 ^ n9486;
  assign n9491 = n9487 & ~n9490;
  assign n9492 = n9491 ^ x84;
  assign n9493 = n9492 ^ x85;
  assign n9494 = n9137 ^ x84;
  assign n9495 = n9328 & n9494;
  assign n9496 = n9495 ^ n8989;
  assign n9497 = n9496 ^ n9492;
  assign n9498 = n9493 & ~n9497;
  assign n9499 = n9498 ^ x85;
  assign n9500 = n9499 ^ x86;
  assign n9501 = n9137 ^ n8989;
  assign n9502 = n9494 & ~n9501;
  assign n9503 = n9502 ^ x84;
  assign n9504 = n9503 ^ x85;
  assign n9505 = n9328 & n9504;
  assign n9506 = n9505 ^ n8992;
  assign n9507 = n9506 ^ n9499;
  assign n9508 = n9500 & ~n9507;
  assign n9509 = n9508 ^ x86;
  assign n9510 = n9509 ^ x87;
  assign n9511 = ~n9145 & n9328;
  assign n9512 = n9511 ^ n9148;
  assign n9513 = n9512 ^ n9509;
  assign n9514 = n9510 & ~n9513;
  assign n9515 = n9514 ^ x87;
  assign n9516 = n9515 ^ x88;
  assign n9517 = n9152 & n9328;
  assign n9518 = n9517 ^ n9156;
  assign n9519 = n9518 ^ n9515;
  assign n9520 = n9516 & ~n9519;
  assign n9521 = n9520 ^ x88;
  assign n9522 = n9521 ^ x89;
  assign n9523 = n9160 & n9328;
  assign n9524 = n9523 ^ n9162;
  assign n9525 = n9524 ^ n9521;
  assign n9526 = n9522 & ~n9525;
  assign n9527 = n9526 ^ x89;
  assign n9528 = n9527 ^ x90;
  assign n9529 = n9166 & n9328;
  assign n9530 = n9529 ^ n9169;
  assign n9531 = n9530 ^ n9527;
  assign n9532 = n9528 & ~n9531;
  assign n9533 = n9532 ^ x90;
  assign n9534 = n9533 ^ x91;
  assign n9535 = n9173 & n9328;
  assign n9536 = n9535 ^ n9179;
  assign n9537 = n9536 ^ n9533;
  assign n9538 = n9534 & ~n9537;
  assign n9539 = n9538 ^ x91;
  assign n9540 = n9539 ^ x92;
  assign n9541 = n9183 & n9328;
  assign n9542 = n9541 ^ n9186;
  assign n9543 = n9542 ^ n9539;
  assign n9544 = n9540 & ~n9543;
  assign n9545 = n9544 ^ x92;
  assign n9546 = n9545 ^ x93;
  assign n9547 = n9190 & n9328;
  assign n9548 = n9547 ^ n9196;
  assign n9549 = n9548 ^ n9545;
  assign n9550 = n9546 & ~n9549;
  assign n9551 = n9550 ^ x93;
  assign n9552 = n9551 ^ x94;
  assign n9553 = n9200 & n9328;
  assign n9554 = n9553 ^ n9202;
  assign n9555 = n9554 ^ n9551;
  assign n9556 = n9552 & ~n9555;
  assign n9557 = n9556 ^ x94;
  assign n9558 = n9557 ^ x95;
  assign n9559 = n9206 & n9328;
  assign n9560 = n9559 ^ n9208;
  assign n9561 = n9560 ^ n9557;
  assign n9562 = n9558 & ~n9561;
  assign n9563 = n9562 ^ x95;
  assign n9564 = n9563 ^ x96;
  assign n9565 = n9212 & n9328;
  assign n9566 = n9565 ^ n9214;
  assign n9567 = n9566 ^ n9563;
  assign n9568 = n9564 & ~n9567;
  assign n9569 = n9568 ^ x96;
  assign n9570 = n9569 ^ x97;
  assign n9571 = n9217 ^ x96;
  assign n9572 = n9328 & n9571;
  assign n9573 = n9572 ^ n8986;
  assign n9574 = n9573 ^ n9569;
  assign n9575 = n9570 & ~n9574;
  assign n9576 = n9575 ^ x97;
  assign n9577 = n9576 ^ x98;
  assign n9578 = ~n9218 & ~n9222;
  assign n9579 = n9578 ^ x97;
  assign n9580 = n9328 & ~n9579;
  assign n9581 = n9580 ^ n9220;
  assign n9582 = n9581 ^ n9576;
  assign n9583 = n9577 & ~n9582;
  assign n9584 = n9583 ^ x98;
  assign n9585 = n9584 ^ x99;
  assign n9586 = n9227 & n9328;
  assign n9587 = n9586 ^ n9229;
  assign n9588 = n9587 ^ n9584;
  assign n9589 = n9585 & ~n9588;
  assign n9590 = n9589 ^ x99;
  assign n9591 = n9340 & n9590;
  assign n9592 = n9338 ^ x101;
  assign n9593 = x100 & n9335;
  assign n9594 = n9593 ^ n9338;
  assign n9595 = n9592 & ~n9594;
  assign n9596 = n9595 ^ x101;
  assign n9597 = ~n9591 & ~n9596;
  assign n9598 = n9597 ^ x102;
  assign n9599 = n9245 & n9328;
  assign n9600 = n9599 ^ n9247;
  assign n9601 = n9600 ^ n9597;
  assign n9602 = ~n9598 & n9601;
  assign n9603 = n9602 ^ x102;
  assign n9604 = n9603 ^ x103;
  assign n9605 = n9251 & n9328;
  assign n9606 = n9605 ^ n9253;
  assign n9607 = n9606 ^ n9603;
  assign n9608 = n9604 & ~n9607;
  assign n9609 = n9608 ^ x103;
  assign n9610 = n9609 ^ x104;
  assign n9611 = n9257 & n9328;
  assign n9612 = n9611 ^ n9259;
  assign n9613 = n9612 ^ n9609;
  assign n9614 = n9610 & ~n9613;
  assign n9615 = n9614 ^ x104;
  assign n9616 = n9615 ^ x105;
  assign n9617 = n9263 & n9328;
  assign n9618 = n9617 ^ n9265;
  assign n9619 = n9618 ^ n9615;
  assign n9620 = n9616 & ~n9619;
  assign n9621 = n9620 ^ x105;
  assign n9622 = n9621 ^ x106;
  assign n9623 = n9269 & n9328;
  assign n9624 = n9623 ^ n9271;
  assign n9625 = n9624 ^ n9621;
  assign n9626 = n9622 & ~n9625;
  assign n9627 = n9626 ^ x106;
  assign n9628 = n9627 ^ x107;
  assign n9629 = n9274 ^ x106;
  assign n9630 = n9328 & n9629;
  assign n9631 = n9630 ^ n8979;
  assign n9632 = n9631 ^ n9627;
  assign n9633 = n9628 & ~n9632;
  assign n9634 = n9633 ^ x107;
  assign n9635 = n9634 ^ x108;
  assign n9636 = n9274 ^ n8979;
  assign n9637 = n9629 & ~n9636;
  assign n9638 = n9637 ^ x106;
  assign n9639 = n9638 ^ x107;
  assign n9640 = n9328 & n9639;
  assign n9641 = n9640 ^ n8982;
  assign n9642 = n9641 ^ n9634;
  assign n9643 = n9635 & ~n9642;
  assign n9644 = n9643 ^ x108;
  assign n9645 = n9644 ^ x109;
  assign n9646 = ~n9282 & n9328;
  assign n9647 = n9646 ^ n9284;
  assign n9648 = n9647 ^ n9644;
  assign n9649 = n9645 & ~n9648;
  assign n9650 = n9649 ^ x109;
  assign n9651 = n9650 ^ x110;
  assign n9652 = n9288 & n9328;
  assign n9653 = n9652 ^ n9290;
  assign n9654 = n9653 ^ n9650;
  assign n9655 = n9651 & ~n9654;
  assign n9656 = n9655 ^ x110;
  assign n9657 = n9656 ^ x111;
  assign n9658 = n9294 & n9328;
  assign n9659 = n9658 ^ n9296;
  assign n9660 = n9659 ^ n9656;
  assign n9661 = n9657 & ~n9660;
  assign n9662 = n9661 ^ x111;
  assign n9663 = n9662 ^ x112;
  assign n9664 = n9300 & n9328;
  assign n9665 = n9664 ^ n9302;
  assign n9666 = n9665 ^ n9662;
  assign n9667 = n9663 & ~n9666;
  assign n9668 = n9667 ^ x112;
  assign n9669 = n9668 ^ x113;
  assign n9670 = n9306 & n9328;
  assign n9671 = n9670 ^ n9308;
  assign n9672 = n9671 ^ n9668;
  assign n9673 = n9669 & ~n9672;
  assign n9674 = n9673 ^ x113;
  assign n9675 = n9333 & n9674;
  assign n9676 = x114 & ~n9330;
  assign n9677 = ~n9332 & n9676;
  assign n9678 = x115 & ~n9320;
  assign n9679 = n140 & ~n9678;
  assign n9680 = ~n9677 & n9679;
  assign n9681 = ~n9675 & n9680;
  assign n9682 = n9674 ^ x114;
  assign n9683 = n9681 & n9682;
  assign n9684 = n9683 ^ n9330;
  assign n9685 = x115 & ~n9684;
  assign n9686 = n9585 & n9681;
  assign n9687 = n9686 ^ n9587;
  assign n9688 = ~x100 & ~n9687;
  assign n9689 = n9590 ^ x100;
  assign n9690 = n9681 & n9689;
  assign n9691 = n9690 ^ n9335;
  assign n9692 = ~x101 & ~n9691;
  assign n9693 = ~n9688 & ~n9692;
  assign n9694 = n9437 ^ x75;
  assign n9695 = n9681 & n9694;
  assign n9696 = n9695 ^ n9342;
  assign n9697 = n9414 & n9681;
  assign n9698 = n9697 ^ n9416;
  assign n9699 = ~x72 & ~n9698;
  assign n9700 = n293 & ~n9328;
  assign n9701 = n9700 ^ x65;
  assign n9702 = ~x12 & n9701;
  assign n9703 = ~x65 & ~n9702;
  assign n9704 = n9681 & ~n9703;
  assign n9705 = ~n9364 & ~n9704;
  assign n9706 = x65 & n9328;
  assign n9707 = x12 & ~n9706;
  assign n9708 = ~n202 & ~n9707;
  assign n9709 = ~n9702 & n9708;
  assign n9710 = n9681 & n9709;
  assign n9711 = ~n9705 & ~n9710;
  assign n9712 = n9711 ^ x13;
  assign n9713 = n9712 ^ x66;
  assign n9714 = ~x11 & x64;
  assign n9715 = ~x65 & ~n9714;
  assign n9716 = ~x12 & ~n9715;
  assign n9717 = ~n9681 & n9716;
  assign n9718 = x12 ^ x11;
  assign n9719 = ~x64 & n9718;
  assign n9720 = n9719 ^ x11;
  assign n9721 = x65 & ~n9720;
  assign n9722 = ~n9717 & ~n9721;
  assign n9723 = x11 & ~x65;
  assign n9724 = n9372 & ~n9723;
  assign n9725 = n9681 & n9724;
  assign n9726 = n9722 & ~n9725;
  assign n9727 = n9726 ^ n9712;
  assign n9728 = ~n9713 & ~n9727;
  assign n9729 = n9728 ^ x66;
  assign n9730 = n9729 ^ x67;
  assign n9731 = n9377 ^ x66;
  assign n9732 = n9681 & ~n9731;
  assign n9733 = n9732 ^ n9362;
  assign n9734 = n9733 ^ n9729;
  assign n9735 = n9730 & ~n9734;
  assign n9736 = n9735 ^ x67;
  assign n9737 = n9736 ^ x68;
  assign n9738 = n9381 & n9681;
  assign n9739 = n9738 ^ n9392;
  assign n9740 = n9739 ^ n9736;
  assign n9741 = n9737 & n9740;
  assign n9742 = n9741 ^ x68;
  assign n9743 = n9742 ^ x69;
  assign n9744 = n9396 & n9681;
  assign n9745 = n9744 ^ n9398;
  assign n9746 = n9745 ^ n9742;
  assign n9747 = n9743 & n9746;
  assign n9748 = n9747 ^ x69;
  assign n9749 = n9748 ^ x70;
  assign n9750 = n9402 & n9681;
  assign n9751 = n9750 ^ n9404;
  assign n9752 = n9751 ^ n9748;
  assign n9753 = n9749 & ~n9752;
  assign n9754 = n9753 ^ x70;
  assign n9755 = n9754 ^ x71;
  assign n9756 = n9408 & n9681;
  assign n9757 = n9756 ^ n9410;
  assign n9758 = n9757 ^ n9754;
  assign n9759 = n9755 & n9758;
  assign n9760 = n9759 ^ x71;
  assign n9761 = ~n9699 & n9760;
  assign n9762 = n9420 & n9681;
  assign n9763 = n9762 ^ n9422;
  assign n9764 = x73 & n9763;
  assign n9765 = x72 & n9698;
  assign n9766 = ~n9764 & ~n9765;
  assign n9767 = ~n9761 & n9766;
  assign n9768 = ~x73 & ~n9763;
  assign n9769 = ~n9767 & ~n9768;
  assign n9770 = n9769 ^ x74;
  assign n9771 = n9426 & n9681;
  assign n9772 = n9771 ^ n9428;
  assign n9773 = n9772 ^ n9769;
  assign n9774 = n9770 & n9773;
  assign n9775 = n9774 ^ x74;
  assign n9776 = n9775 ^ x75;
  assign n9777 = n9432 & n9681;
  assign n9778 = n9777 ^ n9434;
  assign n9779 = n9778 ^ n9775;
  assign n9780 = n9776 & ~n9779;
  assign n9781 = n9780 ^ x75;
  assign n9782 = ~n9696 & n9781;
  assign n9783 = x76 & n9781;
  assign n9784 = ~n9782 & ~n9783;
  assign n9785 = n9437 ^ n9342;
  assign n9786 = n9694 & n9785;
  assign n9787 = n9786 ^ x75;
  assign n9788 = n9787 ^ x76;
  assign n9789 = n9681 & n9788;
  assign n9790 = n9789 ^ n9345;
  assign n9791 = x76 & x77;
  assign n9792 = ~n9790 & ~n9791;
  assign n9793 = ~n9784 & ~n9792;
  assign n9794 = x77 & n9782;
  assign n9795 = ~n9696 & n9791;
  assign n9796 = ~n9790 & ~n9795;
  assign n9797 = x76 & ~n9696;
  assign n9798 = ~x77 & ~n9797;
  assign n9799 = ~n9796 & ~n9798;
  assign n9800 = ~n9794 & ~n9799;
  assign n9801 = ~n9793 & n9800;
  assign n9802 = ~n9445 & n9681;
  assign n9803 = n9802 ^ n9447;
  assign n9804 = ~x78 & n9803;
  assign n9805 = n9451 & n9681;
  assign n9806 = n9805 ^ n9453;
  assign n9807 = ~x79 & ~n9806;
  assign n9808 = ~n9804 & ~n9807;
  assign n9809 = ~n9801 & n9808;
  assign n9810 = n9806 ^ x79;
  assign n9811 = x78 & ~n9803;
  assign n9812 = n9811 ^ n9806;
  assign n9813 = n9810 & ~n9812;
  assign n9814 = n9813 ^ x79;
  assign n9815 = ~n9809 & ~n9814;
  assign n9816 = n9815 ^ x80;
  assign n9817 = n9457 & n9681;
  assign n9818 = n9817 ^ n9459;
  assign n9819 = n9818 ^ n9815;
  assign n9820 = ~n9816 & n9819;
  assign n9821 = n9820 ^ x80;
  assign n9822 = n9821 ^ x81;
  assign n9823 = n9463 & n9681;
  assign n9824 = n9823 ^ n9465;
  assign n9825 = n9824 ^ n9821;
  assign n9826 = n9822 & ~n9825;
  assign n9827 = n9826 ^ x81;
  assign n9828 = n9827 ^ x82;
  assign n9829 = n9469 & n9681;
  assign n9830 = n9829 ^ n9471;
  assign n9831 = n9830 ^ n9827;
  assign n9832 = n9828 & ~n9831;
  assign n9833 = n9832 ^ x82;
  assign n9834 = n9833 ^ x83;
  assign n9835 = n9475 & n9681;
  assign n9836 = n9835 ^ n9477;
  assign n9837 = n9836 ^ n9833;
  assign n9838 = n9834 & ~n9837;
  assign n9839 = n9838 ^ x83;
  assign n9840 = n9839 ^ x84;
  assign n9841 = n9481 & n9681;
  assign n9842 = n9841 ^ n9483;
  assign n9843 = n9842 ^ n9839;
  assign n9844 = n9840 & ~n9843;
  assign n9845 = n9844 ^ x84;
  assign n9846 = n9845 ^ x85;
  assign n9847 = n9487 & n9681;
  assign n9848 = n9847 ^ n9489;
  assign n9849 = n9848 ^ n9845;
  assign n9850 = n9846 & ~n9849;
  assign n9851 = n9850 ^ x85;
  assign n9852 = n9851 ^ x86;
  assign n9853 = n9493 & n9681;
  assign n9854 = n9853 ^ n9496;
  assign n9855 = n9854 ^ n9851;
  assign n9856 = n9852 & ~n9855;
  assign n9857 = n9856 ^ x86;
  assign n9858 = n9857 ^ x87;
  assign n9859 = n9500 & n9681;
  assign n9860 = n9859 ^ n9506;
  assign n9861 = n9860 ^ n9857;
  assign n9862 = n9858 & ~n9861;
  assign n9863 = n9862 ^ x87;
  assign n9864 = n9863 ^ x88;
  assign n9865 = n9510 & n9681;
  assign n9866 = n9865 ^ n9512;
  assign n9867 = n9866 ^ n9863;
  assign n9868 = n9864 & ~n9867;
  assign n9869 = n9868 ^ x88;
  assign n9870 = n9869 ^ x89;
  assign n9871 = n9516 & n9681;
  assign n9872 = n9871 ^ n9518;
  assign n9873 = n9872 ^ n9869;
  assign n9874 = n9870 & ~n9873;
  assign n9875 = n9874 ^ x89;
  assign n9876 = n9875 ^ x90;
  assign n9877 = n9522 & n9681;
  assign n9878 = n9877 ^ n9524;
  assign n9879 = n9878 ^ n9875;
  assign n9880 = n9876 & ~n9879;
  assign n9881 = n9880 ^ x90;
  assign n9882 = n9881 ^ x91;
  assign n9883 = n9528 & n9681;
  assign n9884 = n9883 ^ n9530;
  assign n9885 = n9884 ^ n9881;
  assign n9886 = n9882 & ~n9885;
  assign n9887 = n9886 ^ x91;
  assign n9888 = n9887 ^ x92;
  assign n9889 = n9534 & n9681;
  assign n9890 = n9889 ^ n9536;
  assign n9891 = n9890 ^ n9887;
  assign n9892 = n9888 & ~n9891;
  assign n9893 = n9892 ^ x92;
  assign n9894 = n9893 ^ x93;
  assign n9895 = n9540 & n9681;
  assign n9896 = n9895 ^ n9542;
  assign n9897 = n9896 ^ n9893;
  assign n9898 = n9894 & ~n9897;
  assign n9899 = n9898 ^ x93;
  assign n9900 = n9899 ^ x94;
  assign n9901 = n9546 & n9681;
  assign n9902 = n9901 ^ n9548;
  assign n9903 = n9902 ^ n9899;
  assign n9904 = n9900 & ~n9903;
  assign n9905 = n9904 ^ x94;
  assign n9906 = n9905 ^ x95;
  assign n9907 = n9552 & n9681;
  assign n9908 = n9907 ^ n9554;
  assign n9909 = n9908 ^ n9905;
  assign n9910 = n9906 & ~n9909;
  assign n9911 = n9910 ^ x95;
  assign n9912 = n9911 ^ x96;
  assign n9913 = n9558 & n9681;
  assign n9914 = n9913 ^ n9560;
  assign n9915 = n9914 ^ n9911;
  assign n9916 = n9912 & ~n9915;
  assign n9917 = n9916 ^ x96;
  assign n9918 = n9917 ^ x97;
  assign n9919 = n9564 & n9681;
  assign n9920 = n9919 ^ n9566;
  assign n9921 = n9920 ^ n9917;
  assign n9922 = n9918 & ~n9921;
  assign n9923 = n9922 ^ x97;
  assign n9924 = n9923 ^ x98;
  assign n9925 = n9570 & n9681;
  assign n9926 = n9925 ^ n9573;
  assign n9927 = n9926 ^ n9923;
  assign n9928 = n9924 & ~n9927;
  assign n9929 = n9928 ^ x98;
  assign n9930 = n9929 ^ x99;
  assign n9931 = n9577 & n9681;
  assign n9932 = n9931 ^ n9581;
  assign n9933 = n9932 ^ n9929;
  assign n9934 = n9930 & ~n9933;
  assign n9935 = n9934 ^ x99;
  assign n9936 = n9693 & n9935;
  assign n9937 = n9691 ^ x101;
  assign n9938 = x100 & n9687;
  assign n9939 = n9938 ^ n9691;
  assign n9940 = n9937 & ~n9939;
  assign n9941 = n9940 ^ x101;
  assign n9942 = ~n9936 & ~n9941;
  assign n9943 = n9942 ^ x102;
  assign n9944 = n9590 ^ n9335;
  assign n9945 = n9689 & ~n9944;
  assign n9946 = n9945 ^ x100;
  assign n9947 = n9946 ^ x101;
  assign n9948 = n9681 & n9947;
  assign n9949 = n9948 ^ n9338;
  assign n9950 = n9949 ^ n9942;
  assign n9951 = ~n9943 & n9950;
  assign n9952 = n9951 ^ x102;
  assign n9953 = n9952 ^ x103;
  assign n9954 = ~n9598 & n9681;
  assign n9955 = n9954 ^ n9600;
  assign n9956 = n9955 ^ n9952;
  assign n9957 = n9953 & ~n9956;
  assign n9958 = n9957 ^ x103;
  assign n9959 = n9958 ^ x104;
  assign n9960 = n9604 & n9681;
  assign n9961 = n9960 ^ n9606;
  assign n9962 = n9961 ^ n9958;
  assign n9963 = n9959 & ~n9962;
  assign n9964 = n9963 ^ x104;
  assign n9965 = n9964 ^ x105;
  assign n9966 = n9610 & n9681;
  assign n9967 = n9966 ^ n9612;
  assign n9968 = n9967 ^ n9964;
  assign n9969 = n9965 & ~n9968;
  assign n9970 = n9969 ^ x105;
  assign n9971 = n9970 ^ x106;
  assign n9972 = n9616 & n9681;
  assign n9973 = n9972 ^ n9618;
  assign n9974 = n9973 ^ n9970;
  assign n9975 = n9971 & ~n9974;
  assign n9976 = n9975 ^ x106;
  assign n9977 = n9976 ^ x107;
  assign n9978 = n9622 & n9681;
  assign n9979 = n9978 ^ n9624;
  assign n9980 = n9979 ^ n9976;
  assign n9981 = n9977 & ~n9980;
  assign n9982 = n9981 ^ x107;
  assign n9983 = n9982 ^ x108;
  assign n9984 = n9628 & n9681;
  assign n9985 = n9984 ^ n9631;
  assign n9986 = n9985 ^ n9982;
  assign n9987 = n9983 & ~n9986;
  assign n9988 = n9987 ^ x108;
  assign n9989 = n9988 ^ x109;
  assign n9990 = n9635 & n9681;
  assign n9991 = n9990 ^ n9641;
  assign n9992 = n9991 ^ n9988;
  assign n9993 = n9989 & ~n9992;
  assign n9994 = n9993 ^ x109;
  assign n9995 = n9994 ^ x110;
  assign n9996 = n9645 & n9681;
  assign n9997 = n9996 ^ n9647;
  assign n9998 = n9997 ^ n9994;
  assign n9999 = n9995 & ~n9998;
  assign n10000 = n9999 ^ x110;
  assign n10001 = n10000 ^ x111;
  assign n10002 = n9651 & n9681;
  assign n10003 = n10002 ^ n9653;
  assign n10004 = n10003 ^ n10000;
  assign n10005 = n10001 & ~n10004;
  assign n10006 = n10005 ^ x111;
  assign n10007 = n10006 ^ x112;
  assign n10008 = n9657 & n9681;
  assign n10009 = n10008 ^ n9659;
  assign n10010 = n10009 ^ n10006;
  assign n10011 = n10007 & ~n10010;
  assign n10012 = n10011 ^ x112;
  assign n10013 = n10012 ^ x113;
  assign n10014 = n9663 & n9681;
  assign n10015 = n10014 ^ n9665;
  assign n10016 = n10015 ^ n10012;
  assign n10017 = n10013 & ~n10016;
  assign n10018 = n10017 ^ x113;
  assign n10019 = n10018 ^ x114;
  assign n10020 = n9669 & n9681;
  assign n10021 = n10020 ^ n9671;
  assign n10022 = n10021 ^ n10018;
  assign n10023 = n10019 & ~n10022;
  assign n10024 = n10023 ^ x114;
  assign n10025 = ~n9685 & ~n10024;
  assign n10026 = ~x115 & n9684;
  assign n10027 = ~n10025 & ~n10026;
  assign n10028 = n10027 ^ x116;
  assign n10029 = n9674 ^ n9330;
  assign n10030 = n9682 & n10029;
  assign n10031 = n10030 ^ x114;
  assign n10032 = n10031 ^ x115;
  assign n10033 = ~n10027 & n10032;
  assign n10034 = ~n10028 & n10033;
  assign n10035 = n10034 ^ n10028;
  assign n10036 = n9324 & n10035;
  assign n10037 = n9320 & ~n10036;
  assign n10038 = ~x117 & n10037;
  assign n10039 = n9320 & ~n10032;
  assign n10040 = ~n10026 & ~n10039;
  assign n10041 = ~n10025 & n10040;
  assign n10042 = ~x116 & ~n10041;
  assign n10043 = n9320 & ~n10027;
  assign n10044 = ~n10042 & ~n10043;
  assign n10045 = n9324 & ~n10044;
  assign n10046 = n10001 & n10045;
  assign n10047 = n10046 ^ n10003;
  assign n10048 = ~x112 & ~n10047;
  assign n10049 = n10007 & n10045;
  assign n10050 = n10049 ^ n10009;
  assign n10051 = ~x113 & ~n10050;
  assign n10052 = ~n10048 & ~n10051;
  assign n10053 = n9776 & n10045;
  assign n10054 = n10053 ^ n9778;
  assign n10055 = ~x76 & ~n10054;
  assign n10056 = n9781 ^ x76;
  assign n10057 = n10045 & n10056;
  assign n10058 = n10057 ^ n9696;
  assign n10059 = ~x77 & n10058;
  assign n10060 = ~n10055 & ~n10059;
  assign n10061 = n9737 & n10045;
  assign n10062 = n10061 ^ n9739;
  assign n10063 = ~x69 & n10062;
  assign n10064 = x65 & ~n9681;
  assign n10065 = n10045 & n10064;
  assign n10066 = ~x65 & n9681;
  assign n10067 = x64 & n10066;
  assign n10068 = ~n10065 & ~n10067;
  assign n10069 = x11 & ~n10068;
  assign n10071 = n9714 & ~n10064;
  assign n10072 = ~n202 & ~n10071;
  assign n10073 = ~n10066 & ~n10072;
  assign n10070 = x64 & n9681;
  assign n10074 = n10073 ^ n10070;
  assign n10075 = ~n10045 & n10074;
  assign n10076 = n10075 ^ n10073;
  assign n10077 = ~n10069 & ~n10076;
  assign n10078 = n10077 ^ x12;
  assign n10079 = n10078 ^ x66;
  assign n10080 = x64 & n10045;
  assign n10081 = x11 & n10080;
  assign n10082 = x10 & ~x65;
  assign n10083 = n10081 & ~n10082;
  assign n10084 = ~x10 & x64;
  assign n10085 = ~x65 & ~n10084;
  assign n10086 = ~x11 & ~n10085;
  assign n10087 = ~n10045 & n10086;
  assign n10088 = ~x11 & n202;
  assign n10089 = ~x10 & x65;
  assign n10090 = x64 & n10089;
  assign n10091 = ~n10088 & ~n10090;
  assign n10092 = ~n10087 & n10091;
  assign n10093 = ~n10083 & n10092;
  assign n10094 = n10093 ^ n10078;
  assign n10095 = n10079 & n10094;
  assign n10096 = n10095 ^ x66;
  assign n10097 = n10096 ^ x67;
  assign n10098 = n9726 ^ x66;
  assign n10099 = n10045 & ~n10098;
  assign n10100 = n10099 ^ n9712;
  assign n10101 = n10100 ^ n10096;
  assign n10102 = n10097 & n10101;
  assign n10103 = n10102 ^ x67;
  assign n10104 = n10103 ^ x68;
  assign n10105 = n9730 & n10045;
  assign n10106 = n10105 ^ n9733;
  assign n10107 = n10106 ^ n10103;
  assign n10108 = n10104 & ~n10107;
  assign n10109 = n10108 ^ x68;
  assign n10110 = ~n10063 & n10109;
  assign n10111 = n9743 & n10045;
  assign n10112 = n10111 ^ n9745;
  assign n10113 = x70 & ~n10112;
  assign n10114 = x69 & ~n10062;
  assign n10115 = ~n10113 & ~n10114;
  assign n10116 = ~n10110 & n10115;
  assign n10117 = ~x70 & n10112;
  assign n10118 = ~n10116 & ~n10117;
  assign n10119 = n10118 ^ x71;
  assign n10120 = n9749 & n10045;
  assign n10121 = n10120 ^ n9751;
  assign n10122 = n10121 ^ n10118;
  assign n10123 = n10119 & ~n10122;
  assign n10124 = n10123 ^ x71;
  assign n10125 = n10124 ^ x72;
  assign n10126 = n9755 & n10045;
  assign n10127 = n10126 ^ n9757;
  assign n10128 = n10127 ^ n10124;
  assign n10129 = n10125 & n10128;
  assign n10130 = n10129 ^ x72;
  assign n10131 = n10130 ^ x73;
  assign n10132 = n9760 ^ x72;
  assign n10133 = n10045 & n10132;
  assign n10134 = n10133 ^ n9698;
  assign n10135 = n10134 ^ n10130;
  assign n10136 = n10131 & ~n10135;
  assign n10137 = n10136 ^ x73;
  assign n10138 = n10137 ^ x74;
  assign n10139 = ~n9761 & ~n9765;
  assign n10140 = n10139 ^ x73;
  assign n10141 = n10045 & ~n10140;
  assign n10142 = n10141 ^ n9763;
  assign n10143 = n10142 ^ n10137;
  assign n10144 = n10138 & ~n10143;
  assign n10145 = n10144 ^ x74;
  assign n10146 = n10145 ^ x75;
  assign n10147 = n9770 & n10045;
  assign n10148 = n10147 ^ n9772;
  assign n10149 = n10148 ^ n10145;
  assign n10150 = n10146 & n10149;
  assign n10151 = n10150 ^ x75;
  assign n10152 = n10060 & n10151;
  assign n10153 = n10058 ^ x77;
  assign n10154 = x76 & n10054;
  assign n10155 = n10154 ^ n10058;
  assign n10156 = ~n10153 & n10155;
  assign n10157 = n10156 ^ x77;
  assign n10158 = ~n10152 & ~n10157;
  assign n10159 = n10158 ^ x78;
  assign n10160 = n9781 ^ n9696;
  assign n10161 = n10056 & n10160;
  assign n10162 = n10161 ^ x76;
  assign n10163 = n10162 ^ x77;
  assign n10164 = n10045 & n10163;
  assign n10165 = n10164 ^ n9790;
  assign n10166 = n10165 ^ n10158;
  assign n10167 = ~n10159 & n10166;
  assign n10168 = n10167 ^ x78;
  assign n10169 = n10168 ^ x79;
  assign n10170 = n9801 ^ x78;
  assign n10171 = n10045 & ~n10170;
  assign n10172 = n10171 ^ n9803;
  assign n10173 = n10172 ^ n10168;
  assign n10174 = n10169 & n10173;
  assign n10175 = n10174 ^ x79;
  assign n10176 = n10175 ^ x80;
  assign n10177 = n9803 ^ n9801;
  assign n10178 = ~n10170 & ~n10177;
  assign n10179 = n10178 ^ x78;
  assign n10180 = n10179 ^ x79;
  assign n10181 = n10045 & n10180;
  assign n10182 = n10181 ^ n9806;
  assign n10183 = n10182 ^ n10175;
  assign n10184 = n10176 & ~n10183;
  assign n10185 = n10184 ^ x80;
  assign n10186 = n10185 ^ x81;
  assign n10187 = ~n9816 & n10045;
  assign n10188 = n10187 ^ n9818;
  assign n10189 = n10188 ^ n10185;
  assign n10190 = n10186 & ~n10189;
  assign n10191 = n10190 ^ x81;
  assign n10192 = n10191 ^ x82;
  assign n10193 = n9822 & n10045;
  assign n10194 = n10193 ^ n9824;
  assign n10195 = n10194 ^ n10191;
  assign n10196 = n10192 & ~n10195;
  assign n10197 = n10196 ^ x82;
  assign n10198 = n10197 ^ x83;
  assign n10199 = n9828 & n10045;
  assign n10200 = n10199 ^ n9830;
  assign n10201 = n10200 ^ n10197;
  assign n10202 = n10198 & ~n10201;
  assign n10203 = n10202 ^ x83;
  assign n10204 = n10203 ^ x84;
  assign n10205 = n9834 & n10045;
  assign n10206 = n10205 ^ n9836;
  assign n10207 = n10206 ^ n10203;
  assign n10208 = n10204 & ~n10207;
  assign n10209 = n10208 ^ x84;
  assign n10210 = n10209 ^ x85;
  assign n10211 = n9840 & n10045;
  assign n10212 = n10211 ^ n9842;
  assign n10213 = n10212 ^ n10209;
  assign n10214 = n10210 & ~n10213;
  assign n10215 = n10214 ^ x85;
  assign n10216 = n10215 ^ x86;
  assign n10217 = n9846 & n10045;
  assign n10218 = n10217 ^ n9848;
  assign n10219 = n10218 ^ n10215;
  assign n10220 = n10216 & ~n10219;
  assign n10221 = n10220 ^ x86;
  assign n10222 = n10221 ^ x87;
  assign n10223 = n9852 & n10045;
  assign n10224 = n10223 ^ n9854;
  assign n10225 = n10224 ^ n10221;
  assign n10226 = n10222 & ~n10225;
  assign n10227 = n10226 ^ x87;
  assign n10228 = n10227 ^ x88;
  assign n10229 = n9858 & n10045;
  assign n10230 = n10229 ^ n9860;
  assign n10231 = n10230 ^ n10227;
  assign n10232 = n10228 & ~n10231;
  assign n10233 = n10232 ^ x88;
  assign n10234 = n10233 ^ x89;
  assign n10235 = n9864 & n10045;
  assign n10236 = n10235 ^ n9866;
  assign n10237 = n10236 ^ n10233;
  assign n10238 = n10234 & ~n10237;
  assign n10239 = n10238 ^ x89;
  assign n10240 = n10239 ^ x90;
  assign n10241 = n9870 & n10045;
  assign n10242 = n10241 ^ n9872;
  assign n10243 = n10242 ^ n10239;
  assign n10244 = n10240 & ~n10243;
  assign n10245 = n10244 ^ x90;
  assign n10246 = n10245 ^ x91;
  assign n10247 = n9876 & n10045;
  assign n10248 = n10247 ^ n9878;
  assign n10249 = n10248 ^ n10245;
  assign n10250 = n10246 & ~n10249;
  assign n10251 = n10250 ^ x91;
  assign n10252 = n10251 ^ x92;
  assign n10253 = n9882 & n10045;
  assign n10254 = n10253 ^ n9884;
  assign n10255 = n10254 ^ n10251;
  assign n10256 = n10252 & ~n10255;
  assign n10257 = n10256 ^ x92;
  assign n10258 = n10257 ^ x93;
  assign n10259 = n9888 & n10045;
  assign n10260 = n10259 ^ n9890;
  assign n10261 = n10260 ^ n10257;
  assign n10262 = n10258 & ~n10261;
  assign n10263 = n10262 ^ x93;
  assign n10264 = n10263 ^ x94;
  assign n10265 = n9894 & n10045;
  assign n10266 = n10265 ^ n9896;
  assign n10267 = n10266 ^ n10263;
  assign n10268 = n10264 & ~n10267;
  assign n10269 = n10268 ^ x94;
  assign n10270 = n10269 ^ x95;
  assign n10271 = n9900 & n10045;
  assign n10272 = n10271 ^ n9902;
  assign n10273 = n10272 ^ n10269;
  assign n10274 = n10270 & ~n10273;
  assign n10275 = n10274 ^ x95;
  assign n10276 = n10275 ^ x96;
  assign n10277 = n9906 & n10045;
  assign n10278 = n10277 ^ n9908;
  assign n10279 = n10278 ^ n10275;
  assign n10280 = n10276 & ~n10279;
  assign n10281 = n10280 ^ x96;
  assign n10282 = n10281 ^ x97;
  assign n10283 = n9912 & n10045;
  assign n10284 = n10283 ^ n9914;
  assign n10285 = n10284 ^ n10281;
  assign n10286 = n10282 & ~n10285;
  assign n10287 = n10286 ^ x97;
  assign n10288 = n10287 ^ x98;
  assign n10289 = n9918 & n10045;
  assign n10290 = n10289 ^ n9920;
  assign n10291 = n10290 ^ n10287;
  assign n10292 = n10288 & ~n10291;
  assign n10293 = n10292 ^ x98;
  assign n10294 = n10293 ^ x99;
  assign n10295 = n9924 & n10045;
  assign n10296 = n10295 ^ n9926;
  assign n10297 = n10296 ^ n10293;
  assign n10298 = n10294 & ~n10297;
  assign n10299 = n10298 ^ x99;
  assign n10300 = n10299 ^ x100;
  assign n10301 = n9930 & n10045;
  assign n10302 = n10301 ^ n9932;
  assign n10303 = n10302 ^ n10299;
  assign n10304 = n10300 & ~n10303;
  assign n10305 = n10304 ^ x100;
  assign n10306 = n10305 ^ x101;
  assign n10307 = n9935 ^ x100;
  assign n10308 = n10045 & n10307;
  assign n10309 = n10308 ^ n9687;
  assign n10310 = n10309 ^ n10305;
  assign n10311 = n10306 & ~n10310;
  assign n10312 = n10311 ^ x101;
  assign n10313 = n10312 ^ x102;
  assign n10314 = n9935 ^ n9687;
  assign n10315 = n10307 & ~n10314;
  assign n10316 = n10315 ^ x100;
  assign n10317 = n10316 ^ x101;
  assign n10318 = n10045 & n10317;
  assign n10319 = n10318 ^ n9691;
  assign n10320 = n10319 ^ n10312;
  assign n10321 = n10313 & ~n10320;
  assign n10322 = n10321 ^ x102;
  assign n10323 = n10322 ^ x103;
  assign n10324 = ~n9943 & n10045;
  assign n10325 = n10324 ^ n9949;
  assign n10326 = n10325 ^ n10322;
  assign n10327 = n10323 & ~n10326;
  assign n10328 = n10327 ^ x103;
  assign n10329 = n10328 ^ x104;
  assign n10330 = n9953 & n10045;
  assign n10331 = n10330 ^ n9955;
  assign n10332 = n10331 ^ n10328;
  assign n10333 = n10329 & ~n10332;
  assign n10334 = n10333 ^ x104;
  assign n10335 = n10334 ^ x105;
  assign n10336 = n9959 & n10045;
  assign n10337 = n10336 ^ n9961;
  assign n10338 = n10337 ^ n10334;
  assign n10339 = n10335 & ~n10338;
  assign n10340 = n10339 ^ x105;
  assign n10341 = n10340 ^ x106;
  assign n10342 = n9965 & n10045;
  assign n10343 = n10342 ^ n9967;
  assign n10344 = n10343 ^ n10340;
  assign n10345 = n10341 & ~n10344;
  assign n10346 = n10345 ^ x106;
  assign n10347 = n10346 ^ x107;
  assign n10348 = n9971 & n10045;
  assign n10349 = n10348 ^ n9973;
  assign n10350 = n10349 ^ n10346;
  assign n10351 = n10347 & ~n10350;
  assign n10352 = n10351 ^ x107;
  assign n10353 = n10352 ^ x108;
  assign n10354 = n9977 & n10045;
  assign n10355 = n10354 ^ n9979;
  assign n10356 = n10355 ^ n10352;
  assign n10357 = n10353 & ~n10356;
  assign n10358 = n10357 ^ x108;
  assign n10359 = n10358 ^ x109;
  assign n10360 = n9983 & n10045;
  assign n10361 = n10360 ^ n9985;
  assign n10362 = n10361 ^ n10358;
  assign n10363 = n10359 & ~n10362;
  assign n10364 = n10363 ^ x109;
  assign n10365 = n10364 ^ x110;
  assign n10366 = n9989 & n10045;
  assign n10367 = n10366 ^ n9991;
  assign n10368 = n10367 ^ n10364;
  assign n10369 = n10365 & ~n10368;
  assign n10370 = n10369 ^ x110;
  assign n10371 = n10370 ^ x111;
  assign n10372 = n9995 & n10045;
  assign n10373 = n10372 ^ n9997;
  assign n10374 = n10373 ^ n10370;
  assign n10375 = n10371 & ~n10374;
  assign n10376 = n10375 ^ x111;
  assign n10377 = n10052 & n10376;
  assign n10378 = n10050 ^ x113;
  assign n10379 = x112 & n10047;
  assign n10380 = n10379 ^ n10050;
  assign n10381 = n10378 & ~n10380;
  assign n10382 = n10381 ^ x113;
  assign n10383 = ~n10377 & ~n10382;
  assign n10384 = n10383 ^ x114;
  assign n10385 = n10013 & n10045;
  assign n10386 = n10385 ^ n10015;
  assign n10387 = n10386 ^ n10383;
  assign n10388 = ~n10384 & n10387;
  assign n10389 = n10388 ^ x114;
  assign n10390 = n10389 ^ x115;
  assign n10391 = n10019 & n10045;
  assign n10392 = n10391 ^ n10021;
  assign n10393 = n10392 ^ n10389;
  assign n10394 = n10390 & ~n10393;
  assign n10395 = n10394 ^ x115;
  assign n10396 = n10395 ^ x116;
  assign n10397 = n10024 ^ x115;
  assign n10398 = n10045 & n10397;
  assign n10399 = n10398 ^ n9684;
  assign n10400 = n10399 ^ n10395;
  assign n10401 = n10396 & n10400;
  assign n10402 = n10401 ^ x116;
  assign n10403 = ~n10038 & n10402;
  assign n10404 = x117 & ~n10037;
  assign n10405 = n9323 & ~n10404;
  assign n10406 = ~n10403 & n10405;
  assign n10407 = n10080 ^ x11;
  assign n10408 = ~n10406 & ~n10407;
  assign n10409 = ~x9 & ~n10082;
  assign n10410 = n10408 & n10409;
  assign n10411 = n10407 ^ x65;
  assign n10412 = x9 & n10082;
  assign n10413 = n10412 ^ x10;
  assign n10414 = ~n10411 & n10413;
  assign n10415 = n10406 & n10414;
  assign n10416 = ~x9 & n10089;
  assign n10417 = ~n10407 & n10416;
  assign n10418 = ~n10415 & ~n10417;
  assign n10419 = ~n10410 & n10418;
  assign n10420 = x64 & ~n10419;
  assign n10421 = x64 & n10406;
  assign n10422 = n10089 & ~n10421;
  assign n10423 = n10407 ^ n10406;
  assign n10424 = n10422 & ~n10423;
  assign n10425 = ~x66 & ~n10424;
  assign n10426 = ~n10420 & n10425;
  assign n10427 = ~x9 & x64;
  assign n10428 = n10085 & ~n10427;
  assign n10429 = n10406 & ~n10428;
  assign n10430 = ~n10082 & n10427;
  assign n10431 = ~n10089 & ~n10430;
  assign n10432 = n10407 & n10431;
  assign n10433 = ~n10429 & n10432;
  assign n10434 = ~x9 & x65;
  assign n10435 = n10084 & ~n10434;
  assign n10436 = ~n10411 & n10435;
  assign n10437 = x10 & n10088;
  assign n10438 = ~n10436 & ~n10437;
  assign n10439 = n10406 & ~n10438;
  assign n10440 = ~n10433 & ~n10439;
  assign n10441 = ~n10426 & n10440;
  assign n10442 = n10441 ^ x67;
  assign n10443 = n10093 ^ x66;
  assign n10444 = n10406 & ~n10443;
  assign n10445 = n10444 ^ n10078;
  assign n10446 = n10445 ^ n10441;
  assign n10447 = n10442 & ~n10446;
  assign n10448 = n10447 ^ x67;
  assign n10449 = n10448 ^ x68;
  assign n10450 = n10097 & n10406;
  assign n10451 = n10450 ^ n10100;
  assign n10452 = n10451 ^ n10448;
  assign n10453 = n10449 & n10452;
  assign n10454 = n10453 ^ x68;
  assign n10455 = n10454 ^ x69;
  assign n10456 = n10104 & n10406;
  assign n10457 = n10456 ^ n10106;
  assign n10458 = n10457 ^ n10454;
  assign n10459 = n10455 & ~n10458;
  assign n10460 = n10459 ^ x69;
  assign n10461 = ~x70 & ~n10460;
  assign n10462 = ~n10110 & ~n10114;
  assign n10463 = n10462 ^ x70;
  assign n10464 = n10406 & ~n10463;
  assign n10465 = n10464 ^ n10112;
  assign n10466 = n10109 ^ x69;
  assign n10467 = n10406 & n10466;
  assign n10468 = n10467 ^ n10062;
  assign n10469 = ~n10465 & ~n10468;
  assign n10470 = ~n10461 & n10469;
  assign n10471 = x70 & ~n10465;
  assign n10472 = ~x71 & ~n10471;
  assign n10473 = ~x70 & n10468;
  assign n10474 = ~n10472 & ~n10473;
  assign n10475 = n10460 & n10474;
  assign n10476 = x70 & ~n10468;
  assign n10477 = n10465 & ~n10476;
  assign n10478 = x71 & ~n10477;
  assign n10479 = ~n10475 & ~n10478;
  assign n10480 = ~n10470 & n10479;
  assign n10481 = n10480 ^ x72;
  assign n10482 = n10119 & n10406;
  assign n10483 = n10482 ^ n10121;
  assign n10484 = n10483 ^ n10480;
  assign n10485 = ~n10481 & n10484;
  assign n10486 = n10485 ^ x72;
  assign n10487 = n10486 ^ x73;
  assign n10488 = n10125 & n10406;
  assign n10489 = n10488 ^ n10127;
  assign n10490 = n10489 ^ n10486;
  assign n10491 = n10487 & n10490;
  assign n10492 = n10491 ^ x73;
  assign n10493 = n10492 ^ x74;
  assign n10494 = n10131 & n10406;
  assign n10495 = n10494 ^ n10134;
  assign n10496 = n10495 ^ n10492;
  assign n10497 = n10493 & ~n10496;
  assign n10498 = n10497 ^ x74;
  assign n10499 = n10498 ^ x75;
  assign n10500 = n10138 & n10406;
  assign n10501 = n10500 ^ n10142;
  assign n10502 = n10501 ^ n10498;
  assign n10503 = n10499 & ~n10502;
  assign n10504 = n10503 ^ x75;
  assign n10505 = n10504 ^ x76;
  assign n10506 = n10146 & n10406;
  assign n10507 = n10506 ^ n10148;
  assign n10508 = n10507 ^ n10504;
  assign n10509 = n10505 & n10508;
  assign n10510 = n10509 ^ x76;
  assign n10511 = n10510 ^ x77;
  assign n10512 = n10151 ^ x76;
  assign n10513 = n10406 & n10512;
  assign n10514 = n10513 ^ n10054;
  assign n10515 = n10514 ^ n10510;
  assign n10516 = n10511 & ~n10515;
  assign n10517 = n10516 ^ x77;
  assign n10518 = n10517 ^ x78;
  assign n10519 = n10151 ^ n10054;
  assign n10520 = n10512 & ~n10519;
  assign n10521 = n10520 ^ x76;
  assign n10522 = n10521 ^ x77;
  assign n10523 = n10406 & n10522;
  assign n10524 = n10523 ^ n10058;
  assign n10525 = n10524 ^ n10517;
  assign n10526 = n10518 & n10525;
  assign n10527 = n10526 ^ x78;
  assign n10528 = n10527 ^ x79;
  assign n10529 = ~n10159 & n10406;
  assign n10530 = n10529 ^ n10165;
  assign n10531 = n10530 ^ n10527;
  assign n10532 = n10528 & ~n10531;
  assign n10533 = n10532 ^ x79;
  assign n10534 = n10533 ^ x80;
  assign n10535 = n10169 & n10406;
  assign n10536 = n10535 ^ n10172;
  assign n10537 = n10536 ^ n10533;
  assign n10538 = n10534 & n10537;
  assign n10539 = n10538 ^ x80;
  assign n10540 = n10539 ^ x81;
  assign n10541 = n10176 & n10406;
  assign n10542 = n10541 ^ n10182;
  assign n10543 = n10542 ^ n10539;
  assign n10544 = n10540 & ~n10543;
  assign n10545 = n10544 ^ x81;
  assign n10546 = n10545 ^ x82;
  assign n10547 = n10186 & n10406;
  assign n10548 = n10547 ^ n10188;
  assign n10549 = n10548 ^ n10545;
  assign n10550 = n10546 & ~n10549;
  assign n10551 = n10550 ^ x82;
  assign n10552 = n10551 ^ x83;
  assign n10553 = n10192 & n10406;
  assign n10554 = n10553 ^ n10194;
  assign n10555 = n10554 ^ n10551;
  assign n10556 = n10552 & ~n10555;
  assign n10557 = n10556 ^ x83;
  assign n10558 = n10557 ^ x84;
  assign n10559 = n10198 & n10406;
  assign n10560 = n10559 ^ n10200;
  assign n10561 = n10560 ^ n10557;
  assign n10562 = n10558 & ~n10561;
  assign n10563 = n10562 ^ x84;
  assign n10564 = n10563 ^ x85;
  assign n10565 = n10204 & n10406;
  assign n10566 = n10565 ^ n10206;
  assign n10567 = n10566 ^ n10563;
  assign n10568 = n10564 & ~n10567;
  assign n10569 = n10568 ^ x85;
  assign n10570 = n10569 ^ x86;
  assign n10571 = n10210 & n10406;
  assign n10572 = n10571 ^ n10212;
  assign n10573 = n10572 ^ n10569;
  assign n10574 = n10570 & ~n10573;
  assign n10575 = n10574 ^ x86;
  assign n10576 = n10575 ^ x87;
  assign n10577 = n10216 & n10406;
  assign n10578 = n10577 ^ n10218;
  assign n10579 = n10578 ^ n10575;
  assign n10580 = n10576 & ~n10579;
  assign n10581 = n10580 ^ x87;
  assign n10582 = n10581 ^ x88;
  assign n10583 = n10222 & n10406;
  assign n10584 = n10583 ^ n10224;
  assign n10585 = n10584 ^ n10581;
  assign n10586 = n10582 & ~n10585;
  assign n10587 = n10586 ^ x88;
  assign n10588 = n10587 ^ x89;
  assign n10589 = n10228 & n10406;
  assign n10590 = n10589 ^ n10230;
  assign n10591 = n10590 ^ n10587;
  assign n10592 = n10588 & ~n10591;
  assign n10593 = n10592 ^ x89;
  assign n10594 = n10593 ^ x90;
  assign n10595 = n10234 & n10406;
  assign n10596 = n10595 ^ n10236;
  assign n10597 = n10596 ^ n10593;
  assign n10598 = n10594 & ~n10597;
  assign n10599 = n10598 ^ x90;
  assign n10600 = n10599 ^ x91;
  assign n10601 = n10240 & n10406;
  assign n10602 = n10601 ^ n10242;
  assign n10603 = n10602 ^ n10599;
  assign n10604 = n10600 & ~n10603;
  assign n10605 = n10604 ^ x91;
  assign n10606 = n10605 ^ x92;
  assign n10607 = n10246 & n10406;
  assign n10608 = n10607 ^ n10248;
  assign n10609 = n10608 ^ n10605;
  assign n10610 = n10606 & ~n10609;
  assign n10611 = n10610 ^ x92;
  assign n10612 = n10611 ^ x93;
  assign n10613 = n10402 ^ x117;
  assign n10614 = n10406 & n10613;
  assign n10615 = n10037 & ~n10614;
  assign n10616 = n10376 ^ x112;
  assign n10617 = n10376 ^ n10047;
  assign n10618 = n10616 & ~n10617;
  assign n10619 = n10618 ^ x112;
  assign n10620 = n10619 ^ x113;
  assign n10621 = n10406 & n10620;
  assign n10622 = n10621 ^ n10050;
  assign n10623 = ~x114 & ~n10622;
  assign n10624 = n10406 & n10616;
  assign n10625 = n10624 ^ n10047;
  assign n10626 = ~x113 & ~n10625;
  assign n10627 = ~n10623 & ~n10626;
  assign n10628 = n10341 & n10406;
  assign n10629 = n10628 ^ n10343;
  assign n10630 = ~x107 & ~n10629;
  assign n10631 = n10347 & n10406;
  assign n10632 = n10631 ^ n10349;
  assign n10633 = ~x108 & ~n10632;
  assign n10634 = ~n10630 & ~n10633;
  assign n10635 = n10252 & n10406;
  assign n10636 = n10635 ^ n10254;
  assign n10637 = n10636 ^ n10611;
  assign n10638 = n10612 & ~n10637;
  assign n10639 = n10638 ^ x93;
  assign n10640 = n10639 ^ x94;
  assign n10641 = n10258 & n10406;
  assign n10642 = n10641 ^ n10260;
  assign n10643 = n10642 ^ n10639;
  assign n10644 = n10640 & ~n10643;
  assign n10645 = n10644 ^ x94;
  assign n10646 = n10645 ^ x95;
  assign n10647 = n10264 & n10406;
  assign n10648 = n10647 ^ n10266;
  assign n10649 = n10648 ^ n10645;
  assign n10650 = n10646 & ~n10649;
  assign n10651 = n10650 ^ x95;
  assign n10652 = n10651 ^ x96;
  assign n10653 = n10270 & n10406;
  assign n10654 = n10653 ^ n10272;
  assign n10655 = n10654 ^ n10651;
  assign n10656 = n10652 & ~n10655;
  assign n10657 = n10656 ^ x96;
  assign n10658 = n10657 ^ x97;
  assign n10659 = n10276 & n10406;
  assign n10660 = n10659 ^ n10278;
  assign n10661 = n10660 ^ n10657;
  assign n10662 = n10658 & ~n10661;
  assign n10663 = n10662 ^ x97;
  assign n10664 = n10663 ^ x98;
  assign n10665 = n10282 & n10406;
  assign n10666 = n10665 ^ n10284;
  assign n10667 = n10666 ^ n10663;
  assign n10668 = n10664 & ~n10667;
  assign n10669 = n10668 ^ x98;
  assign n10670 = n10669 ^ x99;
  assign n10671 = n10288 & n10406;
  assign n10672 = n10671 ^ n10290;
  assign n10673 = n10672 ^ n10669;
  assign n10674 = n10670 & ~n10673;
  assign n10675 = n10674 ^ x99;
  assign n10676 = n10675 ^ x100;
  assign n10677 = n10294 & n10406;
  assign n10678 = n10677 ^ n10296;
  assign n10679 = n10678 ^ n10675;
  assign n10680 = n10676 & ~n10679;
  assign n10681 = n10680 ^ x100;
  assign n10682 = n10681 ^ x101;
  assign n10683 = n10300 & n10406;
  assign n10684 = n10683 ^ n10302;
  assign n10685 = n10684 ^ n10681;
  assign n10686 = n10682 & ~n10685;
  assign n10687 = n10686 ^ x101;
  assign n10688 = n10687 ^ x102;
  assign n10689 = n10306 & n10406;
  assign n10690 = n10689 ^ n10309;
  assign n10691 = n10690 ^ n10687;
  assign n10692 = n10688 & ~n10691;
  assign n10693 = n10692 ^ x102;
  assign n10694 = n10693 ^ x103;
  assign n10695 = n10313 & n10406;
  assign n10696 = n10695 ^ n10319;
  assign n10697 = n10696 ^ n10693;
  assign n10698 = n10694 & ~n10697;
  assign n10699 = n10698 ^ x103;
  assign n10700 = n10699 ^ x104;
  assign n10701 = n10323 & n10406;
  assign n10702 = n10701 ^ n10325;
  assign n10703 = n10702 ^ n10699;
  assign n10704 = n10700 & ~n10703;
  assign n10705 = n10704 ^ x104;
  assign n10706 = n10705 ^ x105;
  assign n10707 = n10329 & n10406;
  assign n10708 = n10707 ^ n10331;
  assign n10709 = n10708 ^ n10705;
  assign n10710 = n10706 & ~n10709;
  assign n10711 = n10710 ^ x105;
  assign n10712 = n10711 ^ x106;
  assign n10713 = n10335 & n10406;
  assign n10714 = n10713 ^ n10337;
  assign n10715 = n10714 ^ n10711;
  assign n10716 = n10712 & ~n10715;
  assign n10717 = n10716 ^ x106;
  assign n10718 = n10634 & n10717;
  assign n10719 = n10632 ^ x108;
  assign n10720 = x107 & n10629;
  assign n10721 = n10720 ^ n10632;
  assign n10722 = n10719 & ~n10721;
  assign n10723 = n10722 ^ x108;
  assign n10724 = ~n10718 & ~n10723;
  assign n10725 = n10724 ^ x109;
  assign n10726 = n10353 & n10406;
  assign n10727 = n10726 ^ n10355;
  assign n10728 = n10727 ^ n10724;
  assign n10729 = ~n10725 & n10728;
  assign n10730 = n10729 ^ x109;
  assign n10731 = n10730 ^ x110;
  assign n10732 = n10359 & n10406;
  assign n10733 = n10732 ^ n10361;
  assign n10734 = n10733 ^ n10730;
  assign n10735 = n10731 & ~n10734;
  assign n10736 = n10735 ^ x110;
  assign n10737 = n10736 ^ x111;
  assign n10738 = n10365 & n10406;
  assign n10739 = n10738 ^ n10367;
  assign n10740 = n10739 ^ n10736;
  assign n10741 = n10737 & ~n10740;
  assign n10742 = n10741 ^ x111;
  assign n10743 = n10742 ^ x112;
  assign n10744 = n10371 & n10406;
  assign n10745 = n10744 ^ n10373;
  assign n10746 = n10745 ^ n10742;
  assign n10747 = n10743 & ~n10746;
  assign n10748 = n10747 ^ x112;
  assign n10749 = n10627 & n10748;
  assign n10750 = n10622 ^ x114;
  assign n10751 = x113 & n10625;
  assign n10752 = n10751 ^ n10622;
  assign n10753 = n10750 & ~n10752;
  assign n10754 = n10753 ^ x114;
  assign n10755 = ~n10749 & ~n10754;
  assign n10756 = ~n10384 & n10406;
  assign n10757 = n10756 ^ n10386;
  assign n10758 = ~x115 & ~n10757;
  assign n10759 = n10390 & n10406;
  assign n10760 = n10759 ^ n10392;
  assign n10761 = ~x116 & ~n10760;
  assign n10762 = ~n10758 & ~n10761;
  assign n10763 = ~n10755 & n10762;
  assign n10764 = n10760 ^ x116;
  assign n10765 = x115 & n10757;
  assign n10766 = n10765 ^ n10760;
  assign n10767 = n10764 & ~n10766;
  assign n10768 = n10767 ^ x116;
  assign n10769 = ~n10763 & ~n10768;
  assign n10770 = x117 & ~n10769;
  assign n10771 = ~n10615 & n10770;
  assign n10772 = n10396 & n10406;
  assign n10773 = n10772 ^ n10399;
  assign n10774 = ~x118 & n10615;
  assign n10775 = ~n10773 & ~n10774;
  assign n10776 = x117 & x118;
  assign n10777 = ~n10775 & ~n10776;
  assign n10778 = ~n10769 & ~n10777;
  assign n10779 = x117 & n10775;
  assign n10780 = x118 & ~n10615;
  assign n10781 = n9322 & ~n10780;
  assign n10782 = ~n10779 & n10781;
  assign n10783 = ~n10778 & n10782;
  assign n10784 = ~n10771 & n10783;
  assign n10785 = n10612 & n10784;
  assign n10786 = n10785 ^ n10636;
  assign n10787 = ~x94 & ~n10786;
  assign n10788 = n10606 & n10784;
  assign n10789 = n10788 ^ n10608;
  assign n10790 = ~x93 & ~n10789;
  assign n10791 = ~n10787 & ~n10790;
  assign n10792 = x65 & n10406;
  assign n10793 = x9 & ~n10792;
  assign n10794 = n10784 & ~n10793;
  assign n10795 = n10421 & ~n10794;
  assign n10796 = n10406 ^ x65;
  assign n10797 = n10427 & ~n10796;
  assign n10798 = ~n202 & ~n10797;
  assign n10799 = x65 & n10793;
  assign n10800 = n10798 & ~n10799;
  assign n10801 = n10784 & ~n10800;
  assign n10802 = ~n10795 & ~n10801;
  assign n10803 = n10802 ^ x10;
  assign n10804 = n10803 ^ x66;
  assign n10805 = x64 & n10784;
  assign n10806 = x9 & ~x65;
  assign n10807 = x8 & n10806;
  assign n10808 = n10807 ^ x9;
  assign n10809 = n10805 & n10808;
  assign n10810 = ~x8 & n10427;
  assign n10811 = ~n10434 & ~n10810;
  assign n10812 = ~n10784 & ~n10811;
  assign n10813 = x8 & x64;
  assign n10814 = x65 & ~n10813;
  assign n10815 = x9 & ~x64;
  assign n10816 = n10814 & ~n10815;
  assign n10817 = ~n10812 & ~n10816;
  assign n10818 = ~n10809 & n10817;
  assign n10819 = n10818 ^ n10803;
  assign n10820 = n10804 & n10819;
  assign n10821 = n10820 ^ x66;
  assign n10822 = n10821 ^ x67;
  assign n10826 = ~x65 & n10406;
  assign n10827 = n10430 & ~n10826;
  assign n10828 = ~n10422 & ~n10827;
  assign n10829 = n10413 & n10421;
  assign n10830 = n10828 & ~n10829;
  assign n10831 = n10830 ^ x66;
  assign n10832 = n10784 & ~n10831;
  assign n10823 = n10084 ^ x65;
  assign n10824 = n10406 & n10823;
  assign n10825 = n10824 ^ n10407;
  assign n10833 = n10832 ^ n10825;
  assign n10834 = n10833 ^ n10821;
  assign n10835 = n10822 & n10834;
  assign n10836 = n10835 ^ x67;
  assign n10837 = n10836 ^ x68;
  assign n10838 = n10442 & n10784;
  assign n10839 = n10838 ^ n10445;
  assign n10840 = n10839 ^ n10836;
  assign n10841 = n10837 & ~n10840;
  assign n10842 = n10841 ^ x68;
  assign n10843 = n10842 ^ x69;
  assign n10844 = n10449 & n10784;
  assign n10845 = n10844 ^ n10451;
  assign n10846 = n10845 ^ n10842;
  assign n10847 = n10843 & n10846;
  assign n10848 = n10847 ^ x69;
  assign n10849 = n10848 ^ x70;
  assign n10850 = n10455 & n10784;
  assign n10851 = n10850 ^ n10457;
  assign n10852 = n10851 ^ n10848;
  assign n10853 = n10849 & ~n10852;
  assign n10854 = n10853 ^ x70;
  assign n10855 = n10854 ^ x71;
  assign n10856 = n10460 ^ x70;
  assign n10857 = n10784 & n10856;
  assign n10858 = n10857 ^ n10468;
  assign n10859 = n10858 ^ n10854;
  assign n10860 = n10855 & n10859;
  assign n10861 = n10860 ^ x71;
  assign n10862 = n10861 ^ x72;
  assign n10863 = n10468 ^ n10460;
  assign n10864 = n10856 & n10863;
  assign n10865 = n10864 ^ x70;
  assign n10866 = n10865 ^ x71;
  assign n10867 = n10784 & n10866;
  assign n10868 = n10867 ^ n10465;
  assign n10869 = n10868 ^ n10861;
  assign n10870 = n10862 & n10869;
  assign n10871 = n10870 ^ x72;
  assign n10872 = n10871 ^ x73;
  assign n10873 = ~n10481 & n10784;
  assign n10874 = n10873 ^ n10483;
  assign n10875 = n10874 ^ n10871;
  assign n10876 = n10872 & ~n10875;
  assign n10877 = n10876 ^ x73;
  assign n10878 = n10877 ^ x74;
  assign n10879 = n10487 & n10784;
  assign n10880 = n10879 ^ n10489;
  assign n10881 = n10880 ^ n10877;
  assign n10882 = n10878 & n10881;
  assign n10883 = n10882 ^ x74;
  assign n10884 = n10883 ^ x75;
  assign n10885 = n10493 & n10784;
  assign n10886 = n10885 ^ n10495;
  assign n10887 = n10886 ^ n10883;
  assign n10888 = n10884 & ~n10887;
  assign n10889 = n10888 ^ x75;
  assign n10890 = n10889 ^ x76;
  assign n10891 = n10499 & n10784;
  assign n10892 = n10891 ^ n10501;
  assign n10893 = n10892 ^ n10889;
  assign n10894 = n10890 & ~n10893;
  assign n10895 = n10894 ^ x76;
  assign n10896 = n10895 ^ x77;
  assign n10897 = n10505 & n10784;
  assign n10898 = n10897 ^ n10507;
  assign n10899 = n10898 ^ n10895;
  assign n10900 = n10896 & n10899;
  assign n10901 = n10900 ^ x77;
  assign n10902 = n10901 ^ x78;
  assign n10903 = n10511 & n10784;
  assign n10904 = n10903 ^ n10514;
  assign n10905 = n10904 ^ n10901;
  assign n10906 = n10902 & ~n10905;
  assign n10907 = n10906 ^ x78;
  assign n10908 = n10907 ^ x79;
  assign n10909 = n10518 & n10784;
  assign n10910 = n10909 ^ n10524;
  assign n10911 = n10910 ^ n10907;
  assign n10912 = n10908 & n10911;
  assign n10913 = n10912 ^ x79;
  assign n10914 = n10913 ^ x80;
  assign n10915 = n10528 & n10784;
  assign n10916 = n10915 ^ n10530;
  assign n10917 = n10916 ^ n10913;
  assign n10918 = n10914 & ~n10917;
  assign n10919 = n10918 ^ x80;
  assign n10920 = n10919 ^ x81;
  assign n10921 = n10534 & n10784;
  assign n10922 = n10921 ^ n10536;
  assign n10923 = n10922 ^ n10919;
  assign n10924 = n10920 & n10923;
  assign n10925 = n10924 ^ x81;
  assign n10926 = n10925 ^ x82;
  assign n10927 = n10540 & n10784;
  assign n10928 = n10927 ^ n10542;
  assign n10929 = n10928 ^ n10925;
  assign n10930 = n10926 & ~n10929;
  assign n10931 = n10930 ^ x82;
  assign n10932 = n10931 ^ x83;
  assign n10933 = n10546 & n10784;
  assign n10934 = n10933 ^ n10548;
  assign n10935 = n10934 ^ n10931;
  assign n10936 = n10932 & ~n10935;
  assign n10937 = n10936 ^ x83;
  assign n10938 = n10937 ^ x84;
  assign n10939 = n10552 & n10784;
  assign n10940 = n10939 ^ n10554;
  assign n10941 = n10940 ^ n10937;
  assign n10942 = n10938 & ~n10941;
  assign n10943 = n10942 ^ x84;
  assign n10944 = n10943 ^ x85;
  assign n10945 = n10558 & n10784;
  assign n10946 = n10945 ^ n10560;
  assign n10947 = n10946 ^ n10943;
  assign n10948 = n10944 & ~n10947;
  assign n10949 = n10948 ^ x85;
  assign n10950 = n10949 ^ x86;
  assign n10951 = n10564 & n10784;
  assign n10952 = n10951 ^ n10566;
  assign n10953 = n10952 ^ n10949;
  assign n10954 = n10950 & ~n10953;
  assign n10955 = n10954 ^ x86;
  assign n10956 = n10955 ^ x87;
  assign n10957 = n10570 & n10784;
  assign n10958 = n10957 ^ n10572;
  assign n10959 = n10958 ^ n10955;
  assign n10960 = n10956 & ~n10959;
  assign n10961 = n10960 ^ x87;
  assign n10962 = n10961 ^ x88;
  assign n10963 = n10576 & n10784;
  assign n10964 = n10963 ^ n10578;
  assign n10965 = n10964 ^ n10961;
  assign n10966 = n10962 & ~n10965;
  assign n10967 = n10966 ^ x88;
  assign n10968 = n10967 ^ x89;
  assign n10969 = n10582 & n10784;
  assign n10970 = n10969 ^ n10584;
  assign n10971 = n10970 ^ n10967;
  assign n10972 = n10968 & ~n10971;
  assign n10973 = n10972 ^ x89;
  assign n10974 = n10973 ^ x90;
  assign n10975 = n10588 & n10784;
  assign n10976 = n10975 ^ n10590;
  assign n10977 = n10976 ^ n10973;
  assign n10978 = n10974 & ~n10977;
  assign n10979 = n10978 ^ x90;
  assign n10980 = n10979 ^ x91;
  assign n10981 = n10594 & n10784;
  assign n10982 = n10981 ^ n10596;
  assign n10983 = n10982 ^ n10979;
  assign n10984 = n10980 & ~n10983;
  assign n10985 = n10984 ^ x91;
  assign n10986 = n10985 ^ x92;
  assign n10987 = n10600 & n10784;
  assign n10988 = n10987 ^ n10602;
  assign n10989 = n10988 ^ n10985;
  assign n10990 = n10986 & ~n10989;
  assign n10991 = n10990 ^ x92;
  assign n10992 = n10791 & n10991;
  assign n10993 = n10786 ^ x94;
  assign n10994 = x93 & n10789;
  assign n10995 = n10994 ^ n10786;
  assign n10996 = n10993 & ~n10995;
  assign n10997 = n10996 ^ x94;
  assign n10998 = ~n10992 & ~n10997;
  assign n10999 = n10998 ^ x95;
  assign n11000 = n10640 & n10784;
  assign n11001 = n11000 ^ n10642;
  assign n11002 = n11001 ^ n10998;
  assign n11003 = ~n10999 & n11002;
  assign n11004 = n11003 ^ x95;
  assign n11005 = n11004 ^ x96;
  assign n11006 = n10646 & n10784;
  assign n11007 = n11006 ^ n10648;
  assign n11008 = n11007 ^ n11004;
  assign n11009 = n11005 & ~n11008;
  assign n11010 = n11009 ^ x96;
  assign n11011 = n11010 ^ x97;
  assign n11012 = n10652 & n10784;
  assign n11013 = n11012 ^ n10654;
  assign n11014 = n11013 ^ n11010;
  assign n11015 = n11011 & ~n11014;
  assign n11016 = n11015 ^ x97;
  assign n11017 = n11016 ^ x98;
  assign n11018 = n10658 & n10784;
  assign n11019 = n11018 ^ n10660;
  assign n11020 = n11019 ^ n11016;
  assign n11021 = n11017 & ~n11020;
  assign n11022 = n11021 ^ x98;
  assign n11023 = n11022 ^ x99;
  assign n11024 = n10664 & n10784;
  assign n11025 = n11024 ^ n10666;
  assign n11026 = n11025 ^ n11022;
  assign n11027 = n11023 & ~n11026;
  assign n11028 = n11027 ^ x99;
  assign n11029 = n11028 ^ x100;
  assign n11030 = n10670 & n10784;
  assign n11031 = n11030 ^ n10672;
  assign n11032 = n11031 ^ n11028;
  assign n11033 = n11029 & ~n11032;
  assign n11034 = n11033 ^ x100;
  assign n11035 = n11034 ^ x101;
  assign n11036 = n10676 & n10784;
  assign n11037 = n11036 ^ n10678;
  assign n11038 = n11037 ^ n11034;
  assign n11039 = n11035 & ~n11038;
  assign n11040 = n11039 ^ x101;
  assign n11041 = n11040 ^ x102;
  assign n11042 = n10682 & n10784;
  assign n11043 = n11042 ^ n10684;
  assign n11044 = n11043 ^ n11040;
  assign n11045 = n11041 & ~n11044;
  assign n11046 = n11045 ^ x102;
  assign n11047 = n11046 ^ x103;
  assign n11048 = n10688 & n10784;
  assign n11049 = n11048 ^ n10690;
  assign n11050 = n11049 ^ n11046;
  assign n11051 = n11047 & ~n11050;
  assign n11052 = n11051 ^ x103;
  assign n11053 = n11052 ^ x104;
  assign n11054 = n10694 & n10784;
  assign n11055 = n11054 ^ n10696;
  assign n11056 = n11055 ^ n11052;
  assign n11057 = n11053 & ~n11056;
  assign n11058 = n11057 ^ x104;
  assign n11059 = n11058 ^ x105;
  assign n11060 = n10700 & n10784;
  assign n11061 = n11060 ^ n10702;
  assign n11062 = n11061 ^ n11058;
  assign n11063 = n11059 & ~n11062;
  assign n11064 = n11063 ^ x105;
  assign n11065 = n11064 ^ x106;
  assign n11066 = n10706 & n10784;
  assign n11067 = n11066 ^ n10708;
  assign n11068 = n11067 ^ n11064;
  assign n11069 = n11065 & ~n11068;
  assign n11070 = n11069 ^ x106;
  assign n11071 = n11070 ^ x107;
  assign n11072 = n10755 ^ x115;
  assign n11073 = n10757 ^ n10755;
  assign n11074 = ~n11072 & n11073;
  assign n11075 = n11074 ^ x115;
  assign n11076 = n11075 ^ x116;
  assign n11077 = n10784 & n11076;
  assign n11078 = n11077 ^ n10760;
  assign n11079 = ~x117 & ~n11078;
  assign n11080 = n10769 ^ x117;
  assign n11081 = n10783 & ~n11080;
  assign n11082 = n11081 ^ n10773;
  assign n11083 = ~x118 & n11082;
  assign n11084 = ~n11079 & ~n11083;
  assign n11085 = n10712 & n10784;
  assign n11086 = n11085 ^ n10714;
  assign n11087 = n11086 ^ n11070;
  assign n11088 = n11071 & ~n11087;
  assign n11089 = n11088 ^ x107;
  assign n11090 = n11089 ^ x108;
  assign n11091 = n10717 ^ x107;
  assign n11092 = n10784 & n11091;
  assign n11093 = n11092 ^ n10629;
  assign n11094 = n11093 ^ n11089;
  assign n11095 = n11090 & ~n11094;
  assign n11096 = n11095 ^ x108;
  assign n11097 = n11096 ^ x109;
  assign n11098 = n10717 ^ n10629;
  assign n11099 = n11091 & ~n11098;
  assign n11100 = n11099 ^ x107;
  assign n11101 = n11100 ^ x108;
  assign n11102 = n10784 & n11101;
  assign n11103 = n11102 ^ n10632;
  assign n11104 = n11103 ^ n11096;
  assign n11105 = n11097 & ~n11104;
  assign n11106 = n11105 ^ x109;
  assign n11107 = n11106 ^ x110;
  assign n11108 = ~n10725 & n10784;
  assign n11109 = n11108 ^ n10727;
  assign n11110 = n11109 ^ n11106;
  assign n11111 = n11107 & ~n11110;
  assign n11112 = n11111 ^ x110;
  assign n11113 = n11112 ^ x111;
  assign n11114 = n10731 & n10784;
  assign n11115 = n11114 ^ n10733;
  assign n11116 = n11115 ^ n11112;
  assign n11117 = n11113 & ~n11116;
  assign n11118 = n11117 ^ x111;
  assign n11119 = n11118 ^ x112;
  assign n11120 = n10737 & n10784;
  assign n11121 = n11120 ^ n10739;
  assign n11122 = n11121 ^ n11118;
  assign n11123 = n11119 & ~n11122;
  assign n11124 = n11123 ^ x112;
  assign n11125 = n11124 ^ x113;
  assign n11126 = n10743 & n10784;
  assign n11127 = n11126 ^ n10745;
  assign n11128 = n11127 ^ n11124;
  assign n11129 = n11125 & ~n11128;
  assign n11130 = n11129 ^ x113;
  assign n11131 = n11130 ^ x114;
  assign n11132 = n10748 ^ x113;
  assign n11133 = n10784 & n11132;
  assign n11134 = n11133 ^ n10625;
  assign n11135 = n11134 ^ n11130;
  assign n11136 = n11131 & ~n11135;
  assign n11137 = n11136 ^ x114;
  assign n11138 = n11137 ^ x115;
  assign n11139 = n10748 ^ n10625;
  assign n11140 = n11132 & ~n11139;
  assign n11141 = n11140 ^ x113;
  assign n11142 = n11141 ^ x114;
  assign n11143 = n10784 & n11142;
  assign n11144 = n11143 ^ n10622;
  assign n11145 = n11144 ^ n11137;
  assign n11146 = n11138 & ~n11145;
  assign n11147 = n11146 ^ x115;
  assign n11148 = n11147 ^ x116;
  assign n11149 = n10784 & ~n11072;
  assign n11150 = n11149 ^ n10757;
  assign n11151 = n11150 ^ n11147;
  assign n11152 = n11148 & ~n11151;
  assign n11153 = n11152 ^ x116;
  assign n11154 = n11084 & n11153;
  assign n11155 = n11082 ^ x118;
  assign n11156 = x117 & n11078;
  assign n11157 = n11156 ^ n11082;
  assign n11158 = ~n11155 & n11157;
  assign n11159 = n11158 ^ x118;
  assign n11160 = ~n11154 & ~n11159;
  assign n11161 = x119 & ~n10037;
  assign n11162 = n9321 & ~n11161;
  assign n11163 = n11160 & n11162;
  assign n11164 = n10773 ^ n10769;
  assign n11165 = ~n11080 & ~n11164;
  assign n11166 = n11165 ^ x117;
  assign n11167 = n11166 ^ x118;
  assign n11168 = n9322 & n11167;
  assign n11169 = n10615 & ~n11168;
  assign n11170 = n9322 & n11169;
  assign n11171 = ~n11163 & ~n11170;
  assign n11172 = n11071 & ~n11171;
  assign n11173 = n11172 ^ n11086;
  assign n11174 = ~x108 & ~n11173;
  assign n11175 = n11065 & ~n11171;
  assign n11176 = n11175 ^ n11067;
  assign n11177 = ~x107 & ~n11176;
  assign n11178 = ~n11174 & ~n11177;
  assign n11179 = n11005 & ~n11171;
  assign n11180 = n11179 ^ n11007;
  assign n11181 = ~x97 & ~n11180;
  assign n11182 = n10902 & ~n11171;
  assign n11183 = n11182 ^ n10904;
  assign n11184 = ~x79 & ~n11183;
  assign n11185 = n10908 & ~n11171;
  assign n11186 = n11185 ^ n10910;
  assign n11187 = ~x80 & n11186;
  assign n11188 = ~n11184 & ~n11187;
  assign n11189 = n10855 & ~n11171;
  assign n11190 = n11189 ^ n10858;
  assign n11191 = ~x72 & n11190;
  assign n11192 = ~x65 & n11171;
  assign n11193 = ~x7 & x64;
  assign n11194 = n11192 & ~n11193;
  assign n11195 = x7 & ~x65;
  assign n11196 = n10813 & ~n11195;
  assign n11197 = n11196 ^ x8;
  assign n11198 = ~n11171 & ~n11197;
  assign n11199 = n11198 ^ x8;
  assign n11200 = ~n11194 & ~n11199;
  assign n11201 = x8 ^ x7;
  assign n11202 = ~x64 & n11201;
  assign n11203 = n11202 ^ x7;
  assign n11204 = x65 & ~n11203;
  assign n11205 = ~n11200 & ~n11204;
  assign n11206 = n11205 ^ x66;
  assign n11207 = x65 & n10784;
  assign n11208 = x8 & ~n11207;
  assign n11209 = ~n11171 & ~n11208;
  assign n11210 = n10805 & ~n11209;
  assign n11211 = n293 & ~n10784;
  assign n11212 = n11211 ^ x65;
  assign n11213 = ~x8 & n11212;
  assign n11214 = ~n202 & ~n11213;
  assign n11215 = x65 & n11208;
  assign n11216 = n11214 & ~n11215;
  assign n11217 = ~n11171 & ~n11216;
  assign n11218 = ~n11210 & ~n11217;
  assign n11219 = n11218 ^ x9;
  assign n11220 = n11219 ^ n11205;
  assign n11221 = ~n11206 & n11220;
  assign n11222 = n11221 ^ x66;
  assign n11223 = n11222 ^ x67;
  assign n11224 = n10818 ^ x66;
  assign n11225 = ~n11171 & ~n11224;
  assign n11226 = n11225 ^ n10803;
  assign n11227 = n11226 ^ n11222;
  assign n11228 = n11223 & ~n11227;
  assign n11229 = n11228 ^ x67;
  assign n11230 = n11229 ^ x68;
  assign n11231 = n10822 & ~n11171;
  assign n11232 = n11231 ^ n10833;
  assign n11233 = n11232 ^ n11229;
  assign n11234 = n11230 & n11233;
  assign n11235 = n11234 ^ x68;
  assign n11236 = n11235 ^ x69;
  assign n11237 = n10837 & ~n11171;
  assign n11238 = n11237 ^ n10839;
  assign n11239 = n11238 ^ n11235;
  assign n11240 = n11236 & ~n11239;
  assign n11241 = n11240 ^ x69;
  assign n11242 = n11241 ^ x70;
  assign n11243 = n10843 & ~n11171;
  assign n11244 = n11243 ^ n10845;
  assign n11245 = n11244 ^ n11241;
  assign n11246 = n11242 & n11245;
  assign n11247 = n11246 ^ x70;
  assign n11248 = n11247 ^ x71;
  assign n11249 = n10849 & ~n11171;
  assign n11250 = n11249 ^ n10851;
  assign n11251 = n11250 ^ n11247;
  assign n11252 = n11248 & ~n11251;
  assign n11253 = n11252 ^ x71;
  assign n11254 = ~n11191 & n11253;
  assign n11255 = n10862 & ~n11171;
  assign n11256 = n11255 ^ n10868;
  assign n11257 = x73 & ~n11256;
  assign n11258 = x72 & ~n11190;
  assign n11259 = ~n11257 & ~n11258;
  assign n11260 = ~n11254 & n11259;
  assign n11261 = ~x73 & n11256;
  assign n11262 = ~n11260 & ~n11261;
  assign n11263 = n11262 ^ x74;
  assign n11264 = n10872 & ~n11171;
  assign n11265 = n11264 ^ n10874;
  assign n11266 = n11265 ^ n11262;
  assign n11267 = n11263 & ~n11266;
  assign n11268 = n11267 ^ x74;
  assign n11269 = n11268 ^ x75;
  assign n11270 = n10878 & ~n11171;
  assign n11271 = n11270 ^ n10880;
  assign n11272 = n11271 ^ n11268;
  assign n11273 = n11269 & n11272;
  assign n11274 = n11273 ^ x75;
  assign n11275 = n11274 ^ x76;
  assign n11276 = n10884 & ~n11171;
  assign n11277 = n11276 ^ n10886;
  assign n11278 = n11277 ^ n11274;
  assign n11279 = n11275 & ~n11278;
  assign n11280 = n11279 ^ x76;
  assign n11281 = n11280 ^ x77;
  assign n11282 = n10890 & ~n11171;
  assign n11283 = n11282 ^ n10892;
  assign n11284 = n11283 ^ n11280;
  assign n11285 = n11281 & ~n11284;
  assign n11286 = n11285 ^ x77;
  assign n11287 = n11286 ^ x78;
  assign n11288 = n10896 & ~n11171;
  assign n11289 = n11288 ^ n10898;
  assign n11290 = n11289 ^ n11286;
  assign n11291 = n11287 & n11290;
  assign n11292 = n11291 ^ x78;
  assign n11293 = n11188 & n11292;
  assign n11294 = n11186 ^ x80;
  assign n11295 = x79 & n11183;
  assign n11296 = n11295 ^ n11186;
  assign n11297 = ~n11294 & n11296;
  assign n11298 = n11297 ^ x80;
  assign n11299 = ~n11293 & ~n11298;
  assign n11300 = n11299 ^ x81;
  assign n11301 = n10914 & ~n11171;
  assign n11302 = n11301 ^ n10916;
  assign n11303 = n11302 ^ n11299;
  assign n11304 = ~n11300 & n11303;
  assign n11305 = n11304 ^ x81;
  assign n11306 = n11305 ^ x82;
  assign n11307 = n10920 & ~n11171;
  assign n11308 = n11307 ^ n10922;
  assign n11309 = n11308 ^ n11305;
  assign n11310 = n11306 & n11309;
  assign n11311 = n11310 ^ x82;
  assign n11312 = n11311 ^ x83;
  assign n11313 = n10926 & ~n11171;
  assign n11314 = n11313 ^ n10928;
  assign n11315 = n11314 ^ n11311;
  assign n11316 = n11312 & ~n11315;
  assign n11317 = n11316 ^ x83;
  assign n11318 = n11317 ^ x84;
  assign n11319 = n10932 & ~n11171;
  assign n11320 = n11319 ^ n10934;
  assign n11321 = n11320 ^ n11317;
  assign n11322 = n11318 & ~n11321;
  assign n11323 = n11322 ^ x84;
  assign n11324 = n11323 ^ x85;
  assign n11325 = n10938 & ~n11171;
  assign n11326 = n11325 ^ n10940;
  assign n11327 = n11326 ^ n11323;
  assign n11328 = n11324 & ~n11327;
  assign n11329 = n11328 ^ x85;
  assign n11330 = n11329 ^ x86;
  assign n11331 = n10944 & ~n11171;
  assign n11332 = n11331 ^ n10946;
  assign n11333 = n11332 ^ n11329;
  assign n11334 = n11330 & ~n11333;
  assign n11335 = n11334 ^ x86;
  assign n11336 = n11335 ^ x87;
  assign n11337 = n10950 & ~n11171;
  assign n11338 = n11337 ^ n10952;
  assign n11339 = n11338 ^ n11335;
  assign n11340 = n11336 & ~n11339;
  assign n11341 = n11340 ^ x87;
  assign n11342 = n11341 ^ x88;
  assign n11343 = n10956 & ~n11171;
  assign n11344 = n11343 ^ n10958;
  assign n11345 = n11344 ^ n11341;
  assign n11346 = n11342 & ~n11345;
  assign n11347 = n11346 ^ x88;
  assign n11348 = n11347 ^ x89;
  assign n11349 = n10962 & ~n11171;
  assign n11350 = n11349 ^ n10964;
  assign n11351 = n11350 ^ n11347;
  assign n11352 = n11348 & ~n11351;
  assign n11353 = n11352 ^ x89;
  assign n11354 = n11353 ^ x90;
  assign n11355 = n10968 & ~n11171;
  assign n11356 = n11355 ^ n10970;
  assign n11357 = n11356 ^ n11353;
  assign n11358 = n11354 & ~n11357;
  assign n11359 = n11358 ^ x90;
  assign n11360 = n11359 ^ x91;
  assign n11361 = n10974 & ~n11171;
  assign n11362 = n11361 ^ n10976;
  assign n11363 = n11362 ^ n11359;
  assign n11364 = n11360 & ~n11363;
  assign n11365 = n11364 ^ x91;
  assign n11366 = n11365 ^ x92;
  assign n11367 = n10980 & ~n11171;
  assign n11368 = n11367 ^ n10982;
  assign n11369 = n11368 ^ n11365;
  assign n11370 = n11366 & ~n11369;
  assign n11371 = n11370 ^ x92;
  assign n11372 = n11371 ^ x93;
  assign n11373 = n10986 & ~n11171;
  assign n11374 = n11373 ^ n10988;
  assign n11375 = n11374 ^ n11371;
  assign n11376 = n11372 & ~n11375;
  assign n11377 = n11376 ^ x93;
  assign n11378 = n11377 ^ x94;
  assign n11379 = n10991 ^ x93;
  assign n11380 = ~n11171 & n11379;
  assign n11381 = n11380 ^ n10789;
  assign n11382 = n11381 ^ n11377;
  assign n11383 = n11378 & ~n11382;
  assign n11384 = n11383 ^ x94;
  assign n11385 = n11384 ^ x95;
  assign n11386 = n10991 ^ n10789;
  assign n11387 = n11379 & ~n11386;
  assign n11388 = n11387 ^ x93;
  assign n11389 = n11388 ^ x94;
  assign n11390 = ~n11171 & n11389;
  assign n11391 = n11390 ^ n10786;
  assign n11392 = n11391 ^ n11384;
  assign n11393 = n11385 & ~n11392;
  assign n11394 = n11393 ^ x95;
  assign n11395 = n11394 ^ x96;
  assign n11396 = ~n10999 & ~n11171;
  assign n11397 = n11396 ^ n11001;
  assign n11398 = n11397 ^ n11394;
  assign n11399 = n11395 & ~n11398;
  assign n11400 = n11399 ^ x96;
  assign n11401 = ~n11181 & n11400;
  assign n11402 = n11011 & ~n11171;
  assign n11403 = n11402 ^ n11013;
  assign n11404 = x98 & n11403;
  assign n11405 = x97 & n11180;
  assign n11406 = ~n11404 & ~n11405;
  assign n11407 = ~n11401 & n11406;
  assign n11408 = ~x98 & ~n11403;
  assign n11409 = ~n11407 & ~n11408;
  assign n11410 = n11409 ^ x99;
  assign n11411 = n11017 & ~n11171;
  assign n11412 = n11411 ^ n11019;
  assign n11413 = n11412 ^ n11409;
  assign n11414 = n11410 & ~n11413;
  assign n11415 = n11414 ^ x99;
  assign n11416 = n11415 ^ x100;
  assign n11417 = n11023 & ~n11171;
  assign n11418 = n11417 ^ n11025;
  assign n11419 = n11418 ^ n11415;
  assign n11420 = n11416 & ~n11419;
  assign n11421 = n11420 ^ x100;
  assign n11422 = n11421 ^ x101;
  assign n11423 = n11029 & ~n11171;
  assign n11424 = n11423 ^ n11031;
  assign n11425 = n11424 ^ n11421;
  assign n11426 = n11422 & ~n11425;
  assign n11427 = n11426 ^ x101;
  assign n11428 = n11427 ^ x102;
  assign n11429 = n11035 & ~n11171;
  assign n11430 = n11429 ^ n11037;
  assign n11431 = n11430 ^ n11427;
  assign n11432 = n11428 & ~n11431;
  assign n11433 = n11432 ^ x102;
  assign n11434 = n11433 ^ x103;
  assign n11435 = n11041 & ~n11171;
  assign n11436 = n11435 ^ n11043;
  assign n11437 = n11436 ^ n11433;
  assign n11438 = n11434 & ~n11437;
  assign n11439 = n11438 ^ x103;
  assign n11440 = n11439 ^ x104;
  assign n11441 = n11047 & ~n11171;
  assign n11442 = n11441 ^ n11049;
  assign n11443 = n11442 ^ n11439;
  assign n11444 = n11440 & ~n11443;
  assign n11445 = n11444 ^ x104;
  assign n11446 = n11445 ^ x105;
  assign n11447 = n11053 & ~n11171;
  assign n11448 = n11447 ^ n11055;
  assign n11449 = n11448 ^ n11445;
  assign n11450 = n11446 & ~n11449;
  assign n11451 = n11450 ^ x105;
  assign n11452 = n11451 ^ x106;
  assign n11453 = n11059 & ~n11171;
  assign n11454 = n11453 ^ n11061;
  assign n11455 = n11454 ^ n11451;
  assign n11456 = n11452 & ~n11455;
  assign n11457 = n11456 ^ x106;
  assign n11458 = n11178 & n11457;
  assign n11459 = n11173 ^ x108;
  assign n11460 = x107 & n11176;
  assign n11461 = n11460 ^ n11173;
  assign n11462 = n11459 & ~n11461;
  assign n11463 = n11462 ^ x108;
  assign n11464 = ~n11458 & ~n11463;
  assign n11465 = n11464 ^ x109;
  assign n11466 = n11093 ^ x108;
  assign n11467 = n11466 ^ n11089;
  assign n11468 = n11467 ^ n11093;
  assign n11469 = ~n11171 & n11468;
  assign n11470 = n11469 ^ n11093;
  assign n11471 = n11470 ^ n11464;
  assign n11472 = ~n11465 & n11471;
  assign n11473 = n11472 ^ x109;
  assign n11474 = n11473 ^ x110;
  assign n11475 = n11097 & ~n11171;
  assign n11476 = n11475 ^ n11103;
  assign n11477 = n11476 ^ n11473;
  assign n11478 = n11474 & ~n11477;
  assign n11479 = n11478 ^ x110;
  assign n11480 = n11479 ^ x111;
  assign n11481 = n11107 & ~n11171;
  assign n11482 = n11481 ^ n11109;
  assign n11483 = n11482 ^ n11479;
  assign n11484 = n11480 & ~n11483;
  assign n11485 = n11484 ^ x111;
  assign n11486 = n11485 ^ x112;
  assign n11487 = n11153 ^ x117;
  assign n11488 = ~n11171 & n11487;
  assign n11489 = n11488 ^ n11078;
  assign n11490 = ~x118 & ~n11489;
  assign n11491 = n11153 ^ n11078;
  assign n11492 = n11487 & ~n11491;
  assign n11493 = n11492 ^ x117;
  assign n11494 = n11493 ^ x118;
  assign n11495 = ~n11171 & n11494;
  assign n11496 = n11495 ^ n11082;
  assign n11497 = ~x119 & n11496;
  assign n11498 = ~n11490 & ~n11497;
  assign n11499 = n11113 & ~n11171;
  assign n11500 = n11499 ^ n11115;
  assign n11501 = n11500 ^ n11485;
  assign n11502 = n11486 & ~n11501;
  assign n11503 = n11502 ^ x112;
  assign n11504 = n11503 ^ x113;
  assign n11505 = n11119 & ~n11171;
  assign n11506 = n11505 ^ n11121;
  assign n11507 = n11506 ^ n11503;
  assign n11508 = n11504 & ~n11507;
  assign n11509 = n11508 ^ x113;
  assign n11510 = n11509 ^ x114;
  assign n11511 = n11125 & ~n11171;
  assign n11512 = n11511 ^ n11127;
  assign n11513 = n11512 ^ n11509;
  assign n11514 = n11510 & ~n11513;
  assign n11515 = n11514 ^ x114;
  assign n11516 = n11515 ^ x115;
  assign n11517 = n11131 & ~n11171;
  assign n11518 = n11517 ^ n11134;
  assign n11519 = n11518 ^ n11515;
  assign n11520 = n11516 & ~n11519;
  assign n11521 = n11520 ^ x115;
  assign n11522 = n11521 ^ x116;
  assign n11523 = n11138 & ~n11171;
  assign n11524 = n11523 ^ n11144;
  assign n11525 = n11524 ^ n11521;
  assign n11526 = n11522 & ~n11525;
  assign n11527 = n11526 ^ x116;
  assign n11528 = n11527 ^ x117;
  assign n11529 = n11148 & ~n11171;
  assign n11530 = n11529 ^ n11150;
  assign n11531 = n11530 ^ n11527;
  assign n11532 = n11528 & ~n11531;
  assign n11533 = n11532 ^ x117;
  assign n11534 = n11498 & n11533;
  assign n11535 = n11496 ^ x119;
  assign n11536 = x118 & n11489;
  assign n11537 = n11536 ^ n11496;
  assign n11538 = ~n11535 & n11537;
  assign n11539 = n11538 ^ x119;
  assign n11540 = ~n11534 & ~n11539;
  assign n11541 = n11160 ^ x119;
  assign n11542 = n9321 & ~n11541;
  assign n11543 = n11169 & ~n11542;
  assign n11544 = ~x120 & n11543;
  assign n11545 = ~n11540 & ~n11544;
  assign n11546 = x120 & ~n10615;
  assign n11547 = n135 & ~n11546;
  assign n11548 = ~n11545 & n11547;
  assign n11549 = n11486 & n11548;
  assign n11550 = n11549 ^ n11500;
  assign n11551 = ~x113 & ~n11550;
  assign n11552 = n11480 & n11548;
  assign n11553 = n11552 ^ n11482;
  assign n11554 = ~x112 & ~n11553;
  assign n11555 = ~n11551 & ~n11554;
  assign n11556 = n11457 ^ x107;
  assign n11557 = n11548 & n11556;
  assign n11558 = n11557 ^ n11176;
  assign n11559 = ~x108 & ~n11558;
  assign n11560 = n11457 ^ n11176;
  assign n11561 = n11556 & ~n11560;
  assign n11562 = n11561 ^ x107;
  assign n11563 = n11562 ^ x108;
  assign n11564 = n11548 & n11563;
  assign n11565 = n11564 ^ n11173;
  assign n11566 = ~x109 & ~n11565;
  assign n11567 = ~n11559 & ~n11566;
  assign n11568 = ~n11401 & ~n11405;
  assign n11569 = n11568 ^ x98;
  assign n11570 = n11548 & ~n11569;
  assign n11571 = n11570 ^ n11403;
  assign n11572 = ~x99 & ~n11571;
  assign n11573 = n11378 & n11548;
  assign n11574 = n11573 ^ n11381;
  assign n11575 = ~x95 & ~n11574;
  assign n11576 = n11342 & n11548;
  assign n11577 = n11576 ^ n11344;
  assign n11578 = ~x89 & ~n11577;
  assign n11579 = n11269 & n11548;
  assign n11580 = n11579 ^ n11271;
  assign n11581 = ~x76 & n11580;
  assign n11582 = n11275 & n11548;
  assign n11583 = n11582 ^ n11277;
  assign n11584 = ~x77 & ~n11583;
  assign n11585 = ~n11581 & ~n11584;
  assign n11586 = ~n11195 & n11548;
  assign n11587 = x64 & ~n11171;
  assign n11588 = ~n11586 & n11587;
  assign n11589 = x7 & n11171;
  assign n11590 = ~n11192 & n11589;
  assign n11591 = ~n202 & ~n11590;
  assign n11592 = n11171 ^ x65;
  assign n11593 = n11193 & n11592;
  assign n11594 = n11591 & ~n11593;
  assign n11595 = n11548 & ~n11594;
  assign n11596 = ~n11588 & ~n11595;
  assign n11597 = n11596 ^ x8;
  assign n11598 = n11597 ^ x66;
  assign n11599 = x64 & n11548;
  assign n11600 = x6 & n11195;
  assign n11601 = n11600 ^ x7;
  assign n11602 = n11599 & n11601;
  assign n11603 = ~x6 & n219;
  assign n11604 = n11603 ^ x65;
  assign n11605 = ~x7 & n11604;
  assign n11606 = ~n11548 & n11605;
  assign n11607 = x6 & x64;
  assign n11608 = x65 & ~n11607;
  assign n11609 = x7 & ~x64;
  assign n11610 = n11608 & ~n11609;
  assign n11611 = ~n11606 & ~n11610;
  assign n11612 = ~n11602 & n11611;
  assign n11613 = n11612 ^ n11597;
  assign n11614 = n11598 & n11613;
  assign n11615 = n11614 ^ x66;
  assign n11616 = n11615 ^ x67;
  assign n11617 = ~n11206 & n11548;
  assign n11618 = n11617 ^ n11219;
  assign n11619 = n11618 ^ n11615;
  assign n11620 = n11616 & ~n11619;
  assign n11621 = n11620 ^ x67;
  assign n11622 = n11621 ^ x68;
  assign n11623 = n11223 & n11548;
  assign n11624 = n11623 ^ n11226;
  assign n11625 = n11624 ^ n11621;
  assign n11626 = n11622 & ~n11625;
  assign n11627 = n11626 ^ x68;
  assign n11628 = n11627 ^ x69;
  assign n11629 = n11230 & n11548;
  assign n11630 = n11629 ^ n11232;
  assign n11631 = n11630 ^ n11627;
  assign n11632 = n11628 & n11631;
  assign n11633 = n11632 ^ x69;
  assign n11634 = n11633 ^ x70;
  assign n11635 = n11236 & n11548;
  assign n11636 = n11635 ^ n11238;
  assign n11637 = n11636 ^ n11633;
  assign n11638 = n11634 & ~n11637;
  assign n11639 = n11638 ^ x70;
  assign n11640 = n11639 ^ x71;
  assign n11641 = n11242 & n11548;
  assign n11642 = n11641 ^ n11244;
  assign n11643 = n11642 ^ n11639;
  assign n11644 = n11640 & n11643;
  assign n11645 = n11644 ^ x71;
  assign n11646 = n11645 ^ x72;
  assign n11647 = n11248 & n11548;
  assign n11648 = n11647 ^ n11250;
  assign n11649 = n11648 ^ n11645;
  assign n11650 = n11646 & ~n11649;
  assign n11651 = n11650 ^ x72;
  assign n11652 = n11651 ^ x73;
  assign n11653 = n11253 ^ x72;
  assign n11654 = n11548 & n11653;
  assign n11655 = n11654 ^ n11190;
  assign n11656 = n11655 ^ n11651;
  assign n11657 = n11652 & n11656;
  assign n11658 = n11657 ^ x73;
  assign n11659 = n11658 ^ x74;
  assign n11660 = ~n11254 & ~n11258;
  assign n11661 = n11660 ^ x73;
  assign n11662 = n11548 & ~n11661;
  assign n11663 = n11662 ^ n11256;
  assign n11664 = n11663 ^ n11658;
  assign n11665 = n11659 & n11664;
  assign n11666 = n11665 ^ x74;
  assign n11667 = n11666 ^ x75;
  assign n11668 = n11263 & n11548;
  assign n11669 = n11668 ^ n11265;
  assign n11670 = n11669 ^ n11666;
  assign n11671 = n11667 & ~n11670;
  assign n11672 = n11671 ^ x75;
  assign n11673 = n11585 & n11672;
  assign n11674 = n11583 ^ x77;
  assign n11675 = x76 & ~n11580;
  assign n11676 = n11675 ^ n11583;
  assign n11677 = n11674 & ~n11676;
  assign n11678 = n11677 ^ x77;
  assign n11679 = ~n11673 & ~n11678;
  assign n11680 = n11679 ^ x78;
  assign n11681 = n11281 & n11548;
  assign n11682 = n11681 ^ n11283;
  assign n11683 = n11682 ^ n11679;
  assign n11684 = ~n11680 & n11683;
  assign n11685 = n11684 ^ x78;
  assign n11686 = n11685 ^ x79;
  assign n11687 = n11287 & n11548;
  assign n11688 = n11687 ^ n11289;
  assign n11689 = n11688 ^ n11685;
  assign n11690 = n11686 & n11689;
  assign n11691 = n11690 ^ x79;
  assign n11692 = n11691 ^ x80;
  assign n11693 = n11292 ^ x79;
  assign n11694 = n11548 & n11693;
  assign n11695 = n11694 ^ n11183;
  assign n11696 = n11695 ^ n11691;
  assign n11697 = n11692 & ~n11696;
  assign n11698 = n11697 ^ x80;
  assign n11699 = n11698 ^ x81;
  assign n11700 = n11292 ^ n11183;
  assign n11701 = n11693 & ~n11700;
  assign n11702 = n11701 ^ x79;
  assign n11703 = n11702 ^ x80;
  assign n11704 = n11548 & n11703;
  assign n11705 = n11704 ^ n11186;
  assign n11706 = n11705 ^ n11698;
  assign n11707 = n11699 & n11706;
  assign n11708 = n11707 ^ x81;
  assign n11709 = n11708 ^ x82;
  assign n11710 = ~n11300 & n11548;
  assign n11711 = n11710 ^ n11302;
  assign n11712 = n11711 ^ n11708;
  assign n11713 = n11709 & ~n11712;
  assign n11714 = n11713 ^ x82;
  assign n11715 = n11714 ^ x83;
  assign n11716 = n11306 & n11548;
  assign n11717 = n11716 ^ n11308;
  assign n11718 = n11717 ^ n11714;
  assign n11719 = n11715 & n11718;
  assign n11720 = n11719 ^ x83;
  assign n11721 = n11720 ^ x84;
  assign n11722 = n11312 & n11548;
  assign n11723 = n11722 ^ n11314;
  assign n11724 = n11723 ^ n11720;
  assign n11725 = n11721 & ~n11724;
  assign n11726 = n11725 ^ x84;
  assign n11727 = n11726 ^ x85;
  assign n11728 = n11318 & n11548;
  assign n11729 = n11728 ^ n11320;
  assign n11730 = n11729 ^ n11726;
  assign n11731 = n11727 & ~n11730;
  assign n11732 = n11731 ^ x85;
  assign n11733 = n11732 ^ x86;
  assign n11734 = n11324 & n11548;
  assign n11735 = n11734 ^ n11326;
  assign n11736 = n11735 ^ n11732;
  assign n11737 = n11733 & ~n11736;
  assign n11738 = n11737 ^ x86;
  assign n11739 = n11738 ^ x87;
  assign n11740 = n11330 & n11548;
  assign n11741 = n11740 ^ n11332;
  assign n11742 = n11741 ^ n11738;
  assign n11743 = n11739 & ~n11742;
  assign n11744 = n11743 ^ x87;
  assign n11745 = n11744 ^ x88;
  assign n11746 = n11336 & n11548;
  assign n11747 = n11746 ^ n11338;
  assign n11748 = n11747 ^ n11744;
  assign n11749 = n11745 & ~n11748;
  assign n11750 = n11749 ^ x88;
  assign n11751 = ~n11578 & n11750;
  assign n11752 = n11348 & n11548;
  assign n11753 = n11752 ^ n11350;
  assign n11754 = x90 & n11753;
  assign n11755 = x89 & n11577;
  assign n11756 = ~n11754 & ~n11755;
  assign n11757 = ~n11751 & n11756;
  assign n11758 = ~x90 & ~n11753;
  assign n11759 = ~n11757 & ~n11758;
  assign n11760 = n11759 ^ x91;
  assign n11761 = n11354 & n11548;
  assign n11762 = n11761 ^ n11356;
  assign n11763 = n11762 ^ n11759;
  assign n11764 = n11760 & ~n11763;
  assign n11765 = n11764 ^ x91;
  assign n11766 = n11765 ^ x92;
  assign n11767 = n11360 & n11548;
  assign n11768 = n11767 ^ n11362;
  assign n11769 = n11768 ^ n11765;
  assign n11770 = n11766 & ~n11769;
  assign n11771 = n11770 ^ x92;
  assign n11772 = n11771 ^ x93;
  assign n11773 = n11366 & n11548;
  assign n11774 = n11773 ^ n11368;
  assign n11775 = n11774 ^ n11771;
  assign n11776 = n11772 & ~n11775;
  assign n11777 = n11776 ^ x93;
  assign n11778 = n11777 ^ x94;
  assign n11779 = n11372 & n11548;
  assign n11780 = n11779 ^ n11374;
  assign n11781 = n11780 ^ n11777;
  assign n11782 = n11778 & ~n11781;
  assign n11783 = n11782 ^ x94;
  assign n11784 = ~n11575 & n11783;
  assign n11785 = n11385 & n11548;
  assign n11786 = n11785 ^ n11391;
  assign n11787 = x96 & n11786;
  assign n11788 = x95 & n11574;
  assign n11789 = ~n11787 & ~n11788;
  assign n11790 = ~n11784 & n11789;
  assign n11791 = ~x96 & ~n11786;
  assign n11792 = ~n11790 & ~n11791;
  assign n11793 = n11792 ^ x97;
  assign n11794 = n11395 & n11548;
  assign n11795 = n11794 ^ n11397;
  assign n11796 = n11795 ^ n11792;
  assign n11797 = n11793 & ~n11796;
  assign n11798 = n11797 ^ x97;
  assign n11799 = n11798 ^ x98;
  assign n11800 = n11400 ^ x97;
  assign n11801 = n11548 & n11800;
  assign n11802 = n11801 ^ n11180;
  assign n11803 = n11802 ^ n11798;
  assign n11804 = n11799 & ~n11803;
  assign n11805 = n11804 ^ x98;
  assign n11806 = ~n11572 & n11805;
  assign n11807 = n11410 & n11548;
  assign n11808 = n11807 ^ n11412;
  assign n11809 = x100 & n11808;
  assign n11810 = x99 & n11571;
  assign n11811 = ~n11809 & ~n11810;
  assign n11812 = ~n11806 & n11811;
  assign n11813 = ~x100 & ~n11808;
  assign n11814 = ~n11812 & ~n11813;
  assign n11815 = n11814 ^ x101;
  assign n11816 = n11416 & n11548;
  assign n11817 = n11816 ^ n11418;
  assign n11818 = n11817 ^ n11814;
  assign n11819 = n11815 & ~n11818;
  assign n11820 = n11819 ^ x101;
  assign n11821 = n11820 ^ x102;
  assign n11822 = n11422 & n11548;
  assign n11823 = n11822 ^ n11424;
  assign n11824 = n11823 ^ n11820;
  assign n11825 = n11821 & ~n11824;
  assign n11826 = n11825 ^ x102;
  assign n11827 = n11826 ^ x103;
  assign n11828 = n11428 & n11548;
  assign n11829 = n11828 ^ n11430;
  assign n11830 = n11829 ^ n11826;
  assign n11831 = n11827 & ~n11830;
  assign n11832 = n11831 ^ x103;
  assign n11833 = n11832 ^ x104;
  assign n11834 = n11434 & n11548;
  assign n11835 = n11834 ^ n11436;
  assign n11836 = n11835 ^ n11832;
  assign n11837 = n11833 & ~n11836;
  assign n11838 = n11837 ^ x104;
  assign n11839 = n11838 ^ x105;
  assign n11840 = n11440 & n11548;
  assign n11841 = n11840 ^ n11442;
  assign n11842 = n11841 ^ n11838;
  assign n11843 = n11839 & ~n11842;
  assign n11844 = n11843 ^ x105;
  assign n11845 = n11844 ^ x106;
  assign n11846 = n11446 & n11548;
  assign n11847 = n11846 ^ n11448;
  assign n11848 = n11847 ^ n11844;
  assign n11849 = n11845 & ~n11848;
  assign n11850 = n11849 ^ x106;
  assign n11851 = n11850 ^ x107;
  assign n11852 = n11452 & n11548;
  assign n11853 = n11852 ^ n11454;
  assign n11854 = n11853 ^ n11850;
  assign n11855 = n11851 & ~n11854;
  assign n11856 = n11855 ^ x107;
  assign n11857 = n11567 & n11856;
  assign n11858 = n11565 ^ x109;
  assign n11859 = x108 & n11558;
  assign n11860 = n11859 ^ n11565;
  assign n11861 = n11858 & ~n11860;
  assign n11862 = n11861 ^ x109;
  assign n11863 = ~n11857 & ~n11862;
  assign n11864 = n11863 ^ x110;
  assign n11865 = ~n11465 & n11548;
  assign n11866 = n11865 ^ n11470;
  assign n11867 = n11866 ^ n11863;
  assign n11868 = ~n11864 & n11867;
  assign n11869 = n11868 ^ x110;
  assign n11870 = n11869 ^ x111;
  assign n11871 = n11474 & n11548;
  assign n11872 = n11871 ^ n11476;
  assign n11873 = n11872 ^ n11869;
  assign n11874 = n11870 & ~n11873;
  assign n11875 = n11874 ^ x111;
  assign n11876 = n11555 & n11875;
  assign n11877 = n11550 ^ x113;
  assign n11878 = x112 & n11553;
  assign n11879 = n11878 ^ n11550;
  assign n11880 = n11877 & ~n11879;
  assign n11881 = n11880 ^ x113;
  assign n11882 = ~n11876 & ~n11881;
  assign n11883 = n11882 ^ x114;
  assign n11884 = n11504 & n11548;
  assign n11885 = n11884 ^ n11506;
  assign n11886 = n11885 ^ n11882;
  assign n11887 = ~n11883 & n11886;
  assign n11888 = n11887 ^ x114;
  assign n11889 = n11888 ^ x115;
  assign n11890 = n11510 & n11548;
  assign n11891 = n11890 ^ n11512;
  assign n11892 = n11891 ^ n11888;
  assign n11893 = n11889 & ~n11892;
  assign n11894 = n11893 ^ x115;
  assign n11895 = n11894 ^ x116;
  assign n11896 = n11516 & n11548;
  assign n11897 = n11896 ^ n11518;
  assign n11898 = n11897 ^ n11894;
  assign n11899 = n11895 & ~n11898;
  assign n11900 = n11899 ^ x116;
  assign n11901 = n11900 ^ x117;
  assign n11902 = n11540 ^ x120;
  assign n11903 = n135 & ~n11902;
  assign n11904 = n11543 & ~n11903;
  assign n11905 = ~x121 & n11904;
  assign n11906 = n11522 & n11548;
  assign n11907 = n11906 ^ n11524;
  assign n11908 = n11907 ^ n11900;
  assign n11909 = n11901 & ~n11908;
  assign n11910 = n11909 ^ x117;
  assign n11911 = n11910 ^ x118;
  assign n11912 = n11528 & n11548;
  assign n11913 = n11912 ^ n11530;
  assign n11914 = n11913 ^ n11910;
  assign n11915 = n11911 & ~n11914;
  assign n11916 = n11915 ^ x118;
  assign n11917 = n11916 ^ x119;
  assign n11918 = n11533 ^ x118;
  assign n11919 = n11548 & n11918;
  assign n11920 = n11919 ^ n11489;
  assign n11921 = n11920 ^ n11916;
  assign n11922 = n11917 & ~n11921;
  assign n11923 = n11922 ^ x119;
  assign n11924 = n11923 ^ x120;
  assign n11925 = n11533 ^ n11489;
  assign n11926 = n11918 & ~n11925;
  assign n11927 = n11926 ^ x118;
  assign n11928 = n11927 ^ x119;
  assign n11929 = n11548 & n11928;
  assign n11930 = n11929 ^ n11496;
  assign n11931 = n11930 ^ n11923;
  assign n11932 = n11924 & n11931;
  assign n11933 = n11932 ^ x120;
  assign n11934 = ~n11905 & n11933;
  assign n11935 = x121 & ~n11169;
  assign n11936 = n134 & ~n11935;
  assign n11937 = ~n11934 & n11936;
  assign n11938 = n11901 & n11937;
  assign n11939 = n11938 ^ n11907;
  assign n11940 = ~x118 & ~n11939;
  assign n11941 = n11875 ^ x112;
  assign n11942 = n11875 ^ n11553;
  assign n11943 = n11941 & ~n11942;
  assign n11944 = n11943 ^ x112;
  assign n11945 = n11944 ^ x113;
  assign n11946 = n11937 & n11945;
  assign n11947 = n11946 ^ n11550;
  assign n11948 = ~x114 & ~n11947;
  assign n11949 = n11845 & n11937;
  assign n11950 = n11949 ^ n11847;
  assign n11951 = ~x107 & ~n11950;
  assign n11952 = n11851 & n11937;
  assign n11953 = n11952 ^ n11853;
  assign n11954 = ~x108 & ~n11953;
  assign n11955 = ~n11951 & ~n11954;
  assign n11956 = n11766 & n11937;
  assign n11957 = n11956 ^ n11768;
  assign n11958 = ~x93 & ~n11957;
  assign n11959 = n11733 & n11937;
  assign n11960 = n11959 ^ n11735;
  assign n11961 = ~x87 & ~n11960;
  assign n11962 = n11667 & n11937;
  assign n11963 = n11962 ^ n11669;
  assign n11964 = ~x76 & ~n11963;
  assign n11965 = x65 & ~n11548;
  assign n11966 = n11937 & n11965;
  assign n11967 = n219 & n11548;
  assign n11968 = ~n11966 & ~n11967;
  assign n11969 = x6 & ~n11968;
  assign n11970 = n11548 ^ x65;
  assign n11971 = n341 & ~n11970;
  assign n11972 = x6 & n11971;
  assign n11973 = n11972 ^ n340;
  assign n11974 = n11937 & n11973;
  assign n11975 = n11974 ^ n11599;
  assign n11976 = ~n11969 & ~n11975;
  assign n11977 = n11976 ^ x7;
  assign n11978 = n11977 ^ x66;
  assign n11979 = ~x5 & x64;
  assign n11980 = ~x65 & ~n11979;
  assign n11981 = ~x6 & ~n11980;
  assign n11982 = ~n11937 & n11981;
  assign n11983 = x6 ^ x5;
  assign n11984 = ~x64 & n11983;
  assign n11985 = n11984 ^ x5;
  assign n11986 = x65 & ~n11985;
  assign n11987 = ~n11982 & ~n11986;
  assign n11988 = x5 & ~x65;
  assign n11989 = n11607 & ~n11988;
  assign n11990 = n11937 & n11989;
  assign n11991 = n11987 & ~n11990;
  assign n11992 = n11991 ^ n11977;
  assign n11993 = n11978 & n11992;
  assign n11994 = n11993 ^ x66;
  assign n11995 = n11994 ^ x67;
  assign n11996 = n11612 ^ x66;
  assign n11997 = n11937 & ~n11996;
  assign n11998 = n11997 ^ n11597;
  assign n11999 = n11998 ^ n11994;
  assign n12000 = n11995 & ~n11999;
  assign n12001 = n12000 ^ x67;
  assign n12002 = n12001 ^ x68;
  assign n12003 = n11616 & n11937;
  assign n12004 = n12003 ^ n11618;
  assign n12005 = n12004 ^ n12001;
  assign n12006 = n12002 & ~n12005;
  assign n12007 = n12006 ^ x68;
  assign n12008 = n12007 ^ x69;
  assign n12009 = n11622 & n11937;
  assign n12010 = n12009 ^ n11624;
  assign n12011 = n12010 ^ n12007;
  assign n12012 = n12008 & ~n12011;
  assign n12013 = n12012 ^ x69;
  assign n12014 = n12013 ^ x70;
  assign n12015 = n11628 & n11937;
  assign n12016 = n12015 ^ n11630;
  assign n12017 = n12016 ^ n12013;
  assign n12018 = n12014 & n12017;
  assign n12019 = n12018 ^ x70;
  assign n12020 = n12019 ^ x71;
  assign n12021 = n11634 & n11937;
  assign n12022 = n12021 ^ n11636;
  assign n12023 = n12022 ^ n12019;
  assign n12024 = n12020 & ~n12023;
  assign n12025 = n12024 ^ x71;
  assign n12026 = n12025 ^ x72;
  assign n12027 = n11640 & n11937;
  assign n12028 = n12027 ^ n11642;
  assign n12029 = n12028 ^ n12025;
  assign n12030 = n12026 & n12029;
  assign n12031 = n12030 ^ x72;
  assign n12032 = n12031 ^ x73;
  assign n12033 = n11646 & n11937;
  assign n12034 = n12033 ^ n11648;
  assign n12035 = n12034 ^ n12031;
  assign n12036 = n12032 & ~n12035;
  assign n12037 = n12036 ^ x73;
  assign n12038 = n12037 ^ x74;
  assign n12039 = n11652 & n11937;
  assign n12040 = n12039 ^ n11655;
  assign n12041 = n12040 ^ n12037;
  assign n12042 = n12038 & n12041;
  assign n12043 = n12042 ^ x74;
  assign n12044 = n12043 ^ x75;
  assign n12045 = n11659 & n11937;
  assign n12046 = n12045 ^ n11663;
  assign n12047 = n12046 ^ n12043;
  assign n12048 = n12044 & n12047;
  assign n12049 = n12048 ^ x75;
  assign n12050 = ~n11964 & n12049;
  assign n12051 = n11672 ^ x76;
  assign n12052 = n11937 & n12051;
  assign n12053 = n12052 ^ n11580;
  assign n12054 = x77 & ~n12053;
  assign n12055 = x76 & n11963;
  assign n12056 = ~n12054 & ~n12055;
  assign n12057 = ~n12050 & n12056;
  assign n12058 = ~x77 & n12053;
  assign n12059 = ~n12057 & ~n12058;
  assign n12060 = n12059 ^ x78;
  assign n12061 = n11672 ^ n11580;
  assign n12062 = n12051 & n12061;
  assign n12063 = n12062 ^ x76;
  assign n12064 = n12063 ^ x77;
  assign n12065 = n11937 & n12064;
  assign n12066 = n12065 ^ n11583;
  assign n12067 = n12066 ^ n12059;
  assign n12068 = n12060 & ~n12067;
  assign n12069 = n12068 ^ x78;
  assign n12070 = n12069 ^ x79;
  assign n12071 = ~n11680 & n11937;
  assign n12072 = n12071 ^ n11682;
  assign n12073 = n12072 ^ n12069;
  assign n12074 = n12070 & ~n12073;
  assign n12075 = n12074 ^ x79;
  assign n12076 = n12075 ^ x80;
  assign n12077 = n11686 & n11937;
  assign n12078 = n12077 ^ n11688;
  assign n12079 = n12078 ^ n12075;
  assign n12080 = n12076 & n12079;
  assign n12081 = n12080 ^ x80;
  assign n12082 = n12081 ^ x81;
  assign n12083 = n11692 & n11937;
  assign n12084 = n12083 ^ n11695;
  assign n12085 = n12084 ^ n12081;
  assign n12086 = n12082 & ~n12085;
  assign n12087 = n12086 ^ x81;
  assign n12088 = n12087 ^ x82;
  assign n12089 = n11699 & n11937;
  assign n12090 = n12089 ^ n11705;
  assign n12091 = n12090 ^ n12087;
  assign n12092 = n12088 & n12091;
  assign n12093 = n12092 ^ x82;
  assign n12094 = n12093 ^ x83;
  assign n12095 = n11709 & n11937;
  assign n12096 = n12095 ^ n11711;
  assign n12097 = n12096 ^ n12093;
  assign n12098 = n12094 & ~n12097;
  assign n12099 = n12098 ^ x83;
  assign n12100 = n12099 ^ x84;
  assign n12101 = n11715 & n11937;
  assign n12102 = n12101 ^ n11717;
  assign n12103 = n12102 ^ n12099;
  assign n12104 = n12100 & n12103;
  assign n12105 = n12104 ^ x84;
  assign n12106 = n12105 ^ x85;
  assign n12107 = n11721 & n11937;
  assign n12108 = n12107 ^ n11723;
  assign n12109 = n12108 ^ n12105;
  assign n12110 = n12106 & ~n12109;
  assign n12111 = n12110 ^ x85;
  assign n12112 = n12111 ^ x86;
  assign n12113 = n11727 & n11937;
  assign n12114 = n12113 ^ n11729;
  assign n12115 = n12114 ^ n12111;
  assign n12116 = n12112 & ~n12115;
  assign n12117 = n12116 ^ x86;
  assign n12118 = ~n11961 & n12117;
  assign n12119 = n11739 & n11937;
  assign n12120 = n12119 ^ n11741;
  assign n12121 = x88 & n12120;
  assign n12122 = x87 & n11960;
  assign n12123 = ~n12121 & ~n12122;
  assign n12124 = ~n12118 & n12123;
  assign n12125 = ~x88 & ~n12120;
  assign n12126 = ~n12124 & ~n12125;
  assign n12127 = n12126 ^ x89;
  assign n12128 = n11745 & n11937;
  assign n12129 = n12128 ^ n11747;
  assign n12130 = n12129 ^ n12126;
  assign n12131 = n12127 & ~n12130;
  assign n12132 = n12131 ^ x89;
  assign n12133 = n12132 ^ x90;
  assign n12134 = n11750 ^ x89;
  assign n12135 = n11937 & n12134;
  assign n12136 = n12135 ^ n11577;
  assign n12137 = n12136 ^ n12132;
  assign n12138 = n12133 & ~n12137;
  assign n12139 = n12138 ^ x90;
  assign n12140 = n12139 ^ x91;
  assign n12141 = ~n11751 & ~n11755;
  assign n12142 = n12141 ^ x90;
  assign n12143 = n11937 & ~n12142;
  assign n12144 = n12143 ^ n11753;
  assign n12145 = n12144 ^ n12139;
  assign n12146 = n12140 & ~n12145;
  assign n12147 = n12146 ^ x91;
  assign n12148 = n12147 ^ x92;
  assign n12149 = n11760 & n11937;
  assign n12150 = n12149 ^ n11762;
  assign n12151 = n12150 ^ n12147;
  assign n12152 = n12148 & ~n12151;
  assign n12153 = n12152 ^ x92;
  assign n12154 = ~n11958 & n12153;
  assign n12155 = n11772 & n11937;
  assign n12156 = n12155 ^ n11774;
  assign n12157 = x94 & n12156;
  assign n12158 = x93 & n11957;
  assign n12159 = ~n12157 & ~n12158;
  assign n12160 = ~n12154 & n12159;
  assign n12161 = ~x94 & ~n12156;
  assign n12162 = ~n12160 & ~n12161;
  assign n12163 = n12162 ^ x95;
  assign n12164 = n11778 & n11937;
  assign n12165 = n12164 ^ n11780;
  assign n12166 = n12165 ^ n12162;
  assign n12167 = n12163 & ~n12166;
  assign n12168 = n12167 ^ x95;
  assign n12169 = n12168 ^ x96;
  assign n12170 = n11783 ^ x95;
  assign n12171 = n11937 & n12170;
  assign n12172 = n12171 ^ n11574;
  assign n12173 = n12172 ^ n12168;
  assign n12174 = n12169 & ~n12173;
  assign n12175 = n12174 ^ x96;
  assign n12176 = n12175 ^ x97;
  assign n12177 = ~n11784 & ~n11788;
  assign n12178 = n12177 ^ x96;
  assign n12179 = n11937 & ~n12178;
  assign n12180 = n12179 ^ n11786;
  assign n12181 = n12180 ^ n12175;
  assign n12182 = n12176 & ~n12181;
  assign n12183 = n12182 ^ x97;
  assign n12184 = n12183 ^ x98;
  assign n12185 = n11793 & n11937;
  assign n12186 = n12185 ^ n11795;
  assign n12187 = n12186 ^ n12183;
  assign n12188 = n12184 & ~n12187;
  assign n12189 = n12188 ^ x98;
  assign n12190 = n12189 ^ x99;
  assign n12191 = n11799 & n11937;
  assign n12192 = n12191 ^ n11802;
  assign n12193 = n12192 ^ n12189;
  assign n12194 = n12190 & ~n12193;
  assign n12195 = n12194 ^ x99;
  assign n12196 = n12195 ^ x100;
  assign n12197 = n11805 ^ x99;
  assign n12198 = n11937 & n12197;
  assign n12199 = n12198 ^ n11571;
  assign n12200 = n12199 ^ n12195;
  assign n12201 = n12196 & ~n12200;
  assign n12202 = n12201 ^ x100;
  assign n12203 = n12202 ^ x101;
  assign n12204 = ~n11806 & ~n11810;
  assign n12205 = n12204 ^ x100;
  assign n12206 = n11937 & ~n12205;
  assign n12207 = n12206 ^ n11808;
  assign n12208 = n12207 ^ n12202;
  assign n12209 = n12203 & ~n12208;
  assign n12210 = n12209 ^ x101;
  assign n12211 = n12210 ^ x102;
  assign n12212 = n11815 & n11937;
  assign n12213 = n12212 ^ n11817;
  assign n12214 = n12213 ^ n12210;
  assign n12215 = n12211 & ~n12214;
  assign n12216 = n12215 ^ x102;
  assign n12217 = n12216 ^ x103;
  assign n12218 = n11821 & n11937;
  assign n12219 = n12218 ^ n11823;
  assign n12220 = n12219 ^ n12216;
  assign n12221 = n12217 & ~n12220;
  assign n12222 = n12221 ^ x103;
  assign n12223 = n12222 ^ x104;
  assign n12224 = n11827 & n11937;
  assign n12225 = n12224 ^ n11829;
  assign n12226 = n12225 ^ n12222;
  assign n12227 = n12223 & ~n12226;
  assign n12228 = n12227 ^ x104;
  assign n12229 = n12228 ^ x105;
  assign n12230 = n11833 & n11937;
  assign n12231 = n12230 ^ n11835;
  assign n12232 = n12231 ^ n12228;
  assign n12233 = n12229 & ~n12232;
  assign n12234 = n12233 ^ x105;
  assign n12235 = n12234 ^ x106;
  assign n12236 = n11839 & n11937;
  assign n12237 = n12236 ^ n11841;
  assign n12238 = n12237 ^ n12234;
  assign n12239 = n12235 & ~n12238;
  assign n12240 = n12239 ^ x106;
  assign n12241 = n11955 & n12240;
  assign n12242 = n11953 ^ x108;
  assign n12243 = x107 & n11950;
  assign n12244 = n12243 ^ n11953;
  assign n12245 = n12242 & ~n12244;
  assign n12246 = n12245 ^ x108;
  assign n12247 = ~n12241 & ~n12246;
  assign n12248 = n12247 ^ x109;
  assign n12249 = n11856 ^ x108;
  assign n12250 = n11937 & n12249;
  assign n12251 = n12250 ^ n11558;
  assign n12252 = n12251 ^ n12247;
  assign n12253 = ~n12248 & n12252;
  assign n12254 = n12253 ^ x109;
  assign n12255 = n12254 ^ x110;
  assign n12256 = n11856 ^ n11558;
  assign n12257 = n12249 & ~n12256;
  assign n12258 = n12257 ^ x108;
  assign n12259 = n12258 ^ x109;
  assign n12260 = n11937 & n12259;
  assign n12261 = n12260 ^ n11565;
  assign n12262 = n12261 ^ n12254;
  assign n12263 = n12255 & ~n12262;
  assign n12264 = n12263 ^ x110;
  assign n12265 = n12264 ^ x111;
  assign n12266 = ~n11864 & n11937;
  assign n12267 = n12266 ^ n11866;
  assign n12268 = n12267 ^ n12264;
  assign n12269 = n12265 & ~n12268;
  assign n12270 = n12269 ^ x111;
  assign n12271 = n12270 ^ x112;
  assign n12272 = n11870 & n11937;
  assign n12273 = n12272 ^ n11872;
  assign n12274 = n12273 ^ n12270;
  assign n12275 = n12271 & ~n12274;
  assign n12276 = n12275 ^ x112;
  assign n12277 = n12276 ^ x113;
  assign n12278 = n11937 & n11941;
  assign n12279 = n12278 ^ n11553;
  assign n12280 = n12279 ^ n12276;
  assign n12281 = n12277 & ~n12280;
  assign n12282 = n12281 ^ x113;
  assign n12283 = ~n11948 & n12282;
  assign n12284 = ~n11883 & n11937;
  assign n12285 = n12284 ^ n11885;
  assign n12286 = x115 & n12285;
  assign n12287 = x114 & n11947;
  assign n12288 = ~n12286 & ~n12287;
  assign n12289 = ~n12283 & n12288;
  assign n12290 = ~x115 & ~n12285;
  assign n12291 = ~n12289 & ~n12290;
  assign n12292 = n12291 ^ x116;
  assign n12293 = n11889 & n11937;
  assign n12294 = n12293 ^ n11891;
  assign n12295 = n12294 ^ n12291;
  assign n12296 = n12292 & ~n12295;
  assign n12297 = n12296 ^ x116;
  assign n12298 = n12297 ^ x117;
  assign n12299 = n11895 & n11937;
  assign n12300 = n12299 ^ n11897;
  assign n12301 = n12300 ^ n12297;
  assign n12302 = n12298 & ~n12301;
  assign n12303 = n12302 ^ x117;
  assign n12304 = ~n11940 & n12303;
  assign n12305 = n11911 & n11937;
  assign n12306 = n12305 ^ n11913;
  assign n12307 = x119 & n12306;
  assign n12308 = x118 & n11939;
  assign n12309 = ~n12307 & ~n12308;
  assign n12310 = ~n12304 & n12309;
  assign n12311 = ~x119 & ~n12306;
  assign n12312 = n11917 & n11937;
  assign n12313 = n12312 ^ n11920;
  assign n12314 = ~x120 & ~n12313;
  assign n12315 = ~n12311 & ~n12314;
  assign n12316 = ~n12310 & n12315;
  assign n12317 = x120 & n12313;
  assign n12318 = ~n12316 & ~n12317;
  assign n12319 = n12318 ^ x121;
  assign n12320 = n11924 & n11937;
  assign n12321 = n12320 ^ n11930;
  assign n12322 = n12321 ^ n12318;
  assign n12323 = ~n12319 & ~n12322;
  assign n12324 = n12323 ^ x121;
  assign n12325 = n133 & ~n12324;
  assign n12326 = n11905 & ~n11933;
  assign n12327 = ~n134 & n11904;
  assign n12328 = ~n12326 & ~n12327;
  assign n12329 = ~n12325 & ~n12328;
  assign n12330 = x127 & ~n12329;
  assign n12331 = x122 & ~n11543;
  assign n12332 = n132 & ~n12331;
  assign n12333 = ~n12324 & n12332;
  assign n12334 = n11933 ^ x121;
  assign n12335 = n11904 & ~n12334;
  assign n12336 = n134 & n12335;
  assign n12337 = ~n12333 & ~n12336;
  assign n12338 = n12240 ^ x107;
  assign n12339 = n12240 ^ n11950;
  assign n12340 = n12338 & ~n12339;
  assign n12341 = n12340 ^ x107;
  assign n12342 = n12341 ^ x108;
  assign n12343 = ~n12337 & n12342;
  assign n12344 = n12343 ^ n11953;
  assign n12345 = ~x109 & ~n12344;
  assign n12346 = ~n12337 & n12338;
  assign n12347 = n12346 ^ n11950;
  assign n12348 = ~x108 & ~n12347;
  assign n12349 = ~n12345 & ~n12348;
  assign n12350 = n12190 & ~n12337;
  assign n12351 = n12350 ^ n12192;
  assign n12352 = ~x100 & ~n12351;
  assign n12353 = n12140 & ~n12337;
  assign n12354 = n12353 ^ n12144;
  assign n12355 = ~x92 & ~n12354;
  assign n12356 = n12133 & ~n12337;
  assign n12357 = n12356 ^ n12136;
  assign n12358 = ~x91 & ~n12357;
  assign n12359 = ~n12355 & ~n12358;
  assign n12360 = n12070 & ~n12337;
  assign n12361 = n12360 ^ n12072;
  assign n12362 = x80 & n12361;
  assign n12363 = n12026 & ~n12337;
  assign n12364 = n12363 ^ n12028;
  assign n12365 = ~x73 & n12364;
  assign n12366 = x65 & ~n11937;
  assign n12367 = ~n12337 & n12366;
  assign n12368 = n219 & n11937;
  assign n12369 = ~n12367 & ~n12368;
  assign n12370 = x5 & ~n12369;
  assign n12376 = x64 & n11937;
  assign n12371 = n11937 ^ x65;
  assign n12372 = n341 & ~n12371;
  assign n12373 = x5 & n12372;
  assign n12374 = n12373 ^ n340;
  assign n12375 = ~n12337 & n12374;
  assign n12377 = n12376 ^ n12375;
  assign n12378 = ~n12370 & ~n12377;
  assign n12379 = n12378 ^ x6;
  assign n12380 = n12379 ^ x66;
  assign n12384 = x4 & ~x65;
  assign n12385 = x5 & x64;
  assign n12386 = ~n12384 & n12385;
  assign n12381 = ~x4 & n11979;
  assign n12382 = ~x5 & x65;
  assign n12383 = ~n12381 & ~n12382;
  assign n12387 = n12386 ^ n12383;
  assign n12388 = n12337 & ~n12387;
  assign n12389 = n12388 ^ n12386;
  assign n12390 = ~x4 & x65;
  assign n12391 = n12390 ^ n12382;
  assign n12392 = x64 & n12391;
  assign n12393 = n12392 ^ n12382;
  assign n12394 = ~n12389 & ~n12393;
  assign n12395 = n12394 ^ n12379;
  assign n12396 = n12380 & n12395;
  assign n12397 = n12396 ^ x66;
  assign n12398 = n12397 ^ x67;
  assign n12399 = n11991 ^ x66;
  assign n12400 = ~n12337 & ~n12399;
  assign n12401 = n12400 ^ n11977;
  assign n12402 = n12401 ^ n12397;
  assign n12403 = n12398 & ~n12402;
  assign n12404 = n12403 ^ x67;
  assign n12405 = n12404 ^ x68;
  assign n12406 = n11995 & ~n12337;
  assign n12407 = n12406 ^ n11998;
  assign n12408 = n12407 ^ n12404;
  assign n12409 = n12405 & ~n12408;
  assign n12410 = n12409 ^ x68;
  assign n12411 = n12410 ^ x69;
  assign n12412 = n12002 & ~n12337;
  assign n12413 = n12412 ^ n12004;
  assign n12414 = n12413 ^ n12410;
  assign n12415 = n12411 & ~n12414;
  assign n12416 = n12415 ^ x69;
  assign n12417 = n12416 ^ x70;
  assign n12418 = n12008 & ~n12337;
  assign n12419 = n12418 ^ n12010;
  assign n12420 = n12419 ^ n12416;
  assign n12421 = n12417 & ~n12420;
  assign n12422 = n12421 ^ x70;
  assign n12423 = n12422 ^ x71;
  assign n12424 = n12014 & ~n12337;
  assign n12425 = n12424 ^ n12016;
  assign n12426 = n12425 ^ n12422;
  assign n12427 = n12423 & n12426;
  assign n12428 = n12427 ^ x71;
  assign n12429 = n12428 ^ x72;
  assign n12430 = n12020 & ~n12337;
  assign n12431 = n12430 ^ n12022;
  assign n12432 = n12431 ^ n12428;
  assign n12433 = n12429 & ~n12432;
  assign n12434 = n12433 ^ x72;
  assign n12435 = ~n12365 & n12434;
  assign n12436 = x73 & ~n12364;
  assign n12437 = n12032 & ~n12337;
  assign n12438 = n12437 ^ n12034;
  assign n12439 = x74 & n12438;
  assign n12440 = ~n12436 & ~n12439;
  assign n12441 = ~n12435 & n12440;
  assign n12442 = ~x74 & ~n12438;
  assign n12443 = ~n12441 & ~n12442;
  assign n12444 = n12443 ^ x75;
  assign n12445 = n12038 & ~n12337;
  assign n12446 = n12445 ^ n12040;
  assign n12447 = n12446 ^ n12443;
  assign n12448 = n12444 & n12447;
  assign n12449 = n12448 ^ x75;
  assign n12450 = n12449 ^ x76;
  assign n12451 = n12044 & ~n12337;
  assign n12452 = n12451 ^ n12046;
  assign n12453 = n12452 ^ n12449;
  assign n12454 = n12450 & n12453;
  assign n12455 = n12454 ^ x76;
  assign n12456 = n12455 ^ x77;
  assign n12457 = n12049 ^ x76;
  assign n12458 = ~n12337 & n12457;
  assign n12459 = n12458 ^ n11963;
  assign n12460 = n12459 ^ n12455;
  assign n12461 = n12456 & ~n12460;
  assign n12462 = n12461 ^ x77;
  assign n12463 = n12462 ^ x78;
  assign n12464 = ~n12050 & ~n12055;
  assign n12465 = n12464 ^ x77;
  assign n12466 = ~n12337 & ~n12465;
  assign n12467 = n12466 ^ n12053;
  assign n12468 = n12467 ^ n12462;
  assign n12469 = n12463 & n12468;
  assign n12470 = n12469 ^ x78;
  assign n12471 = n12470 ^ x79;
  assign n12472 = n12060 & ~n12337;
  assign n12473 = n12472 ^ n12066;
  assign n12474 = n12473 ^ n12470;
  assign n12475 = n12471 & ~n12474;
  assign n12476 = n12475 ^ x79;
  assign n12477 = ~n12362 & ~n12476;
  assign n12478 = n12076 & ~n12337;
  assign n12479 = n12478 ^ n12078;
  assign n12480 = ~x81 & n12479;
  assign n12481 = ~x80 & ~n12361;
  assign n12482 = ~n12480 & ~n12481;
  assign n12483 = ~n12477 & n12482;
  assign n12484 = x81 & ~n12479;
  assign n12485 = ~n12483 & ~n12484;
  assign n12486 = n12082 & ~n12337;
  assign n12487 = n12486 ^ n12084;
  assign n12488 = ~x82 & ~n12487;
  assign n12489 = n12088 & ~n12337;
  assign n12490 = n12489 ^ n12090;
  assign n12491 = ~x83 & n12490;
  assign n12492 = ~n12488 & ~n12491;
  assign n12493 = ~n12485 & n12492;
  assign n12494 = n12490 ^ x83;
  assign n12495 = x82 & n12487;
  assign n12496 = n12495 ^ n12490;
  assign n12497 = ~n12494 & n12496;
  assign n12498 = n12497 ^ x83;
  assign n12499 = ~n12493 & ~n12498;
  assign n12500 = n12094 & ~n12337;
  assign n12501 = n12500 ^ n12096;
  assign n12502 = ~x84 & ~n12501;
  assign n12503 = n12100 & ~n12337;
  assign n12504 = n12503 ^ n12102;
  assign n12505 = ~x85 & n12504;
  assign n12506 = ~n12502 & ~n12505;
  assign n12507 = ~n12499 & n12506;
  assign n12508 = n12504 ^ x85;
  assign n12509 = x84 & n12501;
  assign n12510 = n12509 ^ n12504;
  assign n12511 = ~n12508 & n12510;
  assign n12512 = n12511 ^ x85;
  assign n12513 = ~n12507 & ~n12512;
  assign n12514 = n12513 ^ x86;
  assign n12515 = n12106 & ~n12337;
  assign n12516 = n12515 ^ n12108;
  assign n12517 = n12516 ^ n12513;
  assign n12518 = ~n12514 & n12517;
  assign n12519 = n12518 ^ x86;
  assign n12520 = n12519 ^ x87;
  assign n12521 = n12112 & ~n12337;
  assign n12522 = n12521 ^ n12114;
  assign n12523 = n12522 ^ n12519;
  assign n12524 = n12520 & ~n12523;
  assign n12525 = n12524 ^ x87;
  assign n12526 = n12525 ^ x88;
  assign n12527 = n12117 ^ x87;
  assign n12528 = ~n12337 & n12527;
  assign n12529 = n12528 ^ n11960;
  assign n12530 = n12529 ^ n12525;
  assign n12531 = n12526 & ~n12530;
  assign n12532 = n12531 ^ x88;
  assign n12533 = n12532 ^ x89;
  assign n12534 = ~n12118 & ~n12122;
  assign n12535 = n12534 ^ x88;
  assign n12536 = ~n12337 & ~n12535;
  assign n12537 = n12536 ^ n12120;
  assign n12538 = n12537 ^ n12532;
  assign n12539 = n12533 & ~n12538;
  assign n12540 = n12539 ^ x89;
  assign n12541 = n12540 ^ x90;
  assign n12542 = n12127 & ~n12337;
  assign n12543 = n12542 ^ n12129;
  assign n12544 = n12543 ^ n12540;
  assign n12545 = n12541 & ~n12544;
  assign n12546 = n12545 ^ x90;
  assign n12547 = n12359 & n12546;
  assign n12548 = n12354 ^ x92;
  assign n12549 = x91 & n12357;
  assign n12550 = n12549 ^ n12354;
  assign n12551 = n12548 & ~n12550;
  assign n12552 = n12551 ^ x92;
  assign n12553 = ~n12547 & ~n12552;
  assign n12554 = n12553 ^ x93;
  assign n12555 = n12148 & ~n12337;
  assign n12556 = n12555 ^ n12150;
  assign n12557 = n12556 ^ n12553;
  assign n12558 = ~n12554 & n12557;
  assign n12559 = n12558 ^ x93;
  assign n12560 = n12559 ^ x94;
  assign n12561 = n12153 ^ x93;
  assign n12562 = ~n12337 & n12561;
  assign n12563 = n12562 ^ n11957;
  assign n12564 = n12563 ^ n12559;
  assign n12565 = n12560 & ~n12564;
  assign n12566 = n12565 ^ x94;
  assign n12567 = n12566 ^ x95;
  assign n12568 = ~n12154 & ~n12158;
  assign n12569 = n12568 ^ x94;
  assign n12570 = ~n12337 & ~n12569;
  assign n12571 = n12570 ^ n12156;
  assign n12572 = n12571 ^ n12566;
  assign n12573 = n12567 & ~n12572;
  assign n12574 = n12573 ^ x95;
  assign n12575 = n12574 ^ x96;
  assign n12576 = n12163 & ~n12337;
  assign n12577 = n12576 ^ n12165;
  assign n12578 = n12577 ^ n12574;
  assign n12579 = n12575 & ~n12578;
  assign n12580 = n12579 ^ x96;
  assign n12581 = n12580 ^ x97;
  assign n12582 = n12169 & ~n12337;
  assign n12583 = n12582 ^ n12172;
  assign n12584 = n12583 ^ n12580;
  assign n12585 = n12581 & ~n12584;
  assign n12586 = n12585 ^ x97;
  assign n12587 = n12586 ^ x98;
  assign n12588 = n12176 & ~n12337;
  assign n12589 = n12588 ^ n12180;
  assign n12590 = n12589 ^ n12586;
  assign n12591 = n12587 & ~n12590;
  assign n12592 = n12591 ^ x98;
  assign n12593 = n12592 ^ x99;
  assign n12594 = n12184 & ~n12337;
  assign n12595 = n12594 ^ n12186;
  assign n12596 = n12595 ^ n12592;
  assign n12597 = n12593 & ~n12596;
  assign n12598 = n12597 ^ x99;
  assign n12599 = ~n12352 & n12598;
  assign n12600 = n12196 & ~n12337;
  assign n12601 = n12600 ^ n12199;
  assign n12602 = x101 & n12601;
  assign n12603 = x100 & n12351;
  assign n12604 = ~n12602 & ~n12603;
  assign n12605 = ~n12599 & n12604;
  assign n12606 = ~x101 & ~n12601;
  assign n12607 = ~n12605 & ~n12606;
  assign n12608 = n12607 ^ x102;
  assign n12609 = n12203 & ~n12337;
  assign n12610 = n12609 ^ n12207;
  assign n12611 = n12610 ^ n12607;
  assign n12612 = n12608 & ~n12611;
  assign n12613 = n12612 ^ x102;
  assign n12614 = n12613 ^ x103;
  assign n12615 = n12211 & ~n12337;
  assign n12616 = n12615 ^ n12213;
  assign n12617 = n12616 ^ n12613;
  assign n12618 = n12614 & ~n12617;
  assign n12619 = n12618 ^ x103;
  assign n12620 = n12619 ^ x104;
  assign n12621 = n12217 & ~n12337;
  assign n12622 = n12621 ^ n12219;
  assign n12623 = n12622 ^ n12619;
  assign n12624 = n12620 & ~n12623;
  assign n12625 = n12624 ^ x104;
  assign n12626 = n12625 ^ x105;
  assign n12627 = n12223 & ~n12337;
  assign n12628 = n12627 ^ n12225;
  assign n12629 = n12628 ^ n12625;
  assign n12630 = n12626 & ~n12629;
  assign n12631 = n12630 ^ x105;
  assign n12632 = n12631 ^ x106;
  assign n12633 = n12229 & ~n12337;
  assign n12634 = n12633 ^ n12231;
  assign n12635 = n12634 ^ n12631;
  assign n12636 = n12632 & ~n12635;
  assign n12637 = n12636 ^ x106;
  assign n12638 = n12637 ^ x107;
  assign n12639 = n12235 & ~n12337;
  assign n12640 = n12639 ^ n12237;
  assign n12641 = n12640 ^ n12637;
  assign n12642 = n12638 & ~n12641;
  assign n12643 = n12642 ^ x107;
  assign n12644 = n12349 & n12643;
  assign n12645 = n12344 ^ x109;
  assign n12646 = x108 & n12347;
  assign n12647 = n12646 ^ n12344;
  assign n12648 = n12645 & ~n12647;
  assign n12649 = n12648 ^ x109;
  assign n12650 = ~n12644 & ~n12649;
  assign n12651 = n12650 ^ x110;
  assign n12652 = ~n12248 & ~n12337;
  assign n12653 = n12652 ^ n12251;
  assign n12654 = n12653 ^ n12650;
  assign n12655 = ~n12651 & n12654;
  assign n12656 = n12655 ^ x110;
  assign n12657 = n12656 ^ x111;
  assign n12658 = ~n12319 & ~n12337;
  assign n12659 = n12658 ^ n12321;
  assign n12660 = n12659 ^ x122;
  assign n12661 = n12277 & ~n12337;
  assign n12662 = n12661 ^ n12279;
  assign n12663 = x114 & n12662;
  assign n12664 = n12255 & ~n12337;
  assign n12665 = n12664 ^ n12261;
  assign n12666 = n12665 ^ n12656;
  assign n12667 = n12657 & ~n12666;
  assign n12668 = n12667 ^ x111;
  assign n12669 = n12668 ^ x112;
  assign n12670 = n12265 & ~n12337;
  assign n12671 = n12670 ^ n12267;
  assign n12672 = n12671 ^ n12668;
  assign n12673 = n12669 & ~n12672;
  assign n12674 = n12673 ^ x112;
  assign n12675 = n12674 ^ x113;
  assign n12676 = n12271 & ~n12337;
  assign n12677 = n12676 ^ n12273;
  assign n12678 = n12677 ^ n12674;
  assign n12679 = n12675 & ~n12678;
  assign n12680 = n12679 ^ x113;
  assign n12681 = ~n12663 & ~n12680;
  assign n12682 = ~x114 & ~n12662;
  assign n12683 = n12282 ^ x114;
  assign n12684 = ~n12337 & n12683;
  assign n12685 = n12684 ^ n11947;
  assign n12686 = ~n12682 & n12685;
  assign n12687 = ~n12681 & n12686;
  assign n12688 = ~x115 & ~n12687;
  assign n12689 = ~n12681 & ~n12682;
  assign n12690 = ~n12685 & ~n12689;
  assign n12691 = ~n12688 & ~n12690;
  assign n12692 = n12691 ^ x116;
  assign n12693 = ~n12283 & ~n12287;
  assign n12694 = n12693 ^ x115;
  assign n12695 = ~n12337 & ~n12694;
  assign n12696 = n12695 ^ n12285;
  assign n12697 = n12696 ^ n12691;
  assign n12698 = n12692 & ~n12697;
  assign n12699 = n12698 ^ x116;
  assign n12700 = n12699 ^ x117;
  assign n12701 = n12292 & ~n12337;
  assign n12702 = n12701 ^ n12294;
  assign n12703 = n12702 ^ n12699;
  assign n12704 = n12700 & ~n12703;
  assign n12705 = n12704 ^ x117;
  assign n12706 = n12705 ^ x118;
  assign n12707 = n12298 & ~n12337;
  assign n12708 = n12707 ^ n12300;
  assign n12709 = n12708 ^ n12705;
  assign n12710 = n12706 & ~n12709;
  assign n12711 = n12710 ^ x118;
  assign n12712 = n12711 ^ x119;
  assign n12713 = n12303 ^ x118;
  assign n12714 = ~n12337 & n12713;
  assign n12715 = n12714 ^ n11939;
  assign n12716 = n12715 ^ n12711;
  assign n12717 = n12712 & ~n12716;
  assign n12718 = n12717 ^ x119;
  assign n12719 = n12718 ^ x120;
  assign n12720 = ~n12304 & ~n12308;
  assign n12721 = n12720 ^ x119;
  assign n12722 = ~n12337 & ~n12721;
  assign n12723 = n12722 ^ n12306;
  assign n12724 = n12723 ^ n12718;
  assign n12725 = n12719 & ~n12724;
  assign n12726 = n12725 ^ x120;
  assign n12727 = n12726 ^ x121;
  assign n12728 = ~n12310 & ~n12311;
  assign n12729 = n12728 ^ x120;
  assign n12730 = ~n12337 & n12729;
  assign n12731 = n12730 ^ n12313;
  assign n12732 = n12731 ^ n12726;
  assign n12733 = n12727 & ~n12732;
  assign n12734 = n12733 ^ x121;
  assign n12735 = n12734 ^ n12659;
  assign n12736 = ~n12660 & n12735;
  assign n12737 = n12736 ^ x122;
  assign n12738 = n11543 & ~n12737;
  assign n12739 = ~n12329 & n12737;
  assign n12740 = ~x123 & ~n12739;
  assign n12741 = ~n12738 & ~n12740;
  assign n12742 = n131 & ~n12741;
  assign n12743 = n12657 & n12742;
  assign n12744 = n12743 ^ n12665;
  assign n12745 = ~x112 & ~n12744;
  assign n12746 = n12560 & n12742;
  assign n12747 = n12746 ^ n12563;
  assign n12748 = ~x95 & ~n12747;
  assign n12749 = n12567 & n12742;
  assign n12750 = n12749 ^ n12571;
  assign n12751 = ~x96 & ~n12750;
  assign n12752 = ~n12748 & ~n12751;
  assign n12753 = n12520 & n12742;
  assign n12754 = n12753 ^ n12522;
  assign n12755 = ~x88 & ~n12754;
  assign n12756 = n12526 & n12742;
  assign n12757 = n12756 ^ n12529;
  assign n12758 = ~x89 & ~n12757;
  assign n12759 = ~n12755 & ~n12758;
  assign n12760 = n12434 ^ x73;
  assign n12761 = n12742 & n12760;
  assign n12762 = n12761 ^ n12364;
  assign n12763 = ~x74 & n12762;
  assign n12764 = ~n12435 & ~n12436;
  assign n12765 = n12764 ^ x74;
  assign n12766 = n12742 & ~n12765;
  assign n12767 = n12766 ^ n12438;
  assign n12768 = ~x75 & ~n12767;
  assign n12769 = ~n12763 & ~n12768;
  assign n12770 = x64 & n12742;
  assign n12771 = x4 & n12770;
  assign n12772 = x3 & ~x65;
  assign n12773 = n12771 & ~n12772;
  assign n12774 = ~x3 & x64;
  assign n12775 = ~x65 & ~n12774;
  assign n12776 = ~x4 & ~n12775;
  assign n12777 = ~n12742 & n12776;
  assign n12778 = ~x3 & x65;
  assign n12779 = x64 & n12778;
  assign n12780 = ~x64 & n12390;
  assign n12781 = ~n12779 & ~n12780;
  assign n12782 = ~n12777 & n12781;
  assign n12783 = ~n12773 & n12782;
  assign n12784 = n12783 ^ x66;
  assign n12785 = x65 & n131;
  assign n12786 = n12337 & n12785;
  assign n12787 = ~n12741 & n12786;
  assign n12788 = n219 & ~n12337;
  assign n12789 = ~n12787 & ~n12788;
  assign n12790 = x4 & ~n12789;
  assign n12791 = ~x4 & n219;
  assign n12792 = n12337 & n12791;
  assign n12793 = ~n202 & ~n12792;
  assign n12794 = n12742 & ~n12793;
  assign n12795 = ~n12390 & ~n12741;
  assign n12796 = x64 & ~n12337;
  assign n12797 = ~n12795 & n12796;
  assign n12798 = ~n12794 & ~n12797;
  assign n12799 = ~n12790 & n12798;
  assign n12800 = n12799 ^ x5;
  assign n12801 = n12800 ^ n12783;
  assign n12802 = ~n12784 & n12801;
  assign n12803 = n12802 ^ x66;
  assign n12804 = ~x67 & ~n12803;
  assign n12805 = ~x66 & ~n12800;
  assign n12806 = x67 & ~n12783;
  assign n12807 = ~n12805 & n12806;
  assign n12808 = n1724 & n12800;
  assign n12809 = n12394 ^ x66;
  assign n12810 = n12742 & ~n12809;
  assign n12811 = n12810 ^ n12379;
  assign n12812 = ~n12808 & ~n12811;
  assign n12813 = ~n12807 & n12812;
  assign n12814 = ~n12804 & ~n12813;
  assign n12815 = n12814 ^ x68;
  assign n12816 = n12398 & n12742;
  assign n12817 = n12816 ^ n12401;
  assign n12818 = n12817 ^ n12814;
  assign n12819 = n12815 & ~n12818;
  assign n12820 = n12819 ^ x68;
  assign n12821 = n12820 ^ x69;
  assign n12822 = n12405 & n12742;
  assign n12823 = n12822 ^ n12407;
  assign n12824 = n12823 ^ n12820;
  assign n12825 = n12821 & ~n12824;
  assign n12826 = n12825 ^ x69;
  assign n12827 = n12826 ^ x70;
  assign n12828 = n12411 & n12742;
  assign n12829 = n12828 ^ n12413;
  assign n12830 = n12829 ^ n12826;
  assign n12831 = n12827 & ~n12830;
  assign n12832 = n12831 ^ x70;
  assign n12833 = n12832 ^ x71;
  assign n12834 = n12417 & n12742;
  assign n12835 = n12834 ^ n12419;
  assign n12836 = n12835 ^ n12832;
  assign n12837 = n12833 & ~n12836;
  assign n12838 = n12837 ^ x71;
  assign n12839 = n12838 ^ x72;
  assign n12840 = n12423 & n12742;
  assign n12841 = n12840 ^ n12425;
  assign n12842 = n12841 ^ n12838;
  assign n12843 = n12839 & n12842;
  assign n12844 = n12843 ^ x72;
  assign n12845 = n12844 ^ x73;
  assign n12846 = n12429 & n12742;
  assign n12847 = n12846 ^ n12431;
  assign n12848 = n12847 ^ n12844;
  assign n12849 = n12845 & ~n12848;
  assign n12850 = n12849 ^ x73;
  assign n12851 = n12769 & n12850;
  assign n12852 = n12767 ^ x75;
  assign n12853 = x74 & ~n12762;
  assign n12854 = n12853 ^ n12767;
  assign n12855 = n12852 & ~n12854;
  assign n12856 = n12855 ^ x75;
  assign n12857 = ~n12851 & ~n12856;
  assign n12858 = n12857 ^ x76;
  assign n12859 = n12444 & n12742;
  assign n12860 = n12859 ^ n12446;
  assign n12861 = n12860 ^ n12857;
  assign n12862 = ~n12858 & ~n12861;
  assign n12863 = n12862 ^ x76;
  assign n12864 = n12863 ^ x77;
  assign n12865 = n12450 & n12742;
  assign n12866 = n12865 ^ n12452;
  assign n12867 = n12866 ^ n12863;
  assign n12868 = n12864 & n12867;
  assign n12869 = n12868 ^ x77;
  assign n12870 = n12869 ^ x78;
  assign n12871 = n12456 & n12742;
  assign n12872 = n12871 ^ n12459;
  assign n12873 = n12872 ^ n12869;
  assign n12874 = n12870 & ~n12873;
  assign n12875 = n12874 ^ x78;
  assign n12876 = n12875 ^ x79;
  assign n12877 = n12463 & n12742;
  assign n12878 = n12877 ^ n12467;
  assign n12879 = n12878 ^ n12875;
  assign n12880 = n12876 & n12879;
  assign n12881 = n12880 ^ x79;
  assign n12882 = n12881 ^ x80;
  assign n12883 = n12471 & n12742;
  assign n12884 = n12883 ^ n12473;
  assign n12885 = n12884 ^ n12881;
  assign n12886 = n12882 & ~n12885;
  assign n12887 = n12886 ^ x80;
  assign n12888 = n12887 ^ x81;
  assign n12889 = n12476 ^ x80;
  assign n12890 = n12742 & n12889;
  assign n12891 = n12890 ^ n12361;
  assign n12892 = n12891 ^ n12887;
  assign n12893 = n12888 & ~n12892;
  assign n12894 = n12893 ^ x81;
  assign n12895 = n12894 ^ x82;
  assign n12896 = ~n12477 & ~n12481;
  assign n12897 = n12896 ^ x81;
  assign n12898 = n12742 & n12897;
  assign n12899 = n12898 ^ n12479;
  assign n12900 = n12899 ^ n12894;
  assign n12901 = n12895 & n12900;
  assign n12902 = n12901 ^ x82;
  assign n12903 = n12902 ^ x83;
  assign n12904 = n12485 ^ x82;
  assign n12905 = n12742 & ~n12904;
  assign n12906 = n12905 ^ n12487;
  assign n12907 = n12906 ^ n12902;
  assign n12908 = n12903 & ~n12907;
  assign n12909 = n12908 ^ x83;
  assign n12910 = n12909 ^ x84;
  assign n12911 = n12487 ^ n12485;
  assign n12912 = ~n12904 & n12911;
  assign n12913 = n12912 ^ x82;
  assign n12914 = n12913 ^ x83;
  assign n12915 = n12742 & n12914;
  assign n12916 = n12915 ^ n12490;
  assign n12917 = n12916 ^ n12909;
  assign n12918 = n12910 & n12917;
  assign n12919 = n12918 ^ x84;
  assign n12920 = n12919 ^ x85;
  assign n12921 = n12499 ^ x84;
  assign n12922 = n12742 & ~n12921;
  assign n12923 = n12922 ^ n12501;
  assign n12924 = n12923 ^ n12919;
  assign n12925 = n12920 & ~n12924;
  assign n12926 = n12925 ^ x85;
  assign n12927 = n12926 ^ x86;
  assign n12928 = n12501 ^ n12499;
  assign n12929 = ~n12921 & n12928;
  assign n12930 = n12929 ^ x84;
  assign n12931 = n12930 ^ x85;
  assign n12932 = n12742 & n12931;
  assign n12933 = n12932 ^ n12504;
  assign n12934 = n12933 ^ n12926;
  assign n12935 = n12927 & n12934;
  assign n12936 = n12935 ^ x86;
  assign n12937 = n12936 ^ x87;
  assign n12938 = ~n12514 & n12742;
  assign n12939 = n12938 ^ n12516;
  assign n12940 = n12939 ^ n12936;
  assign n12941 = n12937 & ~n12940;
  assign n12942 = n12941 ^ x87;
  assign n12943 = n12759 & n12942;
  assign n12944 = n12757 ^ x89;
  assign n12945 = x88 & n12754;
  assign n12946 = n12945 ^ n12757;
  assign n12947 = n12944 & ~n12946;
  assign n12948 = n12947 ^ x89;
  assign n12949 = ~n12943 & ~n12948;
  assign n12950 = n12949 ^ x90;
  assign n12951 = n12533 & n12742;
  assign n12952 = n12951 ^ n12537;
  assign n12953 = n12952 ^ n12949;
  assign n12954 = ~n12950 & n12953;
  assign n12955 = n12954 ^ x90;
  assign n12956 = n12955 ^ x91;
  assign n12957 = n12541 & n12742;
  assign n12958 = n12957 ^ n12543;
  assign n12959 = n12958 ^ n12955;
  assign n12960 = n12956 & ~n12959;
  assign n12961 = n12960 ^ x91;
  assign n12962 = n12961 ^ x92;
  assign n12963 = n12546 ^ x91;
  assign n12964 = n12742 & n12963;
  assign n12965 = n12964 ^ n12357;
  assign n12966 = n12965 ^ n12961;
  assign n12967 = n12962 & ~n12966;
  assign n12968 = n12967 ^ x92;
  assign n12969 = n12968 ^ x93;
  assign n12970 = n12546 ^ n12357;
  assign n12971 = n12963 & ~n12970;
  assign n12972 = n12971 ^ x91;
  assign n12973 = n12972 ^ x92;
  assign n12974 = n12742 & n12973;
  assign n12975 = n12974 ^ n12354;
  assign n12976 = n12975 ^ n12968;
  assign n12977 = n12969 & ~n12976;
  assign n12978 = n12977 ^ x93;
  assign n12979 = n12978 ^ x94;
  assign n12980 = ~n12554 & n12742;
  assign n12981 = n12980 ^ n12556;
  assign n12982 = n12981 ^ n12978;
  assign n12983 = n12979 & ~n12982;
  assign n12984 = n12983 ^ x94;
  assign n12985 = n12752 & n12984;
  assign n12986 = n12750 ^ x96;
  assign n12987 = x95 & n12747;
  assign n12988 = n12987 ^ n12750;
  assign n12989 = n12986 & ~n12988;
  assign n12990 = n12989 ^ x96;
  assign n12991 = ~n12985 & ~n12990;
  assign n12992 = n12991 ^ x97;
  assign n12993 = n12575 & n12742;
  assign n12994 = n12993 ^ n12577;
  assign n12995 = n12994 ^ n12991;
  assign n12996 = ~n12992 & n12995;
  assign n12997 = n12996 ^ x97;
  assign n12998 = n12997 ^ x98;
  assign n12999 = n12581 & n12742;
  assign n13000 = n12999 ^ n12583;
  assign n13001 = n13000 ^ n12997;
  assign n13002 = n12998 & ~n13001;
  assign n13003 = n13002 ^ x98;
  assign n13004 = n13003 ^ x99;
  assign n13005 = n12587 & n12742;
  assign n13006 = n13005 ^ n12589;
  assign n13007 = n13006 ^ n13003;
  assign n13008 = n13004 & ~n13007;
  assign n13009 = n13008 ^ x99;
  assign n13010 = n13009 ^ x100;
  assign n13011 = n12593 & n12742;
  assign n13012 = n13011 ^ n12595;
  assign n13013 = n13012 ^ n13009;
  assign n13014 = n13010 & ~n13013;
  assign n13015 = n13014 ^ x100;
  assign n13016 = n13015 ^ x101;
  assign n13017 = n12598 ^ x100;
  assign n13018 = n12742 & n13017;
  assign n13019 = n13018 ^ n12351;
  assign n13020 = n13019 ^ n13015;
  assign n13021 = n13016 & ~n13020;
  assign n13022 = n13021 ^ x101;
  assign n13023 = n13022 ^ x102;
  assign n13024 = ~n12599 & ~n12603;
  assign n13025 = n13024 ^ x101;
  assign n13026 = n12742 & ~n13025;
  assign n13027 = n13026 ^ n12601;
  assign n13028 = n13027 ^ n13022;
  assign n13029 = n13023 & ~n13028;
  assign n13030 = n13029 ^ x102;
  assign n13031 = n13030 ^ x103;
  assign n13032 = n12608 & n12742;
  assign n13033 = n13032 ^ n12610;
  assign n13034 = n13033 ^ n13030;
  assign n13035 = n13031 & ~n13034;
  assign n13036 = n13035 ^ x103;
  assign n13037 = n13036 ^ x104;
  assign n13038 = n12614 & n12742;
  assign n13039 = n13038 ^ n12616;
  assign n13040 = n13039 ^ n13036;
  assign n13041 = n13037 & ~n13040;
  assign n13042 = n13041 ^ x104;
  assign n13043 = n13042 ^ x105;
  assign n13044 = n12620 & n12742;
  assign n13045 = n13044 ^ n12622;
  assign n13046 = n13045 ^ n13042;
  assign n13047 = n13043 & ~n13046;
  assign n13048 = n13047 ^ x105;
  assign n13049 = n13048 ^ x106;
  assign n13050 = n12626 & n12742;
  assign n13051 = n13050 ^ n12628;
  assign n13052 = n13051 ^ n13048;
  assign n13053 = n13049 & ~n13052;
  assign n13054 = n13053 ^ x106;
  assign n13055 = n13054 ^ x107;
  assign n13056 = n12632 & n12742;
  assign n13057 = n13056 ^ n12634;
  assign n13058 = n13057 ^ n13054;
  assign n13059 = n13055 & ~n13058;
  assign n13060 = n13059 ^ x107;
  assign n13061 = n13060 ^ x108;
  assign n13062 = n12638 & n12742;
  assign n13063 = n13062 ^ n12640;
  assign n13064 = n13063 ^ n13060;
  assign n13065 = n13061 & ~n13064;
  assign n13066 = n13065 ^ x108;
  assign n13067 = n13066 ^ x109;
  assign n13068 = n12643 ^ x108;
  assign n13069 = n12742 & n13068;
  assign n13070 = n13069 ^ n12347;
  assign n13071 = n13070 ^ n13066;
  assign n13072 = n13067 & ~n13071;
  assign n13073 = n13072 ^ x109;
  assign n13074 = n13073 ^ x110;
  assign n13075 = n12643 ^ n12347;
  assign n13076 = n13068 & ~n13075;
  assign n13077 = n13076 ^ x108;
  assign n13078 = n13077 ^ x109;
  assign n13079 = n12742 & n13078;
  assign n13080 = n13079 ^ n12344;
  assign n13081 = n13080 ^ n13073;
  assign n13082 = n13074 & ~n13081;
  assign n13083 = n13082 ^ x110;
  assign n13084 = n13083 ^ x111;
  assign n13085 = ~n12651 & n12742;
  assign n13086 = n13085 ^ n12653;
  assign n13087 = n13086 ^ n13083;
  assign n13088 = n13084 & ~n13087;
  assign n13089 = n13088 ^ x111;
  assign n13090 = ~n12745 & n13089;
  assign n13091 = n12669 & n12742;
  assign n13092 = n13091 ^ n12671;
  assign n13093 = x113 & n13092;
  assign n13094 = x112 & n12744;
  assign n13095 = ~n13093 & ~n13094;
  assign n13096 = ~n13090 & n13095;
  assign n13097 = ~x113 & ~n13092;
  assign n13098 = ~n13096 & ~n13097;
  assign n13099 = n13098 ^ x114;
  assign n13100 = n12675 & n12742;
  assign n13101 = n13100 ^ n12677;
  assign n13102 = n13101 ^ n13098;
  assign n13103 = n13099 & ~n13102;
  assign n13104 = n13103 ^ x114;
  assign n13105 = n13104 ^ x115;
  assign n13106 = n12680 ^ x114;
  assign n13107 = n12742 & n13106;
  assign n13108 = n13107 ^ n12662;
  assign n13109 = n13108 ^ n13104;
  assign n13110 = n13105 & ~n13109;
  assign n13111 = n13110 ^ x115;
  assign n13112 = n13111 ^ x116;
  assign n13113 = n12689 ^ x115;
  assign n13114 = n12742 & n13113;
  assign n13115 = n13114 ^ n12685;
  assign n13116 = n13115 ^ n13111;
  assign n13117 = n13112 & ~n13116;
  assign n13118 = n13117 ^ x116;
  assign n13119 = n13118 ^ x117;
  assign n13120 = n12692 & n12742;
  assign n13121 = n13120 ^ n12696;
  assign n13122 = n13121 ^ n13118;
  assign n13123 = n13119 & ~n13122;
  assign n13124 = n13123 ^ x117;
  assign n13125 = n13124 ^ x118;
  assign n13126 = n12700 & n12742;
  assign n13127 = n13126 ^ n12702;
  assign n13128 = n13127 ^ n13124;
  assign n13129 = n13125 & ~n13128;
  assign n13130 = n13129 ^ x118;
  assign n13131 = n13130 ^ x119;
  assign n13132 = n12706 & n12742;
  assign n13133 = n13132 ^ n12708;
  assign n13134 = n13133 ^ n13130;
  assign n13135 = n13131 & ~n13134;
  assign n13136 = n13135 ^ x119;
  assign n13137 = n13136 ^ x120;
  assign n13138 = n12712 & n12742;
  assign n13139 = n13138 ^ n12715;
  assign n13140 = n13139 ^ n13136;
  assign n13141 = n13137 & ~n13140;
  assign n13142 = n13141 ^ x120;
  assign n13143 = n13142 ^ x121;
  assign n13144 = n12719 & n12742;
  assign n13145 = n13144 ^ n12723;
  assign n13146 = n13145 ^ n13142;
  assign n13147 = n13143 & ~n13146;
  assign n13148 = n13147 ^ x121;
  assign n13149 = n13148 ^ x122;
  assign n13150 = n12727 & n12742;
  assign n13151 = n13150 ^ n12731;
  assign n13152 = n13151 ^ n13148;
  assign n13153 = n13149 & ~n13152;
  assign n13154 = n13153 ^ x122;
  assign n13155 = n13154 ^ x123;
  assign n13156 = n12734 ^ x122;
  assign n13157 = n12742 & n13156;
  assign n13158 = n13157 ^ n12659;
  assign n13159 = n13158 ^ n13154;
  assign n13160 = n13155 & n13159;
  assign n13161 = n13160 ^ x123;
  assign n13162 = n12737 ^ x123;
  assign n13163 = n12329 & n13162;
  assign n13164 = n131 & n13163;
  assign n13165 = n13164 ^ n12329;
  assign n13166 = ~x124 & n13165;
  assign n13167 = n13161 & ~n13166;
  assign n13168 = x124 & ~n11904;
  assign n13169 = n130 & ~n13168;
  assign n13170 = ~n13167 & n13169;
  assign n13171 = ~x2 & ~x3;
  assign n13172 = ~n13170 & n13171;
  assign n13173 = ~x2 & x65;
  assign n13174 = ~n13172 & ~n13173;
  assign n13175 = n12770 ^ x4;
  assign n13176 = ~n13174 & ~n13175;
  assign n13177 = x3 & n13170;
  assign n13178 = ~n13176 & ~n13177;
  assign n13179 = n13175 ^ x65;
  assign n13180 = x2 & ~x65;
  assign n13181 = ~n13179 & ~n13180;
  assign n13182 = n13177 & ~n13181;
  assign n13183 = x64 & ~n13182;
  assign n13184 = ~n13178 & n13183;
  assign n13185 = x64 & n13170;
  assign n13186 = n12778 & ~n13185;
  assign n13187 = n13175 ^ n13170;
  assign n13188 = n13186 & ~n13187;
  assign n13189 = ~x66 & ~n13188;
  assign n13190 = ~n13184 & n13189;
  assign n13191 = n12772 & ~n13170;
  assign n13192 = ~x2 & x64;
  assign n13193 = ~n13191 & n13192;
  assign n13194 = ~n12775 & n13170;
  assign n13195 = ~n12778 & n13175;
  assign n13196 = ~n13194 & n13195;
  assign n13197 = ~n13193 & n13196;
  assign n13198 = n12774 & ~n13173;
  assign n13199 = ~n13179 & n13198;
  assign n13200 = x3 & n12780;
  assign n13201 = ~n13199 & ~n13200;
  assign n13202 = n13170 & ~n13201;
  assign n13203 = ~n13197 & ~n13202;
  assign n13204 = ~n13190 & n13203;
  assign n13205 = n13204 ^ x67;
  assign n13206 = ~n12784 & n13170;
  assign n13207 = n13206 ^ n12800;
  assign n13208 = n13207 ^ n13204;
  assign n13209 = n13205 & ~n13208;
  assign n13210 = n13209 ^ x67;
  assign n13211 = n13210 ^ x68;
  assign n13212 = n13161 ^ x124;
  assign n13213 = n13165 & n13212;
  assign n13214 = n130 & n13213;
  assign n13215 = n13214 ^ n13165;
  assign n13216 = ~x125 & n13215;
  assign n13217 = n13099 & n13170;
  assign n13218 = n13217 ^ n13101;
  assign n13219 = ~x115 & ~n13218;
  assign n13220 = n13105 & n13170;
  assign n13221 = n13220 ^ n13108;
  assign n13222 = ~x116 & ~n13221;
  assign n13223 = ~n13219 & ~n13222;
  assign n13224 = n13016 & n13170;
  assign n13225 = n13224 ^ n13019;
  assign n13226 = ~x102 & ~n13225;
  assign n13227 = n13023 & n13170;
  assign n13228 = n13227 ^ n13027;
  assign n13229 = ~x103 & ~n13228;
  assign n13230 = ~n13226 & ~n13229;
  assign n13231 = n12998 & n13170;
  assign n13232 = n13231 ^ n13000;
  assign n13233 = ~x99 & ~n13232;
  assign n13234 = n13004 & n13170;
  assign n13235 = n13234 ^ n13006;
  assign n13236 = ~x100 & ~n13235;
  assign n13237 = ~n13233 & ~n13236;
  assign n13238 = n12962 & n13170;
  assign n13239 = n13238 ^ n12965;
  assign n13240 = x93 & n13239;
  assign n13241 = n12821 & n13170;
  assign n13242 = n13241 ^ n12823;
  assign n13243 = n12803 ^ x67;
  assign n13244 = n13170 & n13243;
  assign n13245 = n13244 ^ n12811;
  assign n13246 = n13245 ^ n13210;
  assign n13247 = n13211 & ~n13246;
  assign n13248 = n13247 ^ x68;
  assign n13249 = n13248 ^ x69;
  assign n13250 = n12815 & n13170;
  assign n13251 = n13250 ^ n12817;
  assign n13252 = n13251 ^ n13248;
  assign n13253 = n13249 & ~n13252;
  assign n13254 = n13253 ^ x69;
  assign n13255 = n13242 & n13254;
  assign n13256 = x70 & n13254;
  assign n13257 = ~n13255 & ~n13256;
  assign n13258 = n12827 & n13170;
  assign n13259 = n13258 ^ n12829;
  assign n13260 = ~n579 & ~n13259;
  assign n13261 = ~n13257 & ~n13260;
  assign n13262 = x71 & n13255;
  assign n13263 = n13259 ^ x71;
  assign n13264 = x70 & n13242;
  assign n13265 = n13264 ^ n13259;
  assign n13266 = n13263 & ~n13265;
  assign n13267 = n13266 ^ x71;
  assign n13268 = ~n13262 & ~n13267;
  assign n13269 = ~n13261 & n13268;
  assign n13270 = n13269 ^ x72;
  assign n13271 = n12833 & n13170;
  assign n13272 = n13271 ^ n12835;
  assign n13273 = n13272 ^ n13269;
  assign n13274 = ~n13270 & n13273;
  assign n13275 = n13274 ^ x72;
  assign n13276 = n13275 ^ x73;
  assign n13277 = n12839 & n13170;
  assign n13278 = n13277 ^ n12841;
  assign n13279 = n13278 ^ n13275;
  assign n13280 = n13276 & n13279;
  assign n13281 = n13280 ^ x73;
  assign n13282 = n13281 ^ x74;
  assign n13283 = n12845 & n13170;
  assign n13284 = n13283 ^ n12847;
  assign n13285 = n13284 ^ n13281;
  assign n13286 = n13282 & ~n13285;
  assign n13287 = n13286 ^ x74;
  assign n13288 = n13287 ^ x75;
  assign n13289 = n12850 ^ x74;
  assign n13290 = n13170 & n13289;
  assign n13291 = n13290 ^ n12762;
  assign n13292 = n13291 ^ n13287;
  assign n13293 = n13288 & n13292;
  assign n13294 = n13293 ^ x75;
  assign n13295 = n13294 ^ x76;
  assign n13296 = n12850 ^ n12762;
  assign n13297 = n13289 & n13296;
  assign n13298 = n13297 ^ x74;
  assign n13299 = n13298 ^ x75;
  assign n13300 = n13170 & n13299;
  assign n13301 = n13300 ^ n12767;
  assign n13302 = n13301 ^ n13294;
  assign n13303 = n13295 & ~n13302;
  assign n13304 = n13303 ^ x76;
  assign n13305 = n13304 ^ x77;
  assign n13306 = ~n12858 & n13170;
  assign n13307 = n13306 ^ n12860;
  assign n13308 = n13307 ^ n13304;
  assign n13309 = n13305 & n13308;
  assign n13310 = n13309 ^ x77;
  assign n13311 = n13310 ^ x78;
  assign n13312 = n12864 & n13170;
  assign n13313 = n13312 ^ n12866;
  assign n13314 = n13313 ^ n13310;
  assign n13315 = n13311 & n13314;
  assign n13316 = n13315 ^ x78;
  assign n13317 = n13316 ^ x79;
  assign n13318 = n12870 & n13170;
  assign n13319 = n13318 ^ n12872;
  assign n13320 = n13319 ^ n13316;
  assign n13321 = n13317 & ~n13320;
  assign n13322 = n13321 ^ x79;
  assign n13323 = n13322 ^ x80;
  assign n13324 = n12876 & n13170;
  assign n13325 = n13324 ^ n12878;
  assign n13326 = n13325 ^ n13322;
  assign n13327 = n13323 & n13326;
  assign n13328 = n13327 ^ x80;
  assign n13329 = n13328 ^ x81;
  assign n13330 = n12882 & n13170;
  assign n13331 = n13330 ^ n12884;
  assign n13332 = n13331 ^ n13328;
  assign n13333 = n13329 & ~n13332;
  assign n13334 = n13333 ^ x81;
  assign n13335 = n13334 ^ x82;
  assign n13336 = n12888 & n13170;
  assign n13337 = n13336 ^ n12891;
  assign n13338 = n13337 ^ n13334;
  assign n13339 = n13335 & ~n13338;
  assign n13340 = n13339 ^ x82;
  assign n13341 = n13340 ^ x83;
  assign n13342 = n12895 & n13170;
  assign n13343 = n13342 ^ n12899;
  assign n13344 = n13343 ^ n13340;
  assign n13345 = n13341 & n13344;
  assign n13346 = n13345 ^ x83;
  assign n13347 = n13346 ^ x84;
  assign n13348 = n12903 & n13170;
  assign n13349 = n13348 ^ n12906;
  assign n13350 = n13349 ^ n13346;
  assign n13351 = n13347 & ~n13350;
  assign n13352 = n13351 ^ x84;
  assign n13353 = n13352 ^ x85;
  assign n13354 = n12910 & n13170;
  assign n13355 = n13354 ^ n12916;
  assign n13356 = n13355 ^ n13352;
  assign n13357 = n13353 & n13356;
  assign n13358 = n13357 ^ x85;
  assign n13359 = n13358 ^ x86;
  assign n13360 = n12920 & n13170;
  assign n13361 = n13360 ^ n12923;
  assign n13362 = n13361 ^ n13358;
  assign n13363 = n13359 & ~n13362;
  assign n13364 = n13363 ^ x86;
  assign n13365 = n13364 ^ x87;
  assign n13366 = n12927 & n13170;
  assign n13367 = n13366 ^ n12933;
  assign n13368 = n13367 ^ n13364;
  assign n13369 = n13365 & n13368;
  assign n13370 = n13369 ^ x87;
  assign n13371 = n13370 ^ x88;
  assign n13372 = n12937 & n13170;
  assign n13373 = n13372 ^ n12939;
  assign n13374 = n13373 ^ n13370;
  assign n13375 = n13371 & ~n13374;
  assign n13376 = n13375 ^ x88;
  assign n13377 = n13376 ^ x89;
  assign n13378 = n12942 ^ x88;
  assign n13379 = n13170 & n13378;
  assign n13380 = n13379 ^ n12754;
  assign n13381 = n13380 ^ n13376;
  assign n13382 = n13377 & ~n13381;
  assign n13383 = n13382 ^ x89;
  assign n13384 = n13383 ^ x90;
  assign n13385 = n12942 ^ n12754;
  assign n13386 = n13378 & ~n13385;
  assign n13387 = n13386 ^ x88;
  assign n13388 = n13387 ^ x89;
  assign n13389 = n13170 & n13388;
  assign n13390 = n13389 ^ n12757;
  assign n13391 = n13390 ^ n13383;
  assign n13392 = n13384 & ~n13391;
  assign n13393 = n13392 ^ x90;
  assign n13394 = n13393 ^ x91;
  assign n13395 = ~n12950 & n13170;
  assign n13396 = n13395 ^ n12952;
  assign n13397 = n13396 ^ n13393;
  assign n13398 = n13394 & ~n13397;
  assign n13399 = n13398 ^ x91;
  assign n13400 = n13399 ^ x92;
  assign n13401 = n12956 & n13170;
  assign n13402 = n13401 ^ n12958;
  assign n13403 = n13402 ^ n13399;
  assign n13404 = n13400 & ~n13403;
  assign n13405 = n13404 ^ x92;
  assign n13406 = ~n13240 & ~n13405;
  assign n13407 = ~x93 & ~n13239;
  assign n13408 = n12969 & n13170;
  assign n13409 = n13408 ^ n12975;
  assign n13410 = ~n13407 & n13409;
  assign n13411 = ~n13406 & n13410;
  assign n13412 = ~x94 & ~n13411;
  assign n13413 = ~n13406 & ~n13407;
  assign n13414 = ~n13409 & ~n13413;
  assign n13415 = ~n13412 & ~n13414;
  assign n13416 = n13415 ^ x95;
  assign n13417 = n12979 & n13170;
  assign n13418 = n13417 ^ n12981;
  assign n13419 = n13418 ^ n13415;
  assign n13420 = n13416 & ~n13419;
  assign n13421 = n13420 ^ x95;
  assign n13422 = n13421 ^ x96;
  assign n13423 = n12984 ^ x95;
  assign n13424 = n13170 & n13423;
  assign n13425 = n13424 ^ n12747;
  assign n13426 = n13425 ^ n13421;
  assign n13427 = n13422 & ~n13426;
  assign n13428 = n13427 ^ x96;
  assign n13429 = n13428 ^ x97;
  assign n13430 = n12984 ^ n12747;
  assign n13431 = n13423 & ~n13430;
  assign n13432 = n13431 ^ x95;
  assign n13433 = n13432 ^ x96;
  assign n13434 = n13170 & n13433;
  assign n13435 = n13434 ^ n12750;
  assign n13436 = n13435 ^ n13428;
  assign n13437 = n13429 & ~n13436;
  assign n13438 = n13437 ^ x97;
  assign n13439 = n13438 ^ x98;
  assign n13440 = ~n12992 & n13170;
  assign n13441 = n13440 ^ n12994;
  assign n13442 = n13441 ^ n13438;
  assign n13443 = n13439 & ~n13442;
  assign n13444 = n13443 ^ x98;
  assign n13445 = n13237 & n13444;
  assign n13446 = n13235 ^ x100;
  assign n13447 = x99 & n13232;
  assign n13448 = n13447 ^ n13235;
  assign n13449 = n13446 & ~n13448;
  assign n13450 = n13449 ^ x100;
  assign n13451 = ~n13445 & ~n13450;
  assign n13452 = n13451 ^ x101;
  assign n13453 = n13010 & n13170;
  assign n13454 = n13453 ^ n13012;
  assign n13455 = n13454 ^ n13451;
  assign n13456 = ~n13452 & n13455;
  assign n13457 = n13456 ^ x101;
  assign n13458 = n13230 & n13457;
  assign n13459 = n13228 ^ x103;
  assign n13460 = x102 & n13225;
  assign n13461 = n13460 ^ n13228;
  assign n13462 = n13459 & ~n13461;
  assign n13463 = n13462 ^ x103;
  assign n13464 = ~n13458 & ~n13463;
  assign n13465 = n13464 ^ x104;
  assign n13466 = n13031 & n13170;
  assign n13467 = n13466 ^ n13033;
  assign n13468 = n13467 ^ n13464;
  assign n13469 = ~n13465 & n13468;
  assign n13470 = n13469 ^ x104;
  assign n13471 = n13470 ^ x105;
  assign n13472 = n13037 & n13170;
  assign n13473 = n13472 ^ n13039;
  assign n13474 = n13473 ^ n13470;
  assign n13475 = n13471 & ~n13474;
  assign n13476 = n13475 ^ x105;
  assign n13477 = n13476 ^ x106;
  assign n13478 = n13043 & n13170;
  assign n13479 = n13478 ^ n13045;
  assign n13480 = n13479 ^ n13476;
  assign n13481 = n13477 & ~n13480;
  assign n13482 = n13481 ^ x106;
  assign n13483 = n13482 ^ x107;
  assign n13484 = n13049 & n13170;
  assign n13485 = n13484 ^ n13051;
  assign n13486 = n13485 ^ n13482;
  assign n13487 = n13483 & ~n13486;
  assign n13488 = n13487 ^ x107;
  assign n13489 = n13488 ^ x108;
  assign n13490 = n13055 & n13170;
  assign n13491 = n13490 ^ n13057;
  assign n13492 = n13491 ^ n13488;
  assign n13493 = n13489 & ~n13492;
  assign n13494 = n13493 ^ x108;
  assign n13495 = n13494 ^ x109;
  assign n13496 = n13061 & n13170;
  assign n13497 = n13496 ^ n13063;
  assign n13498 = n13497 ^ n13494;
  assign n13499 = n13495 & ~n13498;
  assign n13500 = n13499 ^ x109;
  assign n13501 = n13500 ^ x110;
  assign n13502 = n13067 & n13170;
  assign n13503 = n13502 ^ n13070;
  assign n13504 = n13503 ^ n13500;
  assign n13505 = n13501 & ~n13504;
  assign n13506 = n13505 ^ x110;
  assign n13507 = n13506 ^ x111;
  assign n13508 = n13074 & n13170;
  assign n13509 = n13508 ^ n13080;
  assign n13510 = n13509 ^ n13506;
  assign n13511 = n13507 & ~n13510;
  assign n13512 = n13511 ^ x111;
  assign n13513 = n13512 ^ x112;
  assign n13514 = n13084 & n13170;
  assign n13515 = n13514 ^ n13086;
  assign n13516 = n13515 ^ n13512;
  assign n13517 = n13513 & ~n13516;
  assign n13518 = n13517 ^ x112;
  assign n13519 = n13518 ^ x113;
  assign n13520 = n13089 ^ x112;
  assign n13521 = n13170 & n13520;
  assign n13522 = n13521 ^ n12744;
  assign n13523 = n13522 ^ n13518;
  assign n13524 = n13519 & ~n13523;
  assign n13525 = n13524 ^ x113;
  assign n13526 = n13525 ^ x114;
  assign n13527 = ~n13090 & ~n13094;
  assign n13528 = n13527 ^ x113;
  assign n13529 = n13170 & ~n13528;
  assign n13530 = n13529 ^ n13092;
  assign n13531 = n13530 ^ n13525;
  assign n13532 = n13526 & ~n13531;
  assign n13533 = n13532 ^ x114;
  assign n13534 = n13223 & n13533;
  assign n13535 = n13221 ^ x116;
  assign n13536 = x115 & n13218;
  assign n13537 = n13536 ^ n13221;
  assign n13538 = n13535 & ~n13537;
  assign n13539 = n13538 ^ x116;
  assign n13540 = ~n13534 & ~n13539;
  assign n13541 = n13540 ^ x117;
  assign n13542 = n13112 & n13170;
  assign n13543 = n13542 ^ n13115;
  assign n13544 = n13543 ^ n13540;
  assign n13545 = ~n13541 & n13544;
  assign n13546 = n13545 ^ x117;
  assign n13547 = n13546 ^ x118;
  assign n13548 = n13119 & n13170;
  assign n13549 = n13548 ^ n13121;
  assign n13550 = n13549 ^ n13546;
  assign n13551 = n13547 & ~n13550;
  assign n13552 = n13551 ^ x118;
  assign n13553 = n13552 ^ x119;
  assign n13554 = n13125 & n13170;
  assign n13555 = n13554 ^ n13127;
  assign n13556 = n13555 ^ n13552;
  assign n13557 = n13553 & ~n13556;
  assign n13558 = n13557 ^ x119;
  assign n13559 = n13558 ^ x120;
  assign n13560 = n13131 & n13170;
  assign n13561 = n13560 ^ n13133;
  assign n13562 = n13561 ^ n13558;
  assign n13563 = n13559 & ~n13562;
  assign n13564 = n13563 ^ x120;
  assign n13565 = n13564 ^ x121;
  assign n13566 = n13137 & n13170;
  assign n13567 = n13566 ^ n13139;
  assign n13568 = n13567 ^ n13564;
  assign n13569 = n13565 & ~n13568;
  assign n13570 = n13569 ^ x121;
  assign n13571 = n13570 ^ x122;
  assign n13572 = n13143 & n13170;
  assign n13573 = n13572 ^ n13145;
  assign n13574 = n13573 ^ n13570;
  assign n13575 = n13571 & ~n13574;
  assign n13576 = n13575 ^ x122;
  assign n13577 = n13576 ^ x123;
  assign n13578 = n13149 & n13170;
  assign n13579 = n13578 ^ n13151;
  assign n13580 = n13579 ^ n13576;
  assign n13581 = n13577 & ~n13580;
  assign n13582 = n13581 ^ x123;
  assign n13583 = n13582 ^ x124;
  assign n13584 = n13155 & n13170;
  assign n13585 = n13584 ^ n13158;
  assign n13586 = n13585 ^ n13582;
  assign n13587 = n13583 & n13586;
  assign n13588 = n13587 ^ x124;
  assign n13589 = ~n13216 & n13588;
  assign n13590 = x125 & ~n11904;
  assign n13591 = ~n13589 & ~n13590;
  assign n13592 = n129 & n13591;
  assign n13593 = n13211 & n13592;
  assign n13594 = n13593 ^ n13245;
  assign n13595 = ~x69 & ~n13594;
  assign n13596 = n13205 & n13592;
  assign n13597 = n13596 ^ n13207;
  assign n13598 = ~x68 & ~n13597;
  assign n13599 = ~n13595 & ~n13598;
  assign n13600 = x64 & n13592;
  assign n13601 = x1 & n13180;
  assign n13602 = n13601 ^ x2;
  assign n13603 = n13600 & n13602;
  assign n13604 = ~x1 & n13192;
  assign n13605 = ~n13173 & ~n13604;
  assign n13606 = ~n13592 & ~n13605;
  assign n13607 = ~x1 & x65;
  assign n13608 = n13607 ^ n13173;
  assign n13609 = x64 & n13608;
  assign n13610 = n13609 ^ n13173;
  assign n13611 = ~n13606 & ~n13610;
  assign n13612 = ~n13603 & n13611;
  assign n13613 = n13612 ^ x66;
  assign n13614 = x65 & n13592;
  assign n13615 = ~n13185 & ~n13192;
  assign n13616 = n13614 & n13615;
  assign n13617 = ~x65 & n13192;
  assign n13618 = ~n13170 & n13617;
  assign n13619 = n13592 & n13618;
  assign n13620 = x65 ^ x2;
  assign n13621 = n13591 & ~n13620;
  assign n13622 = n13185 & ~n13621;
  assign n13623 = ~n13619 & ~n13622;
  assign n13624 = ~n13616 & n13623;
  assign n13625 = n13624 ^ x3;
  assign n13626 = n13625 ^ n13612;
  assign n13627 = ~n13613 & n13626;
  assign n13628 = n13627 ^ x66;
  assign n13629 = n13628 ^ x67;
  assign n13632 = n13177 & ~n13180;
  assign n13633 = n13174 & ~n13632;
  assign n13634 = x64 & ~n13633;
  assign n13635 = ~n13186 & ~n13634;
  assign n13636 = n13635 ^ x66;
  assign n13637 = n13592 & ~n13636;
  assign n13630 = ~n12779 & n13194;
  assign n13631 = n13630 ^ n13175;
  assign n13638 = n13637 ^ n13631;
  assign n13639 = n13638 ^ n13628;
  assign n13640 = n13629 & n13639;
  assign n13641 = n13640 ^ x67;
  assign n13642 = n13599 & n13641;
  assign n13643 = n13594 ^ x69;
  assign n13644 = x68 & n13597;
  assign n13645 = n13644 ^ n13594;
  assign n13646 = n13643 & ~n13645;
  assign n13647 = n13646 ^ x69;
  assign n13648 = ~n13642 & ~n13647;
  assign n13649 = n13648 ^ x70;
  assign n13650 = n13249 & n13592;
  assign n13651 = n13650 ^ n13251;
  assign n13652 = n13651 ^ n13648;
  assign n13653 = ~n13649 & n13652;
  assign n13654 = n13653 ^ x70;
  assign n13655 = n13654 ^ x71;
  assign n13656 = n13254 ^ x70;
  assign n13657 = n13592 & n13656;
  assign n13658 = n13657 ^ n13242;
  assign n13659 = n13658 ^ n13654;
  assign n13660 = n13655 & ~n13659;
  assign n13661 = n13660 ^ x71;
  assign n13662 = n13661 ^ x72;
  assign n13663 = n13257 & ~n13264;
  assign n13664 = n13663 ^ x71;
  assign n13665 = n13592 & ~n13664;
  assign n13666 = n13665 ^ n13259;
  assign n13667 = n13666 ^ n13661;
  assign n13668 = n13662 & ~n13667;
  assign n13669 = n13668 ^ x72;
  assign n13670 = n13669 ^ x73;
  assign n13671 = ~n13270 & n13592;
  assign n13672 = n13671 ^ n13272;
  assign n13673 = n13672 ^ n13669;
  assign n13674 = n13670 & ~n13673;
  assign n13675 = n13674 ^ x73;
  assign n13676 = n13675 ^ x74;
  assign n13677 = n13276 & n13592;
  assign n13678 = n13677 ^ n13278;
  assign n13679 = n13678 ^ n13675;
  assign n13680 = n13676 & n13679;
  assign n13681 = n13680 ^ x74;
  assign n13682 = n13681 ^ x75;
  assign n13683 = n13282 & n13592;
  assign n13684 = n13683 ^ n13284;
  assign n13685 = n13684 ^ n13681;
  assign n13686 = n13682 & ~n13685;
  assign n13687 = n13686 ^ x75;
  assign n13688 = n13687 ^ x76;
  assign n13689 = n13288 & n13592;
  assign n13690 = n13689 ^ n13291;
  assign n13691 = n13690 ^ n13687;
  assign n13692 = n13688 & n13691;
  assign n13693 = n13692 ^ x76;
  assign n13694 = n13693 ^ x77;
  assign n13695 = n13295 & n13592;
  assign n13696 = n13695 ^ n13301;
  assign n13697 = n13696 ^ n13693;
  assign n13698 = n13694 & ~n13697;
  assign n13699 = n13698 ^ x77;
  assign n13700 = n13699 ^ x78;
  assign n13701 = n13305 & n13592;
  assign n13702 = n13701 ^ n13307;
  assign n13703 = n13702 ^ n13699;
  assign n13704 = n13700 & n13703;
  assign n13705 = n13704 ^ x78;
  assign n13706 = n13705 ^ x79;
  assign n13707 = n13311 & n13592;
  assign n13708 = n13707 ^ n13313;
  assign n13709 = n13708 ^ n13705;
  assign n13710 = n13706 & n13709;
  assign n13711 = n13710 ^ x79;
  assign n13712 = n13711 ^ x80;
  assign n13713 = n13317 & n13592;
  assign n13714 = n13713 ^ n13319;
  assign n13715 = n13714 ^ n13711;
  assign n13716 = n13712 & ~n13715;
  assign n13717 = n13716 ^ x80;
  assign n13718 = n13717 ^ x81;
  assign n13719 = n13323 & n13592;
  assign n13720 = n13719 ^ n13325;
  assign n13721 = n13720 ^ n13717;
  assign n13722 = n13718 & n13721;
  assign n13723 = n13722 ^ x81;
  assign n13724 = n13723 ^ x82;
  assign n13725 = n13329 & n13592;
  assign n13726 = n13725 ^ n13331;
  assign n13727 = n13726 ^ n13723;
  assign n13728 = n13724 & ~n13727;
  assign n13729 = n13728 ^ x82;
  assign n13730 = n13729 ^ x83;
  assign n13731 = n13335 & n13592;
  assign n13732 = n13731 ^ n13337;
  assign n13733 = n13732 ^ n13729;
  assign n13734 = n13730 & ~n13733;
  assign n13735 = n13734 ^ x83;
  assign n13736 = n13735 ^ x84;
  assign n13737 = n13341 & n13592;
  assign n13738 = n13737 ^ n13343;
  assign n13739 = n13738 ^ n13735;
  assign n13740 = n13736 & n13739;
  assign n13741 = n13740 ^ x84;
  assign n13742 = n13741 ^ x85;
  assign n13743 = ~n13541 & n13592;
  assign n13744 = n13743 ^ n13543;
  assign n13745 = ~x118 & ~n13744;
  assign n13746 = n13547 & n13592;
  assign n13747 = n13746 ^ n13549;
  assign n13748 = ~x119 & ~n13747;
  assign n13749 = ~n13745 & ~n13748;
  assign n13750 = n13513 & n13592;
  assign n13751 = n13750 ^ n13515;
  assign n13752 = ~x113 & ~n13751;
  assign n13753 = n13519 & n13592;
  assign n13754 = n13753 ^ n13522;
  assign n13755 = ~x114 & ~n13754;
  assign n13756 = ~n13752 & ~n13755;
  assign n13757 = n13457 ^ x102;
  assign n13758 = n13592 & n13757;
  assign n13759 = n13758 ^ n13225;
  assign n13760 = ~x103 & ~n13759;
  assign n13761 = n13347 & n13592;
  assign n13762 = n13761 ^ n13349;
  assign n13763 = n13762 ^ n13741;
  assign n13764 = n13742 & ~n13763;
  assign n13765 = n13764 ^ x85;
  assign n13766 = n13765 ^ x86;
  assign n13767 = n13353 & n13592;
  assign n13768 = n13767 ^ n13355;
  assign n13769 = n13768 ^ n13765;
  assign n13770 = n13766 & n13769;
  assign n13771 = n13770 ^ x86;
  assign n13772 = n13771 ^ x87;
  assign n13773 = n13359 & n13592;
  assign n13774 = n13773 ^ n13361;
  assign n13775 = n13774 ^ n13771;
  assign n13776 = n13772 & ~n13775;
  assign n13777 = n13776 ^ x87;
  assign n13778 = n13777 ^ x88;
  assign n13779 = n13365 & n13592;
  assign n13780 = n13779 ^ n13367;
  assign n13781 = n13780 ^ n13777;
  assign n13782 = n13778 & n13781;
  assign n13783 = n13782 ^ x88;
  assign n13784 = n13783 ^ x89;
  assign n13785 = n13371 & n13592;
  assign n13786 = n13785 ^ n13373;
  assign n13787 = n13786 ^ n13783;
  assign n13788 = n13784 & ~n13787;
  assign n13789 = n13788 ^ x89;
  assign n13790 = n13789 ^ x90;
  assign n13791 = n13377 & n13592;
  assign n13792 = n13791 ^ n13380;
  assign n13793 = n13792 ^ n13789;
  assign n13794 = n13790 & ~n13793;
  assign n13795 = n13794 ^ x90;
  assign n13796 = n13795 ^ x91;
  assign n13797 = n13384 & n13592;
  assign n13798 = n13797 ^ n13390;
  assign n13799 = n13798 ^ n13795;
  assign n13800 = n13796 & ~n13799;
  assign n13801 = n13800 ^ x91;
  assign n13802 = n13801 ^ x92;
  assign n13803 = n13394 & n13592;
  assign n13804 = n13803 ^ n13396;
  assign n13805 = n13804 ^ n13801;
  assign n13806 = n13802 & ~n13805;
  assign n13807 = n13806 ^ x92;
  assign n13808 = n13807 ^ x93;
  assign n13809 = n13400 & n13592;
  assign n13810 = n13809 ^ n13402;
  assign n13811 = n13810 ^ n13807;
  assign n13812 = n13808 & ~n13811;
  assign n13813 = n13812 ^ x93;
  assign n13814 = n13813 ^ x94;
  assign n13815 = n13405 ^ x93;
  assign n13816 = n13592 & n13815;
  assign n13817 = n13816 ^ n13239;
  assign n13818 = n13817 ^ n13813;
  assign n13819 = n13814 & ~n13818;
  assign n13820 = n13819 ^ x94;
  assign n13821 = n13820 ^ x95;
  assign n13822 = n13413 ^ x94;
  assign n13823 = n13592 & n13822;
  assign n13824 = n13823 ^ n13409;
  assign n13825 = n13824 ^ n13820;
  assign n13826 = n13821 & ~n13825;
  assign n13827 = n13826 ^ x95;
  assign n13828 = n13827 ^ x96;
  assign n13829 = n13416 & n13592;
  assign n13830 = n13829 ^ n13418;
  assign n13831 = n13830 ^ n13827;
  assign n13832 = n13828 & ~n13831;
  assign n13833 = n13832 ^ x96;
  assign n13834 = n13833 ^ x97;
  assign n13835 = n13422 & n13592;
  assign n13836 = n13835 ^ n13425;
  assign n13837 = n13836 ^ n13833;
  assign n13838 = n13834 & ~n13837;
  assign n13839 = n13838 ^ x97;
  assign n13840 = n13839 ^ x98;
  assign n13841 = n13429 & n13592;
  assign n13842 = n13841 ^ n13435;
  assign n13843 = n13842 ^ n13839;
  assign n13844 = n13840 & ~n13843;
  assign n13845 = n13844 ^ x98;
  assign n13846 = n13845 ^ x99;
  assign n13847 = n13439 & n13592;
  assign n13848 = n13847 ^ n13441;
  assign n13849 = n13848 ^ n13845;
  assign n13850 = n13846 & ~n13849;
  assign n13851 = n13850 ^ x99;
  assign n13852 = n13851 ^ x100;
  assign n13853 = n13444 ^ x99;
  assign n13854 = n13592 & n13853;
  assign n13855 = n13854 ^ n13232;
  assign n13856 = n13855 ^ n13851;
  assign n13857 = n13852 & ~n13856;
  assign n13858 = n13857 ^ x100;
  assign n13859 = n13858 ^ x101;
  assign n13860 = n13444 ^ n13232;
  assign n13861 = n13853 & ~n13860;
  assign n13862 = n13861 ^ x99;
  assign n13863 = n13862 ^ x100;
  assign n13864 = n13592 & n13863;
  assign n13865 = n13864 ^ n13235;
  assign n13866 = n13865 ^ n13858;
  assign n13867 = n13859 & ~n13866;
  assign n13868 = n13867 ^ x101;
  assign n13869 = n13868 ^ x102;
  assign n13870 = ~n13452 & n13592;
  assign n13871 = n13870 ^ n13454;
  assign n13872 = n13871 ^ n13868;
  assign n13873 = n13869 & ~n13872;
  assign n13874 = n13873 ^ x102;
  assign n13875 = ~n13760 & n13874;
  assign n13876 = x103 & n13759;
  assign n13877 = n13457 ^ n13225;
  assign n13878 = n13757 & ~n13877;
  assign n13879 = n13878 ^ x102;
  assign n13880 = n13879 ^ x103;
  assign n13881 = n13592 & n13880;
  assign n13882 = n13881 ^ n13228;
  assign n13883 = x104 & n13882;
  assign n13884 = ~n13876 & ~n13883;
  assign n13885 = ~n13875 & n13884;
  assign n13886 = ~x104 & ~n13882;
  assign n13887 = ~n13885 & ~n13886;
  assign n13888 = n13887 ^ x105;
  assign n13889 = ~n13465 & n13592;
  assign n13890 = n13889 ^ n13467;
  assign n13891 = n13890 ^ n13887;
  assign n13892 = n13888 & ~n13891;
  assign n13893 = n13892 ^ x105;
  assign n13894 = n13893 ^ x106;
  assign n13895 = n13471 & n13592;
  assign n13896 = n13895 ^ n13473;
  assign n13897 = n13896 ^ n13893;
  assign n13898 = n13894 & ~n13897;
  assign n13899 = n13898 ^ x106;
  assign n13900 = n13899 ^ x107;
  assign n13901 = n13477 & n13592;
  assign n13902 = n13901 ^ n13479;
  assign n13903 = n13902 ^ n13899;
  assign n13904 = n13900 & ~n13903;
  assign n13905 = n13904 ^ x107;
  assign n13906 = n13905 ^ x108;
  assign n13907 = n13483 & n13592;
  assign n13908 = n13907 ^ n13485;
  assign n13909 = n13908 ^ n13905;
  assign n13910 = n13906 & ~n13909;
  assign n13911 = n13910 ^ x108;
  assign n13912 = n13911 ^ x109;
  assign n13913 = n13489 & n13592;
  assign n13914 = n13913 ^ n13491;
  assign n13915 = n13914 ^ n13911;
  assign n13916 = n13912 & ~n13915;
  assign n13917 = n13916 ^ x109;
  assign n13918 = n13917 ^ x110;
  assign n13919 = n13495 & n13592;
  assign n13920 = n13919 ^ n13497;
  assign n13921 = n13920 ^ n13917;
  assign n13922 = n13918 & ~n13921;
  assign n13923 = n13922 ^ x110;
  assign n13924 = n13923 ^ x111;
  assign n13925 = n13501 & n13592;
  assign n13926 = n13925 ^ n13503;
  assign n13927 = n13926 ^ n13923;
  assign n13928 = n13924 & ~n13927;
  assign n13929 = n13928 ^ x111;
  assign n13930 = n13929 ^ x112;
  assign n13931 = n13507 & n13592;
  assign n13932 = n13931 ^ n13509;
  assign n13933 = n13932 ^ n13929;
  assign n13934 = n13930 & ~n13933;
  assign n13935 = n13934 ^ x112;
  assign n13936 = n13756 & n13935;
  assign n13937 = n13754 ^ x114;
  assign n13938 = x113 & n13751;
  assign n13939 = n13938 ^ n13754;
  assign n13940 = n13937 & ~n13939;
  assign n13941 = n13940 ^ x114;
  assign n13942 = ~n13936 & ~n13941;
  assign n13943 = n13942 ^ x115;
  assign n13944 = n13526 & n13592;
  assign n13945 = n13944 ^ n13530;
  assign n13946 = n13945 ^ n13942;
  assign n13947 = ~n13943 & n13946;
  assign n13948 = n13947 ^ x115;
  assign n13949 = n13948 ^ x116;
  assign n13950 = n13533 ^ x115;
  assign n13951 = n13592 & n13950;
  assign n13952 = n13951 ^ n13218;
  assign n13953 = n13952 ^ n13948;
  assign n13954 = n13949 & ~n13953;
  assign n13955 = n13954 ^ x116;
  assign n13956 = n13955 ^ x117;
  assign n13957 = n13533 ^ n13218;
  assign n13958 = n13950 & ~n13957;
  assign n13959 = n13958 ^ x115;
  assign n13960 = n13959 ^ x116;
  assign n13961 = n13592 & n13960;
  assign n13962 = n13961 ^ n13221;
  assign n13963 = n13962 ^ n13955;
  assign n13964 = n13956 & ~n13963;
  assign n13965 = n13964 ^ x117;
  assign n13966 = n13749 & n13965;
  assign n13967 = n13747 ^ x119;
  assign n13968 = x118 & n13744;
  assign n13969 = n13968 ^ n13747;
  assign n13970 = n13967 & ~n13969;
  assign n13971 = n13970 ^ x119;
  assign n13972 = ~n13966 & ~n13971;
  assign n13973 = n13972 ^ x120;
  assign n13974 = n13553 & n13592;
  assign n13975 = n13974 ^ n13555;
  assign n13976 = n13975 ^ n13972;
  assign n13977 = ~n13973 & n13976;
  assign n13978 = n13977 ^ x120;
  assign n13979 = n13978 ^ x121;
  assign n13980 = n13559 & n13592;
  assign n13981 = n13980 ^ n13561;
  assign n13982 = n13981 ^ n13978;
  assign n13983 = n13979 & ~n13982;
  assign n13984 = n13983 ^ x121;
  assign n13985 = n13984 ^ x122;
  assign n13986 = n13565 & n13592;
  assign n13987 = n13986 ^ n13567;
  assign n13988 = n13987 ^ n13984;
  assign n13989 = n13985 & ~n13988;
  assign n13990 = n13989 ^ x122;
  assign n13991 = n13990 ^ x123;
  assign n13992 = n13571 & n13592;
  assign n13993 = n13992 ^ n13573;
  assign n13994 = n13993 ^ n13990;
  assign n13995 = n13991 & ~n13994;
  assign n13996 = n13995 ^ x123;
  assign n13997 = n13996 ^ x124;
  assign n13998 = n13577 & n13592;
  assign n13999 = n13998 ^ n13579;
  assign n14000 = n13999 ^ n13996;
  assign n14001 = n13997 & ~n14000;
  assign n14002 = n14001 ^ x124;
  assign n14003 = n14002 ^ x125;
  assign n14004 = n13583 & n13592;
  assign n14005 = n14004 ^ n13585;
  assign n14006 = n14005 ^ n14002;
  assign n14007 = n14003 & n14006;
  assign n14008 = n14007 ^ x125;
  assign n14009 = n14008 ^ x126;
  assign n14010 = n13588 ^ x125;
  assign n14011 = n13215 & n14010;
  assign n14012 = n129 & n14011;
  assign n14013 = n14012 ^ n13215;
  assign n14014 = n14013 ^ n14008;
  assign n14015 = n14009 & n14014;
  assign n14016 = n14015 ^ x126;
  assign n14017 = ~x127 & ~n14016;
  assign n14018 = n13742 & n14017;
  assign n14019 = n14018 ^ n13762;
  assign n14020 = ~x86 & ~n14019;
  assign n14021 = n13766 & n14017;
  assign n14022 = n14021 ^ n13768;
  assign n14023 = ~x87 & n14022;
  assign n14024 = ~n14020 & ~n14023;
  assign n14025 = n13682 & n14017;
  assign n14026 = n14025 ^ n13684;
  assign n14027 = ~x76 & ~n14026;
  assign n14028 = n13688 & n14017;
  assign n14029 = n14028 ^ n13690;
  assign n14030 = ~x77 & n14029;
  assign n14031 = ~n14027 & ~n14030;
  assign n14032 = ~n13649 & n14017;
  assign n14033 = n14032 ^ n13651;
  assign n14034 = x71 & n14033;
  assign n14035 = x64 & n14017;
  assign n14036 = x0 & ~x65;
  assign n14037 = x1 & ~n14036;
  assign n14038 = n14035 & n14037;
  assign n14039 = ~x0 & x64;
  assign n14040 = ~x1 & n14039;
  assign n14041 = ~n13607 & ~n14040;
  assign n14042 = ~n14017 & ~n14041;
  assign n14043 = x1 ^ x0;
  assign n14044 = ~x64 & n14043;
  assign n14045 = n14044 ^ x0;
  assign n14046 = x65 & ~n14045;
  assign n14047 = ~n14042 & ~n14046;
  assign n14048 = ~n14038 & n14047;
  assign n14049 = n14048 ^ x66;
  assign n14050 = x65 & ~x127;
  assign n14051 = ~n13592 & n14050;
  assign n14052 = ~n14016 & n14051;
  assign n14053 = n219 & n13592;
  assign n14054 = ~n14052 & ~n14053;
  assign n14055 = x1 & ~n14054;
  assign n14056 = n13592 ^ x65;
  assign n14057 = n341 & ~n14056;
  assign n14058 = x1 & n14057;
  assign n14059 = n14058 ^ n340;
  assign n14060 = n14017 & n14059;
  assign n14061 = n14060 ^ n13600;
  assign n14062 = ~n14055 & ~n14061;
  assign n14063 = n14062 ^ x2;
  assign n14064 = n14063 ^ n14048;
  assign n14065 = ~n14049 & n14064;
  assign n14066 = n14065 ^ x66;
  assign n14067 = n14066 ^ x67;
  assign n14068 = ~n13613 & n14017;
  assign n14069 = n14068 ^ n13625;
  assign n14070 = n14069 ^ n14066;
  assign n14071 = n14067 & ~n14070;
  assign n14072 = n14071 ^ x67;
  assign n14073 = n14072 ^ x68;
  assign n14074 = n13629 & n14017;
  assign n14075 = n14074 ^ n13638;
  assign n14076 = n14075 ^ n14072;
  assign n14077 = n14073 & n14076;
  assign n14078 = n14077 ^ x68;
  assign n14079 = n14078 ^ x69;
  assign n14080 = n13641 ^ x68;
  assign n14081 = n14017 & n14080;
  assign n14082 = n14081 ^ n13597;
  assign n14083 = n14082 ^ n14078;
  assign n14084 = n14079 & ~n14083;
  assign n14085 = n14084 ^ x69;
  assign n14086 = n14085 ^ x70;
  assign n14087 = n13641 ^ n13597;
  assign n14088 = n14080 & ~n14087;
  assign n14089 = n14088 ^ x68;
  assign n14090 = n14089 ^ x69;
  assign n14091 = n14017 & n14090;
  assign n14092 = n14091 ^ n13594;
  assign n14093 = n14092 ^ n14085;
  assign n14094 = n14086 & ~n14093;
  assign n14095 = n14094 ^ x70;
  assign n14096 = ~n14034 & ~n14095;
  assign n14097 = ~x71 & ~n14033;
  assign n14098 = n13655 & n14017;
  assign n14099 = n14098 ^ n13658;
  assign n14100 = ~n14097 & n14099;
  assign n14101 = ~n14096 & n14100;
  assign n14102 = ~x72 & ~n14101;
  assign n14103 = ~n14096 & ~n14097;
  assign n14104 = ~n14099 & ~n14103;
  assign n14105 = ~n14102 & ~n14104;
  assign n14106 = n14105 ^ x73;
  assign n14107 = n13662 & n14017;
  assign n14108 = n14107 ^ n13666;
  assign n14109 = n14108 ^ n14105;
  assign n14110 = n14106 & ~n14109;
  assign n14111 = n14110 ^ x73;
  assign n14112 = n14111 ^ x74;
  assign n14113 = n13670 & n14017;
  assign n14114 = n14113 ^ n13672;
  assign n14115 = n14114 ^ n14111;
  assign n14116 = n14112 & ~n14115;
  assign n14117 = n14116 ^ x74;
  assign n14118 = n14117 ^ x75;
  assign n14119 = n13676 & n14017;
  assign n14120 = n14119 ^ n13678;
  assign n14121 = n14120 ^ n14117;
  assign n14122 = n14118 & n14121;
  assign n14123 = n14122 ^ x75;
  assign n14124 = n14031 & n14123;
  assign n14125 = n14029 ^ x77;
  assign n14126 = x76 & n14026;
  assign n14127 = n14126 ^ n14029;
  assign n14128 = ~n14125 & n14127;
  assign n14129 = n14128 ^ x77;
  assign n14130 = ~n14124 & ~n14129;
  assign n14131 = n14130 ^ x78;
  assign n14132 = n13694 & n14017;
  assign n14133 = n14132 ^ n13696;
  assign n14134 = n14133 ^ n14130;
  assign n14135 = ~n14131 & n14134;
  assign n14136 = n14135 ^ x78;
  assign n14137 = n14136 ^ x79;
  assign n14138 = n13700 & n14017;
  assign n14139 = n14138 ^ n13702;
  assign n14140 = n14139 ^ n14136;
  assign n14141 = n14137 & n14140;
  assign n14142 = n14141 ^ x79;
  assign n14143 = n14142 ^ x80;
  assign n14144 = n13706 & n14017;
  assign n14145 = n14144 ^ n13708;
  assign n14146 = n14145 ^ n14142;
  assign n14147 = n14143 & n14146;
  assign n14148 = n14147 ^ x80;
  assign n14149 = n14148 ^ x81;
  assign n14150 = n13712 & n14017;
  assign n14151 = n14150 ^ n13714;
  assign n14152 = n14151 ^ n14148;
  assign n14153 = n14149 & ~n14152;
  assign n14154 = n14153 ^ x81;
  assign n14155 = n14154 ^ x82;
  assign n14156 = n13718 & n14017;
  assign n14157 = n14156 ^ n13720;
  assign n14158 = n14157 ^ n14154;
  assign n14159 = n14155 & n14158;
  assign n14160 = n14159 ^ x82;
  assign n14161 = n14160 ^ x83;
  assign n14162 = n13724 & n14017;
  assign n14163 = n14162 ^ n13726;
  assign n14164 = n14163 ^ n14160;
  assign n14165 = n14161 & ~n14164;
  assign n14166 = n14165 ^ x83;
  assign n14167 = n14166 ^ x84;
  assign n14168 = n13730 & n14017;
  assign n14169 = n14168 ^ n13732;
  assign n14170 = n14169 ^ n14166;
  assign n14171 = n14167 & ~n14170;
  assign n14172 = n14171 ^ x84;
  assign n14173 = n14172 ^ x85;
  assign n14174 = n13736 & n14017;
  assign n14175 = n14174 ^ n13738;
  assign n14176 = n14175 ^ n14172;
  assign n14177 = n14173 & n14176;
  assign n14178 = n14177 ^ x85;
  assign n14179 = n14024 & n14178;
  assign n14180 = n14022 ^ x87;
  assign n14181 = x86 & n14019;
  assign n14182 = n14181 ^ n14022;
  assign n14183 = ~n14180 & n14182;
  assign n14184 = n14183 ^ x87;
  assign n14185 = ~n14179 & ~n14184;
  assign n14186 = n14185 ^ x88;
  assign n14187 = n13772 & n14017;
  assign n14188 = n14187 ^ n13774;
  assign n14189 = n14188 ^ n14185;
  assign n14190 = ~n14186 & n14189;
  assign n14191 = n14190 ^ x88;
  assign n14192 = n14191 ^ x89;
  assign n14193 = n13778 & n14017;
  assign n14194 = n14193 ^ n13780;
  assign n14195 = n14194 ^ n14191;
  assign n14196 = n14192 & n14195;
  assign n14197 = n14196 ^ x89;
  assign n14198 = n14197 ^ x90;
  assign n14199 = n13784 & n14017;
  assign n14200 = n14199 ^ n13786;
  assign n14201 = n14200 ^ n14197;
  assign n14202 = n14198 & ~n14201;
  assign n14203 = n14202 ^ x90;
  assign n14204 = n14203 ^ x91;
  assign n14205 = n13790 & n14017;
  assign n14206 = n14205 ^ n13792;
  assign n14207 = n14206 ^ n14203;
  assign n14208 = n14204 & ~n14207;
  assign n14209 = n14208 ^ x91;
  assign n14210 = n14209 ^ x92;
  assign n14211 = n13796 & n14017;
  assign n14212 = n14211 ^ n13798;
  assign n14213 = n14212 ^ n14209;
  assign n14214 = n14210 & ~n14213;
  assign n14215 = n14214 ^ x92;
  assign n14216 = n14215 ^ x93;
  assign n14217 = n13802 & n14017;
  assign n14218 = n14217 ^ n13804;
  assign n14219 = n14218 ^ n14215;
  assign n14220 = n14216 & ~n14219;
  assign n14221 = n14220 ^ x93;
  assign n14222 = n14221 ^ x94;
  assign n14223 = n13808 & n14017;
  assign n14224 = n14223 ^ n13810;
  assign n14225 = n14224 ^ n14221;
  assign n14226 = n14222 & ~n14225;
  assign n14227 = n14226 ^ x94;
  assign n14228 = n14227 ^ x95;
  assign n14229 = n13814 & n14017;
  assign n14230 = n14229 ^ n13817;
  assign n14231 = n14230 ^ n14227;
  assign n14232 = n14228 & ~n14231;
  assign n14233 = n14232 ^ x95;
  assign n14234 = n14233 ^ x96;
  assign n14235 = n13821 & n14017;
  assign n14236 = n14235 ^ n13824;
  assign n14237 = n14236 ^ n14233;
  assign n14238 = n14234 & ~n14237;
  assign n14239 = n14238 ^ x96;
  assign n14240 = n14239 ^ x97;
  assign n14241 = n13828 & n14017;
  assign n14242 = n14241 ^ n13830;
  assign n14243 = n14242 ^ n14239;
  assign n14244 = n14240 & ~n14243;
  assign n14245 = n14244 ^ x97;
  assign n14246 = n14245 ^ x98;
  assign n14247 = n13834 & n14017;
  assign n14248 = n14247 ^ n13836;
  assign n14249 = n14248 ^ n14245;
  assign n14250 = n14246 & ~n14249;
  assign n14251 = n14250 ^ x98;
  assign n14252 = n14251 ^ x99;
  assign n14253 = n13840 & n14017;
  assign n14254 = n14253 ^ n13842;
  assign n14255 = n14254 ^ n14251;
  assign n14256 = n14252 & ~n14255;
  assign n14257 = n14256 ^ x99;
  assign n14258 = n14257 ^ x100;
  assign n14259 = n13846 & n14017;
  assign n14260 = n14259 ^ n13848;
  assign n14261 = n14260 ^ n14257;
  assign n14262 = n14258 & ~n14261;
  assign n14263 = n14262 ^ x100;
  assign n14264 = n14263 ^ x101;
  assign n14265 = n13852 & n14017;
  assign n14266 = n14265 ^ n13855;
  assign n14267 = n14266 ^ n14263;
  assign n14268 = n14264 & ~n14267;
  assign n14269 = n14268 ^ x101;
  assign n14270 = n14269 ^ x102;
  assign n14271 = n13859 & n14017;
  assign n14272 = n14271 ^ n13865;
  assign n14273 = n14272 ^ n14269;
  assign n14274 = n14270 & ~n14273;
  assign n14275 = n14274 ^ x102;
  assign n14276 = n14275 ^ x103;
  assign n14277 = n13869 & n14017;
  assign n14278 = n14277 ^ n13871;
  assign n14279 = n14278 ^ n14275;
  assign n14280 = n14276 & ~n14279;
  assign n14281 = n14280 ^ x103;
  assign n14282 = n14281 ^ x104;
  assign n14283 = n13874 ^ x103;
  assign n14284 = n14017 & n14283;
  assign n14285 = n14284 ^ n13759;
  assign n14286 = n14285 ^ n14281;
  assign n14287 = n14282 & ~n14286;
  assign n14288 = n14287 ^ x104;
  assign n14289 = n14288 ^ x105;
  assign n14290 = ~n13875 & ~n13876;
  assign n14291 = n14290 ^ x104;
  assign n14292 = n14017 & ~n14291;
  assign n14293 = n14292 ^ n13882;
  assign n14294 = n14293 ^ n14288;
  assign n14295 = n14289 & ~n14294;
  assign n14296 = n14295 ^ x105;
  assign n14297 = n14296 ^ x106;
  assign n14298 = n13888 & n14017;
  assign n14299 = n14298 ^ n13890;
  assign n14300 = n14299 ^ n14296;
  assign n14301 = n14297 & ~n14300;
  assign n14302 = n14301 ^ x106;
  assign n14303 = n14302 ^ x107;
  assign n14304 = n13894 & n14017;
  assign n14305 = n14304 ^ n13896;
  assign n14306 = n14305 ^ n14302;
  assign n14307 = n14303 & ~n14306;
  assign n14308 = n14307 ^ x107;
  assign n14309 = n14308 ^ x108;
  assign n14310 = n13900 & n14017;
  assign n14311 = n14310 ^ n13902;
  assign n14312 = n14311 ^ n14308;
  assign n14313 = n14309 & ~n14312;
  assign n14314 = n14313 ^ x108;
  assign n14315 = n14314 ^ x109;
  assign n14316 = n13906 & n14017;
  assign n14317 = n14316 ^ n13908;
  assign n14318 = n14317 ^ n14314;
  assign n14319 = n14315 & ~n14318;
  assign n14320 = n14319 ^ x109;
  assign n14321 = n14320 ^ x110;
  assign n14322 = n13912 & n14017;
  assign n14323 = n14322 ^ n13914;
  assign n14324 = n14323 ^ n14320;
  assign n14325 = n14321 & ~n14324;
  assign n14326 = n14325 ^ x110;
  assign n14327 = n14326 ^ x111;
  assign n14328 = n13918 & n14017;
  assign n14329 = n14328 ^ n13920;
  assign n14330 = n14329 ^ n14326;
  assign n14331 = n14327 & ~n14330;
  assign n14332 = n14331 ^ x111;
  assign n14333 = n14332 ^ x112;
  assign n14334 = n13924 & n14017;
  assign n14335 = n14334 ^ n13926;
  assign n14336 = n14335 ^ n14332;
  assign n14337 = n14333 & ~n14336;
  assign n14338 = n14337 ^ x112;
  assign n14339 = n14338 ^ x113;
  assign n14340 = n13930 & n14017;
  assign n14341 = n14340 ^ n13932;
  assign n14342 = n14341 ^ n14338;
  assign n14343 = n14339 & ~n14342;
  assign n14344 = n14343 ^ x113;
  assign n14345 = n14344 ^ x114;
  assign n14346 = n13935 ^ x113;
  assign n14347 = n14017 & n14346;
  assign n14348 = n14347 ^ n13751;
  assign n14349 = n14348 ^ n14344;
  assign n14350 = n14345 & ~n14349;
  assign n14351 = n14350 ^ x114;
  assign n14352 = n14351 ^ x115;
  assign n14353 = n13935 ^ n13751;
  assign n14354 = n14346 & ~n14353;
  assign n14355 = n14354 ^ x113;
  assign n14356 = n14355 ^ x114;
  assign n14357 = n14017 & n14356;
  assign n14358 = n14357 ^ n13754;
  assign n14359 = n14358 ^ n14351;
  assign n14360 = n14352 & ~n14359;
  assign n14361 = n14360 ^ x115;
  assign n14362 = n14361 ^ x116;
  assign n14363 = ~n13943 & n14017;
  assign n14364 = n14363 ^ n13945;
  assign n14365 = n14364 ^ n14361;
  assign n14366 = n14362 & ~n14365;
  assign n14367 = n14366 ^ x116;
  assign n14368 = n14367 ^ x117;
  assign n14369 = n13949 & n14017;
  assign n14370 = n14369 ^ n13952;
  assign n14371 = n14370 ^ n14367;
  assign n14372 = n14368 & ~n14371;
  assign n14373 = n14372 ^ x117;
  assign n14374 = n14373 ^ x118;
  assign n14375 = n13956 & n14017;
  assign n14376 = n14375 ^ n13962;
  assign n14377 = n14376 ^ n14373;
  assign n14378 = n14374 & ~n14377;
  assign n14379 = n14378 ^ x118;
  assign n14380 = n14379 ^ x119;
  assign n14381 = n13965 ^ x118;
  assign n14382 = n14017 & n14381;
  assign n14383 = n14382 ^ n13744;
  assign n14384 = n14383 ^ n14379;
  assign n14385 = n14380 & ~n14384;
  assign n14386 = n14385 ^ x119;
  assign n14387 = n14386 ^ x120;
  assign n14388 = n13965 ^ n13744;
  assign n14389 = n14381 & ~n14388;
  assign n14390 = n14389 ^ x118;
  assign n14391 = n14390 ^ x119;
  assign n14392 = n14017 & n14391;
  assign n14393 = n14392 ^ n13747;
  assign n14394 = n14393 ^ n14386;
  assign n14395 = n14387 & ~n14394;
  assign n14396 = n14395 ^ x120;
  assign n14397 = n14396 ^ x121;
  assign n14398 = ~n13973 & n14017;
  assign n14399 = n14398 ^ n13975;
  assign n14400 = n14399 ^ n14396;
  assign n14401 = n14397 & ~n14400;
  assign n14402 = n14401 ^ x121;
  assign n14403 = n14402 ^ x122;
  assign n14404 = n13979 & n14017;
  assign n14405 = n14404 ^ n13981;
  assign n14406 = n14405 ^ n14402;
  assign n14407 = n14403 & ~n14406;
  assign n14408 = n14407 ^ x122;
  assign n14409 = n14408 ^ x123;
  assign n14410 = n13985 & n14017;
  assign n14411 = n14410 ^ n13987;
  assign n14412 = n14411 ^ n14408;
  assign n14413 = n14409 & ~n14412;
  assign n14414 = n14413 ^ x123;
  assign n14415 = n14414 ^ x124;
  assign n14416 = n13991 & n14017;
  assign n14417 = n14416 ^ n13993;
  assign n14418 = n14417 ^ n14414;
  assign n14419 = n14415 & ~n14418;
  assign n14420 = n14419 ^ x124;
  assign n14421 = n14420 ^ x125;
  assign n14422 = n13997 & n14017;
  assign n14423 = n14422 ^ n13999;
  assign n14424 = n14423 ^ n14420;
  assign n14425 = n14421 & ~n14424;
  assign n14426 = n14425 ^ x125;
  assign n14427 = n14426 ^ x126;
  assign n14428 = n14003 & n14017;
  assign n14429 = n14428 ^ n14005;
  assign n14430 = n14429 ^ n14426;
  assign n14431 = n14427 & n14430;
  assign n14432 = n14431 ^ x126;
  assign n14433 = ~n12330 & ~n14432;
  assign n14434 = ~x127 & ~n14009;
  assign n14435 = n14013 & n14434;
  assign n14436 = ~n14433 & ~n14435;
  assign n14437 = ~x62 & n228;
  assign n14438 = n14437 ^ n192;
  assign n14439 = ~x63 & x64;
  assign n14440 = ~x65 & ~x66;
  assign n14441 = ~n14439 & n14440;
  assign n14442 = n189 & n14441;
  assign n14443 = x64 & ~n14436;
  assign n14444 = n14443 ^ x0;
  assign n14445 = ~n14036 & ~n14436;
  assign n14446 = n14035 & ~n14445;
  assign n14447 = ~n14017 & n14039;
  assign n14448 = ~x65 & ~n14447;
  assign n14449 = n14039 ^ n14017;
  assign n14450 = n960 & n14449;
  assign n14451 = ~n14448 & ~n14450;
  assign n14452 = ~n14436 & n14451;
  assign n14453 = ~n14446 & ~n14452;
  assign n14454 = n14453 ^ x1;
  assign n14455 = ~n14049 & ~n14436;
  assign n14456 = n14455 ^ n14063;
  assign n14457 = n14067 & ~n14436;
  assign n14458 = n14457 ^ n14069;
  assign n14459 = n14073 & ~n14436;
  assign n14460 = n14459 ^ n14075;
  assign n14461 = n14079 & ~n14436;
  assign n14462 = n14461 ^ n14082;
  assign n14463 = n14086 & ~n14436;
  assign n14464 = n14463 ^ n14092;
  assign n14465 = n14095 ^ x71;
  assign n14466 = ~n14436 & n14465;
  assign n14467 = n14466 ^ n14033;
  assign n14468 = n14103 ^ x72;
  assign n14469 = ~n14436 & n14468;
  assign n14470 = n14469 ^ n14099;
  assign n14471 = n14106 & ~n14436;
  assign n14472 = n14471 ^ n14108;
  assign n14473 = n14112 & ~n14436;
  assign n14474 = n14473 ^ n14114;
  assign n14475 = n14118 & ~n14436;
  assign n14476 = n14475 ^ n14120;
  assign n14477 = n14123 ^ x76;
  assign n14478 = ~n14436 & n14477;
  assign n14479 = n14478 ^ n14026;
  assign n14480 = n14123 ^ n14026;
  assign n14481 = n14477 & ~n14480;
  assign n14482 = n14481 ^ x76;
  assign n14483 = n14482 ^ x77;
  assign n14484 = ~n14436 & n14483;
  assign n14485 = n14484 ^ n14029;
  assign n14486 = ~n14131 & ~n14436;
  assign n14487 = n14486 ^ n14133;
  assign n14488 = n14137 & ~n14436;
  assign n14489 = n14488 ^ n14139;
  assign n14490 = n14143 & ~n14436;
  assign n14491 = n14490 ^ n14145;
  assign n14492 = n14149 & ~n14436;
  assign n14493 = n14492 ^ n14151;
  assign n14494 = n14155 & ~n14436;
  assign n14495 = n14494 ^ n14157;
  assign n14496 = n14161 & ~n14436;
  assign n14497 = n14496 ^ n14163;
  assign n14498 = n14167 & ~n14436;
  assign n14499 = n14498 ^ n14169;
  assign n14500 = n14173 & ~n14436;
  assign n14501 = n14500 ^ n14175;
  assign n14502 = n14178 ^ x86;
  assign n14503 = ~n14436 & n14502;
  assign n14504 = n14503 ^ n14019;
  assign n14505 = n14178 ^ n14019;
  assign n14506 = n14502 & ~n14505;
  assign n14507 = n14506 ^ x86;
  assign n14508 = n14507 ^ x87;
  assign n14509 = ~n14436 & n14508;
  assign n14510 = n14509 ^ n14022;
  assign n14511 = ~n14186 & ~n14436;
  assign n14512 = n14511 ^ n14188;
  assign n14513 = n14192 & ~n14436;
  assign n14514 = n14513 ^ n14194;
  assign n14515 = n14198 & ~n14436;
  assign n14516 = n14515 ^ n14200;
  assign n14517 = n14204 & ~n14436;
  assign n14518 = n14517 ^ n14206;
  assign n14519 = n14210 & ~n14436;
  assign n14520 = n14519 ^ n14212;
  assign n14521 = n14216 & ~n14436;
  assign n14522 = n14521 ^ n14218;
  assign n14523 = n14222 & ~n14436;
  assign n14524 = n14523 ^ n14224;
  assign n14525 = n14228 & ~n14436;
  assign n14526 = n14525 ^ n14230;
  assign n14527 = n14234 & ~n14436;
  assign n14528 = n14527 ^ n14236;
  assign n14529 = n14240 & ~n14436;
  assign n14530 = n14529 ^ n14242;
  assign n14531 = n14246 & ~n14436;
  assign n14532 = n14531 ^ n14248;
  assign n14533 = n14252 & ~n14436;
  assign n14534 = n14533 ^ n14254;
  assign n14535 = n14258 & ~n14436;
  assign n14536 = n14535 ^ n14260;
  assign n14537 = n14264 & ~n14436;
  assign n14538 = n14537 ^ n14266;
  assign n14539 = n14270 & ~n14436;
  assign n14540 = n14539 ^ n14272;
  assign n14541 = n14276 & ~n14436;
  assign n14542 = n14541 ^ n14278;
  assign n14543 = n14282 & ~n14436;
  assign n14544 = n14543 ^ n14285;
  assign n14545 = n14289 & ~n14436;
  assign n14546 = n14545 ^ n14293;
  assign n14547 = n14297 & ~n14436;
  assign n14548 = n14547 ^ n14299;
  assign n14549 = n14303 & ~n14436;
  assign n14550 = n14549 ^ n14305;
  assign n14551 = n14309 & ~n14436;
  assign n14552 = n14551 ^ n14311;
  assign n14553 = n14315 & ~n14436;
  assign n14554 = n14553 ^ n14317;
  assign n14555 = n14321 & ~n14436;
  assign n14556 = n14555 ^ n14323;
  assign n14557 = n14327 & ~n14436;
  assign n14558 = n14557 ^ n14329;
  assign n14559 = n14333 & ~n14436;
  assign n14560 = n14559 ^ n14335;
  assign n14561 = n14339 & ~n14436;
  assign n14562 = n14561 ^ n14341;
  assign n14563 = n14345 & ~n14436;
  assign n14564 = n14563 ^ n14348;
  assign n14565 = n14352 & ~n14436;
  assign n14566 = n14565 ^ n14358;
  assign n14567 = n14362 & ~n14436;
  assign n14568 = n14567 ^ n14364;
  assign n14569 = n14368 & ~n14436;
  assign n14570 = n14569 ^ n14370;
  assign n14571 = n14374 & ~n14436;
  assign n14572 = n14571 ^ n14376;
  assign n14573 = n14380 & ~n14436;
  assign n14574 = n14573 ^ n14383;
  assign n14575 = n14387 & ~n14436;
  assign n14576 = n14575 ^ n14393;
  assign n14577 = n14397 & ~n14436;
  assign n14578 = n14577 ^ n14399;
  assign n14579 = n14403 & ~n14436;
  assign n14580 = n14579 ^ n14405;
  assign n14581 = n14409 & ~n14436;
  assign n14582 = n14581 ^ n14411;
  assign n14583 = n14415 & ~n14436;
  assign n14584 = n14583 ^ n14417;
  assign n14585 = n14421 & ~n14436;
  assign n14586 = n14585 ^ n14423;
  assign n14587 = n14427 & ~n14436;
  assign n14588 = n14587 ^ n14429;
  assign n14589 = ~x127 & n14432;
  assign n14590 = n14013 & ~n14589;
  assign n14591 = ~n14432 & ~n14434;
  assign n14592 = n14590 & ~n14591;
  assign y0 = ~n14436;
  assign y1 = n14017;
  assign y2 = n13592;
  assign y3 = n13170;
  assign y4 = n12742;
  assign y5 = ~n12337;
  assign y6 = n11937;
  assign y7 = n11548;
  assign y8 = ~n11171;
  assign y9 = n10784;
  assign y10 = n10406;
  assign y11 = n10045;
  assign y12 = n9681;
  assign y13 = n9328;
  assign y14 = n8977;
  assign y15 = ~n8648;
  assign y16 = n8301;
  assign y17 = ~n7987;
  assign y18 = n7671;
  assign y19 = ~n7365;
  assign y20 = n7049;
  assign y21 = n6742;
  assign y22 = ~n6433;
  assign y23 = n6143;
  assign y24 = n5863;
  assign y25 = n5597;
  assign y26 = n5322;
  assign y27 = ~n5046;
  assign y28 = n4786;
  assign y29 = n4546;
  assign y30 = n4318;
  assign y31 = n4086;
  assign y32 = ~n3862;
  assign y33 = n3646;
  assign y34 = n3435;
  assign y35 = n3225;
  assign y36 = n3025;
  assign y37 = n2835;
  assign y38 = n2655;
  assign y39 = n2477;
  assign y40 = n2306;
  assign y41 = ~n2140;
  assign y42 = n1990;
  assign y43 = n1832;
  assign y44 = n1681;
  assign y45 = n1540;
  assign y46 = ~n1415;
  assign y47 = n1288;
  assign y48 = n1170;
  assign y49 = ~n1063;
  assign y50 = n957;
  assign y51 = n860;
  assign y52 = n773;
  assign y53 = ~n689;
  assign y54 = n605;
  assign y55 = ~n525;
  assign y56 = n453;
  assign y57 = n392;
  assign y58 = n334;
  assign y59 = n285;
  assign y60 = ~n247;
  assign y61 = n215;
  assign y62 = n14438;
  assign y63 = n14442;
  assign y64 = n14444;
  assign y65 = ~n14454;
  assign y66 = ~n14456;
  assign y67 = ~n14458;
  assign y68 = n14460;
  assign y69 = ~n14462;
  assign y70 = ~n14464;
  assign y71 = ~n14467;
  assign y72 = ~n14470;
  assign y73 = ~n14472;
  assign y74 = ~n14474;
  assign y75 = n14476;
  assign y76 = ~n14479;
  assign y77 = n14485;
  assign y78 = ~n14487;
  assign y79 = n14489;
  assign y80 = n14491;
  assign y81 = ~n14493;
  assign y82 = n14495;
  assign y83 = ~n14497;
  assign y84 = ~n14499;
  assign y85 = n14501;
  assign y86 = ~n14504;
  assign y87 = n14510;
  assign y88 = ~n14512;
  assign y89 = n14514;
  assign y90 = ~n14516;
  assign y91 = ~n14518;
  assign y92 = ~n14520;
  assign y93 = ~n14522;
  assign y94 = ~n14524;
  assign y95 = ~n14526;
  assign y96 = ~n14528;
  assign y97 = ~n14530;
  assign y98 = ~n14532;
  assign y99 = ~n14534;
  assign y100 = ~n14536;
  assign y101 = ~n14538;
  assign y102 = ~n14540;
  assign y103 = ~n14542;
  assign y104 = ~n14544;
  assign y105 = ~n14546;
  assign y106 = ~n14548;
  assign y107 = ~n14550;
  assign y108 = ~n14552;
  assign y109 = ~n14554;
  assign y110 = ~n14556;
  assign y111 = ~n14558;
  assign y112 = ~n14560;
  assign y113 = ~n14562;
  assign y114 = ~n14564;
  assign y115 = ~n14566;
  assign y116 = ~n14568;
  assign y117 = ~n14570;
  assign y118 = ~n14572;
  assign y119 = ~n14574;
  assign y120 = ~n14576;
  assign y121 = ~n14578;
  assign y122 = ~n14580;
  assign y123 = ~n14582;
  assign y124 = ~n14584;
  assign y125 = ~n14586;
  assign y126 = n14588;
  assign y127 = n14592;
endmodule
