module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63;
  wire n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673;
  assign n65 = x0 & x32;
  assign n74 = x33 & ~n65;
  assign n66 = x32 & ~x33;
  assign n67 = x1 & n66;
  assign n68 = x32 & x33;
  assign n69 = ~x1 & n68;
  assign n70 = ~x32 & x33;
  assign n71 = ~x0 & n70;
  assign n72 = ~n69 & ~n71;
  assign n73 = ~n67 & n72;
  assign n75 = n74 ^ n73;
  assign n84 = ~n73 & n74;
  assign n81 = x34 ^ x33;
  assign n82 = x0 & n81;
  assign n76 = x2 & n66;
  assign n77 = ~x2 & n68;
  assign n78 = ~x1 & n70;
  assign n79 = ~n77 & ~n78;
  assign n80 = ~n76 & n79;
  assign n83 = n82 ^ n80;
  assign n85 = n84 ^ n83;
  assign n110 = ~n80 & n82;
  assign n111 = n80 & ~n82;
  assign n112 = n84 & ~n111;
  assign n113 = ~n110 & ~n112;
  assign n96 = x35 & n81;
  assign n97 = ~x1 & n96;
  assign n98 = x35 ^ x34;
  assign n99 = ~n81 & n98;
  assign n100 = x35 & n99;
  assign n101 = ~x0 & n100;
  assign n102 = ~n97 & ~n101;
  assign n103 = ~x35 & n81;
  assign n104 = x1 & n103;
  assign n105 = ~x35 & n99;
  assign n106 = x0 & n105;
  assign n107 = ~n104 & ~n106;
  assign n108 = n102 & n107;
  assign n90 = x3 & n66;
  assign n91 = ~x3 & n68;
  assign n92 = ~x2 & n70;
  assign n93 = ~n91 & ~n92;
  assign n94 = ~n90 & n93;
  assign n86 = x33 ^ x0;
  assign n87 = ~n81 & n86;
  assign n88 = n87 ^ x0;
  assign n89 = x35 & ~n88;
  assign n95 = n94 ^ n89;
  assign n109 = n108 ^ n95;
  assign n114 = n113 ^ n109;
  assign n133 = ~n95 & ~n108;
  assign n134 = n95 & n108;
  assign n135 = ~n113 & ~n134;
  assign n136 = ~n133 & ~n135;
  assign n131 = n89 & ~n94;
  assign n125 = x4 & n66;
  assign n126 = ~x4 & n68;
  assign n127 = ~x3 & n70;
  assign n128 = ~n126 & ~n127;
  assign n129 = ~n125 & n128;
  assign n122 = x36 ^ x35;
  assign n123 = x0 & n122;
  assign n115 = x2 & n103;
  assign n116 = x1 & n105;
  assign n117 = ~n115 & ~n116;
  assign n118 = ~x2 & n96;
  assign n119 = ~x1 & n100;
  assign n120 = ~n118 & ~n119;
  assign n121 = n117 & n120;
  assign n124 = n123 ^ n121;
  assign n130 = n129 ^ n124;
  assign n132 = n131 ^ n130;
  assign n137 = n136 ^ n132;
  assign n175 = n130 & n131;
  assign n176 = ~n130 & ~n131;
  assign n177 = ~n136 & ~n176;
  assign n178 = ~n175 & ~n177;
  assign n167 = x5 & n66;
  assign n168 = ~x5 & n68;
  assign n169 = ~x4 & n70;
  assign n170 = ~n168 & ~n169;
  assign n171 = ~n167 & n170;
  assign n163 = x35 ^ x0;
  assign n164 = ~n122 & n163;
  assign n165 = n164 ^ x0;
  assign n166 = x37 & ~n165;
  assign n172 = n171 ^ n166;
  assign n155 = x3 & n103;
  assign n156 = x2 & n105;
  assign n157 = ~n155 & ~n156;
  assign n158 = ~x3 & n96;
  assign n159 = ~x2 & n100;
  assign n160 = ~n158 & ~n159;
  assign n161 = n157 & n160;
  assign n142 = x37 & n122;
  assign n143 = ~x1 & n142;
  assign n144 = x37 ^ x36;
  assign n145 = ~n122 & n144;
  assign n146 = x37 & n145;
  assign n147 = ~x0 & n146;
  assign n148 = ~n143 & ~n147;
  assign n149 = ~x37 & n122;
  assign n150 = x1 & n149;
  assign n151 = ~x37 & n145;
  assign n152 = x0 & n151;
  assign n153 = ~n150 & ~n152;
  assign n154 = n148 & n153;
  assign n162 = n161 ^ n154;
  assign n173 = n172 ^ n162;
  assign n138 = n129 ^ n123;
  assign n139 = n129 ^ n121;
  assign n140 = ~n138 & ~n139;
  assign n141 = n140 ^ n123;
  assign n174 = n173 ^ n141;
  assign n179 = n178 ^ n174;
  assign n210 = n141 & ~n173;
  assign n211 = ~n141 & n173;
  assign n212 = ~n178 & ~n211;
  assign n213 = ~n210 & ~n212;
  assign n204 = x38 ^ x37;
  assign n205 = x0 & n204;
  assign n199 = x6 & n66;
  assign n200 = ~x6 & n68;
  assign n201 = ~x5 & n70;
  assign n202 = ~n200 & ~n201;
  assign n203 = ~n199 & n202;
  assign n206 = n205 ^ n203;
  assign n192 = ~x4 & n96;
  assign n193 = ~x3 & n100;
  assign n194 = ~n192 & ~n193;
  assign n195 = x4 & n103;
  assign n196 = x3 & n105;
  assign n197 = ~n195 & ~n196;
  assign n198 = n194 & n197;
  assign n207 = n206 ^ n198;
  assign n184 = ~x2 & n142;
  assign n185 = ~x1 & n146;
  assign n186 = ~n184 & ~n185;
  assign n187 = x2 & n149;
  assign n188 = x1 & n151;
  assign n189 = ~n187 & ~n188;
  assign n190 = n186 & n189;
  assign n183 = n166 & ~n171;
  assign n191 = n190 ^ n183;
  assign n208 = n207 ^ n191;
  assign n180 = n172 ^ n154;
  assign n181 = n162 & ~n180;
  assign n182 = n181 ^ n161;
  assign n209 = n208 ^ n182;
  assign n214 = n213 ^ n209;
  assign n263 = ~n182 & ~n208;
  assign n264 = n182 & n208;
  assign n265 = ~n213 & ~n264;
  assign n266 = ~n263 & ~n265;
  assign n253 = x3 & n149;
  assign n254 = x2 & n151;
  assign n255 = ~n253 & ~n254;
  assign n256 = ~x3 & n142;
  assign n257 = ~x2 & n146;
  assign n258 = ~n256 & ~n257;
  assign n259 = n255 & n258;
  assign n239 = x39 & n204;
  assign n240 = ~x1 & n239;
  assign n241 = x39 ^ x38;
  assign n242 = ~n204 & n241;
  assign n243 = x39 & n242;
  assign n244 = ~x0 & n243;
  assign n245 = ~n240 & ~n244;
  assign n246 = ~x39 & n204;
  assign n247 = x1 & n246;
  assign n248 = ~x39 & n242;
  assign n249 = x0 & n248;
  assign n250 = ~n247 & ~n249;
  assign n251 = n245 & n250;
  assign n232 = x5 & n103;
  assign n233 = x4 & n105;
  assign n234 = ~n232 & ~n233;
  assign n235 = ~x5 & n96;
  assign n236 = ~x4 & n100;
  assign n237 = ~n235 & ~n236;
  assign n238 = n234 & n237;
  assign n252 = n251 ^ n238;
  assign n260 = n259 ^ n252;
  assign n225 = x7 & n66;
  assign n226 = ~x7 & n68;
  assign n227 = ~x6 & n70;
  assign n228 = ~n226 & ~n227;
  assign n229 = ~n225 & n228;
  assign n221 = x37 ^ x0;
  assign n222 = ~n204 & n221;
  assign n223 = n222 ^ x0;
  assign n224 = x39 & ~n223;
  assign n230 = n229 ^ n224;
  assign n218 = n203 ^ n198;
  assign n219 = ~n206 & ~n218;
  assign n220 = n219 ^ n205;
  assign n231 = n230 ^ n220;
  assign n261 = n260 ^ n231;
  assign n215 = n207 ^ n183;
  assign n216 = ~n191 & ~n215;
  assign n217 = n216 ^ n190;
  assign n262 = n261 ^ n217;
  assign n267 = n266 ^ n262;
  assign n312 = ~n217 & n261;
  assign n313 = n217 & ~n261;
  assign n314 = ~n266 & ~n313;
  assign n315 = ~n312 & ~n314;
  assign n308 = n224 & ~n229;
  assign n300 = ~x6 & n96;
  assign n301 = ~x5 & n100;
  assign n302 = ~n300 & ~n301;
  assign n303 = x6 & n103;
  assign n304 = x5 & n105;
  assign n305 = ~n303 & ~n304;
  assign n306 = n302 & n305;
  assign n293 = ~x4 & n142;
  assign n294 = ~x3 & n146;
  assign n295 = ~n293 & ~n294;
  assign n296 = x4 & n149;
  assign n297 = x3 & n151;
  assign n298 = ~n296 & ~n297;
  assign n299 = n295 & n298;
  assign n307 = n306 ^ n299;
  assign n309 = n308 ^ n307;
  assign n288 = x40 ^ x39;
  assign n289 = x0 & n288;
  assign n283 = x8 & n66;
  assign n284 = ~x8 & n68;
  assign n285 = ~x7 & n70;
  assign n286 = ~n284 & ~n285;
  assign n287 = ~n283 & n286;
  assign n290 = n289 ^ n287;
  assign n276 = ~x2 & n239;
  assign n277 = ~x1 & n243;
  assign n278 = ~n276 & ~n277;
  assign n279 = x2 & n246;
  assign n280 = x1 & n248;
  assign n281 = ~n279 & ~n280;
  assign n282 = n278 & n281;
  assign n291 = n290 ^ n282;
  assign n272 = n259 ^ n251;
  assign n273 = n259 ^ n238;
  assign n274 = n272 & ~n273;
  assign n275 = n274 ^ n251;
  assign n292 = n291 ^ n275;
  assign n310 = n309 ^ n292;
  assign n268 = n260 ^ n230;
  assign n269 = n260 ^ n220;
  assign n270 = n268 & n269;
  assign n271 = n270 ^ n230;
  assign n311 = n310 ^ n271;
  assign n316 = n315 ^ n311;
  assign n378 = ~n271 & ~n310;
  assign n379 = n271 & n310;
  assign n380 = ~n315 & ~n379;
  assign n381 = ~n378 & ~n380;
  assign n367 = x5 & n149;
  assign n368 = x4 & n151;
  assign n369 = ~n367 & ~n368;
  assign n370 = ~x5 & n142;
  assign n371 = ~x4 & n146;
  assign n372 = ~n370 & ~n371;
  assign n373 = n369 & n372;
  assign n362 = x39 ^ x0;
  assign n363 = ~n288 & n362;
  assign n364 = n363 ^ x0;
  assign n365 = x41 & ~n364;
  assign n355 = ~x7 & n96;
  assign n356 = ~x6 & n100;
  assign n357 = ~n355 & ~n356;
  assign n358 = x7 & n103;
  assign n359 = x6 & n105;
  assign n360 = ~n358 & ~n359;
  assign n361 = n357 & n360;
  assign n366 = n365 ^ n361;
  assign n374 = n373 ^ n366;
  assign n352 = n287 ^ n282;
  assign n353 = ~n290 & ~n352;
  assign n354 = n353 ^ n289;
  assign n375 = n374 ^ n354;
  assign n345 = x9 & n66;
  assign n346 = ~x9 & n68;
  assign n347 = ~x8 & n70;
  assign n348 = ~n346 & ~n347;
  assign n349 = ~n345 & n348;
  assign n331 = x41 & n288;
  assign n332 = ~x1 & n331;
  assign n333 = x41 ^ x40;
  assign n334 = ~n288 & n333;
  assign n335 = x41 & n334;
  assign n336 = ~x0 & n335;
  assign n337 = ~n332 & ~n336;
  assign n338 = ~x41 & n288;
  assign n339 = x1 & n338;
  assign n340 = ~x41 & n334;
  assign n341 = x0 & n340;
  assign n342 = ~n339 & ~n341;
  assign n343 = n337 & n342;
  assign n324 = ~x3 & n239;
  assign n325 = ~x2 & n243;
  assign n326 = ~n324 & ~n325;
  assign n327 = x3 & n246;
  assign n328 = x2 & n248;
  assign n329 = ~n327 & ~n328;
  assign n330 = n326 & n329;
  assign n344 = n343 ^ n330;
  assign n350 = n349 ^ n344;
  assign n321 = n308 ^ n299;
  assign n322 = n307 & n321;
  assign n323 = n322 ^ n306;
  assign n351 = n350 ^ n323;
  assign n376 = n375 ^ n351;
  assign n317 = n309 ^ n291;
  assign n318 = n309 ^ n275;
  assign n319 = n317 & n318;
  assign n320 = n319 ^ n291;
  assign n377 = n376 ^ n320;
  assign n382 = n381 ^ n377;
  assign n438 = n320 & n376;
  assign n439 = ~n320 & ~n376;
  assign n440 = ~n381 & ~n439;
  assign n441 = ~n438 & ~n440;
  assign n427 = x4 & n246;
  assign n428 = x3 & n248;
  assign n429 = ~n427 & ~n428;
  assign n430 = ~x4 & n239;
  assign n431 = ~x3 & n243;
  assign n432 = ~n430 & ~n431;
  assign n433 = n429 & n432;
  assign n424 = x42 ^ x41;
  assign n425 = x0 & n424;
  assign n417 = ~x8 & n96;
  assign n418 = ~x7 & n100;
  assign n419 = ~n417 & ~n418;
  assign n420 = x8 & n103;
  assign n421 = x7 & n105;
  assign n422 = ~n420 & ~n421;
  assign n423 = n419 & n422;
  assign n426 = n425 ^ n423;
  assign n434 = n433 ^ n426;
  assign n415 = ~n361 & n365;
  assign n412 = n349 ^ n343;
  assign n413 = ~n344 & n412;
  assign n414 = n413 ^ n349;
  assign n416 = n415 ^ n414;
  assign n435 = n434 ^ n416;
  assign n403 = ~x6 & n142;
  assign n404 = ~x5 & n146;
  assign n405 = ~n403 & ~n404;
  assign n406 = x6 & n149;
  assign n407 = x5 & n151;
  assign n408 = ~n406 & ~n407;
  assign n409 = n405 & n408;
  assign n397 = x10 & n66;
  assign n398 = ~x10 & n68;
  assign n399 = ~x9 & n70;
  assign n400 = ~n398 & ~n399;
  assign n401 = ~n397 & n400;
  assign n390 = ~x2 & n331;
  assign n391 = ~x1 & n335;
  assign n392 = ~n390 & ~n391;
  assign n393 = x2 & n338;
  assign n394 = x1 & n340;
  assign n395 = ~n393 & ~n394;
  assign n396 = n392 & n395;
  assign n402 = n401 ^ n396;
  assign n410 = n409 ^ n402;
  assign n387 = n366 ^ n354;
  assign n388 = n374 & n387;
  assign n389 = n388 ^ n373;
  assign n411 = n410 ^ n389;
  assign n436 = n435 ^ n411;
  assign n383 = n375 ^ n350;
  assign n384 = n375 ^ n323;
  assign n385 = ~n383 & n384;
  assign n386 = n385 ^ n350;
  assign n437 = n436 ^ n386;
  assign n442 = n441 ^ n437;
  assign n516 = ~n386 & ~n436;
  assign n517 = n386 & n436;
  assign n518 = ~n441 & ~n517;
  assign n519 = ~n516 & ~n518;
  assign n504 = ~x7 & n142;
  assign n505 = ~x6 & n146;
  assign n506 = ~n504 & ~n505;
  assign n507 = x7 & n149;
  assign n508 = x6 & n151;
  assign n509 = ~n507 & ~n508;
  assign n510 = n506 & n509;
  assign n491 = ~x43 & n424;
  assign n492 = x1 & n491;
  assign n493 = x43 ^ x42;
  assign n494 = ~n424 & n493;
  assign n495 = ~x43 & n494;
  assign n496 = x0 & n495;
  assign n497 = ~n492 & ~n496;
  assign n498 = x43 & n424;
  assign n499 = ~x1 & n498;
  assign n500 = x43 & n494;
  assign n501 = ~x0 & n500;
  assign n502 = ~n499 & ~n501;
  assign n503 = n497 & n502;
  assign n511 = n510 ^ n503;
  assign n486 = x41 ^ x0;
  assign n487 = ~n424 & n486;
  assign n488 = n487 ^ x0;
  assign n489 = x43 & ~n488;
  assign n479 = x9 & n103;
  assign n480 = x8 & n105;
  assign n481 = ~n479 & ~n480;
  assign n482 = ~x9 & n96;
  assign n483 = ~x8 & n100;
  assign n484 = ~n482 & ~n483;
  assign n485 = n481 & n484;
  assign n490 = n489 ^ n485;
  assign n512 = n511 ^ n490;
  assign n472 = x11 & n66;
  assign n473 = ~x11 & n68;
  assign n474 = ~x10 & n70;
  assign n475 = ~n473 & ~n474;
  assign n476 = ~n472 & n475;
  assign n464 = ~x5 & n239;
  assign n465 = ~x4 & n243;
  assign n466 = ~n464 & ~n465;
  assign n467 = x5 & n246;
  assign n468 = x4 & n248;
  assign n469 = ~n467 & ~n468;
  assign n470 = n466 & n469;
  assign n457 = ~x3 & n331;
  assign n458 = ~x2 & n335;
  assign n459 = ~n457 & ~n458;
  assign n460 = x3 & n338;
  assign n461 = x2 & n340;
  assign n462 = ~n460 & ~n461;
  assign n463 = n459 & n462;
  assign n471 = n470 ^ n463;
  assign n477 = n476 ^ n471;
  assign n453 = n409 ^ n396;
  assign n454 = n402 & ~n453;
  assign n455 = n454 ^ n401;
  assign n450 = n433 ^ n423;
  assign n451 = ~n426 & ~n450;
  assign n452 = n451 ^ n425;
  assign n456 = n455 ^ n452;
  assign n478 = n477 ^ n456;
  assign n513 = n512 ^ n478;
  assign n447 = n434 ^ n415;
  assign n448 = n416 & n447;
  assign n449 = n448 ^ n434;
  assign n514 = n513 ^ n449;
  assign n443 = n435 ^ n410;
  assign n444 = n435 ^ n389;
  assign n445 = n443 & ~n444;
  assign n446 = n445 ^ n410;
  assign n515 = n514 ^ n446;
  assign n520 = n519 ^ n515;
  assign n587 = ~n446 & ~n514;
  assign n588 = n446 & n514;
  assign n589 = ~n519 & ~n588;
  assign n590 = ~n587 & ~n589;
  assign n575 = ~x6 & n239;
  assign n576 = ~x5 & n243;
  assign n577 = ~n575 & ~n576;
  assign n578 = x6 & n246;
  assign n579 = x5 & n248;
  assign n580 = ~n578 & ~n579;
  assign n581 = n577 & n580;
  assign n572 = x44 ^ x43;
  assign n573 = x0 & n572;
  assign n565 = x10 & n103;
  assign n566 = x9 & n105;
  assign n567 = ~n565 & ~n566;
  assign n568 = ~x10 & n96;
  assign n569 = ~x9 & n100;
  assign n570 = ~n568 & ~n569;
  assign n571 = n567 & n570;
  assign n574 = n573 ^ n571;
  assign n582 = n581 ^ n574;
  assign n557 = x2 & n491;
  assign n558 = x1 & n495;
  assign n559 = ~n557 & ~n558;
  assign n560 = ~x2 & n498;
  assign n561 = ~x1 & n500;
  assign n562 = ~n560 & ~n561;
  assign n563 = n559 & n562;
  assign n551 = x12 & n66;
  assign n552 = ~x12 & n68;
  assign n553 = ~x11 & n70;
  assign n554 = ~n552 & ~n553;
  assign n555 = ~n551 & n554;
  assign n544 = ~x4 & n331;
  assign n545 = ~x3 & n335;
  assign n546 = ~n544 & ~n545;
  assign n547 = x4 & n338;
  assign n548 = x3 & n340;
  assign n549 = ~n547 & ~n548;
  assign n550 = n546 & n549;
  assign n556 = n555 ^ n550;
  assign n564 = n563 ^ n556;
  assign n583 = n582 ^ n564;
  assign n541 = n503 ^ n490;
  assign n542 = n511 & ~n541;
  assign n543 = n542 ^ n510;
  assign n584 = n583 ^ n543;
  assign n531 = ~x8 & n142;
  assign n532 = ~x7 & n146;
  assign n533 = ~n531 & ~n532;
  assign n534 = x8 & n149;
  assign n535 = x7 & n151;
  assign n536 = ~n534 & ~n535;
  assign n537 = n533 & n536;
  assign n530 = ~n485 & n489;
  assign n538 = n537 ^ n530;
  assign n527 = n476 ^ n470;
  assign n528 = ~n471 & n527;
  assign n529 = n528 ^ n476;
  assign n539 = n538 ^ n529;
  assign n524 = n477 ^ n455;
  assign n525 = n456 & n524;
  assign n526 = n525 ^ n477;
  assign n540 = n539 ^ n526;
  assign n585 = n584 ^ n540;
  assign n521 = n478 ^ n449;
  assign n522 = ~n513 & ~n521;
  assign n523 = n522 ^ n512;
  assign n586 = n585 ^ n523;
  assign n591 = n590 ^ n586;
  assign n677 = ~n523 & ~n585;
  assign n678 = n523 & n585;
  assign n679 = ~n590 & ~n678;
  assign n680 = ~n677 & ~n679;
  assign n665 = x5 & n338;
  assign n666 = x4 & n340;
  assign n667 = ~n665 & ~n666;
  assign n668 = ~x5 & n331;
  assign n669 = ~x4 & n335;
  assign n670 = ~n668 & ~n669;
  assign n671 = n667 & n670;
  assign n657 = x7 & n246;
  assign n658 = x6 & n248;
  assign n659 = ~n657 & ~n658;
  assign n660 = ~x7 & n239;
  assign n661 = ~x6 & n243;
  assign n662 = ~n660 & ~n661;
  assign n663 = n659 & n662;
  assign n650 = ~x11 & n96;
  assign n651 = ~x10 & n100;
  assign n652 = ~n650 & ~n651;
  assign n653 = x11 & n103;
  assign n654 = x10 & n105;
  assign n655 = ~n653 & ~n654;
  assign n656 = n652 & n655;
  assign n664 = n663 ^ n656;
  assign n672 = n671 ^ n664;
  assign n636 = x45 & n572;
  assign n637 = ~x1 & n636;
  assign n638 = x45 ^ x44;
  assign n639 = ~n572 & n638;
  assign n640 = x45 & n639;
  assign n641 = ~x0 & n640;
  assign n642 = ~n637 & ~n641;
  assign n643 = ~x45 & n572;
  assign n644 = x1 & n643;
  assign n645 = ~x45 & n639;
  assign n646 = x0 & n645;
  assign n647 = ~n644 & ~n646;
  assign n648 = n642 & n647;
  assign n628 = ~x9 & n142;
  assign n629 = ~x8 & n146;
  assign n630 = ~n628 & ~n629;
  assign n631 = x9 & n149;
  assign n632 = x8 & n151;
  assign n633 = ~n631 & ~n632;
  assign n634 = n630 & n633;
  assign n621 = x3 & n491;
  assign n622 = x2 & n495;
  assign n623 = ~n621 & ~n622;
  assign n624 = ~x3 & n498;
  assign n625 = ~x2 & n500;
  assign n626 = ~n624 & ~n625;
  assign n627 = n623 & n626;
  assign n635 = n634 ^ n627;
  assign n649 = n648 ^ n635;
  assign n673 = n672 ^ n649;
  assign n618 = n530 ^ n529;
  assign n619 = ~n538 & n618;
  assign n620 = n619 ^ n537;
  assign n674 = n673 ^ n620;
  assign n609 = x13 & n66;
  assign n610 = ~x13 & n68;
  assign n611 = ~x12 & n70;
  assign n612 = ~n610 & ~n611;
  assign n613 = ~n609 & n612;
  assign n605 = x43 ^ x0;
  assign n606 = ~n572 & n605;
  assign n607 = n606 ^ x0;
  assign n608 = x45 & ~n607;
  assign n614 = n613 ^ n608;
  assign n601 = n581 ^ n573;
  assign n602 = n581 ^ n571;
  assign n603 = ~n601 & ~n602;
  assign n604 = n603 ^ n573;
  assign n615 = n614 ^ n604;
  assign n598 = n563 ^ n550;
  assign n599 = n556 & ~n598;
  assign n600 = n599 ^ n555;
  assign n616 = n615 ^ n600;
  assign n595 = n564 ^ n543;
  assign n596 = ~n583 & ~n595;
  assign n597 = n596 ^ n582;
  assign n617 = n616 ^ n597;
  assign n675 = n674 ^ n617;
  assign n592 = n584 ^ n539;
  assign n593 = n540 & n592;
  assign n594 = n593 ^ n584;
  assign n676 = n675 ^ n594;
  assign n681 = n680 ^ n676;
  assign n760 = n594 & ~n675;
  assign n761 = ~n594 & n675;
  assign n762 = ~n680 & ~n761;
  assign n763 = ~n760 & ~n762;
  assign n752 = x46 ^ x45;
  assign n753 = x0 & n752;
  assign n747 = x14 & n66;
  assign n748 = ~x14 & n68;
  assign n749 = ~x13 & n70;
  assign n750 = ~n748 & ~n749;
  assign n751 = ~n747 & n750;
  assign n754 = n753 ^ n751;
  assign n740 = ~x12 & n96;
  assign n741 = ~x11 & n100;
  assign n742 = ~n740 & ~n741;
  assign n743 = x12 & n103;
  assign n744 = x11 & n105;
  assign n745 = ~n743 & ~n744;
  assign n746 = n742 & n745;
  assign n755 = n754 ^ n746;
  assign n736 = n671 ^ n656;
  assign n737 = n664 & ~n736;
  assign n738 = n737 ^ n663;
  assign n733 = n648 ^ n627;
  assign n734 = n635 & ~n733;
  assign n735 = n734 ^ n634;
  assign n739 = n738 ^ n735;
  assign n756 = n755 ^ n739;
  assign n723 = x10 & n149;
  assign n724 = x9 & n151;
  assign n725 = ~n723 & ~n724;
  assign n726 = ~x10 & n142;
  assign n727 = ~x9 & n146;
  assign n728 = ~n726 & ~n727;
  assign n729 = n725 & n728;
  assign n715 = x8 & n246;
  assign n716 = x7 & n248;
  assign n717 = ~n715 & ~n716;
  assign n718 = ~x8 & n239;
  assign n719 = ~x7 & n243;
  assign n720 = ~n718 & ~n719;
  assign n721 = n717 & n720;
  assign n708 = ~x6 & n331;
  assign n709 = ~x5 & n335;
  assign n710 = ~n708 & ~n709;
  assign n711 = x6 & n338;
  assign n712 = x5 & n340;
  assign n713 = ~n711 & ~n712;
  assign n714 = n710 & n713;
  assign n722 = n721 ^ n714;
  assign n730 = n729 ^ n722;
  assign n706 = n608 & ~n613;
  assign n698 = x4 & n491;
  assign n699 = x3 & n495;
  assign n700 = ~n698 & ~n699;
  assign n701 = ~x4 & n498;
  assign n702 = ~x3 & n500;
  assign n703 = ~n701 & ~n702;
  assign n704 = n700 & n703;
  assign n691 = x2 & n643;
  assign n692 = x1 & n645;
  assign n693 = ~n691 & ~n692;
  assign n694 = ~x2 & n636;
  assign n695 = ~x1 & n640;
  assign n696 = ~n694 & ~n695;
  assign n697 = n693 & n696;
  assign n705 = n704 ^ n697;
  assign n707 = n706 ^ n705;
  assign n731 = n730 ^ n707;
  assign n688 = n604 ^ n600;
  assign n689 = ~n615 & n688;
  assign n690 = n689 ^ n614;
  assign n732 = n731 ^ n690;
  assign n757 = n756 ^ n732;
  assign n685 = n649 ^ n620;
  assign n686 = n673 & ~n685;
  assign n687 = n686 ^ n672;
  assign n758 = n757 ^ n687;
  assign n682 = n674 ^ n597;
  assign n683 = n617 & n682;
  assign n684 = n683 ^ n616;
  assign n759 = n758 ^ n684;
  assign n764 = n763 ^ n759;
  assign n862 = n684 & ~n758;
  assign n863 = ~n684 & n758;
  assign n864 = ~n763 & ~n863;
  assign n865 = ~n862 & ~n864;
  assign n849 = ~x3 & n636;
  assign n850 = ~x2 & n640;
  assign n851 = ~n849 & ~n850;
  assign n852 = x3 & n643;
  assign n853 = x2 & n645;
  assign n854 = ~n852 & ~n853;
  assign n855 = n851 & n854;
  assign n843 = x15 & n66;
  assign n844 = ~x15 & n68;
  assign n845 = ~x14 & n70;
  assign n846 = ~n844 & ~n845;
  assign n847 = ~n843 & n846;
  assign n839 = x45 ^ x0;
  assign n840 = ~n752 & n839;
  assign n841 = n840 ^ x0;
  assign n842 = x47 & ~n841;
  assign n848 = n847 ^ n842;
  assign n856 = n855 ^ n848;
  assign n836 = n751 ^ n746;
  assign n837 = ~n754 & ~n836;
  assign n838 = n837 ^ n753;
  assign n857 = n856 ^ n838;
  assign n833 = n706 ^ n697;
  assign n834 = n705 & n833;
  assign n835 = n834 ^ n704;
  assign n858 = n857 ^ n835;
  assign n830 = n755 ^ n738;
  assign n831 = ~n739 & ~n830;
  assign n832 = n831 ^ n755;
  assign n859 = n858 ^ n832;
  assign n820 = x9 & n246;
  assign n821 = x8 & n248;
  assign n822 = ~n820 & ~n821;
  assign n823 = ~x9 & n239;
  assign n824 = ~x8 & n243;
  assign n825 = ~n823 & ~n824;
  assign n826 = n822 & n825;
  assign n812 = ~x13 & n96;
  assign n813 = ~x12 & n100;
  assign n814 = ~n812 & ~n813;
  assign n815 = x13 & n103;
  assign n816 = x12 & n105;
  assign n817 = ~n815 & ~n816;
  assign n818 = n814 & n817;
  assign n799 = ~x47 & n752;
  assign n800 = x1 & n799;
  assign n801 = x47 ^ x46;
  assign n802 = ~n752 & n801;
  assign n803 = ~x47 & n802;
  assign n804 = x0 & n803;
  assign n805 = ~n800 & ~n804;
  assign n806 = x47 & n752;
  assign n807 = ~x1 & n806;
  assign n808 = x47 & n802;
  assign n809 = ~x0 & n808;
  assign n810 = ~n807 & ~n809;
  assign n811 = n805 & n810;
  assign n819 = n818 ^ n811;
  assign n827 = n826 ^ n819;
  assign n790 = x5 & n491;
  assign n791 = x4 & n495;
  assign n792 = ~n790 & ~n791;
  assign n793 = ~x5 & n498;
  assign n794 = ~x4 & n500;
  assign n795 = ~n793 & ~n794;
  assign n796 = n792 & n795;
  assign n782 = ~x7 & n331;
  assign n783 = ~x6 & n335;
  assign n784 = ~n782 & ~n783;
  assign n785 = x7 & n338;
  assign n786 = x6 & n340;
  assign n787 = ~n785 & ~n786;
  assign n788 = n784 & n787;
  assign n775 = ~x11 & n142;
  assign n776 = ~x10 & n146;
  assign n777 = ~n775 & ~n776;
  assign n778 = x11 & n149;
  assign n779 = x10 & n151;
  assign n780 = ~n778 & ~n779;
  assign n781 = n777 & n780;
  assign n789 = n788 ^ n781;
  assign n797 = n796 ^ n789;
  assign n771 = n729 ^ n721;
  assign n772 = n729 ^ n714;
  assign n773 = n771 & ~n772;
  assign n774 = n773 ^ n721;
  assign n798 = n797 ^ n774;
  assign n828 = n827 ^ n798;
  assign n768 = n707 ^ n690;
  assign n769 = ~n731 & n768;
  assign n770 = n769 ^ n730;
  assign n829 = n828 ^ n770;
  assign n860 = n859 ^ n829;
  assign n765 = n732 ^ n687;
  assign n766 = n757 & n765;
  assign n767 = n766 ^ n756;
  assign n861 = n860 ^ n767;
  assign n866 = n865 ^ n861;
  assign n960 = n767 & ~n860;
  assign n961 = ~n767 & n860;
  assign n962 = ~n865 & ~n961;
  assign n963 = ~n960 & ~n962;
  assign n953 = n842 & ~n847;
  assign n950 = n826 ^ n811;
  assign n951 = n819 & ~n950;
  assign n952 = n951 ^ n818;
  assign n954 = n953 ^ n952;
  assign n946 = n796 ^ n788;
  assign n947 = n796 ^ n781;
  assign n948 = n946 & ~n947;
  assign n949 = n948 ^ n788;
  assign n955 = n954 ^ n949;
  assign n943 = n848 ^ n838;
  assign n944 = n856 & n943;
  assign n945 = n944 ^ n855;
  assign n956 = n955 ^ n945;
  assign n939 = n827 ^ n797;
  assign n940 = n827 ^ n774;
  assign n941 = n939 & ~n940;
  assign n942 = n941 ^ n797;
  assign n957 = n956 ^ n942;
  assign n929 = x8 & n338;
  assign n930 = x7 & n340;
  assign n931 = ~n929 & ~n930;
  assign n932 = ~x8 & n331;
  assign n933 = ~x7 & n335;
  assign n934 = ~n932 & ~n933;
  assign n935 = n931 & n934;
  assign n921 = ~x2 & n806;
  assign n922 = ~x1 & n808;
  assign n923 = ~n921 & ~n922;
  assign n924 = x2 & n799;
  assign n925 = x1 & n803;
  assign n926 = ~n924 & ~n925;
  assign n927 = n923 & n926;
  assign n914 = x10 & n246;
  assign n915 = x9 & n248;
  assign n916 = ~n914 & ~n915;
  assign n917 = ~x10 & n239;
  assign n918 = ~x9 & n243;
  assign n919 = ~n917 & ~n918;
  assign n920 = n916 & n919;
  assign n928 = n927 ^ n920;
  assign n936 = n935 ^ n928;
  assign n909 = x48 ^ x47;
  assign n910 = x0 & n909;
  assign n904 = x16 & n66;
  assign n905 = ~x16 & n68;
  assign n906 = ~x15 & n70;
  assign n907 = ~n905 & ~n906;
  assign n908 = ~n904 & n907;
  assign n911 = n910 ^ n908;
  assign n897 = ~x14 & n96;
  assign n898 = ~x13 & n100;
  assign n899 = ~n897 & ~n898;
  assign n900 = x14 & n103;
  assign n901 = x13 & n105;
  assign n902 = ~n900 & ~n901;
  assign n903 = n899 & n902;
  assign n912 = n911 ^ n903;
  assign n889 = x4 & n643;
  assign n890 = x3 & n645;
  assign n891 = ~n889 & ~n890;
  assign n892 = ~x4 & n636;
  assign n893 = ~x3 & n640;
  assign n894 = ~n892 & ~n893;
  assign n895 = n891 & n894;
  assign n881 = x12 & n149;
  assign n882 = x11 & n151;
  assign n883 = ~n881 & ~n882;
  assign n884 = ~x12 & n142;
  assign n885 = ~x11 & n146;
  assign n886 = ~n884 & ~n885;
  assign n887 = n883 & n886;
  assign n874 = ~x6 & n498;
  assign n875 = ~x5 & n500;
  assign n876 = ~n874 & ~n875;
  assign n877 = x6 & n491;
  assign n878 = x5 & n495;
  assign n879 = ~n877 & ~n878;
  assign n880 = n876 & n879;
  assign n888 = n887 ^ n880;
  assign n896 = n895 ^ n888;
  assign n913 = n912 ^ n896;
  assign n937 = n936 ^ n913;
  assign n871 = n835 ^ n832;
  assign n872 = ~n858 & n871;
  assign n873 = n872 ^ n857;
  assign n938 = n937 ^ n873;
  assign n958 = n957 ^ n938;
  assign n867 = n859 ^ n828;
  assign n868 = n859 ^ n770;
  assign n869 = n867 & ~n868;
  assign n870 = n869 ^ n828;
  assign n959 = n958 ^ n870;
  assign n964 = n963 ^ n959;
  assign n1074 = ~n870 & n958;
  assign n1075 = n870 & ~n958;
  assign n1076 = ~n963 & ~n1075;
  assign n1077 = ~n1074 & ~n1076;
  assign n1065 = n908 ^ n903;
  assign n1066 = ~n911 & ~n1065;
  assign n1067 = n1066 ^ n910;
  assign n1062 = n895 ^ n887;
  assign n1063 = ~n888 & n1062;
  assign n1064 = n1063 ^ n895;
  assign n1068 = n1067 ^ n1064;
  assign n1059 = n935 ^ n920;
  assign n1060 = n928 & ~n1059;
  assign n1061 = n1060 ^ n927;
  assign n1069 = n1068 ^ n1061;
  assign n1056 = n952 ^ n949;
  assign n1057 = ~n954 & ~n1056;
  assign n1058 = n1057 ^ n953;
  assign n1070 = n1069 ^ n1058;
  assign n1053 = n936 ^ n896;
  assign n1054 = ~n913 & ~n1053;
  assign n1055 = n1054 ^ n912;
  assign n1071 = n1070 ^ n1055;
  assign n1044 = x17 & n66;
  assign n1045 = ~x17 & n68;
  assign n1046 = ~x16 & n70;
  assign n1047 = ~n1045 & ~n1046;
  assign n1048 = ~n1044 & n1047;
  assign n1040 = x47 ^ x0;
  assign n1041 = ~n909 & n1040;
  assign n1042 = n1041 ^ x0;
  assign n1043 = x49 & ~n1042;
  assign n1049 = n1048 ^ n1043;
  assign n1032 = x5 & n643;
  assign n1033 = x4 & n645;
  assign n1034 = ~n1032 & ~n1033;
  assign n1035 = ~x5 & n636;
  assign n1036 = ~x4 & n640;
  assign n1037 = ~n1035 & ~n1036;
  assign n1038 = n1034 & n1037;
  assign n1025 = ~x7 & n498;
  assign n1026 = ~x6 & n500;
  assign n1027 = ~n1025 & ~n1026;
  assign n1028 = x7 & n491;
  assign n1029 = x6 & n495;
  assign n1030 = ~n1028 & ~n1029;
  assign n1031 = n1027 & n1030;
  assign n1039 = n1038 ^ n1031;
  assign n1050 = n1049 ^ n1039;
  assign n1016 = ~x13 & n142;
  assign n1017 = ~x12 & n146;
  assign n1018 = ~n1016 & ~n1017;
  assign n1019 = x13 & n149;
  assign n1020 = x12 & n151;
  assign n1021 = ~n1019 & ~n1020;
  assign n1022 = n1018 & n1021;
  assign n1008 = x15 & n103;
  assign n1009 = x14 & n105;
  assign n1010 = ~n1008 & ~n1009;
  assign n1011 = ~x15 & n96;
  assign n1012 = ~x14 & n100;
  assign n1013 = ~n1011 & ~n1012;
  assign n1014 = n1010 & n1013;
  assign n1001 = x9 & n338;
  assign n1002 = x8 & n340;
  assign n1003 = ~n1001 & ~n1002;
  assign n1004 = ~x9 & n331;
  assign n1005 = ~x8 & n335;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = n1003 & n1006;
  assign n1015 = n1014 ^ n1007;
  assign n1023 = n1022 ^ n1015;
  assign n987 = x49 & n909;
  assign n988 = ~x1 & n987;
  assign n989 = x49 ^ x48;
  assign n990 = ~n909 & n989;
  assign n991 = x49 & n990;
  assign n992 = ~x0 & n991;
  assign n993 = ~n988 & ~n992;
  assign n994 = ~x49 & n909;
  assign n995 = x1 & n994;
  assign n996 = ~x49 & n990;
  assign n997 = x0 & n996;
  assign n998 = ~n995 & ~n997;
  assign n999 = n993 & n998;
  assign n979 = ~x3 & n806;
  assign n980 = ~x2 & n808;
  assign n981 = ~n979 & ~n980;
  assign n982 = x3 & n799;
  assign n983 = x2 & n803;
  assign n984 = ~n982 & ~n983;
  assign n985 = n981 & n984;
  assign n972 = ~x11 & n239;
  assign n973 = ~x10 & n243;
  assign n974 = ~n972 & ~n973;
  assign n975 = x11 & n246;
  assign n976 = x10 & n248;
  assign n977 = ~n975 & ~n976;
  assign n978 = n974 & n977;
  assign n986 = n985 ^ n978;
  assign n1000 = n999 ^ n986;
  assign n1024 = n1023 ^ n1000;
  assign n1051 = n1050 ^ n1024;
  assign n969 = n945 ^ n942;
  assign n970 = ~n956 & ~n969;
  assign n971 = n970 ^ n955;
  assign n1052 = n1051 ^ n971;
  assign n1072 = n1071 ^ n1052;
  assign n965 = n957 ^ n937;
  assign n966 = n957 ^ n873;
  assign n967 = n965 & ~n966;
  assign n968 = n967 ^ n937;
  assign n1073 = n1072 ^ n968;
  assign n1078 = n1077 ^ n1073;
  assign n1182 = n968 & ~n1072;
  assign n1183 = ~n968 & n1072;
  assign n1184 = ~n1077 & ~n1183;
  assign n1185 = ~n1182 & ~n1184;
  assign n1174 = x50 ^ x49;
  assign n1175 = x0 & n1174;
  assign n1169 = x18 & n66;
  assign n1170 = ~x18 & n68;
  assign n1171 = ~x17 & n70;
  assign n1172 = ~n1170 & ~n1171;
  assign n1173 = ~n1169 & n1172;
  assign n1176 = n1175 ^ n1173;
  assign n1162 = ~x12 & n239;
  assign n1163 = ~x11 & n243;
  assign n1164 = ~n1162 & ~n1163;
  assign n1165 = x12 & n246;
  assign n1166 = x11 & n248;
  assign n1167 = ~n1165 & ~n1166;
  assign n1168 = n1164 & n1167;
  assign n1177 = n1176 ^ n1168;
  assign n1153 = ~x8 & n498;
  assign n1154 = ~x7 & n500;
  assign n1155 = ~n1153 & ~n1154;
  assign n1156 = x8 & n491;
  assign n1157 = x7 & n495;
  assign n1158 = ~n1156 & ~n1157;
  assign n1159 = n1155 & n1158;
  assign n1145 = ~x10 & n331;
  assign n1146 = ~x9 & n335;
  assign n1147 = ~n1145 & ~n1146;
  assign n1148 = x10 & n338;
  assign n1149 = x9 & n340;
  assign n1150 = ~n1148 & ~n1149;
  assign n1151 = n1147 & n1150;
  assign n1138 = ~x14 & n142;
  assign n1139 = ~x13 & n146;
  assign n1140 = ~n1138 & ~n1139;
  assign n1141 = x14 & n149;
  assign n1142 = x13 & n151;
  assign n1143 = ~n1141 & ~n1142;
  assign n1144 = n1140 & n1143;
  assign n1152 = n1151 ^ n1144;
  assign n1160 = n1159 ^ n1152;
  assign n1135 = n1022 ^ n1007;
  assign n1136 = n1015 & ~n1135;
  assign n1137 = n1136 ^ n1014;
  assign n1161 = n1160 ^ n1137;
  assign n1178 = n1177 ^ n1161;
  assign n1131 = n1050 ^ n1023;
  assign n1132 = ~n1024 & n1131;
  assign n1133 = n1132 ^ n1050;
  assign n1128 = n1064 ^ n1061;
  assign n1129 = ~n1068 & ~n1128;
  assign n1130 = n1129 ^ n1067;
  assign n1134 = n1133 ^ n1130;
  assign n1179 = n1178 ^ n1134;
  assign n1117 = x6 & n643;
  assign n1118 = x5 & n645;
  assign n1119 = ~n1117 & ~n1118;
  assign n1120 = ~x6 & n636;
  assign n1121 = ~x5 & n640;
  assign n1122 = ~n1120 & ~n1121;
  assign n1123 = n1119 & n1122;
  assign n1116 = n1043 & ~n1048;
  assign n1124 = n1123 ^ n1116;
  assign n1113 = n999 ^ n985;
  assign n1114 = ~n986 & n1113;
  assign n1115 = n1114 ^ n999;
  assign n1125 = n1124 ^ n1115;
  assign n1104 = ~x16 & n96;
  assign n1105 = ~x15 & n100;
  assign n1106 = ~n1104 & ~n1105;
  assign n1107 = x16 & n103;
  assign n1108 = x15 & n105;
  assign n1109 = ~n1107 & ~n1108;
  assign n1110 = n1106 & n1109;
  assign n1096 = x4 & n799;
  assign n1097 = x3 & n803;
  assign n1098 = ~n1096 & ~n1097;
  assign n1099 = ~x4 & n806;
  assign n1100 = ~x3 & n808;
  assign n1101 = ~n1099 & ~n1100;
  assign n1102 = n1098 & n1101;
  assign n1089 = x2 & n994;
  assign n1090 = x1 & n996;
  assign n1091 = ~n1089 & ~n1090;
  assign n1092 = ~x2 & n987;
  assign n1093 = ~x1 & n991;
  assign n1094 = ~n1092 & ~n1093;
  assign n1095 = n1091 & n1094;
  assign n1103 = n1102 ^ n1095;
  assign n1111 = n1110 ^ n1103;
  assign n1086 = n1049 ^ n1031;
  assign n1087 = n1039 & ~n1086;
  assign n1088 = n1087 ^ n1038;
  assign n1112 = n1111 ^ n1088;
  assign n1126 = n1125 ^ n1112;
  assign n1083 = n1069 ^ n1055;
  assign n1084 = ~n1070 & n1083;
  assign n1085 = n1084 ^ n1055;
  assign n1127 = n1126 ^ n1085;
  assign n1180 = n1179 ^ n1127;
  assign n1079 = n1071 ^ n1051;
  assign n1080 = n1071 ^ n971;
  assign n1081 = ~n1079 & ~n1080;
  assign n1082 = n1081 ^ n1051;
  assign n1181 = n1180 ^ n1082;
  assign n1186 = n1185 ^ n1181;
  assign n1308 = ~n1082 & ~n1180;
  assign n1309 = n1082 & n1180;
  assign n1310 = ~n1185 & ~n1309;
  assign n1311 = ~n1308 & ~n1310;
  assign n1295 = ~x3 & n987;
  assign n1296 = ~x2 & n991;
  assign n1297 = ~n1295 & ~n1296;
  assign n1298 = x3 & n994;
  assign n1299 = x2 & n996;
  assign n1300 = ~n1298 & ~n1299;
  assign n1301 = n1297 & n1300;
  assign n1287 = x13 & n246;
  assign n1288 = x12 & n248;
  assign n1289 = ~n1287 & ~n1288;
  assign n1290 = ~x13 & n239;
  assign n1291 = ~x12 & n243;
  assign n1292 = ~n1290 & ~n1291;
  assign n1293 = n1289 & n1292;
  assign n1280 = x5 & n799;
  assign n1281 = x4 & n803;
  assign n1282 = ~n1280 & ~n1281;
  assign n1283 = ~x5 & n806;
  assign n1284 = ~x4 & n808;
  assign n1285 = ~n1283 & ~n1284;
  assign n1286 = n1282 & n1285;
  assign n1294 = n1293 ^ n1286;
  assign n1302 = n1301 ^ n1294;
  assign n1271 = ~x7 & n636;
  assign n1272 = ~x6 & n640;
  assign n1273 = ~n1271 & ~n1272;
  assign n1274 = x7 & n643;
  assign n1275 = x6 & n645;
  assign n1276 = ~n1274 & ~n1275;
  assign n1277 = n1273 & n1276;
  assign n1263 = ~x15 & n142;
  assign n1264 = ~x14 & n146;
  assign n1265 = ~n1263 & ~n1264;
  assign n1266 = x15 & n149;
  assign n1267 = x14 & n151;
  assign n1268 = ~n1266 & ~n1267;
  assign n1269 = n1265 & n1268;
  assign n1256 = ~x9 & n498;
  assign n1257 = ~x8 & n500;
  assign n1258 = ~n1256 & ~n1257;
  assign n1259 = x9 & n491;
  assign n1260 = x8 & n495;
  assign n1261 = ~n1259 & ~n1260;
  assign n1262 = n1258 & n1261;
  assign n1270 = n1269 ^ n1262;
  assign n1278 = n1277 ^ n1270;
  assign n1253 = n1159 ^ n1151;
  assign n1254 = ~n1152 & n1253;
  assign n1255 = n1254 ^ n1159;
  assign n1279 = n1278 ^ n1255;
  assign n1303 = n1302 ^ n1279;
  assign n1250 = n1177 ^ n1160;
  assign n1251 = ~n1161 & ~n1250;
  assign n1252 = n1251 ^ n1177;
  assign n1304 = n1303 ^ n1252;
  assign n1247 = n1125 ^ n1088;
  assign n1248 = n1112 & n1247;
  assign n1249 = n1248 ^ n1111;
  assign n1305 = n1304 ^ n1249;
  assign n1237 = x19 & n66;
  assign n1238 = ~x19 & n68;
  assign n1239 = ~x18 & n70;
  assign n1240 = ~n1238 & ~n1239;
  assign n1241 = ~n1237 & n1240;
  assign n1233 = x49 ^ x0;
  assign n1234 = ~n1174 & n1233;
  assign n1235 = n1234 ^ x0;
  assign n1236 = x51 & ~n1235;
  assign n1242 = n1241 ^ n1236;
  assign n1230 = n1173 ^ n1168;
  assign n1231 = ~n1176 & ~n1230;
  assign n1232 = n1231 ^ n1175;
  assign n1243 = n1242 ^ n1232;
  assign n1227 = n1110 ^ n1102;
  assign n1228 = ~n1103 & n1227;
  assign n1229 = n1228 ^ n1110;
  assign n1244 = n1243 ^ n1229;
  assign n1218 = x11 & n338;
  assign n1219 = x10 & n340;
  assign n1220 = ~n1218 & ~n1219;
  assign n1221 = ~x11 & n331;
  assign n1222 = ~x10 & n335;
  assign n1223 = ~n1221 & ~n1222;
  assign n1224 = n1220 & n1223;
  assign n1204 = ~x51 & n1174;
  assign n1205 = x1 & n1204;
  assign n1206 = x51 ^ x50;
  assign n1207 = ~n1174 & n1206;
  assign n1208 = ~x51 & n1207;
  assign n1209 = x0 & n1208;
  assign n1210 = ~n1205 & ~n1209;
  assign n1211 = x51 & n1174;
  assign n1212 = ~x1 & n1211;
  assign n1213 = x51 & n1207;
  assign n1214 = ~x0 & n1213;
  assign n1215 = ~n1212 & ~n1214;
  assign n1216 = n1210 & n1215;
  assign n1197 = x17 & n103;
  assign n1198 = x16 & n105;
  assign n1199 = ~n1197 & ~n1198;
  assign n1200 = ~x17 & n96;
  assign n1201 = ~x16 & n100;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = n1199 & n1202;
  assign n1217 = n1216 ^ n1203;
  assign n1225 = n1224 ^ n1217;
  assign n1194 = n1116 ^ n1115;
  assign n1195 = ~n1124 & n1194;
  assign n1196 = n1195 ^ n1123;
  assign n1226 = n1225 ^ n1196;
  assign n1245 = n1244 ^ n1226;
  assign n1191 = n1178 ^ n1133;
  assign n1192 = n1134 & ~n1191;
  assign n1193 = n1192 ^ n1178;
  assign n1246 = n1245 ^ n1193;
  assign n1306 = n1305 ^ n1246;
  assign n1187 = n1179 ^ n1126;
  assign n1188 = n1179 ^ n1085;
  assign n1189 = ~n1187 & n1188;
  assign n1190 = n1189 ^ n1126;
  assign n1307 = n1306 ^ n1190;
  assign n1312 = n1311 ^ n1307;
  assign n1431 = n1190 & n1306;
  assign n1432 = ~n1190 & ~n1306;
  assign n1433 = ~n1311 & ~n1432;
  assign n1434 = ~n1431 & ~n1433;
  assign n1418 = x16 & n149;
  assign n1419 = x15 & n151;
  assign n1420 = ~n1418 & ~n1419;
  assign n1421 = ~x16 & n142;
  assign n1422 = ~x15 & n146;
  assign n1423 = ~n1421 & ~n1422;
  assign n1424 = n1420 & n1423;
  assign n1410 = ~x2 & n1211;
  assign n1411 = ~x1 & n1213;
  assign n1412 = ~n1410 & ~n1411;
  assign n1413 = x2 & n1204;
  assign n1414 = x1 & n1208;
  assign n1415 = ~n1413 & ~n1414;
  assign n1416 = n1412 & n1415;
  assign n1403 = ~x12 & n331;
  assign n1404 = ~x11 & n335;
  assign n1405 = ~n1403 & ~n1404;
  assign n1406 = x12 & n338;
  assign n1407 = x11 & n340;
  assign n1408 = ~n1406 & ~n1407;
  assign n1409 = n1405 & n1408;
  assign n1417 = n1416 ^ n1409;
  assign n1425 = n1424 ^ n1417;
  assign n1398 = x52 ^ x51;
  assign n1399 = x0 & n1398;
  assign n1393 = x20 & n66;
  assign n1394 = ~x20 & n68;
  assign n1395 = ~x19 & n70;
  assign n1396 = ~n1394 & ~n1395;
  assign n1397 = ~n1393 & n1396;
  assign n1400 = n1399 ^ n1397;
  assign n1386 = ~x14 & n239;
  assign n1387 = ~x13 & n243;
  assign n1388 = ~n1386 & ~n1387;
  assign n1389 = x14 & n246;
  assign n1390 = x13 & n248;
  assign n1391 = ~n1389 & ~n1390;
  assign n1392 = n1388 & n1391;
  assign n1401 = n1400 ^ n1392;
  assign n1378 = ~x18 & n96;
  assign n1379 = ~x17 & n100;
  assign n1380 = ~n1378 & ~n1379;
  assign n1381 = x18 & n103;
  assign n1382 = x17 & n105;
  assign n1383 = ~n1381 & ~n1382;
  assign n1384 = n1380 & n1383;
  assign n1370 = ~x4 & n987;
  assign n1371 = ~x3 & n991;
  assign n1372 = ~n1370 & ~n1371;
  assign n1373 = x4 & n994;
  assign n1374 = x3 & n996;
  assign n1375 = ~n1373 & ~n1374;
  assign n1376 = n1372 & n1375;
  assign n1363 = ~x6 & n806;
  assign n1364 = ~x5 & n808;
  assign n1365 = ~n1363 & ~n1364;
  assign n1366 = x6 & n799;
  assign n1367 = x5 & n803;
  assign n1368 = ~n1366 & ~n1367;
  assign n1369 = n1365 & n1368;
  assign n1377 = n1376 ^ n1369;
  assign n1385 = n1384 ^ n1377;
  assign n1402 = n1401 ^ n1385;
  assign n1426 = n1425 ^ n1402;
  assign n1358 = n1277 ^ n1262;
  assign n1359 = n1270 & ~n1358;
  assign n1360 = n1359 ^ n1269;
  assign n1355 = n1301 ^ n1286;
  assign n1356 = n1294 & ~n1355;
  assign n1357 = n1356 ^ n1293;
  assign n1361 = n1360 ^ n1357;
  assign n1352 = n1224 ^ n1216;
  assign n1353 = ~n1217 & n1352;
  assign n1354 = n1353 ^ n1224;
  assign n1362 = n1361 ^ n1354;
  assign n1427 = n1426 ^ n1362;
  assign n1348 = n1236 & ~n1241;
  assign n1340 = ~x10 & n498;
  assign n1341 = ~x9 & n500;
  assign n1342 = ~n1340 & ~n1341;
  assign n1343 = x10 & n491;
  assign n1344 = x9 & n495;
  assign n1345 = ~n1343 & ~n1344;
  assign n1346 = n1342 & n1345;
  assign n1333 = ~x8 & n636;
  assign n1334 = ~x7 & n640;
  assign n1335 = ~n1333 & ~n1334;
  assign n1336 = x8 & n643;
  assign n1337 = x7 & n645;
  assign n1338 = ~n1336 & ~n1337;
  assign n1339 = n1335 & n1338;
  assign n1347 = n1346 ^ n1339;
  assign n1349 = n1348 ^ n1347;
  assign n1330 = n1232 ^ n1229;
  assign n1331 = ~n1243 & n1330;
  assign n1332 = n1331 ^ n1242;
  assign n1350 = n1349 ^ n1332;
  assign n1326 = n1302 ^ n1278;
  assign n1327 = n1302 ^ n1255;
  assign n1328 = n1326 & ~n1327;
  assign n1329 = n1328 ^ n1278;
  assign n1351 = n1350 ^ n1329;
  assign n1428 = n1427 ^ n1351;
  assign n1321 = n1244 ^ n1225;
  assign n1322 = n1244 ^ n1196;
  assign n1323 = ~n1321 & n1322;
  assign n1324 = n1323 ^ n1225;
  assign n1317 = n1303 ^ n1249;
  assign n1318 = n1252 ^ n1249;
  assign n1319 = n1317 & n1318;
  assign n1320 = n1319 ^ n1303;
  assign n1325 = n1324 ^ n1320;
  assign n1429 = n1428 ^ n1325;
  assign n1313 = n1305 ^ n1245;
  assign n1314 = n1305 ^ n1193;
  assign n1315 = n1313 & ~n1314;
  assign n1316 = n1315 ^ n1245;
  assign n1430 = n1429 ^ n1316;
  assign n1435 = n1434 ^ n1430;
  assign n1570 = n1316 & ~n1429;
  assign n1571 = ~n1316 & n1429;
  assign n1572 = ~n1434 & ~n1571;
  assign n1573 = ~n1570 & ~n1572;
  assign n1549 = x53 & n1398;
  assign n1550 = ~x1 & n1549;
  assign n1551 = x53 ^ x52;
  assign n1552 = ~n1398 & n1551;
  assign n1553 = x53 & n1552;
  assign n1554 = ~x0 & n1553;
  assign n1555 = ~n1550 & ~n1554;
  assign n1556 = ~x53 & n1398;
  assign n1557 = x1 & n1556;
  assign n1558 = ~x53 & n1552;
  assign n1559 = x0 & n1558;
  assign n1560 = ~n1557 & ~n1559;
  assign n1561 = n1555 & n1560;
  assign n1541 = ~x13 & n331;
  assign n1542 = ~x12 & n335;
  assign n1543 = ~n1541 & ~n1542;
  assign n1544 = x13 & n338;
  assign n1545 = x12 & n340;
  assign n1546 = ~n1544 & ~n1545;
  assign n1547 = n1543 & n1546;
  assign n1534 = x3 & n1204;
  assign n1535 = x2 & n1208;
  assign n1536 = ~n1534 & ~n1535;
  assign n1537 = ~x3 & n1211;
  assign n1538 = ~x2 & n1213;
  assign n1539 = ~n1537 & ~n1538;
  assign n1540 = n1536 & n1539;
  assign n1548 = n1547 ^ n1540;
  assign n1562 = n1561 ^ n1548;
  assign n1526 = ~x5 & n987;
  assign n1527 = ~x4 & n991;
  assign n1528 = ~n1526 & ~n1527;
  assign n1529 = x5 & n994;
  assign n1530 = x4 & n996;
  assign n1531 = ~n1529 & ~n1530;
  assign n1532 = n1528 & n1531;
  assign n1518 = x7 & n799;
  assign n1519 = x6 & n803;
  assign n1520 = ~n1518 & ~n1519;
  assign n1521 = ~x7 & n806;
  assign n1522 = ~x6 & n808;
  assign n1523 = ~n1521 & ~n1522;
  assign n1524 = n1520 & n1523;
  assign n1511 = ~x15 & n239;
  assign n1512 = ~x14 & n243;
  assign n1513 = ~n1511 & ~n1512;
  assign n1514 = x15 & n246;
  assign n1515 = x14 & n248;
  assign n1516 = ~n1514 & ~n1515;
  assign n1517 = n1513 & n1516;
  assign n1525 = n1524 ^ n1517;
  assign n1533 = n1532 ^ n1525;
  assign n1563 = n1562 ^ n1533;
  assign n1508 = n1348 ^ n1339;
  assign n1509 = n1347 & n1508;
  assign n1510 = n1509 ^ n1346;
  assign n1564 = n1563 ^ n1510;
  assign n1505 = n1425 ^ n1385;
  assign n1506 = ~n1402 & ~n1505;
  assign n1507 = n1506 ^ n1401;
  assign n1565 = n1564 ^ n1507;
  assign n1495 = ~x11 & n498;
  assign n1496 = ~x10 & n500;
  assign n1497 = ~n1495 & ~n1496;
  assign n1498 = x11 & n491;
  assign n1499 = x10 & n495;
  assign n1500 = ~n1498 & ~n1499;
  assign n1501 = n1497 & n1500;
  assign n1487 = ~x17 & n142;
  assign n1488 = ~x16 & n146;
  assign n1489 = ~n1487 & ~n1488;
  assign n1490 = x17 & n149;
  assign n1491 = x16 & n151;
  assign n1492 = ~n1490 & ~n1491;
  assign n1493 = n1489 & n1492;
  assign n1482 = ~x20 & n70;
  assign n1483 = x33 ^ x21;
  assign n1484 = ~n1482 & n1483;
  assign n1485 = x32 & n1484;
  assign n1486 = n1485 ^ n1482;
  assign n1494 = n1493 ^ n1486;
  assign n1502 = n1501 ^ n1494;
  assign n1478 = n1397 ^ n1392;
  assign n1479 = ~n1400 & ~n1478;
  assign n1480 = n1479 ^ n1399;
  assign n1475 = n1424 ^ n1409;
  assign n1476 = n1417 & ~n1475;
  assign n1477 = n1476 ^ n1416;
  assign n1481 = n1480 ^ n1477;
  assign n1503 = n1502 ^ n1481;
  assign n1465 = x9 & n643;
  assign n1466 = x8 & n645;
  assign n1467 = ~n1465 & ~n1466;
  assign n1468 = ~x9 & n636;
  assign n1469 = ~x8 & n640;
  assign n1470 = ~n1468 & ~n1469;
  assign n1471 = n1467 & n1470;
  assign n1460 = x51 ^ x0;
  assign n1461 = ~n1398 & n1460;
  assign n1462 = n1461 ^ x0;
  assign n1463 = x53 & ~n1462;
  assign n1453 = x19 & n103;
  assign n1454 = x18 & n105;
  assign n1455 = ~n1453 & ~n1454;
  assign n1456 = ~x19 & n96;
  assign n1457 = ~x18 & n100;
  assign n1458 = ~n1456 & ~n1457;
  assign n1459 = n1455 & n1458;
  assign n1464 = n1463 ^ n1459;
  assign n1472 = n1471 ^ n1464;
  assign n1449 = n1384 ^ n1376;
  assign n1450 = n1384 ^ n1369;
  assign n1451 = n1449 & ~n1450;
  assign n1452 = n1451 ^ n1376;
  assign n1473 = n1472 ^ n1452;
  assign n1446 = n1357 ^ n1354;
  assign n1447 = n1361 & ~n1446;
  assign n1448 = n1447 ^ n1360;
  assign n1474 = n1473 ^ n1448;
  assign n1504 = n1503 ^ n1474;
  assign n1566 = n1565 ^ n1504;
  assign n1442 = n1349 ^ n1329;
  assign n1443 = n1332 ^ n1329;
  assign n1444 = ~n1442 & ~n1443;
  assign n1445 = n1444 ^ n1349;
  assign n1567 = n1566 ^ n1445;
  assign n1439 = n1362 ^ n1351;
  assign n1440 = ~n1427 & n1439;
  assign n1441 = n1440 ^ n1426;
  assign n1568 = n1567 ^ n1441;
  assign n1436 = n1428 ^ n1324;
  assign n1437 = ~n1325 & n1436;
  assign n1438 = n1437 ^ n1428;
  assign n1569 = n1568 ^ n1438;
  assign n1574 = n1573 ^ n1569;
  assign n1703 = ~n1438 & n1568;
  assign n1704 = n1438 & ~n1568;
  assign n1705 = ~n1573 & ~n1704;
  assign n1706 = ~n1703 & ~n1705;
  assign n1695 = ~n1459 & n1463;
  assign n1692 = n1501 ^ n1493;
  assign n1693 = ~n1494 & ~n1692;
  assign n1694 = n1693 ^ n1486;
  assign n1696 = n1695 ^ n1694;
  assign n1689 = n1561 ^ n1547;
  assign n1690 = ~n1548 & n1689;
  assign n1691 = n1690 ^ n1561;
  assign n1697 = n1696 ^ n1691;
  assign n1686 = n1502 ^ n1480;
  assign n1687 = n1481 & n1686;
  assign n1688 = n1687 ^ n1502;
  assign n1698 = n1697 ^ n1688;
  assign n1683 = n1533 ^ n1510;
  assign n1684 = n1563 & ~n1683;
  assign n1685 = n1684 ^ n1562;
  assign n1699 = n1698 ^ n1685;
  assign n1672 = x14 & n338;
  assign n1673 = x13 & n340;
  assign n1674 = ~n1672 & ~n1673;
  assign n1675 = ~x14 & n331;
  assign n1676 = ~x13 & n335;
  assign n1677 = ~n1675 & ~n1676;
  assign n1678 = n1674 & n1677;
  assign n1664 = x8 & n799;
  assign n1665 = x7 & n803;
  assign n1666 = ~n1664 & ~n1665;
  assign n1667 = ~x8 & n806;
  assign n1668 = ~x7 & n808;
  assign n1669 = ~n1667 & ~n1668;
  assign n1670 = n1666 & n1669;
  assign n1657 = ~x6 & n987;
  assign n1658 = ~x5 & n991;
  assign n1659 = ~n1657 & ~n1658;
  assign n1660 = x6 & n994;
  assign n1661 = x5 & n996;
  assign n1662 = ~n1660 & ~n1661;
  assign n1663 = n1659 & n1662;
  assign n1671 = n1670 ^ n1663;
  assign n1679 = n1678 ^ n1671;
  assign n1648 = ~x10 & n636;
  assign n1649 = ~x9 & n640;
  assign n1650 = ~n1648 & ~n1649;
  assign n1651 = x10 & n643;
  assign n1652 = x9 & n645;
  assign n1653 = ~n1651 & ~n1652;
  assign n1654 = n1650 & n1653;
  assign n1640 = ~x18 & n142;
  assign n1641 = ~x17 & n146;
  assign n1642 = ~n1640 & ~n1641;
  assign n1643 = x18 & n149;
  assign n1644 = x17 & n151;
  assign n1645 = ~n1643 & ~n1644;
  assign n1646 = n1642 & n1645;
  assign n1633 = ~x12 & n498;
  assign n1634 = ~x11 & n500;
  assign n1635 = ~n1633 & ~n1634;
  assign n1636 = x12 & n491;
  assign n1637 = x11 & n495;
  assign n1638 = ~n1636 & ~n1637;
  assign n1639 = n1635 & n1638;
  assign n1647 = n1646 ^ n1639;
  assign n1655 = n1654 ^ n1647;
  assign n1630 = n1532 ^ n1517;
  assign n1631 = n1525 & ~n1630;
  assign n1632 = n1631 ^ n1524;
  assign n1656 = n1655 ^ n1632;
  assign n1680 = n1679 ^ n1656;
  assign n1620 = ~x16 & n239;
  assign n1621 = ~x15 & n243;
  assign n1622 = ~n1620 & ~n1621;
  assign n1623 = x16 & n246;
  assign n1624 = x15 & n248;
  assign n1625 = ~n1623 & ~n1624;
  assign n1626 = n1622 & n1625;
  assign n1617 = x54 ^ x53;
  assign n1618 = x0 & n1617;
  assign n1610 = x20 & n103;
  assign n1611 = x19 & n105;
  assign n1612 = ~n1610 & ~n1611;
  assign n1613 = ~x20 & n96;
  assign n1614 = ~x19 & n100;
  assign n1615 = ~n1613 & ~n1614;
  assign n1616 = n1612 & n1615;
  assign n1619 = n1618 ^ n1616;
  assign n1627 = n1626 ^ n1619;
  assign n1604 = x22 & n66;
  assign n1605 = ~x22 & n68;
  assign n1606 = ~x21 & n70;
  assign n1607 = ~n1605 & ~n1606;
  assign n1608 = ~n1604 & n1607;
  assign n1596 = x4 & n1204;
  assign n1597 = x3 & n1208;
  assign n1598 = ~n1596 & ~n1597;
  assign n1599 = ~x4 & n1211;
  assign n1600 = ~x3 & n1213;
  assign n1601 = ~n1599 & ~n1600;
  assign n1602 = n1598 & n1601;
  assign n1589 = x2 & n1556;
  assign n1590 = x1 & n1558;
  assign n1591 = ~n1589 & ~n1590;
  assign n1592 = ~x2 & n1549;
  assign n1593 = ~x1 & n1553;
  assign n1594 = ~n1592 & ~n1593;
  assign n1595 = n1591 & n1594;
  assign n1603 = n1602 ^ n1595;
  assign n1609 = n1608 ^ n1603;
  assign n1628 = n1627 ^ n1609;
  assign n1586 = n1464 ^ n1452;
  assign n1587 = n1472 & ~n1586;
  assign n1588 = n1587 ^ n1471;
  assign n1629 = n1628 ^ n1588;
  assign n1681 = n1680 ^ n1629;
  assign n1582 = n1503 ^ n1473;
  assign n1583 = n1503 ^ n1448;
  assign n1584 = n1582 & ~n1583;
  assign n1585 = n1584 ^ n1473;
  assign n1682 = n1681 ^ n1585;
  assign n1700 = n1699 ^ n1682;
  assign n1579 = n1564 ^ n1504;
  assign n1580 = ~n1565 & ~n1579;
  assign n1581 = n1580 ^ n1507;
  assign n1701 = n1700 ^ n1581;
  assign n1575 = n1566 ^ n1441;
  assign n1576 = n1445 ^ n1441;
  assign n1577 = n1575 & ~n1576;
  assign n1578 = n1577 ^ n1566;
  assign n1702 = n1701 ^ n1578;
  assign n1707 = n1706 ^ n1702;
  assign n1854 = n1578 & n1701;
  assign n1855 = ~n1578 & ~n1701;
  assign n1856 = ~n1706 & ~n1855;
  assign n1857 = ~n1854 & ~n1856;
  assign n1841 = ~x3 & n1549;
  assign n1842 = ~x2 & n1553;
  assign n1843 = ~n1841 & ~n1842;
  assign n1844 = x3 & n1556;
  assign n1845 = x2 & n1558;
  assign n1846 = ~n1844 & ~n1845;
  assign n1847 = n1843 & n1846;
  assign n1833 = x15 & n338;
  assign n1834 = x14 & n340;
  assign n1835 = ~n1833 & ~n1834;
  assign n1836 = ~x15 & n331;
  assign n1837 = ~x14 & n335;
  assign n1838 = ~n1836 & ~n1837;
  assign n1839 = n1835 & n1838;
  assign n1826 = x5 & n1204;
  assign n1827 = x4 & n1208;
  assign n1828 = ~n1826 & ~n1827;
  assign n1829 = ~x5 & n1211;
  assign n1830 = ~x4 & n1213;
  assign n1831 = ~n1829 & ~n1830;
  assign n1832 = n1828 & n1831;
  assign n1840 = n1839 ^ n1832;
  assign n1848 = n1847 ^ n1840;
  assign n1811 = x55 & n1617;
  assign n1812 = ~x1 & n1811;
  assign n1813 = x55 ^ x54;
  assign n1814 = ~n1617 & n1813;
  assign n1815 = x55 & n1814;
  assign n1816 = ~x0 & n1815;
  assign n1817 = ~n1812 & ~n1816;
  assign n1818 = ~x55 & n1617;
  assign n1819 = x1 & n1818;
  assign n1820 = ~x55 & n1814;
  assign n1821 = x0 & n1820;
  assign n1822 = ~n1819 & ~n1821;
  assign n1823 = n1817 & n1822;
  assign n1805 = x23 & n66;
  assign n1806 = ~x23 & n68;
  assign n1807 = ~x22 & n70;
  assign n1808 = ~n1806 & ~n1807;
  assign n1809 = ~n1805 & n1808;
  assign n1798 = x19 & n149;
  assign n1799 = x18 & n151;
  assign n1800 = ~n1798 & ~n1799;
  assign n1801 = ~x19 & n142;
  assign n1802 = ~x18 & n146;
  assign n1803 = ~n1801 & ~n1802;
  assign n1804 = n1800 & n1803;
  assign n1810 = n1809 ^ n1804;
  assign n1824 = n1823 ^ n1810;
  assign n1795 = n1678 ^ n1670;
  assign n1796 = ~n1671 & n1795;
  assign n1797 = n1796 ^ n1678;
  assign n1825 = n1824 ^ n1797;
  assign n1849 = n1848 ^ n1825;
  assign n1789 = n1654 ^ n1639;
  assign n1790 = n1647 & ~n1789;
  assign n1791 = n1790 ^ n1646;
  assign n1786 = n1608 ^ n1602;
  assign n1787 = ~n1603 & n1786;
  assign n1788 = n1787 ^ n1608;
  assign n1792 = n1791 ^ n1788;
  assign n1782 = n1626 ^ n1618;
  assign n1783 = n1626 ^ n1616;
  assign n1784 = ~n1782 & ~n1783;
  assign n1785 = n1784 ^ n1618;
  assign n1793 = n1792 ^ n1785;
  assign n1778 = n1679 ^ n1655;
  assign n1779 = n1679 ^ n1632;
  assign n1780 = n1778 & ~n1779;
  assign n1781 = n1780 ^ n1655;
  assign n1794 = n1793 ^ n1781;
  assign n1850 = n1849 ^ n1794;
  assign n1766 = ~x13 & n498;
  assign n1767 = ~x12 & n500;
  assign n1768 = ~n1766 & ~n1767;
  assign n1769 = x13 & n491;
  assign n1770 = x12 & n495;
  assign n1771 = ~n1769 & ~n1770;
  assign n1772 = n1768 & n1771;
  assign n1759 = ~x11 & n636;
  assign n1760 = ~x10 & n640;
  assign n1761 = ~n1759 & ~n1760;
  assign n1762 = x11 & n643;
  assign n1763 = x10 & n645;
  assign n1764 = ~n1762 & ~n1763;
  assign n1765 = n1761 & n1764;
  assign n1773 = n1772 ^ n1765;
  assign n1754 = x53 ^ x0;
  assign n1755 = ~n1617 & n1754;
  assign n1756 = n1755 ^ x0;
  assign n1757 = x55 & ~n1756;
  assign n1747 = ~x21 & n96;
  assign n1748 = ~x20 & n100;
  assign n1749 = ~n1747 & ~n1748;
  assign n1750 = x21 & n103;
  assign n1751 = x20 & n105;
  assign n1752 = ~n1750 & ~n1751;
  assign n1753 = n1749 & n1752;
  assign n1758 = n1757 ^ n1753;
  assign n1774 = n1773 ^ n1758;
  assign n1739 = ~x7 & n987;
  assign n1740 = ~x6 & n991;
  assign n1741 = ~n1739 & ~n1740;
  assign n1742 = x7 & n994;
  assign n1743 = x6 & n996;
  assign n1744 = ~n1742 & ~n1743;
  assign n1745 = n1741 & n1744;
  assign n1731 = ~x17 & n239;
  assign n1732 = ~x16 & n243;
  assign n1733 = ~n1731 & ~n1732;
  assign n1734 = x17 & n246;
  assign n1735 = x16 & n248;
  assign n1736 = ~n1734 & ~n1735;
  assign n1737 = n1733 & n1736;
  assign n1724 = x9 & n799;
  assign n1725 = x8 & n803;
  assign n1726 = ~n1724 & ~n1725;
  assign n1727 = ~x9 & n806;
  assign n1728 = ~x8 & n808;
  assign n1729 = ~n1727 & ~n1728;
  assign n1730 = n1726 & n1729;
  assign n1738 = n1737 ^ n1730;
  assign n1746 = n1745 ^ n1738;
  assign n1775 = n1774 ^ n1746;
  assign n1721 = n1694 ^ n1691;
  assign n1722 = n1696 & n1721;
  assign n1723 = n1722 ^ n1695;
  assign n1776 = n1775 ^ n1723;
  assign n1718 = n1609 ^ n1588;
  assign n1719 = ~n1628 & ~n1718;
  assign n1720 = n1719 ^ n1627;
  assign n1777 = n1776 ^ n1720;
  assign n1851 = n1850 ^ n1777;
  assign n1714 = n1688 ^ n1685;
  assign n1715 = ~n1698 & n1714;
  assign n1716 = n1715 ^ n1697;
  assign n1711 = n1629 ^ n1585;
  assign n1712 = ~n1681 & n1711;
  assign n1713 = n1712 ^ n1680;
  assign n1717 = n1716 ^ n1713;
  assign n1852 = n1851 ^ n1717;
  assign n1708 = n1682 ^ n1581;
  assign n1709 = n1700 & ~n1708;
  assign n1710 = n1709 ^ n1699;
  assign n1853 = n1852 ^ n1710;
  assign n1858 = n1857 ^ n1853;
  assign n1998 = n1710 & n1852;
  assign n1999 = ~n1710 & ~n1852;
  assign n2000 = ~n1857 & ~n1999;
  assign n2001 = ~n1998 & ~n2000;
  assign n1985 = ~x16 & n331;
  assign n1986 = ~x15 & n335;
  assign n1987 = ~n1985 & ~n1986;
  assign n1988 = x16 & n338;
  assign n1989 = x15 & n340;
  assign n1990 = ~n1988 & ~n1989;
  assign n1991 = n1987 & n1990;
  assign n1977 = x8 & n994;
  assign n1978 = x7 & n996;
  assign n1979 = ~n1977 & ~n1978;
  assign n1980 = ~x8 & n987;
  assign n1981 = ~x7 & n991;
  assign n1982 = ~n1980 & ~n1981;
  assign n1983 = n1979 & n1982;
  assign n1970 = x10 & n799;
  assign n1971 = x9 & n803;
  assign n1972 = ~n1970 & ~n1971;
  assign n1973 = ~x10 & n806;
  assign n1974 = ~x9 & n808;
  assign n1975 = ~n1973 & ~n1974;
  assign n1976 = n1972 & n1975;
  assign n1984 = n1983 ^ n1976;
  assign n1992 = n1991 ^ n1984;
  assign n1961 = ~x18 & n239;
  assign n1962 = ~x17 & n243;
  assign n1963 = ~n1961 & ~n1962;
  assign n1964 = x18 & n246;
  assign n1965 = x17 & n248;
  assign n1966 = ~n1964 & ~n1965;
  assign n1967 = n1963 & n1966;
  assign n1958 = x56 ^ x55;
  assign n1959 = x0 & n1958;
  assign n1951 = ~x22 & n96;
  assign n1952 = ~x21 & n100;
  assign n1953 = ~n1951 & ~n1952;
  assign n1954 = x22 & n103;
  assign n1955 = x21 & n105;
  assign n1956 = ~n1954 & ~n1955;
  assign n1957 = n1953 & n1956;
  assign n1960 = n1959 ^ n1957;
  assign n1968 = n1967 ^ n1960;
  assign n1945 = x24 & n66;
  assign n1946 = ~x24 & n68;
  assign n1947 = ~x23 & n70;
  assign n1948 = ~n1946 & ~n1947;
  assign n1949 = ~n1945 & n1948;
  assign n1937 = ~x6 & n1211;
  assign n1938 = ~x5 & n1213;
  assign n1939 = ~n1937 & ~n1938;
  assign n1940 = x6 & n1204;
  assign n1941 = x5 & n1208;
  assign n1942 = ~n1940 & ~n1941;
  assign n1943 = n1939 & n1942;
  assign n1930 = ~x4 & n1549;
  assign n1931 = ~x3 & n1553;
  assign n1932 = ~n1930 & ~n1931;
  assign n1933 = x4 & n1556;
  assign n1934 = x3 & n1558;
  assign n1935 = ~n1933 & ~n1934;
  assign n1936 = n1932 & n1935;
  assign n1944 = n1943 ^ n1936;
  assign n1950 = n1949 ^ n1944;
  assign n1969 = n1968 ^ n1950;
  assign n1993 = n1992 ^ n1969;
  assign n1920 = ~x14 & n498;
  assign n1921 = ~x13 & n500;
  assign n1922 = ~n1920 & ~n1921;
  assign n1923 = x14 & n491;
  assign n1924 = x13 & n495;
  assign n1925 = ~n1923 & ~n1924;
  assign n1926 = n1922 & n1925;
  assign n1912 = ~x2 & n1811;
  assign n1913 = ~x1 & n1815;
  assign n1914 = ~n1912 & ~n1913;
  assign n1915 = x2 & n1818;
  assign n1916 = x1 & n1820;
  assign n1917 = ~n1915 & ~n1916;
  assign n1918 = n1914 & n1917;
  assign n1905 = ~x20 & n142;
  assign n1906 = ~x19 & n146;
  assign n1907 = ~n1905 & ~n1906;
  assign n1908 = x20 & n149;
  assign n1909 = x19 & n151;
  assign n1910 = ~n1908 & ~n1909;
  assign n1911 = n1907 & n1910;
  assign n1919 = n1918 ^ n1911;
  assign n1927 = n1926 ^ n1919;
  assign n1901 = n1823 ^ n1804;
  assign n1902 = n1810 & ~n1901;
  assign n1903 = n1902 ^ n1809;
  assign n1898 = n1745 ^ n1737;
  assign n1899 = ~n1738 & n1898;
  assign n1900 = n1899 ^ n1745;
  assign n1904 = n1903 ^ n1900;
  assign n1928 = n1927 ^ n1904;
  assign n1895 = n1848 ^ n1824;
  assign n1896 = ~n1825 & n1895;
  assign n1897 = n1896 ^ n1848;
  assign n1929 = n1928 ^ n1897;
  assign n1994 = n1993 ^ n1929;
  assign n1883 = ~x12 & n636;
  assign n1884 = ~x11 & n640;
  assign n1885 = ~n1883 & ~n1884;
  assign n1886 = x12 & n643;
  assign n1887 = x11 & n645;
  assign n1888 = ~n1886 & ~n1887;
  assign n1889 = n1885 & n1888;
  assign n1882 = ~n1753 & n1757;
  assign n1890 = n1889 ^ n1882;
  assign n1879 = n1847 ^ n1839;
  assign n1880 = ~n1840 & n1879;
  assign n1881 = n1880 ^ n1847;
  assign n1891 = n1890 ^ n1881;
  assign n1875 = n1765 ^ n1758;
  assign n1876 = n1773 & ~n1875;
  assign n1877 = n1876 ^ n1772;
  assign n1872 = n1791 ^ n1785;
  assign n1873 = ~n1792 & ~n1872;
  assign n1874 = n1873 ^ n1785;
  assign n1878 = n1877 ^ n1874;
  assign n1892 = n1891 ^ n1878;
  assign n1869 = n1746 ^ n1723;
  assign n1870 = n1775 & n1869;
  assign n1871 = n1870 ^ n1774;
  assign n1893 = n1892 ^ n1871;
  assign n1866 = n1849 ^ n1793;
  assign n1867 = n1794 & ~n1866;
  assign n1868 = n1867 ^ n1849;
  assign n1894 = n1893 ^ n1868;
  assign n1995 = n1994 ^ n1894;
  assign n1862 = n1850 ^ n1776;
  assign n1863 = n1850 ^ n1720;
  assign n1864 = n1862 & ~n1863;
  assign n1865 = n1864 ^ n1776;
  assign n1996 = n1995 ^ n1865;
  assign n1859 = n1851 ^ n1716;
  assign n1860 = ~n1717 & ~n1859;
  assign n1861 = n1860 ^ n1851;
  assign n1997 = n1996 ^ n1861;
  assign n2002 = n2001 ^ n1997;
  assign n2163 = n1861 & ~n1996;
  assign n2164 = ~n1861 & n1996;
  assign n2165 = ~n2001 & ~n2164;
  assign n2166 = ~n2163 & ~n2165;
  assign n2149 = ~x13 & n636;
  assign n2150 = ~x12 & n640;
  assign n2151 = ~n2149 & ~n2150;
  assign n2152 = x13 & n643;
  assign n2153 = x12 & n645;
  assign n2154 = ~n2152 & ~n2153;
  assign n2155 = n2151 & n2154;
  assign n2135 = x57 & n1958;
  assign n2136 = ~x1 & n2135;
  assign n2137 = x57 ^ x56;
  assign n2138 = ~n1958 & n2137;
  assign n2139 = x57 & n2138;
  assign n2140 = ~x0 & n2139;
  assign n2141 = ~n2136 & ~n2140;
  assign n2142 = ~x57 & n1958;
  assign n2143 = x1 & n2142;
  assign n2144 = ~x57 & n2138;
  assign n2145 = x0 & n2144;
  assign n2146 = ~n2143 & ~n2145;
  assign n2147 = n2141 & n2146;
  assign n2128 = ~x21 & n142;
  assign n2129 = ~x20 & n146;
  assign n2130 = ~n2128 & ~n2129;
  assign n2131 = x21 & n149;
  assign n2132 = x20 & n151;
  assign n2133 = ~n2131 & ~n2132;
  assign n2134 = n2130 & n2133;
  assign n2148 = n2147 ^ n2134;
  assign n2156 = n2155 ^ n2148;
  assign n2124 = n1967 ^ n1957;
  assign n2125 = ~n1960 & ~n2124;
  assign n2126 = n2125 ^ n1959;
  assign n2120 = n1926 ^ n1918;
  assign n2121 = n1926 ^ n1911;
  assign n2122 = n2120 & ~n2121;
  assign n2123 = n2122 ^ n1918;
  assign n2127 = n2126 ^ n2123;
  assign n2157 = n2156 ^ n2127;
  assign n2117 = n1882 ^ n1881;
  assign n2118 = ~n1890 & n2117;
  assign n2119 = n2118 ^ n1889;
  assign n2158 = n2157 ^ n2119;
  assign n2113 = n1992 ^ n1968;
  assign n2114 = n1992 ^ n1950;
  assign n2115 = ~n2113 & ~n2114;
  assign n2116 = n2115 ^ n1968;
  assign n2159 = n2158 ^ n2116;
  assign n2109 = n1993 ^ n1928;
  assign n2110 = ~n1929 & ~n2109;
  assign n2111 = n2110 ^ n1993;
  assign n2105 = n1891 ^ n1877;
  assign n2106 = n1891 ^ n1874;
  assign n2107 = ~n2105 & ~n2106;
  assign n2108 = n2107 ^ n1877;
  assign n2112 = n2111 ^ n2108;
  assign n2160 = n2159 ^ n2112;
  assign n2094 = x3 & n1818;
  assign n2095 = x2 & n1820;
  assign n2096 = ~n2094 & ~n2095;
  assign n2097 = ~x3 & n1811;
  assign n2098 = ~x2 & n1815;
  assign n2099 = ~n2097 & ~n2098;
  assign n2100 = n2096 & n2099;
  assign n2088 = x25 & n66;
  assign n2089 = ~x25 & n68;
  assign n2090 = ~x24 & n70;
  assign n2091 = ~n2089 & ~n2090;
  assign n2092 = ~n2088 & n2091;
  assign n2081 = x15 & n491;
  assign n2082 = x14 & n495;
  assign n2083 = ~n2081 & ~n2082;
  assign n2084 = ~x15 & n498;
  assign n2085 = ~x14 & n500;
  assign n2086 = ~n2084 & ~n2085;
  assign n2087 = n2083 & n2086;
  assign n2093 = n2092 ^ n2087;
  assign n2101 = n2100 ^ n2093;
  assign n2072 = ~x9 & n987;
  assign n2073 = ~x8 & n991;
  assign n2074 = ~n2072 & ~n2073;
  assign n2075 = x9 & n994;
  assign n2076 = x8 & n996;
  assign n2077 = ~n2075 & ~n2076;
  assign n2078 = n2074 & n2077;
  assign n2064 = ~x19 & n239;
  assign n2065 = ~x18 & n243;
  assign n2066 = ~n2064 & ~n2065;
  assign n2067 = x19 & n246;
  assign n2068 = x18 & n248;
  assign n2069 = ~n2067 & ~n2068;
  assign n2070 = n2066 & n2069;
  assign n2057 = ~x11 & n806;
  assign n2058 = ~x10 & n808;
  assign n2059 = ~n2057 & ~n2058;
  assign n2060 = x11 & n799;
  assign n2061 = x10 & n803;
  assign n2062 = ~n2060 & ~n2061;
  assign n2063 = n2059 & n2062;
  assign n2071 = n2070 ^ n2063;
  assign n2079 = n2078 ^ n2071;
  assign n2049 = x5 & n1556;
  assign n2050 = x4 & n1558;
  assign n2051 = ~n2049 & ~n2050;
  assign n2052 = ~x5 & n1549;
  assign n2053 = ~x4 & n1553;
  assign n2054 = ~n2052 & ~n2053;
  assign n2055 = n2051 & n2054;
  assign n2041 = ~x17 & n331;
  assign n2042 = ~x16 & n335;
  assign n2043 = ~n2041 & ~n2042;
  assign n2044 = x17 & n338;
  assign n2045 = x16 & n340;
  assign n2046 = ~n2044 & ~n2045;
  assign n2047 = n2043 & n2046;
  assign n2034 = x7 & n1204;
  assign n2035 = x6 & n1208;
  assign n2036 = ~n2034 & ~n2035;
  assign n2037 = ~x7 & n1211;
  assign n2038 = ~x6 & n1213;
  assign n2039 = ~n2037 & ~n2038;
  assign n2040 = n2036 & n2039;
  assign n2048 = n2047 ^ n2040;
  assign n2056 = n2055 ^ n2048;
  assign n2080 = n2079 ^ n2056;
  assign n2102 = n2101 ^ n2080;
  assign n2026 = x55 ^ x0;
  assign n2027 = ~n1958 & n2026;
  assign n2028 = n2027 ^ x0;
  assign n2029 = x57 & ~n2028;
  assign n2019 = x23 & n103;
  assign n2020 = x22 & n105;
  assign n2021 = ~n2019 & ~n2020;
  assign n2022 = ~x23 & n96;
  assign n2023 = ~x22 & n100;
  assign n2024 = ~n2022 & ~n2023;
  assign n2025 = n2021 & n2024;
  assign n2030 = n2029 ^ n2025;
  assign n2015 = n1991 ^ n1983;
  assign n2016 = n1991 ^ n1976;
  assign n2017 = n2015 & ~n2016;
  assign n2018 = n2017 ^ n1983;
  assign n2031 = n2030 ^ n2018;
  assign n2012 = n1949 ^ n1943;
  assign n2013 = ~n1944 & n2012;
  assign n2014 = n2013 ^ n1949;
  assign n2032 = n2031 ^ n2014;
  assign n2009 = n1927 ^ n1903;
  assign n2010 = ~n1904 & n2009;
  assign n2011 = n2010 ^ n1927;
  assign n2033 = n2032 ^ n2011;
  assign n2103 = n2102 ^ n2033;
  assign n2006 = n1871 ^ n1868;
  assign n2007 = n1893 & ~n2006;
  assign n2008 = n2007 ^ n1892;
  assign n2104 = n2103 ^ n2008;
  assign n2161 = n2160 ^ n2104;
  assign n2003 = n1894 ^ n1865;
  assign n2004 = ~n1995 & n2003;
  assign n2005 = n2004 ^ n1994;
  assign n2162 = n2161 ^ n2005;
  assign n2167 = n2166 ^ n2162;
  assign n2322 = n2005 & n2161;
  assign n2323 = ~n2005 & ~n2161;
  assign n2324 = ~n2166 & ~n2323;
  assign n2325 = ~n2322 & ~n2324;
  assign n2313 = n2018 ^ n2014;
  assign n2314 = n2031 & ~n2313;
  assign n2315 = n2314 ^ n2030;
  assign n2310 = n2156 ^ n2126;
  assign n2311 = n2127 & ~n2310;
  assign n2312 = n2311 ^ n2156;
  assign n2316 = n2315 ^ n2312;
  assign n2307 = n2101 ^ n2056;
  assign n2308 = n2080 & ~n2307;
  assign n2309 = n2308 ^ n2079;
  assign n2317 = n2316 ^ n2309;
  assign n2303 = n2157 ^ n2116;
  assign n2304 = n2119 ^ n2116;
  assign n2305 = n2303 & n2304;
  assign n2306 = n2305 ^ n2157;
  assign n2318 = n2317 ^ n2306;
  assign n2300 = n2102 ^ n2032;
  assign n2301 = ~n2033 & n2300;
  assign n2302 = n2301 ^ n2102;
  assign n2319 = n2318 ^ n2302;
  assign n2291 = x26 & n66;
  assign n2292 = ~x26 & n68;
  assign n2293 = ~x25 & n70;
  assign n2294 = ~n2292 & ~n2293;
  assign n2295 = ~n2291 & n2294;
  assign n2283 = ~x6 & n1549;
  assign n2284 = ~x5 & n1553;
  assign n2285 = ~n2283 & ~n2284;
  assign n2286 = x6 & n1556;
  assign n2287 = x5 & n1558;
  assign n2288 = ~n2286 & ~n2287;
  assign n2289 = n2285 & n2288;
  assign n2276 = ~x8 & n1211;
  assign n2277 = ~x7 & n1213;
  assign n2278 = ~n2276 & ~n2277;
  assign n2279 = x8 & n1204;
  assign n2280 = x7 & n1208;
  assign n2281 = ~n2279 & ~n2280;
  assign n2282 = n2278 & n2281;
  assign n2290 = n2289 ^ n2282;
  assign n2296 = n2295 ^ n2290;
  assign n2267 = ~x20 & n239;
  assign n2268 = ~x19 & n243;
  assign n2269 = ~n2267 & ~n2268;
  assign n2270 = x20 & n246;
  assign n2271 = x19 & n248;
  assign n2272 = ~n2270 & ~n2271;
  assign n2273 = n2269 & n2272;
  assign n2264 = x58 ^ x57;
  assign n2265 = x0 & n2264;
  assign n2257 = ~x24 & n96;
  assign n2258 = ~x23 & n100;
  assign n2259 = ~n2257 & ~n2258;
  assign n2260 = x24 & n103;
  assign n2261 = x23 & n105;
  assign n2262 = ~n2260 & ~n2261;
  assign n2263 = n2259 & n2262;
  assign n2266 = n2265 ^ n2263;
  assign n2274 = n2273 ^ n2266;
  assign n2254 = n2155 ^ n2134;
  assign n2255 = n2148 & ~n2254;
  assign n2256 = n2255 ^ n2147;
  assign n2275 = n2274 ^ n2256;
  assign n2297 = n2296 ^ n2275;
  assign n2243 = ~x18 & n331;
  assign n2244 = ~x17 & n335;
  assign n2245 = ~n2243 & ~n2244;
  assign n2246 = x18 & n338;
  assign n2247 = x17 & n340;
  assign n2248 = ~n2246 & ~n2247;
  assign n2249 = n2245 & n2248;
  assign n2235 = x10 & n994;
  assign n2236 = x9 & n996;
  assign n2237 = ~n2235 & ~n2236;
  assign n2238 = ~x10 & n987;
  assign n2239 = ~x9 & n991;
  assign n2240 = ~n2238 & ~n2239;
  assign n2241 = n2237 & n2240;
  assign n2228 = x12 & n799;
  assign n2229 = x11 & n803;
  assign n2230 = ~n2228 & ~n2229;
  assign n2231 = ~x12 & n806;
  assign n2232 = ~x11 & n808;
  assign n2233 = ~n2231 & ~n2232;
  assign n2234 = n2230 & n2233;
  assign n2242 = n2241 ^ n2234;
  assign n2250 = n2249 ^ n2242;
  assign n2220 = ~x2 & n2135;
  assign n2221 = ~x1 & n2139;
  assign n2222 = ~n2220 & ~n2221;
  assign n2223 = x2 & n2142;
  assign n2224 = x1 & n2144;
  assign n2225 = ~n2223 & ~n2224;
  assign n2226 = n2222 & n2225;
  assign n2212 = ~x4 & n1811;
  assign n2213 = ~x3 & n1815;
  assign n2214 = ~n2212 & ~n2213;
  assign n2215 = x4 & n1818;
  assign n2216 = x3 & n1820;
  assign n2217 = ~n2215 & ~n2216;
  assign n2218 = n2214 & n2217;
  assign n2205 = ~x16 & n498;
  assign n2206 = ~x15 & n500;
  assign n2207 = ~n2205 & ~n2206;
  assign n2208 = x16 & n491;
  assign n2209 = x15 & n495;
  assign n2210 = ~n2208 & ~n2209;
  assign n2211 = n2207 & n2210;
  assign n2219 = n2218 ^ n2211;
  assign n2227 = n2226 ^ n2219;
  assign n2251 = n2250 ^ n2227;
  assign n2196 = x22 & n149;
  assign n2197 = x21 & n151;
  assign n2198 = ~n2196 & ~n2197;
  assign n2199 = ~x22 & n142;
  assign n2200 = ~x21 & n146;
  assign n2201 = ~n2199 & ~n2200;
  assign n2202 = n2198 & n2201;
  assign n2189 = ~x14 & n636;
  assign n2190 = ~x13 & n640;
  assign n2191 = ~n2189 & ~n2190;
  assign n2192 = x14 & n643;
  assign n2193 = x13 & n645;
  assign n2194 = ~n2192 & ~n2193;
  assign n2195 = n2191 & n2194;
  assign n2203 = n2202 ^ n2195;
  assign n2188 = ~n2025 & n2029;
  assign n2204 = n2203 ^ n2188;
  assign n2252 = n2251 ^ n2204;
  assign n2183 = n2078 ^ n2063;
  assign n2184 = n2071 & ~n2183;
  assign n2185 = n2184 ^ n2070;
  assign n2179 = n2055 ^ n2047;
  assign n2180 = n2055 ^ n2040;
  assign n2181 = n2179 & ~n2180;
  assign n2182 = n2181 ^ n2047;
  assign n2186 = n2185 ^ n2182;
  assign n2175 = n2100 ^ n2092;
  assign n2176 = n2100 ^ n2087;
  assign n2177 = n2175 & ~n2176;
  assign n2178 = n2177 ^ n2092;
  assign n2187 = n2186 ^ n2178;
  assign n2253 = n2252 ^ n2187;
  assign n2298 = n2297 ^ n2253;
  assign n2172 = n2159 ^ n2111;
  assign n2173 = n2112 & ~n2172;
  assign n2174 = n2173 ^ n2159;
  assign n2299 = n2298 ^ n2174;
  assign n2320 = n2319 ^ n2299;
  assign n2168 = n2160 ^ n2103;
  assign n2169 = n2160 ^ n2008;
  assign n2170 = ~n2168 & n2169;
  assign n2171 = n2170 ^ n2103;
  assign n2321 = n2320 ^ n2171;
  assign n2326 = n2325 ^ n2321;
  assign n2498 = ~n2171 & n2320;
  assign n2499 = n2171 & ~n2320;
  assign n2500 = ~n2325 & ~n2499;
  assign n2501 = ~n2498 & ~n2500;
  assign n2488 = n2249 ^ n2241;
  assign n2489 = n2249 ^ n2234;
  assign n2490 = n2488 & ~n2489;
  assign n2491 = n2490 ^ n2241;
  assign n2485 = n2295 ^ n2289;
  assign n2486 = ~n2290 & n2485;
  assign n2487 = n2486 ^ n2295;
  assign n2492 = n2491 ^ n2487;
  assign n2482 = n2226 ^ n2211;
  assign n2483 = n2219 & ~n2482;
  assign n2484 = n2483 ^ n2218;
  assign n2493 = n2492 ^ n2484;
  assign n2478 = n2296 ^ n2274;
  assign n2479 = n2275 & ~n2478;
  assign n2480 = n2479 ^ n2296;
  assign n2475 = n2182 ^ n2178;
  assign n2476 = n2186 & ~n2475;
  assign n2477 = n2476 ^ n2185;
  assign n2481 = n2480 ^ n2477;
  assign n2494 = n2493 ^ n2481;
  assign n2470 = n2297 ^ n2252;
  assign n2471 = n2297 ^ n2187;
  assign n2472 = n2470 & n2471;
  assign n2473 = n2472 ^ n2252;
  assign n2467 = n2315 ^ n2309;
  assign n2468 = ~n2316 & n2467;
  assign n2469 = n2468 ^ n2309;
  assign n2474 = n2473 ^ n2469;
  assign n2495 = n2494 ^ n2474;
  assign n2455 = x15 & n643;
  assign n2456 = x14 & n645;
  assign n2457 = ~n2455 & ~n2456;
  assign n2458 = ~x15 & n636;
  assign n2459 = ~x14 & n640;
  assign n2460 = ~n2458 & ~n2459;
  assign n2461 = n2457 & n2460;
  assign n2450 = x57 ^ x0;
  assign n2451 = ~n2264 & n2450;
  assign n2452 = n2451 ^ x0;
  assign n2453 = x59 & ~n2452;
  assign n2443 = ~x25 & n96;
  assign n2444 = ~x24 & n100;
  assign n2445 = ~n2443 & ~n2444;
  assign n2446 = x25 & n103;
  assign n2447 = x24 & n105;
  assign n2448 = ~n2446 & ~n2447;
  assign n2449 = n2445 & n2448;
  assign n2454 = n2453 ^ n2449;
  assign n2462 = n2461 ^ n2454;
  assign n2440 = n2273 ^ n2263;
  assign n2441 = ~n2266 & ~n2440;
  assign n2442 = n2441 ^ n2265;
  assign n2463 = n2462 ^ n2442;
  assign n2431 = ~x7 & n1549;
  assign n2432 = ~x6 & n1553;
  assign n2433 = ~n2431 & ~n2432;
  assign n2434 = x7 & n1556;
  assign n2435 = x6 & n1558;
  assign n2436 = ~n2434 & ~n2435;
  assign n2437 = n2433 & n2436;
  assign n2423 = x19 & n338;
  assign n2424 = x18 & n340;
  assign n2425 = ~n2423 & ~n2424;
  assign n2426 = ~x19 & n331;
  assign n2427 = ~x18 & n335;
  assign n2428 = ~n2426 & ~n2427;
  assign n2429 = n2425 & n2428;
  assign n2416 = ~x9 & n1211;
  assign n2417 = ~x8 & n1213;
  assign n2418 = ~n2416 & ~n2417;
  assign n2419 = x9 & n1204;
  assign n2420 = x8 & n1208;
  assign n2421 = ~n2419 & ~n2420;
  assign n2422 = n2418 & n2421;
  assign n2430 = n2429 ^ n2422;
  assign n2438 = n2437 ^ n2430;
  assign n2413 = n2195 ^ n2188;
  assign n2414 = n2203 & n2413;
  assign n2415 = n2414 ^ n2202;
  assign n2439 = n2438 ^ n2415;
  assign n2464 = n2463 ^ n2439;
  assign n2403 = ~x5 & n1811;
  assign n2404 = ~x4 & n1815;
  assign n2405 = ~n2403 & ~n2404;
  assign n2406 = x5 & n1818;
  assign n2407 = x4 & n1820;
  assign n2408 = ~n2406 & ~n2407;
  assign n2409 = n2405 & n2408;
  assign n2397 = x27 & n66;
  assign n2398 = ~x27 & n68;
  assign n2399 = ~x26 & n70;
  assign n2400 = ~n2398 & ~n2399;
  assign n2401 = ~n2397 & n2400;
  assign n2390 = ~x17 & n498;
  assign n2391 = ~x16 & n500;
  assign n2392 = ~n2390 & ~n2391;
  assign n2393 = x17 & n491;
  assign n2394 = x16 & n495;
  assign n2395 = ~n2393 & ~n2394;
  assign n2396 = n2392 & n2395;
  assign n2402 = n2401 ^ n2396;
  assign n2410 = n2409 ^ n2402;
  assign n2381 = ~x11 & n987;
  assign n2382 = ~x10 & n991;
  assign n2383 = ~n2381 & ~n2382;
  assign n2384 = x11 & n994;
  assign n2385 = x10 & n996;
  assign n2386 = ~n2384 & ~n2385;
  assign n2387 = n2383 & n2386;
  assign n2373 = x21 & n246;
  assign n2374 = x20 & n248;
  assign n2375 = ~n2373 & ~n2374;
  assign n2376 = ~x21 & n239;
  assign n2377 = ~x20 & n243;
  assign n2378 = ~n2376 & ~n2377;
  assign n2379 = n2375 & n2378;
  assign n2366 = ~x13 & n806;
  assign n2367 = ~x12 & n808;
  assign n2368 = ~n2366 & ~n2367;
  assign n2369 = x13 & n799;
  assign n2370 = x12 & n803;
  assign n2371 = ~n2369 & ~n2370;
  assign n2372 = n2368 & n2371;
  assign n2380 = n2379 ^ n2372;
  assign n2388 = n2387 ^ n2380;
  assign n2352 = ~x59 & n2264;
  assign n2353 = x1 & n2352;
  assign n2354 = x59 ^ x58;
  assign n2355 = ~n2264 & n2354;
  assign n2356 = ~x59 & n2355;
  assign n2357 = x0 & n2356;
  assign n2358 = ~n2353 & ~n2357;
  assign n2359 = x59 & n2264;
  assign n2360 = ~x1 & n2359;
  assign n2361 = x59 & n2355;
  assign n2362 = ~x0 & n2361;
  assign n2363 = ~n2360 & ~n2362;
  assign n2364 = n2358 & n2363;
  assign n2344 = x3 & n2142;
  assign n2345 = x2 & n2144;
  assign n2346 = ~n2344 & ~n2345;
  assign n2347 = ~x3 & n2135;
  assign n2348 = ~x2 & n2139;
  assign n2349 = ~n2347 & ~n2348;
  assign n2350 = n2346 & n2349;
  assign n2337 = x23 & n149;
  assign n2338 = x22 & n151;
  assign n2339 = ~n2337 & ~n2338;
  assign n2340 = ~x23 & n142;
  assign n2341 = ~x22 & n146;
  assign n2342 = ~n2340 & ~n2341;
  assign n2343 = n2339 & n2342;
  assign n2351 = n2350 ^ n2343;
  assign n2365 = n2364 ^ n2351;
  assign n2389 = n2388 ^ n2365;
  assign n2411 = n2410 ^ n2389;
  assign n2334 = n2227 ^ n2204;
  assign n2335 = n2251 & n2334;
  assign n2336 = n2335 ^ n2250;
  assign n2412 = n2411 ^ n2336;
  assign n2465 = n2464 ^ n2412;
  assign n2331 = n2306 ^ n2302;
  assign n2332 = ~n2318 & n2331;
  assign n2333 = n2332 ^ n2317;
  assign n2466 = n2465 ^ n2333;
  assign n2496 = n2495 ^ n2466;
  assign n2327 = n2319 ^ n2298;
  assign n2328 = n2319 ^ n2174;
  assign n2329 = ~n2327 & n2328;
  assign n2330 = n2329 ^ n2298;
  assign n2497 = n2496 ^ n2330;
  assign n2502 = n2501 ^ n2497;
  assign n2668 = ~n2330 & ~n2496;
  assign n2669 = n2330 & n2496;
  assign n2670 = ~n2501 & ~n2669;
  assign n2671 = ~n2668 & ~n2670;
  assign n2653 = ~x20 & n331;
  assign n2654 = ~x19 & n335;
  assign n2655 = ~n2653 & ~n2654;
  assign n2656 = x20 & n338;
  assign n2657 = x19 & n340;
  assign n2658 = ~n2656 & ~n2657;
  assign n2659 = n2655 & n2658;
  assign n2645 = ~x14 & n806;
  assign n2646 = ~x13 & n808;
  assign n2647 = ~n2645 & ~n2646;
  assign n2648 = x14 & n799;
  assign n2649 = x13 & n803;
  assign n2650 = ~n2648 & ~n2649;
  assign n2651 = n2647 & n2650;
  assign n2638 = ~x12 & n987;
  assign n2639 = ~x11 & n991;
  assign n2640 = ~n2638 & ~n2639;
  assign n2641 = x12 & n994;
  assign n2642 = x11 & n996;
  assign n2643 = ~n2641 & ~n2642;
  assign n2644 = n2640 & n2643;
  assign n2652 = n2651 ^ n2644;
  assign n2660 = n2659 ^ n2652;
  assign n2634 = n2409 ^ n2396;
  assign n2635 = n2402 & ~n2634;
  assign n2636 = n2635 ^ n2401;
  assign n2631 = n2364 ^ n2343;
  assign n2632 = n2351 & ~n2631;
  assign n2633 = n2632 ^ n2350;
  assign n2637 = n2636 ^ n2633;
  assign n2661 = n2660 ^ n2637;
  assign n2628 = ~n2449 & n2453;
  assign n2625 = n2387 ^ n2372;
  assign n2626 = n2380 & ~n2625;
  assign n2627 = n2626 ^ n2379;
  assign n2629 = n2628 ^ n2627;
  assign n2622 = n2437 ^ n2422;
  assign n2623 = n2430 & ~n2622;
  assign n2624 = n2623 ^ n2429;
  assign n2630 = n2629 ^ n2624;
  assign n2662 = n2661 ^ n2630;
  assign n2619 = n2410 ^ n2388;
  assign n2620 = ~n2389 & n2619;
  assign n2621 = n2620 ^ n2410;
  assign n2663 = n2662 ^ n2621;
  assign n2609 = ~x4 & n2135;
  assign n2610 = ~x3 & n2139;
  assign n2611 = ~n2609 & ~n2610;
  assign n2612 = x4 & n2142;
  assign n2613 = x3 & n2144;
  assign n2614 = ~n2612 & ~n2613;
  assign n2615 = n2611 & n2614;
  assign n2601 = x18 & n491;
  assign n2602 = x17 & n495;
  assign n2603 = ~n2601 & ~n2602;
  assign n2604 = ~x18 & n498;
  assign n2605 = ~x17 & n500;
  assign n2606 = ~n2604 & ~n2605;
  assign n2607 = n2603 & n2606;
  assign n2594 = ~x6 & n1811;
  assign n2595 = ~x5 & n1815;
  assign n2596 = ~n2594 & ~n2595;
  assign n2597 = x6 & n1818;
  assign n2598 = x5 & n1820;
  assign n2599 = ~n2597 & ~n2598;
  assign n2600 = n2596 & n2599;
  assign n2608 = n2607 ^ n2600;
  assign n2616 = n2615 ^ n2608;
  assign n2591 = n2491 ^ n2484;
  assign n2592 = ~n2492 & n2591;
  assign n2593 = n2592 ^ n2484;
  assign n2617 = n2616 ^ n2593;
  assign n2588 = n2454 ^ n2442;
  assign n2589 = n2462 & n2588;
  assign n2590 = n2589 ^ n2461;
  assign n2618 = n2617 ^ n2590;
  assign n2664 = n2663 ^ n2618;
  assign n2584 = n2464 ^ n2411;
  assign n2585 = n2464 ^ n2336;
  assign n2586 = ~n2584 & n2585;
  assign n2587 = n2586 ^ n2411;
  assign n2665 = n2664 ^ n2587;
  assign n2574 = x28 & n66;
  assign n2575 = ~x28 & n68;
  assign n2576 = ~x27 & n70;
  assign n2577 = ~n2575 & ~n2576;
  assign n2578 = ~n2574 & n2577;
  assign n2566 = x10 & n1204;
  assign n2567 = x9 & n1208;
  assign n2568 = ~n2566 & ~n2567;
  assign n2569 = ~x10 & n1211;
  assign n2570 = ~x9 & n1213;
  assign n2571 = ~n2569 & ~n2570;
  assign n2572 = n2568 & n2571;
  assign n2559 = x8 & n1556;
  assign n2560 = x7 & n1558;
  assign n2561 = ~n2559 & ~n2560;
  assign n2562 = ~x8 & n1549;
  assign n2563 = ~x7 & n1553;
  assign n2564 = ~n2562 & ~n2563;
  assign n2565 = n2561 & n2564;
  assign n2573 = n2572 ^ n2565;
  assign n2579 = n2578 ^ n2573;
  assign n2550 = x22 & n246;
  assign n2551 = x21 & n248;
  assign n2552 = ~n2550 & ~n2551;
  assign n2553 = ~x22 & n239;
  assign n2554 = ~x21 & n243;
  assign n2555 = ~n2553 & ~n2554;
  assign n2556 = n2552 & n2555;
  assign n2547 = x60 ^ x59;
  assign n2548 = x0 & n2547;
  assign n2540 = ~x26 & n96;
  assign n2541 = ~x25 & n100;
  assign n2542 = ~n2540 & ~n2541;
  assign n2543 = x26 & n103;
  assign n2544 = x25 & n105;
  assign n2545 = ~n2543 & ~n2544;
  assign n2546 = n2542 & n2545;
  assign n2549 = n2548 ^ n2546;
  assign n2557 = n2556 ^ n2549;
  assign n2532 = ~x16 & n636;
  assign n2533 = ~x15 & n640;
  assign n2534 = ~n2532 & ~n2533;
  assign n2535 = x16 & n643;
  assign n2536 = x15 & n645;
  assign n2537 = ~n2535 & ~n2536;
  assign n2538 = n2534 & n2537;
  assign n2524 = x24 & n149;
  assign n2525 = x23 & n151;
  assign n2526 = ~n2524 & ~n2525;
  assign n2527 = ~x24 & n142;
  assign n2528 = ~x23 & n146;
  assign n2529 = ~n2527 & ~n2528;
  assign n2530 = n2526 & n2529;
  assign n2517 = ~x2 & n2359;
  assign n2518 = ~x1 & n2361;
  assign n2519 = ~n2517 & ~n2518;
  assign n2520 = x2 & n2352;
  assign n2521 = x1 & n2356;
  assign n2522 = ~n2520 & ~n2521;
  assign n2523 = n2519 & n2522;
  assign n2531 = n2530 ^ n2523;
  assign n2539 = n2538 ^ n2531;
  assign n2558 = n2557 ^ n2539;
  assign n2580 = n2579 ^ n2558;
  assign n2514 = n2463 ^ n2415;
  assign n2515 = n2439 & n2514;
  assign n2516 = n2515 ^ n2438;
  assign n2581 = n2580 ^ n2516;
  assign n2511 = n2493 ^ n2480;
  assign n2512 = ~n2481 & n2511;
  assign n2513 = n2512 ^ n2493;
  assign n2582 = n2581 ^ n2513;
  assign n2507 = n2494 ^ n2473;
  assign n2508 = n2494 ^ n2469;
  assign n2509 = ~n2507 & ~n2508;
  assign n2510 = n2509 ^ n2473;
  assign n2583 = n2582 ^ n2510;
  assign n2666 = n2665 ^ n2583;
  assign n2503 = n2495 ^ n2465;
  assign n2504 = n2495 ^ n2333;
  assign n2505 = n2503 & n2504;
  assign n2506 = n2505 ^ n2465;
  assign n2667 = n2666 ^ n2506;
  assign n2672 = n2671 ^ n2667;
  assign n2856 = n2506 & n2666;
  assign n2857 = ~n2506 & ~n2666;
  assign n2858 = ~n2671 & ~n2857;
  assign n2859 = ~n2856 & ~n2858;
  assign n2842 = ~x15 & n806;
  assign n2843 = ~x14 & n808;
  assign n2844 = ~n2842 & ~n2843;
  assign n2845 = x15 & n799;
  assign n2846 = x14 & n803;
  assign n2847 = ~n2845 & ~n2846;
  assign n2848 = n2844 & n2847;
  assign n2834 = x27 & n103;
  assign n2835 = x26 & n105;
  assign n2836 = ~n2834 & ~n2835;
  assign n2837 = ~x27 & n96;
  assign n2838 = ~x26 & n100;
  assign n2839 = ~n2837 & ~n2838;
  assign n2840 = n2836 & n2839;
  assign n2827 = ~x23 & n239;
  assign n2828 = ~x22 & n243;
  assign n2829 = ~n2827 & ~n2828;
  assign n2830 = x23 & n246;
  assign n2831 = x22 & n248;
  assign n2832 = ~n2830 & ~n2831;
  assign n2833 = n2829 & n2832;
  assign n2841 = n2840 ^ n2833;
  assign n2849 = n2848 ^ n2841;
  assign n2823 = n2615 ^ n2607;
  assign n2824 = ~n2608 & n2823;
  assign n2825 = n2824 ^ n2615;
  assign n2820 = n2538 ^ n2530;
  assign n2821 = ~n2531 & n2820;
  assign n2822 = n2821 ^ n2538;
  assign n2826 = n2825 ^ n2822;
  assign n2850 = n2849 ^ n2826;
  assign n2813 = n2556 ^ n2548;
  assign n2814 = n2556 ^ n2546;
  assign n2815 = ~n2813 & ~n2814;
  assign n2816 = n2815 ^ n2548;
  assign n2810 = n2578 ^ n2572;
  assign n2811 = ~n2573 & n2810;
  assign n2812 = n2811 ^ n2578;
  assign n2817 = n2816 ^ n2812;
  assign n2807 = n2659 ^ n2644;
  assign n2808 = n2652 & ~n2807;
  assign n2809 = n2808 ^ n2651;
  assign n2818 = n2817 ^ n2809;
  assign n2804 = n2660 ^ n2636;
  assign n2805 = ~n2637 & n2804;
  assign n2806 = n2805 ^ n2660;
  assign n2819 = n2818 ^ n2806;
  assign n2851 = n2850 ^ n2819;
  assign n2795 = x29 & n66;
  assign n2796 = ~x29 & n68;
  assign n2797 = ~x28 & n70;
  assign n2798 = ~n2796 & ~n2797;
  assign n2799 = ~n2795 & n2798;
  assign n2791 = x59 ^ x0;
  assign n2792 = ~n2547 & n2791;
  assign n2793 = n2792 ^ x0;
  assign n2794 = x61 & ~n2793;
  assign n2800 = n2799 ^ n2794;
  assign n2783 = x3 & n2352;
  assign n2784 = x2 & n2356;
  assign n2785 = ~n2783 & ~n2784;
  assign n2786 = ~x3 & n2359;
  assign n2787 = ~x2 & n2361;
  assign n2788 = ~n2786 & ~n2787;
  assign n2789 = n2785 & n2788;
  assign n2770 = x61 & n2547;
  assign n2771 = ~x1 & n2770;
  assign n2772 = x61 ^ x60;
  assign n2773 = ~n2547 & n2772;
  assign n2774 = x61 & n2773;
  assign n2775 = ~x0 & n2774;
  assign n2776 = ~n2771 & ~n2775;
  assign n2777 = ~x61 & n2547;
  assign n2778 = x1 & n2777;
  assign n2779 = ~x61 & n2773;
  assign n2780 = x0 & n2779;
  assign n2781 = ~n2778 & ~n2780;
  assign n2782 = n2776 & n2781;
  assign n2790 = n2789 ^ n2782;
  assign n2801 = n2800 ^ n2790;
  assign n2767 = n2627 ^ n2624;
  assign n2768 = ~n2629 & ~n2767;
  assign n2769 = n2768 ^ n2628;
  assign n2802 = n2801 ^ n2769;
  assign n2763 = n2579 ^ n2557;
  assign n2764 = n2579 ^ n2539;
  assign n2765 = ~n2763 & ~n2764;
  assign n2766 = n2765 ^ n2557;
  assign n2803 = n2802 ^ n2766;
  assign n2852 = n2851 ^ n2803;
  assign n2752 = ~x19 & n498;
  assign n2753 = ~x18 & n500;
  assign n2754 = ~n2752 & ~n2753;
  assign n2755 = x19 & n491;
  assign n2756 = x18 & n495;
  assign n2757 = ~n2755 & ~n2756;
  assign n2758 = n2754 & n2757;
  assign n2744 = ~x9 & n1549;
  assign n2745 = ~x8 & n1553;
  assign n2746 = ~n2744 & ~n2745;
  assign n2747 = x9 & n1556;
  assign n2748 = x8 & n1558;
  assign n2749 = ~n2747 & ~n2748;
  assign n2750 = n2746 & n2749;
  assign n2737 = x25 & n149;
  assign n2738 = x24 & n151;
  assign n2739 = ~n2737 & ~n2738;
  assign n2740 = ~x25 & n142;
  assign n2741 = ~x24 & n146;
  assign n2742 = ~n2740 & ~n2741;
  assign n2743 = n2739 & n2742;
  assign n2751 = n2750 ^ n2743;
  assign n2759 = n2758 ^ n2751;
  assign n2728 = ~x17 & n636;
  assign n2729 = ~x16 & n640;
  assign n2730 = ~n2728 & ~n2729;
  assign n2731 = x17 & n643;
  assign n2732 = x16 & n645;
  assign n2733 = ~n2731 & ~n2732;
  assign n2734 = n2730 & n2733;
  assign n2720 = ~x7 & n1811;
  assign n2721 = ~x6 & n1815;
  assign n2722 = ~n2720 & ~n2721;
  assign n2723 = x7 & n1818;
  assign n2724 = x6 & n1820;
  assign n2725 = ~n2723 & ~n2724;
  assign n2726 = n2722 & n2725;
  assign n2713 = ~x5 & n2135;
  assign n2714 = ~x4 & n2139;
  assign n2715 = ~n2713 & ~n2714;
  assign n2716 = x5 & n2142;
  assign n2717 = x4 & n2144;
  assign n2718 = ~n2716 & ~n2717;
  assign n2719 = n2715 & n2718;
  assign n2727 = n2726 ^ n2719;
  assign n2735 = n2734 ^ n2727;
  assign n2705 = x11 & n1204;
  assign n2706 = x10 & n1208;
  assign n2707 = ~n2705 & ~n2706;
  assign n2708 = ~x11 & n1211;
  assign n2709 = ~x10 & n1213;
  assign n2710 = ~n2708 & ~n2709;
  assign n2711 = n2707 & n2710;
  assign n2697 = ~x13 & n987;
  assign n2698 = ~x12 & n991;
  assign n2699 = ~n2697 & ~n2698;
  assign n2700 = x13 & n994;
  assign n2701 = x12 & n996;
  assign n2702 = ~n2700 & ~n2701;
  assign n2703 = n2699 & n2702;
  assign n2690 = ~x21 & n331;
  assign n2691 = ~x20 & n335;
  assign n2692 = ~n2690 & ~n2691;
  assign n2693 = x21 & n338;
  assign n2694 = x20 & n340;
  assign n2695 = ~n2693 & ~n2694;
  assign n2696 = n2692 & n2695;
  assign n2704 = n2703 ^ n2696;
  assign n2712 = n2711 ^ n2704;
  assign n2736 = n2735 ^ n2712;
  assign n2760 = n2759 ^ n2736;
  assign n2686 = n2616 ^ n2590;
  assign n2687 = n2593 ^ n2590;
  assign n2688 = n2686 & ~n2687;
  assign n2689 = n2688 ^ n2616;
  assign n2761 = n2760 ^ n2689;
  assign n2683 = n2661 ^ n2621;
  assign n2684 = n2662 & n2683;
  assign n2685 = n2684 ^ n2621;
  assign n2762 = n2761 ^ n2685;
  assign n2853 = n2852 ^ n2762;
  assign n2679 = n2618 ^ n2587;
  assign n2680 = ~n2664 & ~n2679;
  assign n2681 = n2680 ^ n2663;
  assign n2676 = n2516 ^ n2513;
  assign n2677 = ~n2581 & ~n2676;
  assign n2678 = n2677 ^ n2580;
  assign n2682 = n2681 ^ n2678;
  assign n2854 = n2853 ^ n2682;
  assign n2673 = n2665 ^ n2582;
  assign n2674 = ~n2583 & n2673;
  assign n2675 = n2674 ^ n2665;
  assign n2855 = n2854 ^ n2675;
  assign n2860 = n2859 ^ n2855;
  assign n3037 = n2675 & n2854;
  assign n3038 = ~n2675 & ~n2854;
  assign n3039 = ~n2859 & ~n3038;
  assign n3040 = ~n3037 & ~n3039;
  assign n3023 = x8 & n1818;
  assign n3024 = x7 & n1820;
  assign n3025 = ~n3023 & ~n3024;
  assign n3026 = ~x8 & n1811;
  assign n3027 = ~x7 & n1815;
  assign n3028 = ~n3026 & ~n3027;
  assign n3029 = n3025 & n3028;
  assign n3015 = ~x26 & n142;
  assign n3016 = ~x25 & n146;
  assign n3017 = ~n3015 & ~n3016;
  assign n3018 = x26 & n149;
  assign n3019 = x25 & n151;
  assign n3020 = ~n3018 & ~n3019;
  assign n3021 = n3017 & n3020;
  assign n3008 = ~x20 & n498;
  assign n3009 = ~x19 & n500;
  assign n3010 = ~n3008 & ~n3009;
  assign n3011 = x20 & n491;
  assign n3012 = x19 & n495;
  assign n3013 = ~n3011 & ~n3012;
  assign n3014 = n3010 & n3013;
  assign n3022 = n3021 ^ n3014;
  assign n3030 = n3029 ^ n3022;
  assign n3003 = x62 ^ x61;
  assign n3004 = x0 & n3003;
  assign n2998 = x30 & n66;
  assign n2999 = ~x30 & n68;
  assign n3000 = ~x29 & n70;
  assign n3001 = ~n2999 & ~n3000;
  assign n3002 = ~n2998 & n3001;
  assign n3005 = n3004 ^ n3002;
  assign n2991 = ~x28 & n96;
  assign n2992 = ~x27 & n100;
  assign n2993 = ~n2991 & ~n2992;
  assign n2994 = x28 & n103;
  assign n2995 = x27 & n105;
  assign n2996 = ~n2994 & ~n2995;
  assign n2997 = n2993 & n2996;
  assign n3006 = n3005 ^ n2997;
  assign n2983 = x4 & n2352;
  assign n2984 = x3 & n2356;
  assign n2985 = ~n2983 & ~n2984;
  assign n2986 = ~x4 & n2359;
  assign n2987 = ~x3 & n2361;
  assign n2988 = ~n2986 & ~n2987;
  assign n2989 = n2985 & n2988;
  assign n2975 = ~x6 & n2135;
  assign n2976 = ~x5 & n2139;
  assign n2977 = ~n2975 & ~n2976;
  assign n2978 = x6 & n2142;
  assign n2979 = x5 & n2144;
  assign n2980 = ~n2978 & ~n2979;
  assign n2981 = n2977 & n2980;
  assign n2968 = ~x18 & n636;
  assign n2969 = ~x17 & n640;
  assign n2970 = ~n2968 & ~n2969;
  assign n2971 = x18 & n643;
  assign n2972 = x17 & n645;
  assign n2973 = ~n2971 & ~n2972;
  assign n2974 = n2970 & n2973;
  assign n2982 = n2981 ^ n2974;
  assign n2990 = n2989 ^ n2982;
  assign n3007 = n3006 ^ n2990;
  assign n3031 = n3030 ^ n3007;
  assign n2965 = n2850 ^ n2818;
  assign n2966 = n2819 & ~n2965;
  assign n2967 = n2966 ^ n2850;
  assign n3032 = n3031 ^ n2967;
  assign n2961 = n2801 ^ n2766;
  assign n2962 = n2769 ^ n2766;
  assign n2963 = ~n2961 & ~n2962;
  assign n2964 = n2963 ^ n2801;
  assign n3033 = n3032 ^ n2964;
  assign n2948 = ~x14 & n987;
  assign n2949 = ~x13 & n991;
  assign n2950 = ~n2948 & ~n2949;
  assign n2951 = x14 & n994;
  assign n2952 = x13 & n996;
  assign n2953 = ~n2951 & ~n2952;
  assign n2954 = n2950 & n2953;
  assign n2940 = x24 & n246;
  assign n2941 = x23 & n248;
  assign n2942 = ~n2940 & ~n2941;
  assign n2943 = ~x24 & n239;
  assign n2944 = ~x23 & n243;
  assign n2945 = ~n2943 & ~n2944;
  assign n2946 = n2942 & n2945;
  assign n2933 = ~x16 & n806;
  assign n2934 = ~x15 & n808;
  assign n2935 = ~n2933 & ~n2934;
  assign n2936 = x16 & n799;
  assign n2937 = x15 & n803;
  assign n2938 = ~n2936 & ~n2937;
  assign n2939 = n2935 & n2938;
  assign n2947 = n2946 ^ n2939;
  assign n2955 = n2954 ^ n2947;
  assign n2925 = ~x10 & n1549;
  assign n2926 = ~x9 & n1553;
  assign n2927 = ~n2925 & ~n2926;
  assign n2928 = x10 & n1556;
  assign n2929 = x9 & n1558;
  assign n2930 = ~n2928 & ~n2929;
  assign n2931 = n2927 & n2930;
  assign n2917 = ~x22 & n331;
  assign n2918 = ~x21 & n335;
  assign n2919 = ~n2917 & ~n2918;
  assign n2920 = x22 & n338;
  assign n2921 = x21 & n340;
  assign n2922 = ~n2920 & ~n2921;
  assign n2923 = n2919 & n2922;
  assign n2910 = ~x12 & n1211;
  assign n2911 = ~x11 & n1213;
  assign n2912 = ~n2910 & ~n2911;
  assign n2913 = x12 & n1204;
  assign n2914 = x11 & n1208;
  assign n2915 = ~n2913 & ~n2914;
  assign n2916 = n2912 & n2915;
  assign n2924 = n2923 ^ n2916;
  assign n2932 = n2931 ^ n2924;
  assign n2956 = n2955 ^ n2932;
  assign n2907 = n2800 ^ n2782;
  assign n2908 = n2790 & ~n2907;
  assign n2909 = n2908 ^ n2789;
  assign n2957 = n2956 ^ n2909;
  assign n2901 = n2758 ^ n2743;
  assign n2902 = n2751 & ~n2901;
  assign n2903 = n2902 ^ n2750;
  assign n2898 = n2711 ^ n2696;
  assign n2899 = n2704 & ~n2898;
  assign n2900 = n2899 ^ n2703;
  assign n2904 = n2903 ^ n2900;
  assign n2895 = n2734 ^ n2719;
  assign n2896 = n2727 & ~n2895;
  assign n2897 = n2896 ^ n2726;
  assign n2905 = n2904 ^ n2897;
  assign n2892 = n2849 ^ n2825;
  assign n2893 = ~n2826 & n2892;
  assign n2894 = n2893 ^ n2849;
  assign n2906 = n2905 ^ n2894;
  assign n2958 = n2957 ^ n2906;
  assign n2881 = ~x2 & n2770;
  assign n2882 = ~x1 & n2774;
  assign n2883 = ~n2881 & ~n2882;
  assign n2884 = x2 & n2777;
  assign n2885 = x1 & n2779;
  assign n2886 = ~n2884 & ~n2885;
  assign n2887 = n2883 & n2886;
  assign n2880 = n2794 & ~n2799;
  assign n2888 = n2887 ^ n2880;
  assign n2877 = n2848 ^ n2833;
  assign n2878 = n2841 & ~n2877;
  assign n2879 = n2878 ^ n2840;
  assign n2889 = n2888 ^ n2879;
  assign n2874 = n2816 ^ n2809;
  assign n2875 = n2817 & ~n2874;
  assign n2876 = n2875 ^ n2809;
  assign n2890 = n2889 ^ n2876;
  assign n2871 = n2759 ^ n2735;
  assign n2872 = ~n2736 & n2871;
  assign n2873 = n2872 ^ n2759;
  assign n2891 = n2890 ^ n2873;
  assign n2959 = n2958 ^ n2891;
  assign n2867 = n2760 ^ n2685;
  assign n2868 = n2689 ^ n2685;
  assign n2869 = n2867 & ~n2868;
  assign n2870 = n2869 ^ n2760;
  assign n2960 = n2959 ^ n2870;
  assign n3034 = n3033 ^ n2960;
  assign n2864 = n2803 ^ n2762;
  assign n2865 = ~n2852 & ~n2864;
  assign n2866 = n2865 ^ n2851;
  assign n3035 = n3034 ^ n2866;
  assign n2861 = n2853 ^ n2681;
  assign n2862 = ~n2682 & n2861;
  assign n2863 = n2862 ^ n2853;
  assign n3036 = n3035 ^ n2863;
  assign n3041 = n3040 ^ n3036;
  assign n3237 = n2863 & n3035;
  assign n3238 = ~n2863 & ~n3035;
  assign n3239 = ~n3040 & ~n3238;
  assign n3240 = ~n3237 & ~n3239;
  assign n3222 = x7 & n2142;
  assign n3223 = x6 & n2144;
  assign n3224 = ~n3222 & ~n3223;
  assign n3225 = ~x7 & n2135;
  assign n3226 = ~x6 & n2139;
  assign n3227 = ~n3225 & ~n3226;
  assign n3228 = n3224 & n3227;
  assign n3214 = ~x9 & n1811;
  assign n3215 = ~x8 & n1815;
  assign n3216 = ~n3214 & ~n3215;
  assign n3217 = x9 & n1818;
  assign n3218 = x8 & n1820;
  assign n3219 = ~n3217 & ~n3218;
  assign n3220 = n3216 & n3219;
  assign n3207 = x21 & n491;
  assign n3208 = x20 & n495;
  assign n3209 = ~n3207 & ~n3208;
  assign n3210 = ~x21 & n498;
  assign n3211 = ~x20 & n500;
  assign n3212 = ~n3210 & ~n3211;
  assign n3213 = n3209 & n3212;
  assign n3221 = n3220 ^ n3213;
  assign n3229 = n3228 ^ n3221;
  assign n3199 = ~x27 & n142;
  assign n3200 = ~x26 & n146;
  assign n3201 = ~n3199 & ~n3200;
  assign n3202 = x27 & n149;
  assign n3203 = x26 & n151;
  assign n3204 = ~n3202 & ~n3203;
  assign n3205 = n3201 & n3204;
  assign n3191 = x13 & n1204;
  assign n3192 = x12 & n1208;
  assign n3193 = ~n3191 & ~n3192;
  assign n3194 = ~x13 & n1211;
  assign n3195 = ~x12 & n1213;
  assign n3196 = ~n3194 & ~n3195;
  assign n3197 = n3193 & n3196;
  assign n3184 = ~x11 & n1549;
  assign n3185 = ~x10 & n1553;
  assign n3186 = ~n3184 & ~n3185;
  assign n3187 = x11 & n1556;
  assign n3188 = x10 & n1558;
  assign n3189 = ~n3187 & ~n3188;
  assign n3190 = n3186 & n3189;
  assign n3198 = n3197 ^ n3190;
  assign n3206 = n3205 ^ n3198;
  assign n3230 = n3229 ^ n3206;
  assign n3181 = n2903 ^ n2897;
  assign n3182 = ~n2904 & n3181;
  assign n3183 = n3182 ^ n2897;
  assign n3231 = n3230 ^ n3183;
  assign n3177 = n2889 ^ n2873;
  assign n3178 = n2876 ^ n2873;
  assign n3179 = ~n3177 & ~n3178;
  assign n3180 = n3179 ^ n2889;
  assign n3232 = n3231 ^ n3180;
  assign n3174 = n2957 ^ n2905;
  assign n3175 = ~n2906 & n3174;
  assign n3176 = n3175 ^ n2957;
  assign n3233 = n3232 ^ n3176;
  assign n3163 = x31 & n66;
  assign n3164 = ~x31 & n68;
  assign n3165 = ~x30 & n70;
  assign n3166 = ~n3164 & ~n3165;
  assign n3167 = ~n3163 & n3166;
  assign n3159 = x61 ^ x0;
  assign n3160 = ~n3003 & n3159;
  assign n3161 = n3160 ^ x0;
  assign n3162 = x63 & ~n3161;
  assign n3168 = n3167 ^ n3162;
  assign n3156 = n3002 ^ n2997;
  assign n3157 = ~n3005 & ~n3156;
  assign n3158 = n3157 ^ n3004;
  assign n3169 = n3168 ^ n3158;
  assign n3153 = n2954 ^ n2939;
  assign n3154 = n2947 & ~n3153;
  assign n3155 = n3154 ^ n2946;
  assign n3170 = n3169 ^ n3155;
  assign n3147 = n2931 ^ n2916;
  assign n3148 = n2924 & ~n3147;
  assign n3149 = n3148 ^ n2923;
  assign n3144 = n3029 ^ n3014;
  assign n3145 = n3022 & ~n3144;
  assign n3146 = n3145 ^ n3021;
  assign n3150 = n3149 ^ n3146;
  assign n3141 = n2989 ^ n2974;
  assign n3142 = n2982 & ~n3141;
  assign n3143 = n3142 ^ n2981;
  assign n3151 = n3150 ^ n3143;
  assign n3138 = n2880 ^ n2879;
  assign n3139 = ~n2888 & n3138;
  assign n3140 = n3139 ^ n2887;
  assign n3152 = n3151 ^ n3140;
  assign n3171 = n3170 ^ n3152;
  assign n3128 = ~x23 & n331;
  assign n3129 = ~x22 & n335;
  assign n3130 = ~n3128 & ~n3129;
  assign n3131 = x23 & n338;
  assign n3132 = x22 & n340;
  assign n3133 = ~n3131 & ~n3132;
  assign n3134 = n3130 & n3133;
  assign n3120 = ~x15 & n987;
  assign n3121 = ~x14 & n991;
  assign n3122 = ~n3120 & ~n3121;
  assign n3123 = x15 & n994;
  assign n3124 = x14 & n996;
  assign n3125 = ~n3123 & ~n3124;
  assign n3126 = n3122 & n3125;
  assign n3113 = x17 & n799;
  assign n3114 = x16 & n803;
  assign n3115 = ~n3113 & ~n3114;
  assign n3116 = ~x17 & n806;
  assign n3117 = ~x16 & n808;
  assign n3118 = ~n3116 & ~n3117;
  assign n3119 = n3115 & n3118;
  assign n3127 = n3126 ^ n3119;
  assign n3135 = n3134 ^ n3127;
  assign n3098 = x63 & n3003;
  assign n3099 = ~x1 & n3098;
  assign n3100 = x63 ^ x62;
  assign n3101 = ~n3003 & n3100;
  assign n3102 = x63 & n3101;
  assign n3103 = ~x0 & n3102;
  assign n3104 = ~n3099 & ~n3103;
  assign n3105 = ~x63 & n3003;
  assign n3106 = x1 & n3105;
  assign n3107 = ~x63 & n3101;
  assign n3108 = x0 & n3107;
  assign n3109 = ~n3106 & ~n3108;
  assign n3110 = n3104 & n3109;
  assign n3090 = ~x29 & n96;
  assign n3091 = ~x28 & n100;
  assign n3092 = ~n3090 & ~n3091;
  assign n3093 = x29 & n103;
  assign n3094 = x28 & n105;
  assign n3095 = ~n3093 & ~n3094;
  assign n3096 = n3092 & n3095;
  assign n3083 = ~x25 & n239;
  assign n3084 = ~x24 & n243;
  assign n3085 = ~n3083 & ~n3084;
  assign n3086 = x25 & n246;
  assign n3087 = x24 & n248;
  assign n3088 = ~n3086 & ~n3087;
  assign n3089 = n3085 & n3088;
  assign n3097 = n3096 ^ n3089;
  assign n3111 = n3110 ^ n3097;
  assign n3075 = ~x3 & n2770;
  assign n3076 = ~x2 & n2774;
  assign n3077 = ~n3075 & ~n3076;
  assign n3078 = x3 & n2777;
  assign n3079 = x2 & n2779;
  assign n3080 = ~n3078 & ~n3079;
  assign n3081 = n3077 & n3080;
  assign n3067 = ~x5 & n2359;
  assign n3068 = ~x4 & n2361;
  assign n3069 = ~n3067 & ~n3068;
  assign n3070 = x5 & n2352;
  assign n3071 = x4 & n2356;
  assign n3072 = ~n3070 & ~n3071;
  assign n3073 = n3069 & n3072;
  assign n3060 = x19 & n643;
  assign n3061 = x18 & n645;
  assign n3062 = ~n3060 & ~n3061;
  assign n3063 = ~x19 & n636;
  assign n3064 = ~x18 & n640;
  assign n3065 = ~n3063 & ~n3064;
  assign n3066 = n3062 & n3065;
  assign n3074 = n3073 ^ n3066;
  assign n3082 = n3081 ^ n3074;
  assign n3112 = n3111 ^ n3082;
  assign n3136 = n3135 ^ n3112;
  assign n3055 = n3030 ^ n3006;
  assign n3056 = n3030 ^ n2990;
  assign n3057 = ~n3055 & ~n3056;
  assign n3058 = n3057 ^ n3006;
  assign n3052 = n2932 ^ n2909;
  assign n3053 = n2956 & ~n3052;
  assign n3054 = n3053 ^ n2955;
  assign n3059 = n3058 ^ n3054;
  assign n3137 = n3136 ^ n3059;
  assign n3172 = n3171 ^ n3137;
  assign n3049 = n2967 ^ n2964;
  assign n3050 = ~n3032 & ~n3049;
  assign n3051 = n3050 ^ n3031;
  assign n3173 = n3172 ^ n3051;
  assign n3234 = n3233 ^ n3173;
  assign n3046 = n2891 ^ n2870;
  assign n3047 = ~n2959 & n3046;
  assign n3048 = n3047 ^ n2958;
  assign n3235 = n3234 ^ n3048;
  assign n3042 = n3033 ^ n2866;
  assign n3043 = n2960 ^ n2866;
  assign n3044 = n3042 & ~n3043;
  assign n3045 = n3044 ^ n3033;
  assign n3236 = n3235 ^ n3045;
  assign n3241 = n3240 ^ n3236;
  assign n3425 = n3045 & ~n3235;
  assign n3426 = ~n3045 & n3235;
  assign n3427 = ~n3240 & ~n3426;
  assign n3428 = ~n3425 & ~n3427;
  assign n3416 = x0 & x63;
  assign n3414 = ~x31 & n70;
  assign n3415 = ~n68 & ~n3414;
  assign n3417 = n3416 ^ n3415;
  assign n3407 = ~x30 & n96;
  assign n3408 = ~x29 & n100;
  assign n3409 = ~n3407 & ~n3408;
  assign n3410 = x30 & n103;
  assign n3411 = x29 & n105;
  assign n3412 = ~n3410 & ~n3411;
  assign n3413 = n3409 & n3412;
  assign n3418 = n3417 ^ n3413;
  assign n3403 = n3228 ^ n3220;
  assign n3404 = ~n3221 & n3403;
  assign n3405 = n3404 ^ n3228;
  assign n3400 = n3081 ^ n3073;
  assign n3401 = ~n3074 & n3400;
  assign n3402 = n3401 ^ n3081;
  assign n3406 = n3405 ^ n3402;
  assign n3419 = n3418 ^ n3406;
  assign n3396 = n3135 ^ n3111;
  assign n3397 = ~n3112 & n3396;
  assign n3398 = n3397 ^ n3135;
  assign n3393 = n3158 ^ n3155;
  assign n3394 = ~n3169 & n3393;
  assign n3395 = n3394 ^ n3168;
  assign n3399 = n3398 ^ n3395;
  assign n3420 = n3419 ^ n3399;
  assign n3382 = x20 & n643;
  assign n3383 = x19 & n645;
  assign n3384 = ~n3382 & ~n3383;
  assign n3385 = ~x20 & n636;
  assign n3386 = ~x19 & n640;
  assign n3387 = ~n3385 & ~n3386;
  assign n3388 = n3384 & n3387;
  assign n3374 = ~x10 & n1811;
  assign n3375 = ~x9 & n1815;
  assign n3376 = ~n3374 & ~n3375;
  assign n3377 = x10 & n1818;
  assign n3378 = x9 & n1820;
  assign n3379 = ~n3377 & ~n3378;
  assign n3380 = n3376 & n3379;
  assign n3367 = x8 & n2142;
  assign n3368 = x7 & n2144;
  assign n3369 = ~n3367 & ~n3368;
  assign n3370 = ~x8 & n2135;
  assign n3371 = ~x7 & n2139;
  assign n3372 = ~n3370 & ~n3371;
  assign n3373 = n3369 & n3372;
  assign n3381 = n3380 ^ n3373;
  assign n3389 = n3388 ^ n3381;
  assign n3358 = ~x14 & n1211;
  assign n3359 = ~x13 & n1213;
  assign n3360 = ~n3358 & ~n3359;
  assign n3361 = x14 & n1204;
  assign n3362 = x13 & n1208;
  assign n3363 = ~n3361 & ~n3362;
  assign n3364 = n3360 & n3363;
  assign n3350 = ~x24 & n331;
  assign n3351 = ~x23 & n335;
  assign n3352 = ~n3350 & ~n3351;
  assign n3353 = x24 & n338;
  assign n3354 = x23 & n340;
  assign n3355 = ~n3353 & ~n3354;
  assign n3356 = n3352 & n3355;
  assign n3343 = ~x16 & n987;
  assign n3344 = ~x15 & n991;
  assign n3345 = ~n3343 & ~n3344;
  assign n3346 = x16 & n994;
  assign n3347 = x15 & n996;
  assign n3348 = ~n3346 & ~n3347;
  assign n3349 = n3345 & n3348;
  assign n3357 = n3356 ^ n3349;
  assign n3365 = n3364 ^ n3357;
  assign n3335 = x22 & n491;
  assign n3336 = x21 & n495;
  assign n3337 = ~n3335 & ~n3336;
  assign n3338 = ~x22 & n498;
  assign n3339 = ~x21 & n500;
  assign n3340 = ~n3338 & ~n3339;
  assign n3341 = n3337 & n3340;
  assign n3327 = x28 & n149;
  assign n3328 = x27 & n151;
  assign n3329 = ~n3327 & ~n3328;
  assign n3330 = ~x28 & n142;
  assign n3331 = ~x27 & n146;
  assign n3332 = ~n3330 & ~n3331;
  assign n3333 = n3329 & n3332;
  assign n3320 = x12 & n1556;
  assign n3321 = x11 & n1558;
  assign n3322 = ~n3320 & ~n3321;
  assign n3323 = ~x12 & n1549;
  assign n3324 = ~x11 & n1553;
  assign n3325 = ~n3323 & ~n3324;
  assign n3326 = n3322 & n3325;
  assign n3334 = n3333 ^ n3326;
  assign n3342 = n3341 ^ n3334;
  assign n3366 = n3365 ^ n3342;
  assign n3390 = n3389 ^ n3366;
  assign n3315 = n3134 ^ n3126;
  assign n3316 = ~n3127 & n3315;
  assign n3317 = n3316 ^ n3134;
  assign n3312 = n3110 ^ n3089;
  assign n3313 = n3097 & ~n3312;
  assign n3314 = n3313 ^ n3096;
  assign n3318 = n3317 ^ n3314;
  assign n3308 = n3205 ^ n3197;
  assign n3309 = n3205 ^ n3190;
  assign n3310 = n3308 & ~n3309;
  assign n3311 = n3310 ^ n3197;
  assign n3319 = n3318 ^ n3311;
  assign n3391 = n3390 ^ n3319;
  assign n3305 = n3206 ^ n3183;
  assign n3306 = n3230 & ~n3305;
  assign n3307 = n3306 ^ n3229;
  assign n3392 = n3391 ^ n3307;
  assign n3421 = n3420 ^ n3392;
  assign n3299 = n3162 & ~n3167;
  assign n3291 = ~x6 & n2359;
  assign n3292 = ~x5 & n2361;
  assign n3293 = ~n3291 & ~n3292;
  assign n3294 = x6 & n2352;
  assign n3295 = x5 & n2356;
  assign n3296 = ~n3294 & ~n3295;
  assign n3297 = n3293 & n3296;
  assign n3284 = ~x4 & n2770;
  assign n3285 = ~x3 & n2774;
  assign n3286 = ~n3284 & ~n3285;
  assign n3287 = x4 & n2777;
  assign n3288 = x3 & n2779;
  assign n3289 = ~n3287 & ~n3288;
  assign n3290 = n3286 & n3289;
  assign n3298 = n3297 ^ n3290;
  assign n3300 = n3299 ^ n3298;
  assign n3276 = x18 & n799;
  assign n3277 = x17 & n803;
  assign n3278 = ~n3276 & ~n3277;
  assign n3279 = ~x18 & n806;
  assign n3280 = ~x17 & n808;
  assign n3281 = ~n3279 & ~n3280;
  assign n3282 = n3278 & n3281;
  assign n3268 = x2 & n3105;
  assign n3269 = x1 & n3107;
  assign n3270 = ~n3268 & ~n3269;
  assign n3271 = ~x2 & n3098;
  assign n3272 = ~x1 & n3102;
  assign n3273 = ~n3271 & ~n3272;
  assign n3274 = n3270 & n3273;
  assign n3261 = ~x26 & n239;
  assign n3262 = ~x25 & n243;
  assign n3263 = ~n3261 & ~n3262;
  assign n3264 = x26 & n246;
  assign n3265 = x25 & n248;
  assign n3266 = ~n3264 & ~n3265;
  assign n3267 = n3263 & n3266;
  assign n3275 = n3274 ^ n3267;
  assign n3283 = n3282 ^ n3275;
  assign n3301 = n3300 ^ n3283;
  assign n3258 = n3146 ^ n3143;
  assign n3259 = n3150 & ~n3258;
  assign n3260 = n3259 ^ n3149;
  assign n3302 = n3301 ^ n3260;
  assign n3255 = n3170 ^ n3151;
  assign n3256 = ~n3152 & ~n3255;
  assign n3257 = n3256 ^ n3170;
  assign n3303 = n3302 ^ n3257;
  assign n3252 = n3136 ^ n3058;
  assign n3253 = n3059 & ~n3252;
  assign n3254 = n3253 ^ n3136;
  assign n3304 = n3303 ^ n3254;
  assign n3422 = n3421 ^ n3304;
  assign n3248 = n3180 ^ n3176;
  assign n3249 = ~n3232 & n3248;
  assign n3250 = n3249 ^ n3231;
  assign n3245 = n3137 ^ n3051;
  assign n3246 = n3172 & ~n3245;
  assign n3247 = n3246 ^ n3171;
  assign n3251 = n3250 ^ n3247;
  assign n3423 = n3422 ^ n3251;
  assign n3242 = n3173 ^ n3048;
  assign n3243 = n3234 & n3242;
  assign n3244 = n3243 ^ n3233;
  assign n3424 = n3423 ^ n3244;
  assign n3429 = n3428 ^ n3424;
  assign n3616 = n3244 & ~n3423;
  assign n3617 = ~n3244 & n3423;
  assign n3618 = ~n3428 & ~n3617;
  assign n3619 = ~n3616 & ~n3618;
  assign n3601 = ~x5 & n2770;
  assign n3602 = ~x4 & n2774;
  assign n3603 = ~n3601 & ~n3602;
  assign n3604 = x5 & n2777;
  assign n3605 = x4 & n2779;
  assign n3606 = ~n3604 & ~n3605;
  assign n3607 = n3603 & n3606;
  assign n3608 = n3607 ^ x33;
  assign n3598 = n3415 ^ n3413;
  assign n3599 = ~n3417 & ~n3598;
  assign n3600 = n3599 ^ n3416;
  assign n3609 = n3608 ^ n3600;
  assign n3592 = n3282 ^ n3274;
  assign n3593 = n3282 ^ n3267;
  assign n3594 = n3592 & ~n3593;
  assign n3595 = n3594 ^ n3274;
  assign n3589 = n3364 ^ n3349;
  assign n3590 = n3357 & ~n3589;
  assign n3591 = n3590 ^ n3356;
  assign n3596 = n3595 ^ n3591;
  assign n3585 = n3388 ^ n3380;
  assign n3586 = n3388 ^ n3373;
  assign n3587 = n3585 & ~n3586;
  assign n3588 = n3587 ^ n3380;
  assign n3597 = n3596 ^ n3588;
  assign n3610 = n3609 ^ n3597;
  assign n3582 = n3389 ^ n3342;
  assign n3583 = n3366 & ~n3582;
  assign n3584 = n3583 ^ n3365;
  assign n3611 = n3610 ^ n3584;
  assign n3576 = n3299 ^ n3290;
  assign n3577 = n3298 & n3576;
  assign n3578 = n3577 ^ n3297;
  assign n3573 = n3314 ^ n3311;
  assign n3574 = n3318 & ~n3573;
  assign n3575 = n3574 ^ n3317;
  assign n3579 = n3578 ^ n3575;
  assign n3570 = n3418 ^ n3405;
  assign n3571 = ~n3406 & ~n3570;
  assign n3572 = n3571 ^ n3418;
  assign n3580 = n3579 ^ n3572;
  assign n3566 = n3419 ^ n3398;
  assign n3567 = n3419 ^ n3395;
  assign n3568 = ~n3566 & n3567;
  assign n3569 = n3568 ^ n3398;
  assign n3581 = n3580 ^ n3569;
  assign n3612 = n3611 ^ n3581;
  assign n3553 = ~x13 & n1549;
  assign n3554 = ~x12 & n1553;
  assign n3555 = ~n3553 & ~n3554;
  assign n3556 = x13 & n1556;
  assign n3557 = x12 & n1558;
  assign n3558 = ~n3556 & ~n3557;
  assign n3559 = n3555 & n3558;
  assign n3545 = x15 & n1204;
  assign n3546 = x14 & n1208;
  assign n3547 = ~n3545 & ~n3546;
  assign n3548 = ~x15 & n1211;
  assign n3549 = ~x14 & n1213;
  assign n3550 = ~n3548 & ~n3549;
  assign n3551 = n3547 & n3550;
  assign n3538 = ~x25 & n331;
  assign n3539 = ~x24 & n335;
  assign n3540 = ~n3538 & ~n3539;
  assign n3541 = x25 & n338;
  assign n3542 = x24 & n340;
  assign n3543 = ~n3541 & ~n3542;
  assign n3544 = n3540 & n3543;
  assign n3552 = n3551 ^ n3544;
  assign n3560 = n3559 ^ n3552;
  assign n3529 = ~x11 & n1811;
  assign n3530 = ~x10 & n1815;
  assign n3531 = ~n3529 & ~n3530;
  assign n3532 = x11 & n1818;
  assign n3533 = x10 & n1820;
  assign n3534 = ~n3532 & ~n3533;
  assign n3535 = n3531 & n3534;
  assign n3521 = ~x29 & n142;
  assign n3522 = ~x28 & n146;
  assign n3523 = ~n3521 & ~n3522;
  assign n3524 = x29 & n149;
  assign n3525 = x28 & n151;
  assign n3526 = ~n3524 & ~n3525;
  assign n3527 = n3523 & n3526;
  assign n3514 = x23 & n491;
  assign n3515 = x22 & n495;
  assign n3516 = ~n3514 & ~n3515;
  assign n3517 = ~x23 & n498;
  assign n3518 = ~x22 & n500;
  assign n3519 = ~n3517 & ~n3518;
  assign n3520 = n3516 & n3519;
  assign n3528 = n3527 ^ n3520;
  assign n3536 = n3535 ^ n3528;
  assign n3506 = x27 & n246;
  assign n3507 = x26 & n248;
  assign n3508 = ~n3506 & ~n3507;
  assign n3509 = ~x27 & n239;
  assign n3510 = ~x26 & n243;
  assign n3511 = ~n3509 & ~n3510;
  assign n3512 = n3508 & n3511;
  assign n3498 = ~x31 & n96;
  assign n3499 = ~x30 & n100;
  assign n3500 = ~n3498 & ~n3499;
  assign n3501 = x31 & n103;
  assign n3502 = x30 & n105;
  assign n3503 = ~n3501 & ~n3502;
  assign n3504 = n3500 & n3503;
  assign n3491 = ~x17 & n987;
  assign n3492 = ~x16 & n991;
  assign n3493 = ~n3491 & ~n3492;
  assign n3494 = x17 & n994;
  assign n3495 = x16 & n996;
  assign n3496 = ~n3494 & ~n3495;
  assign n3497 = n3493 & n3496;
  assign n3505 = n3504 ^ n3497;
  assign n3513 = n3512 ^ n3505;
  assign n3537 = n3536 ^ n3513;
  assign n3561 = n3560 ^ n3537;
  assign n3482 = x7 & n2352;
  assign n3483 = x6 & n2356;
  assign n3484 = ~n3482 & ~n3483;
  assign n3485 = ~x7 & n2359;
  assign n3486 = ~x6 & n2361;
  assign n3487 = ~n3485 & ~n3486;
  assign n3488 = n3484 & n3487;
  assign n3474 = ~x21 & n636;
  assign n3475 = ~x20 & n640;
  assign n3476 = ~n3474 & ~n3475;
  assign n3477 = x21 & n643;
  assign n3478 = x20 & n645;
  assign n3479 = ~n3477 & ~n3478;
  assign n3480 = n3476 & n3479;
  assign n3467 = ~x9 & n2135;
  assign n3468 = ~x8 & n2139;
  assign n3469 = ~n3467 & ~n3468;
  assign n3470 = x9 & n2142;
  assign n3471 = x8 & n2144;
  assign n3472 = ~n3470 & ~n3471;
  assign n3473 = n3469 & n3472;
  assign n3481 = n3480 ^ n3473;
  assign n3489 = n3488 ^ n3481;
  assign n3464 = x1 & x63;
  assign n3456 = ~x19 & n806;
  assign n3457 = ~x18 & n808;
  assign n3458 = ~n3456 & ~n3457;
  assign n3459 = x19 & n799;
  assign n3460 = x18 & n803;
  assign n3461 = ~n3459 & ~n3460;
  assign n3462 = n3458 & n3461;
  assign n3449 = ~x3 & n3098;
  assign n3450 = ~x2 & n3102;
  assign n3451 = ~n3449 & ~n3450;
  assign n3452 = x3 & n3105;
  assign n3453 = x2 & n3107;
  assign n3454 = ~n3452 & ~n3453;
  assign n3455 = n3451 & n3454;
  assign n3463 = n3462 ^ n3455;
  assign n3465 = n3464 ^ n3463;
  assign n3445 = n3341 ^ n3333;
  assign n3446 = n3341 ^ n3326;
  assign n3447 = n3445 & ~n3446;
  assign n3448 = n3447 ^ n3333;
  assign n3466 = n3465 ^ n3448;
  assign n3490 = n3489 ^ n3466;
  assign n3562 = n3561 ^ n3490;
  assign n3442 = n3283 ^ n3260;
  assign n3443 = ~n3301 & ~n3442;
  assign n3444 = n3443 ^ n3300;
  assign n3563 = n3562 ^ n3444;
  assign n3439 = n3319 ^ n3307;
  assign n3440 = n3391 & ~n3439;
  assign n3441 = n3440 ^ n3390;
  assign n3564 = n3563 ^ n3441;
  assign n3436 = n3257 ^ n3254;
  assign n3437 = n3303 & n3436;
  assign n3438 = n3437 ^ n3302;
  assign n3565 = n3564 ^ n3438;
  assign n3613 = n3612 ^ n3565;
  assign n3433 = n3392 ^ n3304;
  assign n3434 = ~n3421 & ~n3433;
  assign n3435 = n3434 ^ n3420;
  assign n3614 = n3613 ^ n3435;
  assign n3430 = n3422 ^ n3250;
  assign n3431 = n3251 & ~n3430;
  assign n3432 = n3431 ^ n3422;
  assign n3615 = n3614 ^ n3432;
  assign n3620 = n3619 ^ n3615;
  assign n3803 = n3432 & n3614;
  assign n3804 = ~n3432 & ~n3614;
  assign n3805 = ~n3619 & ~n3804;
  assign n3806 = ~n3803 & ~n3805;
  assign n3792 = x35 ^ x31;
  assign n3793 = n99 & n3792;
  assign n3794 = ~n96 & ~n3793;
  assign n3795 = n3794 ^ x33;
  assign n3789 = n3464 ^ n3462;
  assign n3790 = ~n3463 & ~n3789;
  assign n3791 = n3790 ^ n3464;
  assign n3796 = n3795 ^ n3791;
  assign n3786 = n3489 ^ n3465;
  assign n3787 = n3466 & ~n3786;
  assign n3788 = n3787 ^ n3489;
  assign n3797 = n3796 ^ n3788;
  assign n3782 = n3560 ^ n3536;
  assign n3783 = n3560 ^ n3513;
  assign n3784 = n3782 & ~n3783;
  assign n3785 = n3784 ^ n3536;
  assign n3798 = n3797 ^ n3785;
  assign n3775 = n3559 ^ n3544;
  assign n3776 = n3552 & ~n3775;
  assign n3777 = n3776 ^ n3551;
  assign n3772 = n3512 ^ n3504;
  assign n3773 = ~n3505 & n3772;
  assign n3774 = n3773 ^ n3512;
  assign n3778 = n3777 ^ n3774;
  assign n3769 = n3535 ^ n3527;
  assign n3770 = ~n3528 & n3769;
  assign n3771 = n3770 ^ n3535;
  assign n3779 = n3778 ^ n3771;
  assign n3765 = n3607 ^ n3600;
  assign n3766 = ~n3608 & n3765;
  assign n3767 = n3766 ^ x33;
  assign n3762 = n3595 ^ n3588;
  assign n3763 = ~n3596 & n3762;
  assign n3764 = n3763 ^ n3588;
  assign n3768 = n3767 ^ n3764;
  assign n3780 = n3779 ^ n3768;
  assign n3758 = n3578 ^ n3572;
  assign n3759 = n3575 ^ n3572;
  assign n3760 = ~n3758 & n3759;
  assign n3761 = n3760 ^ n3578;
  assign n3781 = n3780 ^ n3761;
  assign n3799 = n3798 ^ n3781;
  assign n3745 = ~x8 & n2359;
  assign n3746 = ~x7 & n2361;
  assign n3747 = ~n3745 & ~n3746;
  assign n3748 = x8 & n2352;
  assign n3749 = x7 & n2356;
  assign n3750 = ~n3748 & ~n3749;
  assign n3751 = n3747 & n3750;
  assign n3737 = ~x22 & n636;
  assign n3738 = ~x21 & n640;
  assign n3739 = ~n3737 & ~n3738;
  assign n3740 = x22 & n643;
  assign n3741 = x21 & n645;
  assign n3742 = ~n3740 & ~n3741;
  assign n3743 = n3739 & n3742;
  assign n3730 = ~x10 & n2135;
  assign n3731 = ~x9 & n2139;
  assign n3732 = ~n3730 & ~n3731;
  assign n3733 = x10 & n2142;
  assign n3734 = x9 & n2144;
  assign n3735 = ~n3733 & ~n3734;
  assign n3736 = n3732 & n3735;
  assign n3744 = n3743 ^ n3736;
  assign n3752 = n3751 ^ n3744;
  assign n3727 = x2 & x63;
  assign n3719 = ~x26 & n331;
  assign n3720 = ~x25 & n335;
  assign n3721 = ~n3719 & ~n3720;
  assign n3722 = x26 & n338;
  assign n3723 = x25 & n340;
  assign n3724 = ~n3722 & ~n3723;
  assign n3725 = n3721 & n3724;
  assign n3712 = ~x30 & n142;
  assign n3713 = ~x29 & n146;
  assign n3714 = ~n3712 & ~n3713;
  assign n3715 = x30 & n149;
  assign n3716 = x29 & n151;
  assign n3717 = ~n3715 & ~n3716;
  assign n3718 = n3714 & n3717;
  assign n3726 = n3725 ^ n3718;
  assign n3728 = n3727 ^ n3726;
  assign n3704 = ~x28 & n239;
  assign n3705 = ~x27 & n243;
  assign n3706 = ~n3704 & ~n3705;
  assign n3707 = x28 & n246;
  assign n3708 = x27 & n248;
  assign n3709 = ~n3707 & ~n3708;
  assign n3710 = n3706 & n3709;
  assign n3696 = ~x12 & n1811;
  assign n3697 = ~x11 & n1815;
  assign n3698 = ~n3696 & ~n3697;
  assign n3699 = x12 & n1818;
  assign n3700 = x11 & n1820;
  assign n3701 = ~n3699 & ~n3700;
  assign n3702 = n3698 & n3701;
  assign n3689 = ~x14 & n1549;
  assign n3690 = ~x13 & n1553;
  assign n3691 = ~n3689 & ~n3690;
  assign n3692 = x14 & n1556;
  assign n3693 = x13 & n1558;
  assign n3694 = ~n3692 & ~n3693;
  assign n3695 = n3691 & n3694;
  assign n3703 = n3702 ^ n3695;
  assign n3711 = n3710 ^ n3703;
  assign n3729 = n3728 ^ n3711;
  assign n3753 = n3752 ^ n3729;
  assign n3680 = ~x24 & n498;
  assign n3681 = ~x23 & n500;
  assign n3682 = ~n3680 & ~n3681;
  assign n3683 = x24 & n491;
  assign n3684 = x23 & n495;
  assign n3685 = ~n3683 & ~n3684;
  assign n3686 = n3682 & n3685;
  assign n3672 = ~x18 & n987;
  assign n3673 = ~x17 & n991;
  assign n3674 = ~n3672 & ~n3673;
  assign n3675 = x18 & n994;
  assign n3676 = x17 & n996;
  assign n3677 = ~n3675 & ~n3676;
  assign n3678 = n3674 & n3677;
  assign n3665 = x16 & n1204;
  assign n3666 = x15 & n1208;
  assign n3667 = ~n3665 & ~n3666;
  assign n3668 = ~x16 & n1211;
  assign n3669 = ~x15 & n1213;
  assign n3670 = ~n3668 & ~n3669;
  assign n3671 = n3667 & n3670;
  assign n3679 = n3678 ^ n3671;
  assign n3687 = n3686 ^ n3679;
  assign n3656 = ~x4 & n3098;
  assign n3657 = ~x3 & n3102;
  assign n3658 = ~n3656 & ~n3657;
  assign n3659 = x4 & n3105;
  assign n3660 = x3 & n3107;
  assign n3661 = ~n3659 & ~n3660;
  assign n3662 = n3658 & n3661;
  assign n3648 = ~x6 & n2770;
  assign n3649 = ~x5 & n2774;
  assign n3650 = ~n3648 & ~n3649;
  assign n3651 = x6 & n2777;
  assign n3652 = x5 & n2779;
  assign n3653 = ~n3651 & ~n3652;
  assign n3654 = n3650 & n3653;
  assign n3641 = x20 & n799;
  assign n3642 = x19 & n803;
  assign n3643 = ~n3641 & ~n3642;
  assign n3644 = ~x20 & n806;
  assign n3645 = ~x19 & n808;
  assign n3646 = ~n3644 & ~n3645;
  assign n3647 = n3643 & n3646;
  assign n3655 = n3654 ^ n3647;
  assign n3663 = n3662 ^ n3655;
  assign n3637 = n3488 ^ n3480;
  assign n3638 = n3488 ^ n3473;
  assign n3639 = n3637 & ~n3638;
  assign n3640 = n3639 ^ n3480;
  assign n3664 = n3663 ^ n3640;
  assign n3688 = n3687 ^ n3664;
  assign n3754 = n3753 ^ n3688;
  assign n3633 = n3609 ^ n3584;
  assign n3634 = n3597 ^ n3584;
  assign n3635 = n3633 & ~n3634;
  assign n3636 = n3635 ^ n3609;
  assign n3755 = n3754 ^ n3636;
  assign n3630 = n3490 ^ n3444;
  assign n3631 = ~n3562 & ~n3630;
  assign n3632 = n3631 ^ n3561;
  assign n3756 = n3755 ^ n3632;
  assign n3627 = n3611 ^ n3580;
  assign n3628 = n3581 & ~n3627;
  assign n3629 = n3628 ^ n3611;
  assign n3757 = n3756 ^ n3629;
  assign n3800 = n3799 ^ n3757;
  assign n3624 = n3441 ^ n3438;
  assign n3625 = n3564 & n3624;
  assign n3626 = n3625 ^ n3563;
  assign n3801 = n3800 ^ n3626;
  assign n3621 = n3565 ^ n3435;
  assign n3622 = n3613 & ~n3621;
  assign n3623 = n3622 ^ n3612;
  assign n3802 = n3801 ^ n3623;
  assign n3807 = n3806 ^ n3802;
  assign n3988 = n3623 & ~n3801;
  assign n3989 = ~n3623 & n3801;
  assign n3990 = ~n3806 & ~n3989;
  assign n3991 = ~n3988 & ~n3990;
  assign n3977 = n3710 ^ n3702;
  assign n3978 = ~n3703 & n3977;
  assign n3979 = n3978 ^ n3710;
  assign n3974 = n3686 ^ n3671;
  assign n3975 = n3679 & ~n3974;
  assign n3976 = n3975 ^ n3678;
  assign n3980 = n3979 ^ n3976;
  assign n3971 = n3751 ^ n3736;
  assign n3972 = n3744 & ~n3971;
  assign n3973 = n3972 ^ n3743;
  assign n3981 = n3980 ^ n3973;
  assign n3967 = n3752 ^ n3728;
  assign n3968 = n3752 ^ n3711;
  assign n3969 = ~n3967 & ~n3968;
  assign n3970 = n3969 ^ n3728;
  assign n3982 = n3981 ^ n3970;
  assign n3963 = n3687 ^ n3663;
  assign n3964 = n3687 ^ n3640;
  assign n3965 = n3963 & ~n3964;
  assign n3966 = n3965 ^ n3663;
  assign n3983 = n3982 ^ n3966;
  assign n3958 = n3796 ^ n3785;
  assign n3959 = n3788 ^ n3785;
  assign n3960 = n3958 & ~n3959;
  assign n3961 = n3960 ^ n3796;
  assign n3955 = n3779 ^ n3767;
  assign n3956 = n3768 & ~n3955;
  assign n3957 = n3956 ^ n3779;
  assign n3962 = n3961 ^ n3957;
  assign n3984 = n3983 ^ n3962;
  assign n3942 = x11 & n2142;
  assign n3943 = x10 & n2144;
  assign n3944 = ~n3942 & ~n3943;
  assign n3945 = ~x11 & n2135;
  assign n3946 = ~x10 & n2139;
  assign n3947 = ~n3945 & ~n3946;
  assign n3948 = n3944 & n3947;
  assign n3934 = ~x29 & n239;
  assign n3935 = ~x28 & n243;
  assign n3936 = ~n3934 & ~n3935;
  assign n3937 = x29 & n246;
  assign n3938 = x28 & n248;
  assign n3939 = ~n3937 & ~n3938;
  assign n3940 = n3936 & n3939;
  assign n3927 = x23 & n643;
  assign n3928 = x22 & n645;
  assign n3929 = ~n3927 & ~n3928;
  assign n3930 = ~x23 & n636;
  assign n3931 = ~x22 & n640;
  assign n3932 = ~n3930 & ~n3931;
  assign n3933 = n3929 & n3932;
  assign n3941 = n3940 ^ n3933;
  assign n3949 = n3948 ^ n3941;
  assign n3918 = ~x7 & n2770;
  assign n3919 = ~x6 & n2774;
  assign n3920 = ~n3918 & ~n3919;
  assign n3921 = x7 & n2777;
  assign n3922 = x6 & n2779;
  assign n3923 = ~n3921 & ~n3922;
  assign n3924 = n3920 & n3923;
  assign n3910 = ~x21 & n806;
  assign n3911 = ~x20 & n808;
  assign n3912 = ~n3910 & ~n3911;
  assign n3913 = x21 & n799;
  assign n3914 = x20 & n803;
  assign n3915 = ~n3913 & ~n3914;
  assign n3916 = n3912 & n3915;
  assign n3903 = x9 & n2352;
  assign n3904 = x8 & n2356;
  assign n3905 = ~n3903 & ~n3904;
  assign n3906 = ~x9 & n2359;
  assign n3907 = ~x8 & n2361;
  assign n3908 = ~n3906 & ~n3907;
  assign n3909 = n3905 & n3908;
  assign n3917 = n3916 ^ n3909;
  assign n3925 = n3924 ^ n3917;
  assign n3895 = ~x13 & n1811;
  assign n3896 = ~x12 & n1815;
  assign n3897 = ~n3895 & ~n3896;
  assign n3898 = x13 & n1818;
  assign n3899 = x12 & n1820;
  assign n3900 = ~n3898 & ~n3899;
  assign n3901 = n3897 & n3900;
  assign n3887 = ~x25 & n498;
  assign n3888 = ~x24 & n500;
  assign n3889 = ~n3887 & ~n3888;
  assign n3890 = x25 & n491;
  assign n3891 = x24 & n495;
  assign n3892 = ~n3890 & ~n3891;
  assign n3893 = n3889 & n3892;
  assign n3880 = ~x15 & n1549;
  assign n3881 = ~x14 & n1553;
  assign n3882 = ~n3880 & ~n3881;
  assign n3883 = x15 & n1556;
  assign n3884 = x14 & n1558;
  assign n3885 = ~n3883 & ~n3884;
  assign n3886 = n3882 & n3885;
  assign n3894 = n3893 ^ n3886;
  assign n3902 = n3901 ^ n3894;
  assign n3926 = n3925 ^ n3902;
  assign n3950 = n3949 ^ n3926;
  assign n3871 = x27 & n338;
  assign n3872 = x26 & n340;
  assign n3873 = ~n3871 & ~n3872;
  assign n3874 = ~x27 & n331;
  assign n3875 = ~x26 & n335;
  assign n3876 = ~n3874 & ~n3875;
  assign n3877 = n3873 & n3876;
  assign n3869 = ~n96 & ~n100;
  assign n3862 = x31 & n149;
  assign n3863 = x30 & n151;
  assign n3864 = ~n3862 & ~n3863;
  assign n3865 = ~x31 & n142;
  assign n3866 = ~x30 & n146;
  assign n3867 = ~n3865 & ~n3866;
  assign n3868 = n3864 & n3867;
  assign n3870 = n3869 ^ n3868;
  assign n3878 = n3877 ^ n3870;
  assign n3853 = ~x17 & n1211;
  assign n3854 = ~x16 & n1213;
  assign n3855 = ~n3853 & ~n3854;
  assign n3856 = x17 & n1204;
  assign n3857 = x16 & n1208;
  assign n3858 = ~n3856 & ~n3857;
  assign n3859 = n3855 & n3858;
  assign n3851 = x3 & x63;
  assign n3844 = ~x19 & n987;
  assign n3845 = ~x18 & n991;
  assign n3846 = ~n3844 & ~n3845;
  assign n3847 = x19 & n994;
  assign n3848 = x18 & n996;
  assign n3849 = ~n3847 & ~n3848;
  assign n3850 = n3846 & n3849;
  assign n3852 = n3851 ^ n3850;
  assign n3860 = n3859 ^ n3852;
  assign n3841 = n3662 ^ n3654;
  assign n3842 = ~n3655 & n3841;
  assign n3843 = n3842 ^ n3662;
  assign n3861 = n3860 ^ n3843;
  assign n3879 = n3878 ^ n3861;
  assign n3951 = n3950 ^ n3879;
  assign n3830 = x5 & n3105;
  assign n3831 = x4 & n3107;
  assign n3832 = ~n3830 & ~n3831;
  assign n3833 = ~x5 & n3098;
  assign n3834 = ~x4 & n3102;
  assign n3835 = ~n3833 & ~n3834;
  assign n3836 = n3832 & n3835;
  assign n3837 = n3836 ^ n3794;
  assign n3827 = n3727 ^ n3725;
  assign n3828 = ~n3726 & ~n3827;
  assign n3829 = n3828 ^ n3727;
  assign n3838 = n3837 ^ n3829;
  assign n3824 = n3774 ^ n3771;
  assign n3825 = n3778 & ~n3824;
  assign n3826 = n3825 ^ n3777;
  assign n3839 = n3838 ^ n3826;
  assign n3821 = n3794 ^ n3791;
  assign n3822 = ~n3795 & ~n3821;
  assign n3823 = n3822 ^ x33;
  assign n3840 = n3839 ^ n3823;
  assign n3952 = n3951 ^ n3840;
  assign n3818 = n3688 ^ n3636;
  assign n3819 = ~n3754 & ~n3818;
  assign n3820 = n3819 ^ n3753;
  assign n3953 = n3952 ^ n3820;
  assign n3815 = n3798 ^ n3780;
  assign n3816 = n3781 & ~n3815;
  assign n3817 = n3816 ^ n3798;
  assign n3954 = n3953 ^ n3817;
  assign n3985 = n3984 ^ n3954;
  assign n3811 = n3755 ^ n3629;
  assign n3812 = n3632 ^ n3629;
  assign n3813 = ~n3811 & ~n3812;
  assign n3814 = n3813 ^ n3755;
  assign n3986 = n3985 ^ n3814;
  assign n3808 = n3757 ^ n3626;
  assign n3809 = n3800 & n3808;
  assign n3810 = n3809 ^ n3799;
  assign n3987 = n3986 ^ n3810;
  assign n3992 = n3991 ^ n3987;
  assign n4169 = n3810 & ~n3986;
  assign n4170 = ~n3810 & n3986;
  assign n4171 = ~n3991 & ~n4170;
  assign n4172 = ~n4169 & ~n4171;
  assign n4155 = x18 & n1204;
  assign n4156 = x17 & n1208;
  assign n4157 = ~n4155 & ~n4156;
  assign n4158 = ~x18 & n1211;
  assign n4159 = ~x17 & n1213;
  assign n4160 = ~n4158 & ~n4159;
  assign n4161 = n4157 & n4160;
  assign n4147 = ~x26 & n498;
  assign n4148 = ~x25 & n500;
  assign n4149 = ~n4147 & ~n4148;
  assign n4150 = x26 & n491;
  assign n4151 = x25 & n495;
  assign n4152 = ~n4150 & ~n4151;
  assign n4153 = n4149 & n4152;
  assign n4140 = ~x30 & n239;
  assign n4141 = ~x29 & n243;
  assign n4142 = ~n4140 & ~n4141;
  assign n4143 = x30 & n246;
  assign n4144 = x29 & n248;
  assign n4145 = ~n4143 & ~n4144;
  assign n4146 = n4142 & n4145;
  assign n4154 = n4153 ^ n4146;
  assign n4162 = n4161 ^ n4154;
  assign n4136 = n3948 ^ n3933;
  assign n4137 = n3941 & ~n4136;
  assign n4138 = n4137 ^ n3940;
  assign n4132 = n3924 ^ n3916;
  assign n4133 = n3924 ^ n3909;
  assign n4134 = n4132 & ~n4133;
  assign n4135 = n4134 ^ n3916;
  assign n4139 = n4138 ^ n4135;
  assign n4163 = n4162 ^ n4139;
  assign n4125 = n3877 ^ n3869;
  assign n4126 = n3877 ^ n3868;
  assign n4127 = ~n4125 & ~n4126;
  assign n4128 = n4127 ^ n3869;
  assign n4121 = n3859 ^ n3851;
  assign n4122 = n3859 ^ n3850;
  assign n4123 = ~n4121 & ~n4122;
  assign n4124 = n4123 ^ n3851;
  assign n4129 = n4128 ^ n4124;
  assign n4117 = n3901 ^ n3893;
  assign n4118 = n3901 ^ n3886;
  assign n4119 = n4117 & ~n4118;
  assign n4120 = n4119 ^ n3893;
  assign n4130 = n4129 ^ n4120;
  assign n4113 = n3878 ^ n3860;
  assign n4114 = n3878 ^ n3843;
  assign n4115 = n4113 & n4114;
  assign n4116 = n4115 ^ n3860;
  assign n4131 = n4130 ^ n4116;
  assign n4164 = n4163 ^ n4131;
  assign n4106 = x37 ^ x31;
  assign n4107 = n145 & n4106;
  assign n4108 = ~n142 & ~n4107;
  assign n4104 = x4 & x63;
  assign n4097 = x6 & n3105;
  assign n4098 = x5 & n3107;
  assign n4099 = ~n4097 & ~n4098;
  assign n4100 = ~x6 & n3098;
  assign n4101 = ~x5 & n3102;
  assign n4102 = ~n4100 & ~n4101;
  assign n4103 = n4099 & n4102;
  assign n4105 = n4104 ^ n4103;
  assign n4109 = n4108 ^ n4105;
  assign n4093 = n3979 ^ n3973;
  assign n4094 = n3976 ^ n3973;
  assign n4095 = n4093 & ~n4094;
  assign n4096 = n4095 ^ n3979;
  assign n4110 = n4109 ^ n4096;
  assign n4090 = n3836 ^ n3829;
  assign n4091 = n3837 & n4090;
  assign n4092 = n4091 ^ n3794;
  assign n4111 = n4110 ^ n4092;
  assign n4087 = n3970 ^ n3966;
  assign n4088 = ~n3982 & n4087;
  assign n4089 = n4088 ^ n3981;
  assign n4112 = n4111 ^ n4089;
  assign n4165 = n4164 ^ n4112;
  assign n4074 = x22 & n799;
  assign n4075 = x21 & n803;
  assign n4076 = ~n4074 & ~n4075;
  assign n4077 = ~x22 & n806;
  assign n4078 = ~x21 & n808;
  assign n4079 = ~n4077 & ~n4078;
  assign n4080 = n4076 & n4079;
  assign n4066 = ~x28 & n331;
  assign n4067 = ~x27 & n335;
  assign n4068 = ~n4066 & ~n4067;
  assign n4069 = x28 & n338;
  assign n4070 = x27 & n340;
  assign n4071 = ~n4069 & ~n4070;
  assign n4072 = n4068 & n4071;
  assign n4059 = ~x12 & n2135;
  assign n4060 = ~x11 & n2139;
  assign n4061 = ~n4059 & ~n4060;
  assign n4062 = x12 & n2142;
  assign n4063 = x11 & n2144;
  assign n4064 = ~n4062 & ~n4063;
  assign n4065 = n4061 & n4064;
  assign n4073 = n4072 ^ n4065;
  assign n4081 = n4080 ^ n4073;
  assign n4050 = ~x20 & n987;
  assign n4051 = ~x19 & n991;
  assign n4052 = ~n4050 & ~n4051;
  assign n4053 = x20 & n994;
  assign n4054 = x19 & n996;
  assign n4055 = ~n4053 & ~n4054;
  assign n4056 = n4052 & n4055;
  assign n4042 = x10 & n2352;
  assign n4043 = x9 & n2356;
  assign n4044 = ~n4042 & ~n4043;
  assign n4045 = ~x10 & n2359;
  assign n4046 = ~x9 & n2361;
  assign n4047 = ~n4045 & ~n4046;
  assign n4048 = n4044 & n4047;
  assign n4035 = x8 & n2777;
  assign n4036 = x7 & n2779;
  assign n4037 = ~n4035 & ~n4036;
  assign n4038 = ~x8 & n2770;
  assign n4039 = ~x7 & n2774;
  assign n4040 = ~n4038 & ~n4039;
  assign n4041 = n4037 & n4040;
  assign n4049 = n4048 ^ n4041;
  assign n4057 = n4056 ^ n4049;
  assign n4027 = x14 & n1818;
  assign n4028 = x13 & n1820;
  assign n4029 = ~n4027 & ~n4028;
  assign n4030 = ~x14 & n1811;
  assign n4031 = ~x13 & n1815;
  assign n4032 = ~n4030 & ~n4031;
  assign n4033 = n4029 & n4032;
  assign n4019 = ~x16 & n1549;
  assign n4020 = ~x15 & n1553;
  assign n4021 = ~n4019 & ~n4020;
  assign n4022 = x16 & n1556;
  assign n4023 = x15 & n1558;
  assign n4024 = ~n4022 & ~n4023;
  assign n4025 = n4021 & n4024;
  assign n4012 = ~x24 & n636;
  assign n4013 = ~x23 & n640;
  assign n4014 = ~n4012 & ~n4013;
  assign n4015 = x24 & n643;
  assign n4016 = x23 & n645;
  assign n4017 = ~n4015 & ~n4016;
  assign n4018 = n4014 & n4017;
  assign n4026 = n4025 ^ n4018;
  assign n4034 = n4033 ^ n4026;
  assign n4058 = n4057 ^ n4034;
  assign n4082 = n4081 ^ n4058;
  assign n4009 = n3949 ^ n3925;
  assign n4010 = ~n3926 & n4009;
  assign n4011 = n4010 ^ n3949;
  assign n4083 = n4082 ^ n4011;
  assign n4005 = n3838 ^ n3823;
  assign n4006 = n3826 ^ n3823;
  assign n4007 = ~n4005 & ~n4006;
  assign n4008 = n4007 ^ n3838;
  assign n4084 = n4083 ^ n4008;
  assign n4002 = n3879 ^ n3840;
  assign n4003 = n3951 & n4002;
  assign n4004 = n4003 ^ n3950;
  assign n4085 = n4084 ^ n4004;
  assign n3999 = n3983 ^ n3961;
  assign n4000 = ~n3962 & ~n3999;
  assign n4001 = n4000 ^ n3983;
  assign n4086 = n4085 ^ n4001;
  assign n4166 = n4165 ^ n4086;
  assign n3996 = n3820 ^ n3817;
  assign n3997 = n3953 & n3996;
  assign n3998 = n3997 ^ n3952;
  assign n4167 = n4166 ^ n3998;
  assign n3993 = n3954 ^ n3814;
  assign n3994 = ~n3985 & n3993;
  assign n3995 = n3994 ^ n3984;
  assign n4168 = n4167 ^ n3995;
  assign n4173 = n4172 ^ n4168;
  assign n4344 = n3995 & ~n4167;
  assign n4345 = ~n3995 & n4167;
  assign n4346 = ~n4172 & ~n4345;
  assign n4347 = ~n4344 & ~n4346;
  assign n4329 = ~x25 & n636;
  assign n4330 = ~x24 & n640;
  assign n4331 = ~n4329 & ~n4330;
  assign n4332 = x25 & n643;
  assign n4333 = x24 & n645;
  assign n4334 = ~n4332 & ~n4333;
  assign n4335 = n4331 & n4334;
  assign n4321 = ~x19 & n1211;
  assign n4322 = ~x18 & n1213;
  assign n4323 = ~n4321 & ~n4322;
  assign n4324 = x19 & n1204;
  assign n4325 = x18 & n1208;
  assign n4326 = ~n4324 & ~n4325;
  assign n4327 = n4323 & n4326;
  assign n4314 = x17 & n1556;
  assign n4315 = x16 & n1558;
  assign n4316 = ~n4314 & ~n4315;
  assign n4317 = ~x17 & n1549;
  assign n4318 = ~x16 & n1553;
  assign n4319 = ~n4317 & ~n4318;
  assign n4320 = n4316 & n4319;
  assign n4328 = n4327 ^ n4320;
  assign n4336 = n4335 ^ n4328;
  assign n4310 = n4056 ^ n4048;
  assign n4311 = ~n4049 & n4310;
  assign n4312 = n4311 ^ n4056;
  assign n4306 = n4080 ^ n4072;
  assign n4307 = n4080 ^ n4065;
  assign n4308 = n4306 & ~n4307;
  assign n4309 = n4308 ^ n4072;
  assign n4313 = n4312 ^ n4309;
  assign n4337 = n4336 ^ n4313;
  assign n4301 = n4161 ^ n4146;
  assign n4302 = n4154 & ~n4301;
  assign n4303 = n4302 ^ n4153;
  assign n4304 = n4303 ^ n4108;
  assign n4298 = n4033 ^ n4018;
  assign n4299 = n4026 & ~n4298;
  assign n4300 = n4299 ^ n4025;
  assign n4305 = n4304 ^ n4300;
  assign n4338 = n4337 ^ n4305;
  assign n4295 = n4162 ^ n4138;
  assign n4296 = ~n4139 & n4295;
  assign n4297 = n4296 ^ n4162;
  assign n4339 = n4338 ^ n4297;
  assign n4290 = n4109 ^ n4092;
  assign n4291 = n4096 ^ n4092;
  assign n4292 = n4290 & ~n4291;
  assign n4293 = n4292 ^ n4109;
  assign n4287 = n4163 ^ n4130;
  assign n4288 = n4131 & n4287;
  assign n4289 = n4288 ^ n4163;
  assign n4294 = n4293 ^ n4289;
  assign n4340 = n4339 ^ n4294;
  assign n4274 = ~x9 & n2770;
  assign n4275 = ~x8 & n2774;
  assign n4276 = ~n4274 & ~n4275;
  assign n4277 = x9 & n2777;
  assign n4278 = x8 & n2779;
  assign n4279 = ~n4277 & ~n4278;
  assign n4280 = n4276 & n4279;
  assign n4266 = ~x23 & n806;
  assign n4267 = ~x22 & n808;
  assign n4268 = ~n4266 & ~n4267;
  assign n4269 = x23 & n799;
  assign n4270 = x22 & n803;
  assign n4271 = ~n4269 & ~n4270;
  assign n4272 = n4268 & n4271;
  assign n4259 = ~x11 & n2359;
  assign n4260 = ~x10 & n2361;
  assign n4261 = ~n4259 & ~n4260;
  assign n4262 = x11 & n2352;
  assign n4263 = x10 & n2356;
  assign n4264 = ~n4262 & ~n4263;
  assign n4265 = n4261 & n4264;
  assign n4273 = n4272 ^ n4265;
  assign n4281 = n4280 ^ n4273;
  assign n4250 = ~x27 & n498;
  assign n4251 = ~x26 & n500;
  assign n4252 = ~n4250 & ~n4251;
  assign n4253 = x27 & n491;
  assign n4254 = x26 & n495;
  assign n4255 = ~n4253 & ~n4254;
  assign n4256 = n4252 & n4255;
  assign n4248 = ~n142 & ~n146;
  assign n4241 = ~x31 & n239;
  assign n4242 = ~x30 & n243;
  assign n4243 = ~n4241 & ~n4242;
  assign n4244 = x31 & n246;
  assign n4245 = x30 & n248;
  assign n4246 = ~n4244 & ~n4245;
  assign n4247 = n4243 & n4246;
  assign n4249 = n4248 ^ n4247;
  assign n4257 = n4256 ^ n4249;
  assign n4239 = x5 & x63;
  assign n4231 = ~x21 & n987;
  assign n4232 = ~x20 & n991;
  assign n4233 = ~n4231 & ~n4232;
  assign n4234 = x21 & n994;
  assign n4235 = x20 & n996;
  assign n4236 = ~n4234 & ~n4235;
  assign n4237 = n4233 & n4236;
  assign n4224 = ~x7 & n3098;
  assign n4225 = ~x6 & n3102;
  assign n4226 = ~n4224 & ~n4225;
  assign n4227 = x7 & n3105;
  assign n4228 = x6 & n3107;
  assign n4229 = ~n4227 & ~n4228;
  assign n4230 = n4226 & n4229;
  assign n4238 = n4237 ^ n4230;
  assign n4240 = n4239 ^ n4238;
  assign n4258 = n4257 ^ n4240;
  assign n4282 = n4281 ^ n4258;
  assign n4220 = n4081 ^ n4057;
  assign n4221 = n4081 ^ n4034;
  assign n4222 = n4220 & ~n4221;
  assign n4223 = n4222 ^ n4057;
  assign n4283 = n4282 ^ n4223;
  assign n4210 = ~x29 & n331;
  assign n4211 = ~x28 & n335;
  assign n4212 = ~n4210 & ~n4211;
  assign n4213 = x29 & n338;
  assign n4214 = x28 & n340;
  assign n4215 = ~n4213 & ~n4214;
  assign n4216 = n4212 & n4215;
  assign n4202 = ~x15 & n1811;
  assign n4203 = ~x14 & n1815;
  assign n4204 = ~n4202 & ~n4203;
  assign n4205 = x15 & n1818;
  assign n4206 = x14 & n1820;
  assign n4207 = ~n4205 & ~n4206;
  assign n4208 = n4204 & n4207;
  assign n4195 = x13 & n2142;
  assign n4196 = x12 & n2144;
  assign n4197 = ~n4195 & ~n4196;
  assign n4198 = ~x13 & n2135;
  assign n4199 = ~x12 & n2139;
  assign n4200 = ~n4198 & ~n4199;
  assign n4201 = n4197 & n4200;
  assign n4209 = n4208 ^ n4201;
  assign n4217 = n4216 ^ n4209;
  assign n4191 = n4108 ^ n4104;
  assign n4192 = n4108 ^ n4103;
  assign n4193 = n4191 & n4192;
  assign n4194 = n4193 ^ n4104;
  assign n4218 = n4217 ^ n4194;
  assign n4187 = n4128 ^ n4120;
  assign n4188 = n4124 ^ n4120;
  assign n4189 = ~n4187 & n4188;
  assign n4190 = n4189 ^ n4128;
  assign n4219 = n4218 ^ n4190;
  assign n4284 = n4283 ^ n4219;
  assign n4184 = n4011 ^ n4008;
  assign n4185 = n4083 & n4184;
  assign n4186 = n4185 ^ n4082;
  assign n4285 = n4284 ^ n4186;
  assign n4180 = n4164 ^ n4111;
  assign n4181 = n4164 ^ n4089;
  assign n4182 = ~n4180 & n4181;
  assign n4183 = n4182 ^ n4111;
  assign n4286 = n4285 ^ n4183;
  assign n4341 = n4340 ^ n4286;
  assign n4177 = n4004 ^ n4001;
  assign n4178 = ~n4085 & n4177;
  assign n4179 = n4178 ^ n4084;
  assign n4342 = n4341 ^ n4179;
  assign n4174 = n4086 ^ n3998;
  assign n4175 = ~n4166 & n4174;
  assign n4176 = n4175 ^ n4165;
  assign n4343 = n4342 ^ n4176;
  assign n4348 = n4347 ^ n4343;
  assign n4508 = n4176 & n4342;
  assign n4509 = ~n4176 & ~n4342;
  assign n4510 = ~n4347 & ~n4509;
  assign n4511 = ~n4508 & ~n4510;
  assign n4495 = n4256 ^ n4248;
  assign n4496 = n4256 ^ n4247;
  assign n4497 = ~n4495 & ~n4496;
  assign n4498 = n4497 ^ n4248;
  assign n4492 = n4335 ^ n4327;
  assign n4493 = ~n4328 & n4492;
  assign n4494 = n4493 ^ n4335;
  assign n4499 = n4498 ^ n4494;
  assign n4489 = n4216 ^ n4201;
  assign n4490 = n4209 & ~n4489;
  assign n4491 = n4490 ^ n4208;
  assign n4500 = n4499 ^ n4491;
  assign n4486 = n4303 ^ n4300;
  assign n4487 = n4304 & ~n4486;
  assign n4488 = n4487 ^ n4108;
  assign n4501 = n4500 ^ n4488;
  assign n4483 = n4336 ^ n4312;
  assign n4484 = ~n4313 & n4483;
  assign n4485 = n4484 ^ n4336;
  assign n4502 = n4501 ^ n4485;
  assign n4472 = ~x10 & n2770;
  assign n4473 = ~x9 & n2774;
  assign n4474 = ~n4472 & ~n4473;
  assign n4475 = x10 & n2777;
  assign n4476 = x9 & n2779;
  assign n4477 = ~n4475 & ~n4476;
  assign n4478 = n4474 & n4477;
  assign n4468 = x39 ^ x31;
  assign n4469 = n242 & n4468;
  assign n4470 = ~n239 & ~n4469;
  assign n4461 = ~x22 & n987;
  assign n4462 = ~x21 & n991;
  assign n4463 = ~n4461 & ~n4462;
  assign n4464 = x22 & n994;
  assign n4465 = x21 & n996;
  assign n4466 = ~n4464 & ~n4465;
  assign n4467 = n4463 & n4466;
  assign n4471 = n4470 ^ n4467;
  assign n4479 = n4478 ^ n4471;
  assign n4453 = x12 & n2352;
  assign n4454 = x11 & n2356;
  assign n4455 = ~n4453 & ~n4454;
  assign n4456 = ~x12 & n2359;
  assign n4457 = ~x11 & n2361;
  assign n4458 = ~n4456 & ~n4457;
  assign n4459 = n4455 & n4458;
  assign n4445 = ~x24 & n806;
  assign n4446 = ~x23 & n808;
  assign n4447 = ~n4445 & ~n4446;
  assign n4448 = x24 & n799;
  assign n4449 = x23 & n803;
  assign n4450 = ~n4448 & ~n4449;
  assign n4451 = n4447 & n4450;
  assign n4438 = ~x14 & n2135;
  assign n4439 = ~x13 & n2139;
  assign n4440 = ~n4438 & ~n4439;
  assign n4441 = x14 & n2142;
  assign n4442 = x13 & n2144;
  assign n4443 = ~n4441 & ~n4442;
  assign n4444 = n4440 & n4443;
  assign n4452 = n4451 ^ n4444;
  assign n4460 = n4459 ^ n4452;
  assign n4480 = n4479 ^ n4460;
  assign n4429 = ~x30 & n331;
  assign n4430 = ~x29 & n335;
  assign n4431 = ~n4429 & ~n4430;
  assign n4432 = x30 & n338;
  assign n4433 = x29 & n340;
  assign n4434 = ~n4432 & ~n4433;
  assign n4435 = n4431 & n4434;
  assign n4422 = ~x20 & n1211;
  assign n4423 = ~x19 & n1213;
  assign n4424 = ~n4422 & ~n4423;
  assign n4425 = x20 & n1204;
  assign n4426 = x19 & n1208;
  assign n4427 = ~n4425 & ~n4426;
  assign n4428 = n4424 & n4427;
  assign n4436 = n4435 ^ n4428;
  assign n4419 = n4280 ^ n4272;
  assign n4420 = ~n4273 & n4419;
  assign n4421 = n4420 ^ n4280;
  assign n4437 = n4436 ^ n4421;
  assign n4481 = n4480 ^ n4437;
  assign n4416 = n4305 ^ n4297;
  assign n4417 = n4338 & ~n4416;
  assign n4418 = n4417 ^ n4337;
  assign n4482 = n4481 ^ n4418;
  assign n4503 = n4502 ^ n4482;
  assign n4404 = ~x16 & n1811;
  assign n4405 = ~x15 & n1815;
  assign n4406 = ~n4404 & ~n4405;
  assign n4407 = x16 & n1818;
  assign n4408 = x15 & n1820;
  assign n4409 = ~n4407 & ~n4408;
  assign n4410 = n4406 & n4409;
  assign n4396 = ~x26 & n636;
  assign n4397 = ~x25 & n640;
  assign n4398 = ~n4396 & ~n4397;
  assign n4399 = x26 & n643;
  assign n4400 = x25 & n645;
  assign n4401 = ~n4399 & ~n4400;
  assign n4402 = n4398 & n4401;
  assign n4389 = ~x18 & n1549;
  assign n4390 = ~x17 & n1553;
  assign n4391 = ~n4389 & ~n4390;
  assign n4392 = x18 & n1556;
  assign n4393 = x17 & n1558;
  assign n4394 = ~n4392 & ~n4393;
  assign n4395 = n4391 & n4394;
  assign n4403 = n4402 ^ n4395;
  assign n4411 = n4410 ^ n4403;
  assign n4386 = x6 & x63;
  assign n4378 = ~x28 & n498;
  assign n4379 = ~x27 & n500;
  assign n4380 = ~n4378 & ~n4379;
  assign n4381 = x28 & n491;
  assign n4382 = x27 & n495;
  assign n4383 = ~n4381 & ~n4382;
  assign n4384 = n4380 & n4383;
  assign n4371 = ~x8 & n3098;
  assign n4372 = ~x7 & n3102;
  assign n4373 = ~n4371 & ~n4372;
  assign n4374 = x8 & n3105;
  assign n4375 = x7 & n3107;
  assign n4376 = ~n4374 & ~n4375;
  assign n4377 = n4373 & n4376;
  assign n4385 = n4384 ^ n4377;
  assign n4387 = n4386 ^ n4385;
  assign n4368 = n4239 ^ n4237;
  assign n4369 = ~n4238 & ~n4368;
  assign n4370 = n4369 ^ n4239;
  assign n4388 = n4387 ^ n4370;
  assign n4412 = n4411 ^ n4388;
  assign n4364 = n4281 ^ n4257;
  assign n4365 = n4281 ^ n4240;
  assign n4366 = ~n4364 & n4365;
  assign n4367 = n4366 ^ n4257;
  assign n4413 = n4412 ^ n4367;
  assign n4361 = n4194 ^ n4190;
  assign n4362 = ~n4218 & ~n4361;
  assign n4363 = n4362 ^ n4217;
  assign n4414 = n4413 ^ n4363;
  assign n4358 = n4223 ^ n4219;
  assign n4359 = n4283 & ~n4358;
  assign n4360 = n4359 ^ n4282;
  assign n4415 = n4414 ^ n4360;
  assign n4504 = n4503 ^ n4415;
  assign n4355 = n4339 ^ n4293;
  assign n4356 = ~n4294 & n4355;
  assign n4357 = n4356 ^ n4339;
  assign n4505 = n4504 ^ n4357;
  assign n4352 = n4186 ^ n4183;
  assign n4353 = n4285 & ~n4352;
  assign n4354 = n4353 ^ n4284;
  assign n4506 = n4505 ^ n4354;
  assign n4349 = n4286 ^ n4179;
  assign n4350 = n4341 & n4349;
  assign n4351 = n4350 ^ n4340;
  assign n4507 = n4506 ^ n4351;
  assign n4512 = n4511 ^ n4507;
  assign n4668 = ~n4351 & n4506;
  assign n4669 = n4351 & ~n4506;
  assign n4670 = ~n4511 & ~n4669;
  assign n4671 = ~n4668 & ~n4670;
  assign n4656 = n4459 ^ n4451;
  assign n4657 = ~n4452 & n4656;
  assign n4658 = n4657 ^ n4459;
  assign n4653 = n4410 ^ n4402;
  assign n4654 = ~n4403 & n4653;
  assign n4655 = n4654 ^ n4410;
  assign n4659 = n4658 ^ n4655;
  assign n4650 = n4478 ^ n4467;
  assign n4651 = n4471 & ~n4650;
  assign n4652 = n4651 ^ n4470;
  assign n4660 = n4659 ^ n4652;
  assign n4646 = n4428 ^ n4421;
  assign n4647 = ~n4436 & ~n4646;
  assign n4648 = n4647 ^ n4435;
  assign n4643 = n4494 ^ n4491;
  assign n4644 = ~n4499 & ~n4643;
  assign n4645 = n4644 ^ n4498;
  assign n4649 = n4648 ^ n4645;
  assign n4661 = n4660 ^ n4649;
  assign n4640 = n4460 ^ n4437;
  assign n4641 = n4480 & n4640;
  assign n4642 = n4641 ^ n4479;
  assign n4662 = n4661 ^ n4642;
  assign n4636 = n4500 ^ n4485;
  assign n4637 = n4488 ^ n4485;
  assign n4638 = ~n4636 & ~n4637;
  assign n4639 = n4638 ^ n4500;
  assign n4663 = n4662 ^ n4639;
  assign n4630 = x7 & x63;
  assign n4623 = ~x21 & n1211;
  assign n4624 = ~x20 & n1213;
  assign n4625 = ~n4623 & ~n4624;
  assign n4626 = x21 & n1204;
  assign n4627 = x20 & n1208;
  assign n4628 = ~n4626 & ~n4627;
  assign n4629 = n4625 & n4628;
  assign n4631 = n4630 ^ n4629;
  assign n4632 = n4631 ^ n4435;
  assign n4614 = x9 & n3105;
  assign n4615 = x8 & n3107;
  assign n4616 = ~n4614 & ~n4615;
  assign n4617 = ~x9 & n3098;
  assign n4618 = ~x8 & n3102;
  assign n4619 = ~n4617 & ~n4618;
  assign n4620 = n4616 & n4619;
  assign n4606 = x23 & n994;
  assign n4607 = x22 & n996;
  assign n4608 = ~n4606 & ~n4607;
  assign n4609 = ~x23 & n987;
  assign n4610 = ~x22 & n991;
  assign n4611 = ~n4609 & ~n4610;
  assign n4612 = n4608 & n4611;
  assign n4599 = ~x11 & n2770;
  assign n4600 = ~x10 & n2774;
  assign n4601 = ~n4599 & ~n4600;
  assign n4602 = x11 & n2777;
  assign n4603 = x10 & n2779;
  assign n4604 = ~n4602 & ~n4603;
  assign n4605 = n4601 & n4604;
  assign n4613 = n4612 ^ n4605;
  assign n4621 = n4620 ^ n4613;
  assign n4591 = ~x29 & n498;
  assign n4592 = ~x28 & n500;
  assign n4593 = ~n4591 & ~n4592;
  assign n4594 = x29 & n491;
  assign n4595 = x28 & n495;
  assign n4596 = ~n4594 & ~n4595;
  assign n4597 = n4593 & n4596;
  assign n4583 = x15 & n2142;
  assign n4584 = x14 & n2144;
  assign n4585 = ~n4583 & ~n4584;
  assign n4586 = ~x15 & n2135;
  assign n4587 = ~x14 & n2139;
  assign n4588 = ~n4586 & ~n4587;
  assign n4589 = n4585 & n4588;
  assign n4576 = ~x13 & n2359;
  assign n4577 = ~x12 & n2361;
  assign n4578 = ~n4576 & ~n4577;
  assign n4579 = x13 & n2352;
  assign n4580 = x12 & n2356;
  assign n4581 = ~n4579 & ~n4580;
  assign n4582 = n4578 & n4581;
  assign n4590 = n4589 ^ n4582;
  assign n4598 = n4597 ^ n4590;
  assign n4622 = n4621 ^ n4598;
  assign n4633 = n4632 ^ n4622;
  assign n4566 = x27 & n643;
  assign n4567 = x26 & n645;
  assign n4568 = ~n4566 & ~n4567;
  assign n4569 = ~x27 & n636;
  assign n4570 = ~x26 & n640;
  assign n4571 = ~n4569 & ~n4570;
  assign n4572 = n4568 & n4571;
  assign n4564 = ~n239 & ~n243;
  assign n4557 = ~x31 & n331;
  assign n4558 = ~x30 & n335;
  assign n4559 = ~n4557 & ~n4558;
  assign n4560 = x31 & n338;
  assign n4561 = x30 & n340;
  assign n4562 = ~n4560 & ~n4561;
  assign n4563 = n4559 & n4562;
  assign n4565 = n4564 ^ n4563;
  assign n4573 = n4572 ^ n4565;
  assign n4548 = ~x25 & n806;
  assign n4549 = ~x24 & n808;
  assign n4550 = ~n4548 & ~n4549;
  assign n4551 = x25 & n799;
  assign n4552 = x24 & n803;
  assign n4553 = ~n4551 & ~n4552;
  assign n4554 = n4550 & n4553;
  assign n4540 = ~x19 & n1549;
  assign n4541 = ~x18 & n1553;
  assign n4542 = ~n4540 & ~n4541;
  assign n4543 = x19 & n1556;
  assign n4544 = x18 & n1558;
  assign n4545 = ~n4543 & ~n4544;
  assign n4546 = n4542 & n4545;
  assign n4533 = ~x17 & n1811;
  assign n4534 = ~x16 & n1815;
  assign n4535 = ~n4533 & ~n4534;
  assign n4536 = x17 & n1818;
  assign n4537 = x16 & n1820;
  assign n4538 = ~n4536 & ~n4537;
  assign n4539 = n4535 & n4538;
  assign n4547 = n4546 ^ n4539;
  assign n4555 = n4554 ^ n4547;
  assign n4530 = n4386 ^ n4384;
  assign n4531 = ~n4385 & ~n4530;
  assign n4532 = n4531 ^ n4386;
  assign n4556 = n4555 ^ n4532;
  assign n4574 = n4573 ^ n4556;
  assign n4527 = n4411 ^ n4387;
  assign n4528 = ~n4388 & ~n4527;
  assign n4529 = n4528 ^ n4411;
  assign n4575 = n4574 ^ n4529;
  assign n4634 = n4633 ^ n4575;
  assign n4524 = n4367 ^ n4363;
  assign n4525 = ~n4413 & n4524;
  assign n4526 = n4525 ^ n4412;
  assign n4635 = n4634 ^ n4526;
  assign n4664 = n4663 ^ n4635;
  assign n4520 = n4502 ^ n4481;
  assign n4521 = n4502 ^ n4418;
  assign n4522 = n4520 & n4521;
  assign n4523 = n4522 ^ n4481;
  assign n4665 = n4664 ^ n4523;
  assign n4516 = n4503 ^ n4414;
  assign n4517 = n4503 ^ n4360;
  assign n4518 = ~n4516 & ~n4517;
  assign n4519 = n4518 ^ n4414;
  assign n4666 = n4665 ^ n4519;
  assign n4513 = n4357 ^ n4354;
  assign n4514 = ~n4505 & ~n4513;
  assign n4515 = n4514 ^ n4504;
  assign n4667 = n4666 ^ n4515;
  assign n4672 = n4671 ^ n4667;
  assign n4821 = n4515 & ~n4666;
  assign n4822 = ~n4515 & n4666;
  assign n4823 = ~n4671 & ~n4822;
  assign n4824 = ~n4821 & ~n4823;
  assign n4807 = ~x30 & n498;
  assign n4808 = ~x29 & n500;
  assign n4809 = ~n4807 & ~n4808;
  assign n4810 = x30 & n491;
  assign n4811 = x29 & n495;
  assign n4812 = ~n4810 & ~n4811;
  assign n4813 = n4809 & n4812;
  assign n4804 = n4554 ^ n4546;
  assign n4805 = ~n4547 & n4804;
  assign n4806 = n4805 ^ n4554;
  assign n4814 = n4813 ^ n4806;
  assign n4801 = n4597 ^ n4589;
  assign n4802 = ~n4590 & n4801;
  assign n4803 = n4802 ^ n4597;
  assign n4815 = n4814 ^ n4803;
  assign n4797 = n4629 ^ n4435;
  assign n4798 = ~n4631 & ~n4797;
  assign n4799 = n4798 ^ n4630;
  assign n4794 = n4655 ^ n4652;
  assign n4795 = n4659 & ~n4794;
  assign n4796 = n4795 ^ n4658;
  assign n4800 = n4799 ^ n4796;
  assign n4816 = n4815 ^ n4800;
  assign n4784 = ~x12 & n2770;
  assign n4785 = ~x11 & n2774;
  assign n4786 = ~n4784 & ~n4785;
  assign n4787 = x12 & n2777;
  assign n4788 = x11 & n2779;
  assign n4789 = ~n4787 & ~n4788;
  assign n4790 = n4786 & n4789;
  assign n4776 = ~x24 & n987;
  assign n4777 = ~x23 & n991;
  assign n4778 = ~n4776 & ~n4777;
  assign n4779 = x24 & n994;
  assign n4780 = x23 & n996;
  assign n4781 = ~n4779 & ~n4780;
  assign n4782 = n4778 & n4781;
  assign n4769 = ~x14 & n2359;
  assign n4770 = ~x13 & n2361;
  assign n4771 = ~n4769 & ~n4770;
  assign n4772 = x14 & n2352;
  assign n4773 = x13 & n2356;
  assign n4774 = ~n4772 & ~n4773;
  assign n4775 = n4771 & n4774;
  assign n4783 = n4782 ^ n4775;
  assign n4791 = n4790 ^ n4783;
  assign n4760 = ~x16 & n2135;
  assign n4761 = ~x15 & n2139;
  assign n4762 = ~n4760 & ~n4761;
  assign n4763 = x16 & n2142;
  assign n4764 = x15 & n2144;
  assign n4765 = ~n4763 & ~n4764;
  assign n4766 = n4762 & n4765;
  assign n4752 = ~x18 & n1811;
  assign n4753 = ~x17 & n1815;
  assign n4754 = ~n4752 & ~n4753;
  assign n4755 = x18 & n1818;
  assign n4756 = x17 & n1820;
  assign n4757 = ~n4755 & ~n4756;
  assign n4758 = n4754 & n4757;
  assign n4745 = x26 & n799;
  assign n4746 = x25 & n803;
  assign n4747 = ~n4745 & ~n4746;
  assign n4748 = ~x26 & n806;
  assign n4749 = ~x25 & n808;
  assign n4750 = ~n4748 & ~n4749;
  assign n4751 = n4747 & n4750;
  assign n4759 = n4758 ^ n4751;
  assign n4767 = n4766 ^ n4759;
  assign n4737 = ~x10 & n3098;
  assign n4738 = ~x9 & n3102;
  assign n4739 = ~n4737 & ~n4738;
  assign n4740 = x10 & n3105;
  assign n4741 = x9 & n3107;
  assign n4742 = ~n4740 & ~n4741;
  assign n4743 = n4739 & n4742;
  assign n4733 = x41 ^ x31;
  assign n4734 = n334 & n4733;
  assign n4735 = ~n331 & ~n4734;
  assign n4726 = x22 & n1204;
  assign n4727 = x21 & n1208;
  assign n4728 = ~n4726 & ~n4727;
  assign n4729 = ~x22 & n1211;
  assign n4730 = ~x21 & n1213;
  assign n4731 = ~n4729 & ~n4730;
  assign n4732 = n4728 & n4731;
  assign n4736 = n4735 ^ n4732;
  assign n4744 = n4743 ^ n4736;
  assign n4768 = n4767 ^ n4744;
  assign n4792 = n4791 ^ n4768;
  assign n4723 = n4660 ^ n4648;
  assign n4724 = ~n4649 & ~n4723;
  assign n4725 = n4724 ^ n4660;
  assign n4793 = n4792 ^ n4725;
  assign n4817 = n4816 ^ n4793;
  assign n4710 = ~x20 & n1549;
  assign n4711 = ~x19 & n1553;
  assign n4712 = ~n4710 & ~n4711;
  assign n4713 = x20 & n1556;
  assign n4714 = x19 & n1558;
  assign n4715 = ~n4713 & ~n4714;
  assign n4716 = n4712 & n4715;
  assign n4708 = x8 & x63;
  assign n4701 = x28 & n643;
  assign n4702 = x27 & n645;
  assign n4703 = ~n4701 & ~n4702;
  assign n4704 = ~x28 & n636;
  assign n4705 = ~x27 & n640;
  assign n4706 = ~n4704 & ~n4705;
  assign n4707 = n4703 & n4706;
  assign n4709 = n4708 ^ n4707;
  assign n4717 = n4716 ^ n4709;
  assign n4696 = n4572 ^ n4564;
  assign n4697 = n4572 ^ n4563;
  assign n4698 = ~n4696 & ~n4697;
  assign n4699 = n4698 ^ n4564;
  assign n4693 = n4620 ^ n4605;
  assign n4694 = n4613 & ~n4693;
  assign n4695 = n4694 ^ n4612;
  assign n4700 = n4699 ^ n4695;
  assign n4718 = n4717 ^ n4700;
  assign n4690 = n4573 ^ n4555;
  assign n4691 = n4556 & ~n4690;
  assign n4692 = n4691 ^ n4573;
  assign n4719 = n4718 ^ n4692;
  assign n4687 = n4632 ^ n4621;
  assign n4688 = ~n4622 & ~n4687;
  assign n4689 = n4688 ^ n4632;
  assign n4720 = n4719 ^ n4689;
  assign n4684 = n4633 ^ n4574;
  assign n4685 = ~n4575 & ~n4684;
  assign n4686 = n4685 ^ n4633;
  assign n4721 = n4720 ^ n4686;
  assign n4681 = n4661 ^ n4639;
  assign n4682 = n4662 & n4681;
  assign n4683 = n4682 ^ n4642;
  assign n4722 = n4721 ^ n4683;
  assign n4818 = n4817 ^ n4722;
  assign n4677 = n4663 ^ n4634;
  assign n4678 = n4663 ^ n4526;
  assign n4679 = n4677 & n4678;
  assign n4680 = n4679 ^ n4634;
  assign n4819 = n4818 ^ n4680;
  assign n4673 = n4523 ^ n4519;
  assign n4674 = n4664 ^ n4519;
  assign n4675 = n4673 & n4674;
  assign n4676 = n4675 ^ n4523;
  assign n4820 = n4819 ^ n4676;
  assign n4825 = n4824 ^ n4820;
  assign n4972 = n4676 & ~n4819;
  assign n4973 = ~n4676 & n4819;
  assign n4974 = ~n4824 & ~n4973;
  assign n4975 = ~n4972 & ~n4974;
  assign n4964 = x9 & x63;
  assign n4956 = ~x23 & n1211;
  assign n4957 = ~x22 & n1213;
  assign n4958 = ~n4956 & ~n4957;
  assign n4959 = x23 & n1204;
  assign n4960 = x22 & n1208;
  assign n4961 = ~n4959 & ~n4960;
  assign n4962 = n4958 & n4961;
  assign n4949 = ~x11 & n3098;
  assign n4950 = ~x10 & n3102;
  assign n4951 = ~n4949 & ~n4950;
  assign n4952 = x11 & n3105;
  assign n4953 = x10 & n3107;
  assign n4954 = ~n4952 & ~n4953;
  assign n4955 = n4951 & n4954;
  assign n4963 = n4962 ^ n4955;
  assign n4965 = n4964 ^ n4963;
  assign n4940 = ~x21 & n1549;
  assign n4941 = ~x20 & n1553;
  assign n4942 = ~n4940 & ~n4941;
  assign n4943 = x21 & n1556;
  assign n4944 = x20 & n1558;
  assign n4945 = ~n4943 & ~n4944;
  assign n4946 = n4942 & n4945;
  assign n4947 = n4946 ^ n4813;
  assign n4937 = n4790 ^ n4782;
  assign n4938 = ~n4783 & n4937;
  assign n4939 = n4938 ^ n4790;
  assign n4948 = n4947 ^ n4939;
  assign n4966 = n4965 ^ n4948;
  assign n4934 = n4806 ^ n4803;
  assign n4935 = ~n4814 & ~n4934;
  assign n4936 = n4935 ^ n4813;
  assign n4967 = n4966 ^ n4936;
  assign n4924 = x25 & n994;
  assign n4925 = x24 & n996;
  assign n4926 = ~n4924 & ~n4925;
  assign n4927 = ~x25 & n987;
  assign n4928 = ~x24 & n991;
  assign n4929 = ~n4927 & ~n4928;
  assign n4930 = n4926 & n4929;
  assign n4916 = x19 & n1818;
  assign n4917 = x18 & n1820;
  assign n4918 = ~n4916 & ~n4917;
  assign n4919 = ~x19 & n1811;
  assign n4920 = ~x18 & n1815;
  assign n4921 = ~n4919 & ~n4920;
  assign n4922 = n4918 & n4921;
  assign n4909 = ~x17 & n2135;
  assign n4910 = ~x16 & n2139;
  assign n4911 = ~n4909 & ~n4910;
  assign n4912 = x17 & n2142;
  assign n4913 = x16 & n2144;
  assign n4914 = ~n4912 & ~n4913;
  assign n4915 = n4911 & n4914;
  assign n4923 = n4922 ^ n4915;
  assign n4931 = n4930 ^ n4923;
  assign n4900 = x27 & n799;
  assign n4901 = x26 & n803;
  assign n4902 = ~n4900 & ~n4901;
  assign n4903 = ~x27 & n806;
  assign n4904 = ~x26 & n808;
  assign n4905 = ~n4903 & ~n4904;
  assign n4906 = n4902 & n4905;
  assign n4898 = ~n331 & ~n335;
  assign n4891 = ~x31 & n498;
  assign n4892 = ~x30 & n500;
  assign n4893 = ~n4891 & ~n4892;
  assign n4894 = x31 & n491;
  assign n4895 = x30 & n495;
  assign n4896 = ~n4894 & ~n4895;
  assign n4897 = n4893 & n4896;
  assign n4899 = n4898 ^ n4897;
  assign n4907 = n4906 ^ n4899;
  assign n4883 = ~x29 & n636;
  assign n4884 = ~x28 & n640;
  assign n4885 = ~n4883 & ~n4884;
  assign n4886 = x29 & n643;
  assign n4887 = x28 & n645;
  assign n4888 = ~n4886 & ~n4887;
  assign n4889 = n4885 & n4888;
  assign n4875 = ~x15 & n2359;
  assign n4876 = ~x14 & n2361;
  assign n4877 = ~n4875 & ~n4876;
  assign n4878 = x15 & n2352;
  assign n4879 = x14 & n2356;
  assign n4880 = ~n4878 & ~n4879;
  assign n4881 = n4877 & n4880;
  assign n4868 = ~x13 & n2770;
  assign n4869 = ~x12 & n2774;
  assign n4870 = ~n4868 & ~n4869;
  assign n4871 = x13 & n2777;
  assign n4872 = x12 & n2779;
  assign n4873 = ~n4871 & ~n4872;
  assign n4874 = n4870 & n4873;
  assign n4882 = n4881 ^ n4874;
  assign n4890 = n4889 ^ n4882;
  assign n4908 = n4907 ^ n4890;
  assign n4932 = n4931 ^ n4908;
  assign n4864 = n4815 ^ n4799;
  assign n4865 = n4815 ^ n4796;
  assign n4866 = n4864 & n4865;
  assign n4867 = n4866 ^ n4799;
  assign n4933 = n4932 ^ n4867;
  assign n4968 = n4967 ^ n4933;
  assign n4855 = n4716 ^ n4707;
  assign n4856 = ~n4709 & ~n4855;
  assign n4857 = n4856 ^ n4708;
  assign n4851 = n4743 ^ n4735;
  assign n4852 = n4743 ^ n4732;
  assign n4853 = n4851 & ~n4852;
  assign n4854 = n4853 ^ n4735;
  assign n4858 = n4857 ^ n4854;
  assign n4847 = n4766 ^ n4758;
  assign n4848 = n4766 ^ n4751;
  assign n4849 = n4847 & ~n4848;
  assign n4850 = n4849 ^ n4758;
  assign n4859 = n4858 ^ n4850;
  assign n4844 = n4717 ^ n4699;
  assign n4845 = n4700 & n4844;
  assign n4846 = n4845 ^ n4717;
  assign n4860 = n4859 ^ n4846;
  assign n4840 = n4791 ^ n4767;
  assign n4841 = n4791 ^ n4744;
  assign n4842 = n4840 & ~n4841;
  assign n4843 = n4842 ^ n4767;
  assign n4861 = n4860 ^ n4843;
  assign n4836 = n4718 ^ n4689;
  assign n4837 = n4692 ^ n4689;
  assign n4838 = ~n4836 & ~n4837;
  assign n4839 = n4838 ^ n4718;
  assign n4862 = n4861 ^ n4839;
  assign n4832 = n4816 ^ n4792;
  assign n4833 = n4816 ^ n4725;
  assign n4834 = n4832 & ~n4833;
  assign n4835 = n4834 ^ n4792;
  assign n4863 = n4862 ^ n4835;
  assign n4969 = n4968 ^ n4863;
  assign n4829 = n4686 ^ n4683;
  assign n4830 = ~n4721 & n4829;
  assign n4831 = n4830 ^ n4720;
  assign n4970 = n4969 ^ n4831;
  assign n4826 = n4722 ^ n4680;
  assign n4827 = ~n4818 & ~n4826;
  assign n4828 = n4827 ^ n4817;
  assign n4971 = n4970 ^ n4828;
  assign n4976 = n4975 ^ n4971;
  assign n5112 = ~n4828 & ~n4970;
  assign n5113 = n4828 & n4970;
  assign n5114 = ~n4975 & ~n5113;
  assign n5115 = ~n5112 & ~n5114;
  assign n5098 = ~x30 & n636;
  assign n5099 = ~x29 & n640;
  assign n5100 = ~n5098 & ~n5099;
  assign n5101 = x30 & n643;
  assign n5102 = x29 & n645;
  assign n5103 = ~n5101 & ~n5102;
  assign n5104 = n5100 & n5103;
  assign n5090 = ~x20 & n1811;
  assign n5091 = ~x19 & n1815;
  assign n5092 = ~n5090 & ~n5091;
  assign n5093 = x20 & n1818;
  assign n5094 = x19 & n1820;
  assign n5095 = ~n5093 & ~n5094;
  assign n5096 = n5092 & n5095;
  assign n5083 = x22 & n1556;
  assign n5084 = x21 & n1558;
  assign n5085 = ~n5083 & ~n5084;
  assign n5086 = ~x22 & n1549;
  assign n5087 = ~x21 & n1553;
  assign n5088 = ~n5086 & ~n5087;
  assign n5089 = n5085 & n5088;
  assign n5097 = n5096 ^ n5089;
  assign n5105 = n5104 ^ n5097;
  assign n5075 = ~x12 & n3098;
  assign n5076 = ~x11 & n3102;
  assign n5077 = ~n5075 & ~n5076;
  assign n5078 = x12 & n3105;
  assign n5079 = x11 & n3107;
  assign n5080 = ~n5078 & ~n5079;
  assign n5081 = n5077 & n5080;
  assign n5067 = x14 & n2777;
  assign n5068 = x13 & n2779;
  assign n5069 = ~n5067 & ~n5068;
  assign n5070 = ~x14 & n2770;
  assign n5071 = ~x13 & n2774;
  assign n5072 = ~n5070 & ~n5071;
  assign n5073 = n5069 & n5072;
  assign n5060 = x24 & n1204;
  assign n5061 = x23 & n1208;
  assign n5062 = ~n5060 & ~n5061;
  assign n5063 = ~x24 & n1211;
  assign n5064 = ~x23 & n1213;
  assign n5065 = ~n5063 & ~n5064;
  assign n5066 = n5062 & n5065;
  assign n5074 = n5073 ^ n5066;
  assign n5082 = n5081 ^ n5074;
  assign n5106 = n5105 ^ n5082;
  assign n5056 = n4857 ^ n4850;
  assign n5057 = n4854 ^ n4850;
  assign n5058 = ~n5056 & ~n5057;
  assign n5059 = n5058 ^ n4857;
  assign n5107 = n5106 ^ n5059;
  assign n5046 = ~x16 & n2359;
  assign n5047 = ~x15 & n2361;
  assign n5048 = ~n5046 & ~n5047;
  assign n5049 = x16 & n2352;
  assign n5050 = x15 & n2356;
  assign n5051 = ~n5049 & ~n5050;
  assign n5052 = n5048 & n5051;
  assign n5038 = ~x18 & n2135;
  assign n5039 = ~x17 & n2139;
  assign n5040 = ~n5038 & ~n5039;
  assign n5041 = x18 & n2142;
  assign n5042 = x17 & n2144;
  assign n5043 = ~n5041 & ~n5042;
  assign n5044 = n5040 & n5043;
  assign n5031 = ~x26 & n987;
  assign n5032 = ~x25 & n991;
  assign n5033 = ~n5031 & ~n5032;
  assign n5034 = x26 & n994;
  assign n5035 = x25 & n996;
  assign n5036 = ~n5034 & ~n5035;
  assign n5037 = n5033 & n5036;
  assign n5045 = n5044 ^ n5037;
  assign n5053 = n5052 ^ n5045;
  assign n5028 = x10 & x63;
  assign n5024 = x43 ^ x31;
  assign n5025 = n494 & n5024;
  assign n5026 = ~n498 & ~n5025;
  assign n5017 = ~x28 & n806;
  assign n5018 = ~x27 & n808;
  assign n5019 = ~n5017 & ~n5018;
  assign n5020 = x28 & n799;
  assign n5021 = x27 & n803;
  assign n5022 = ~n5020 & ~n5021;
  assign n5023 = n5019 & n5022;
  assign n5027 = n5026 ^ n5023;
  assign n5029 = n5028 ^ n5027;
  assign n5014 = n4930 ^ n4915;
  assign n5015 = n4923 & ~n5014;
  assign n5016 = n5015 ^ n4922;
  assign n5030 = n5029 ^ n5016;
  assign n5054 = n5053 ^ n5030;
  assign n5011 = n4948 ^ n4936;
  assign n5012 = ~n4966 & n5011;
  assign n5013 = n5012 ^ n4965;
  assign n5055 = n5054 ^ n5013;
  assign n5108 = n5107 ^ n5055;
  assign n5002 = n4889 ^ n4881;
  assign n5003 = ~n4882 & n5002;
  assign n5004 = n5003 ^ n4889;
  assign n4999 = n4964 ^ n4962;
  assign n5000 = ~n4963 & ~n4999;
  assign n5001 = n5000 ^ n4964;
  assign n5005 = n5004 ^ n5001;
  assign n4996 = n4906 ^ n4897;
  assign n4997 = ~n4899 & ~n4996;
  assign n4998 = n4997 ^ n4898;
  assign n5006 = n5005 ^ n4998;
  assign n4993 = n4946 ^ n4939;
  assign n4994 = n4947 & ~n4993;
  assign n4995 = n4994 ^ n4813;
  assign n5007 = n5006 ^ n4995;
  assign n4990 = n4931 ^ n4890;
  assign n4991 = ~n4908 & ~n4990;
  assign n4992 = n4991 ^ n4907;
  assign n5008 = n5007 ^ n4992;
  assign n4987 = n4859 ^ n4843;
  assign n4988 = ~n4860 & ~n4987;
  assign n4989 = n4988 ^ n4843;
  assign n5009 = n5008 ^ n4989;
  assign n4983 = n4967 ^ n4932;
  assign n4984 = n4967 ^ n4867;
  assign n4985 = ~n4983 & n4984;
  assign n4986 = n4985 ^ n4932;
  assign n5010 = n5009 ^ n4986;
  assign n5109 = n5108 ^ n5010;
  assign n4980 = n4839 ^ n4835;
  assign n4981 = n4862 & ~n4980;
  assign n4982 = n4981 ^ n4861;
  assign n5110 = n5109 ^ n4982;
  assign n4977 = n4863 ^ n4831;
  assign n4978 = n4969 & ~n4977;
  assign n4979 = n4978 ^ n4968;
  assign n5111 = n5110 ^ n4979;
  assign n5116 = n5115 ^ n5111;
  assign n5251 = ~n4979 & ~n5110;
  assign n5252 = n4979 & n5110;
  assign n5253 = ~n5115 & ~n5252;
  assign n5254 = ~n5251 & ~n5253;
  assign n5237 = ~x21 & n1811;
  assign n5238 = ~x20 & n1815;
  assign n5239 = ~n5237 & ~n5238;
  assign n5240 = x21 & n1818;
  assign n5241 = x20 & n1820;
  assign n5242 = ~n5240 & ~n5241;
  assign n5243 = n5239 & n5242;
  assign n5235 = x11 & x63;
  assign n5228 = x23 & n1556;
  assign n5229 = x22 & n1558;
  assign n5230 = ~n5228 & ~n5229;
  assign n5231 = ~x23 & n1549;
  assign n5232 = ~x22 & n1553;
  assign n5233 = ~n5231 & ~n5232;
  assign n5234 = n5230 & n5233;
  assign n5236 = n5235 ^ n5234;
  assign n5244 = n5243 ^ n5236;
  assign n5219 = ~x29 & n806;
  assign n5220 = ~x28 & n808;
  assign n5221 = ~n5219 & ~n5220;
  assign n5222 = x29 & n799;
  assign n5223 = x28 & n803;
  assign n5224 = ~n5222 & ~n5223;
  assign n5225 = n5221 & n5224;
  assign n5211 = ~x15 & n2770;
  assign n5212 = ~x14 & n2774;
  assign n5213 = ~n5211 & ~n5212;
  assign n5214 = x15 & n2777;
  assign n5215 = x14 & n2779;
  assign n5216 = ~n5214 & ~n5215;
  assign n5217 = n5213 & n5216;
  assign n5204 = ~x13 & n3098;
  assign n5205 = ~x12 & n3102;
  assign n5206 = ~n5204 & ~n5205;
  assign n5207 = x13 & n3105;
  assign n5208 = x12 & n3107;
  assign n5209 = ~n5207 & ~n5208;
  assign n5210 = n5206 & n5209;
  assign n5218 = n5217 ^ n5210;
  assign n5226 = n5225 ^ n5218;
  assign n5200 = n5081 ^ n5073;
  assign n5201 = n5081 ^ n5066;
  assign n5202 = n5200 & ~n5201;
  assign n5203 = n5202 ^ n5073;
  assign n5227 = n5226 ^ n5203;
  assign n5245 = n5244 ^ n5227;
  assign n5190 = ~x27 & n987;
  assign n5191 = ~x26 & n991;
  assign n5192 = ~n5190 & ~n5191;
  assign n5193 = x27 & n994;
  assign n5194 = x26 & n996;
  assign n5195 = ~n5193 & ~n5194;
  assign n5196 = n5192 & n5195;
  assign n5188 = ~n498 & ~n500;
  assign n5181 = ~x31 & n636;
  assign n5182 = ~x30 & n640;
  assign n5183 = ~n5181 & ~n5182;
  assign n5184 = x31 & n643;
  assign n5185 = x30 & n645;
  assign n5186 = ~n5184 & ~n5185;
  assign n5187 = n5183 & n5186;
  assign n5189 = n5188 ^ n5187;
  assign n5197 = n5196 ^ n5189;
  assign n5173 = ~x25 & n1211;
  assign n5174 = ~x24 & n1213;
  assign n5175 = ~n5173 & ~n5174;
  assign n5176 = x25 & n1204;
  assign n5177 = x24 & n1208;
  assign n5178 = ~n5176 & ~n5177;
  assign n5179 = n5175 & n5178;
  assign n5165 = x19 & n2142;
  assign n5166 = x18 & n2144;
  assign n5167 = ~n5165 & ~n5166;
  assign n5168 = ~x19 & n2135;
  assign n5169 = ~x18 & n2139;
  assign n5170 = ~n5168 & ~n5169;
  assign n5171 = n5167 & n5170;
  assign n5158 = ~x17 & n2359;
  assign n5159 = ~x16 & n2361;
  assign n5160 = ~n5158 & ~n5159;
  assign n5161 = x17 & n2352;
  assign n5162 = x16 & n2356;
  assign n5163 = ~n5161 & ~n5162;
  assign n5164 = n5160 & n5163;
  assign n5172 = n5171 ^ n5164;
  assign n5180 = n5179 ^ n5172;
  assign n5198 = n5197 ^ n5180;
  assign n5154 = n5104 ^ n5096;
  assign n5155 = n5104 ^ n5089;
  assign n5156 = ~n5154 & n5155;
  assign n5157 = n5156 ^ n5096;
  assign n5199 = n5198 ^ n5157;
  assign n5246 = n5245 ^ n5199;
  assign n5151 = n5082 ^ n5059;
  assign n5152 = ~n5106 & n5151;
  assign n5153 = n5152 ^ n5105;
  assign n5247 = n5246 ^ n5153;
  assign n5143 = n5028 ^ n5026;
  assign n5144 = ~n5027 & ~n5143;
  assign n5145 = n5144 ^ n5028;
  assign n5146 = n5145 ^ n5104;
  assign n5140 = n5052 ^ n5037;
  assign n5141 = n5045 & ~n5140;
  assign n5142 = n5141 ^ n5044;
  assign n5147 = n5146 ^ n5142;
  assign n5135 = n5053 ^ n5029;
  assign n5136 = n5053 ^ n5016;
  assign n5137 = ~n5135 & ~n5136;
  assign n5138 = n5137 ^ n5029;
  assign n5131 = n5004 ^ n4998;
  assign n5132 = n5001 ^ n4998;
  assign n5133 = ~n5131 & ~n5132;
  assign n5134 = n5133 ^ n5004;
  assign n5139 = n5138 ^ n5134;
  assign n5148 = n5147 ^ n5139;
  assign n5127 = n5006 ^ n4992;
  assign n5128 = n4995 ^ n4992;
  assign n5129 = ~n5127 & n5128;
  assign n5130 = n5129 ^ n5006;
  assign n5149 = n5148 ^ n5130;
  assign n5123 = n5107 ^ n5054;
  assign n5124 = n5107 ^ n5013;
  assign n5125 = ~n5123 & n5124;
  assign n5126 = n5125 ^ n5054;
  assign n5150 = n5149 ^ n5126;
  assign n5248 = n5247 ^ n5150;
  assign n5120 = n4989 ^ n4986;
  assign n5121 = ~n5009 & n5120;
  assign n5122 = n5121 ^ n5008;
  assign n5249 = n5248 ^ n5122;
  assign n5117 = n5010 ^ n4982;
  assign n5118 = n5109 & ~n5117;
  assign n5119 = n5118 ^ n5108;
  assign n5250 = n5249 ^ n5119;
  assign n5255 = n5254 ^ n5250;
  assign n5378 = ~n5119 & n5249;
  assign n5379 = n5119 & ~n5249;
  assign n5380 = ~n5254 & ~n5379;
  assign n5381 = ~n5378 & ~n5380;
  assign n5365 = ~x16 & n2770;
  assign n5366 = ~x15 & n2774;
  assign n5367 = ~n5365 & ~n5366;
  assign n5368 = x16 & n2777;
  assign n5369 = x15 & n2779;
  assign n5370 = ~n5368 & ~n5369;
  assign n5371 = n5367 & n5370;
  assign n5357 = x18 & n2352;
  assign n5358 = x17 & n2356;
  assign n5359 = ~n5357 & ~n5358;
  assign n5360 = ~x18 & n2359;
  assign n5361 = ~x17 & n2361;
  assign n5362 = ~n5360 & ~n5361;
  assign n5363 = n5359 & n5362;
  assign n5350 = x26 & n1204;
  assign n5351 = x25 & n1208;
  assign n5352 = ~n5350 & ~n5351;
  assign n5353 = ~x26 & n1211;
  assign n5354 = ~x25 & n1213;
  assign n5355 = ~n5353 & ~n5354;
  assign n5356 = n5352 & n5355;
  assign n5364 = n5363 ^ n5356;
  assign n5372 = n5371 ^ n5364;
  assign n5341 = ~x22 & n1811;
  assign n5342 = ~x21 & n1815;
  assign n5343 = ~n5341 & ~n5342;
  assign n5344 = x22 & n1818;
  assign n5345 = x21 & n1820;
  assign n5346 = ~n5344 & ~n5345;
  assign n5347 = n5343 & n5346;
  assign n5337 = x45 ^ x31;
  assign n5338 = n639 & n5337;
  assign n5339 = ~n636 & ~n5338;
  assign n5330 = ~x28 & n987;
  assign n5331 = ~x27 & n991;
  assign n5332 = ~n5330 & ~n5331;
  assign n5333 = x28 & n994;
  assign n5334 = x27 & n996;
  assign n5335 = ~n5333 & ~n5334;
  assign n5336 = n5332 & n5335;
  assign n5340 = n5339 ^ n5336;
  assign n5348 = n5347 ^ n5340;
  assign n5328 = x12 & x63;
  assign n5320 = x24 & n1556;
  assign n5321 = x23 & n1558;
  assign n5322 = ~n5320 & ~n5321;
  assign n5323 = ~x24 & n1549;
  assign n5324 = ~x23 & n1553;
  assign n5325 = ~n5323 & ~n5324;
  assign n5326 = n5322 & n5325;
  assign n5313 = x14 & n3105;
  assign n5314 = x13 & n3107;
  assign n5315 = ~n5313 & ~n5314;
  assign n5316 = ~x14 & n3098;
  assign n5317 = ~x13 & n3102;
  assign n5318 = ~n5316 & ~n5317;
  assign n5319 = n5315 & n5318;
  assign n5327 = n5326 ^ n5319;
  assign n5329 = n5328 ^ n5327;
  assign n5349 = n5348 ^ n5329;
  assign n5373 = n5372 ^ n5349;
  assign n5309 = n5244 ^ n5226;
  assign n5310 = ~n5227 & ~n5309;
  assign n5311 = n5310 ^ n5244;
  assign n5306 = n5180 ^ n5157;
  assign n5307 = ~n5198 & ~n5306;
  assign n5308 = n5307 ^ n5197;
  assign n5312 = n5311 ^ n5308;
  assign n5374 = n5373 ^ n5312;
  assign n5298 = n5243 ^ n5234;
  assign n5299 = ~n5236 & ~n5298;
  assign n5300 = n5299 ^ n5235;
  assign n5295 = n5196 ^ n5187;
  assign n5296 = ~n5189 & ~n5295;
  assign n5297 = n5296 ^ n5188;
  assign n5301 = n5300 ^ n5297;
  assign n5292 = n5179 ^ n5164;
  assign n5293 = n5172 & ~n5292;
  assign n5294 = n5293 ^ n5171;
  assign n5302 = n5301 ^ n5294;
  assign n5282 = ~x30 & n806;
  assign n5283 = ~x29 & n808;
  assign n5284 = ~n5282 & ~n5283;
  assign n5285 = x30 & n799;
  assign n5286 = x29 & n803;
  assign n5287 = ~n5285 & ~n5286;
  assign n5288 = n5284 & n5287;
  assign n5275 = ~x20 & n2135;
  assign n5276 = ~x19 & n2139;
  assign n5277 = ~n5275 & ~n5276;
  assign n5278 = x20 & n2142;
  assign n5279 = x19 & n2144;
  assign n5280 = ~n5278 & ~n5279;
  assign n5281 = n5277 & n5280;
  assign n5289 = n5288 ^ n5281;
  assign n5271 = n5225 ^ n5217;
  assign n5272 = n5225 ^ n5210;
  assign n5273 = n5271 & ~n5272;
  assign n5274 = n5273 ^ n5217;
  assign n5290 = n5289 ^ n5274;
  assign n5268 = n5145 ^ n5142;
  assign n5269 = ~n5146 & n5268;
  assign n5270 = n5269 ^ n5104;
  assign n5291 = n5290 ^ n5270;
  assign n5303 = n5302 ^ n5291;
  assign n5265 = n5147 ^ n5138;
  assign n5266 = n5139 & n5265;
  assign n5267 = n5266 ^ n5147;
  assign n5304 = n5303 ^ n5267;
  assign n5262 = n5199 ^ n5153;
  assign n5263 = n5246 & ~n5262;
  assign n5264 = n5263 ^ n5245;
  assign n5305 = n5304 ^ n5264;
  assign n5375 = n5374 ^ n5305;
  assign n5259 = n5130 ^ n5126;
  assign n5260 = n5149 & n5259;
  assign n5261 = n5260 ^ n5148;
  assign n5376 = n5375 ^ n5261;
  assign n5256 = n5150 ^ n5122;
  assign n5257 = n5248 & ~n5256;
  assign n5258 = n5257 ^ n5247;
  assign n5377 = n5376 ^ n5258;
  assign n5382 = n5381 ^ n5377;
  assign n5504 = n5258 & ~n5376;
  assign n5505 = ~n5258 & n5376;
  assign n5506 = ~n5381 & ~n5505;
  assign n5507 = ~n5504 & ~n5506;
  assign n5490 = x27 & n1204;
  assign n5491 = x26 & n1208;
  assign n5492 = ~n5490 & ~n5491;
  assign n5493 = ~x27 & n1211;
  assign n5494 = ~x26 & n1213;
  assign n5495 = ~n5493 & ~n5494;
  assign n5496 = n5492 & n5495;
  assign n5488 = ~n636 & ~n640;
  assign n5481 = ~x31 & n806;
  assign n5482 = ~x30 & n808;
  assign n5483 = ~n5481 & ~n5482;
  assign n5484 = x31 & n799;
  assign n5485 = x30 & n803;
  assign n5486 = ~n5484 & ~n5485;
  assign n5487 = n5483 & n5486;
  assign n5489 = n5488 ^ n5487;
  assign n5497 = n5496 ^ n5489;
  assign n5472 = ~x25 & n1549;
  assign n5473 = ~x24 & n1553;
  assign n5474 = ~n5472 & ~n5473;
  assign n5475 = x25 & n1556;
  assign n5476 = x24 & n1558;
  assign n5477 = ~n5475 & ~n5476;
  assign n5478 = n5474 & n5477;
  assign n5464 = x19 & n2352;
  assign n5465 = x18 & n2356;
  assign n5466 = ~n5464 & ~n5465;
  assign n5467 = ~x19 & n2359;
  assign n5468 = ~x18 & n2361;
  assign n5469 = ~n5467 & ~n5468;
  assign n5470 = n5466 & n5469;
  assign n5457 = ~x17 & n2770;
  assign n5458 = ~x16 & n2774;
  assign n5459 = ~n5457 & ~n5458;
  assign n5460 = x17 & n2777;
  assign n5461 = x16 & n2779;
  assign n5462 = ~n5460 & ~n5461;
  assign n5463 = n5459 & n5462;
  assign n5471 = n5470 ^ n5463;
  assign n5479 = n5478 ^ n5471;
  assign n5449 = ~x29 & n987;
  assign n5450 = ~x28 & n991;
  assign n5451 = ~n5449 & ~n5450;
  assign n5452 = x29 & n994;
  assign n5453 = x28 & n996;
  assign n5454 = ~n5452 & ~n5453;
  assign n5455 = n5451 & n5454;
  assign n5447 = x13 & x63;
  assign n5440 = x15 & n3105;
  assign n5441 = x14 & n3107;
  assign n5442 = ~n5440 & ~n5441;
  assign n5443 = ~x15 & n3098;
  assign n5444 = ~x14 & n3102;
  assign n5445 = ~n5443 & ~n5444;
  assign n5446 = n5442 & n5445;
  assign n5448 = n5447 ^ n5446;
  assign n5456 = n5455 ^ n5448;
  assign n5480 = n5479 ^ n5456;
  assign n5498 = n5497 ^ n5480;
  assign n5433 = n5347 ^ n5339;
  assign n5434 = n5347 ^ n5336;
  assign n5435 = n5433 & ~n5434;
  assign n5436 = n5435 ^ n5339;
  assign n5429 = n5371 ^ n5363;
  assign n5430 = n5371 ^ n5356;
  assign n5431 = n5429 & ~n5430;
  assign n5432 = n5431 ^ n5363;
  assign n5437 = n5436 ^ n5432;
  assign n5426 = n5328 ^ n5326;
  assign n5427 = ~n5327 & ~n5426;
  assign n5428 = n5427 ^ n5328;
  assign n5438 = n5437 ^ n5428;
  assign n5422 = n5372 ^ n5348;
  assign n5423 = n5372 ^ n5329;
  assign n5424 = n5422 & n5423;
  assign n5425 = n5424 ^ n5348;
  assign n5439 = n5438 ^ n5425;
  assign n5499 = n5498 ^ n5439;
  assign n5410 = ~x21 & n2135;
  assign n5411 = ~x20 & n2139;
  assign n5412 = ~n5410 & ~n5411;
  assign n5413 = x21 & n2142;
  assign n5414 = x20 & n2144;
  assign n5415 = ~n5413 & ~n5414;
  assign n5416 = n5412 & n5415;
  assign n5403 = x23 & n1818;
  assign n5404 = x22 & n1820;
  assign n5405 = ~n5403 & ~n5404;
  assign n5406 = ~x23 & n1811;
  assign n5407 = ~x22 & n1815;
  assign n5408 = ~n5406 & ~n5407;
  assign n5409 = n5405 & n5408;
  assign n5417 = n5416 ^ n5409;
  assign n5418 = n5417 ^ n5288;
  assign n5399 = n5300 ^ n5294;
  assign n5400 = n5297 ^ n5294;
  assign n5401 = ~n5399 & n5400;
  assign n5402 = n5401 ^ n5300;
  assign n5419 = n5418 ^ n5402;
  assign n5396 = n5281 ^ n5274;
  assign n5397 = ~n5289 & ~n5396;
  assign n5398 = n5397 ^ n5288;
  assign n5420 = n5419 ^ n5398;
  assign n5392 = n5302 ^ n5290;
  assign n5393 = n5302 ^ n5270;
  assign n5394 = ~n5392 & ~n5393;
  assign n5395 = n5394 ^ n5290;
  assign n5421 = n5420 ^ n5395;
  assign n5500 = n5499 ^ n5421;
  assign n5389 = n5373 ^ n5311;
  assign n5390 = ~n5312 & n5389;
  assign n5391 = n5390 ^ n5373;
  assign n5501 = n5500 ^ n5391;
  assign n5386 = n5267 ^ n5264;
  assign n5387 = n5304 & ~n5386;
  assign n5388 = n5387 ^ n5303;
  assign n5502 = n5501 ^ n5388;
  assign n5383 = n5305 ^ n5261;
  assign n5384 = n5375 & n5383;
  assign n5385 = n5384 ^ n5374;
  assign n5503 = n5502 ^ n5385;
  assign n5508 = n5507 ^ n5503;
  assign n5621 = n5385 & ~n5502;
  assign n5622 = ~n5385 & n5502;
  assign n5623 = ~n5507 & ~n5622;
  assign n5624 = ~n5621 & ~n5623;
  assign n5608 = ~x24 & n1811;
  assign n5609 = ~x23 & n1815;
  assign n5610 = ~n5608 & ~n5609;
  assign n5611 = x24 & n1818;
  assign n5612 = x23 & n1820;
  assign n5613 = ~n5611 & ~n5612;
  assign n5614 = n5610 & n5613;
  assign n5606 = x14 & x63;
  assign n5599 = ~x30 & n987;
  assign n5600 = ~x29 & n991;
  assign n5601 = ~n5599 & ~n5600;
  assign n5602 = x30 & n994;
  assign n5603 = x29 & n996;
  assign n5604 = ~n5602 & ~n5603;
  assign n5605 = n5601 & n5604;
  assign n5607 = n5606 ^ n5605;
  assign n5615 = n5614 ^ n5607;
  assign n5590 = ~x16 & n3098;
  assign n5591 = ~x15 & n3102;
  assign n5592 = ~n5590 & ~n5591;
  assign n5593 = x16 & n3105;
  assign n5594 = x15 & n3107;
  assign n5595 = ~n5593 & ~n5594;
  assign n5596 = n5592 & n5595;
  assign n5582 = ~x26 & n1549;
  assign n5583 = ~x25 & n1553;
  assign n5584 = ~n5582 & ~n5583;
  assign n5585 = x26 & n1556;
  assign n5586 = x25 & n1558;
  assign n5587 = ~n5585 & ~n5586;
  assign n5588 = n5584 & n5587;
  assign n5575 = ~x18 & n2770;
  assign n5576 = ~x17 & n2774;
  assign n5577 = ~n5575 & ~n5576;
  assign n5578 = x18 & n2777;
  assign n5579 = x17 & n2779;
  assign n5580 = ~n5578 & ~n5579;
  assign n5581 = n5577 & n5580;
  assign n5589 = n5588 ^ n5581;
  assign n5597 = n5596 ^ n5589;
  assign n5571 = n5455 ^ n5447;
  assign n5572 = n5455 ^ n5446;
  assign n5573 = ~n5571 & ~n5572;
  assign n5574 = n5573 ^ n5447;
  assign n5598 = n5597 ^ n5574;
  assign n5616 = n5615 ^ n5598;
  assign n5565 = x47 ^ x31;
  assign n5566 = n802 & n5565;
  assign n5567 = ~n806 & ~n5566;
  assign n5562 = n5496 ^ n5487;
  assign n5563 = ~n5489 & ~n5562;
  assign n5564 = n5563 ^ n5488;
  assign n5568 = n5567 ^ n5564;
  assign n5559 = n5478 ^ n5470;
  assign n5560 = ~n5471 & n5559;
  assign n5561 = n5560 ^ n5478;
  assign n5569 = n5568 ^ n5561;
  assign n5556 = n5497 ^ n5479;
  assign n5557 = n5480 & ~n5556;
  assign n5558 = n5557 ^ n5497;
  assign n5570 = n5569 ^ n5558;
  assign n5617 = n5616 ^ n5570;
  assign n5544 = x20 & n2352;
  assign n5545 = x19 & n2356;
  assign n5546 = ~n5544 & ~n5545;
  assign n5547 = ~x20 & n2359;
  assign n5548 = ~x19 & n2361;
  assign n5549 = ~n5547 & ~n5548;
  assign n5550 = n5546 & n5549;
  assign n5536 = ~x22 & n2135;
  assign n5537 = ~x21 & n2139;
  assign n5538 = ~n5536 & ~n5537;
  assign n5539 = x22 & n2142;
  assign n5540 = x21 & n2144;
  assign n5541 = ~n5539 & ~n5540;
  assign n5542 = n5538 & n5541;
  assign n5529 = ~x28 & n1211;
  assign n5530 = ~x27 & n1213;
  assign n5531 = ~n5529 & ~n5530;
  assign n5532 = x28 & n1204;
  assign n5533 = x27 & n1208;
  assign n5534 = ~n5532 & ~n5533;
  assign n5535 = n5531 & n5534;
  assign n5543 = n5542 ^ n5535;
  assign n5551 = n5550 ^ n5543;
  assign n5525 = n5416 ^ n5288;
  assign n5526 = n5409 ^ n5288;
  assign n5527 = n5525 & ~n5526;
  assign n5528 = n5527 ^ n5416;
  assign n5552 = n5551 ^ n5528;
  assign n5522 = n5432 ^ n5428;
  assign n5523 = n5437 & n5522;
  assign n5524 = n5523 ^ n5436;
  assign n5553 = n5552 ^ n5524;
  assign n5518 = n5418 ^ n5398;
  assign n5519 = n5402 ^ n5398;
  assign n5520 = ~n5518 & ~n5519;
  assign n5521 = n5520 ^ n5418;
  assign n5554 = n5553 ^ n5521;
  assign n5515 = n5498 ^ n5425;
  assign n5516 = n5439 & n5515;
  assign n5517 = n5516 ^ n5498;
  assign n5555 = n5554 ^ n5517;
  assign n5618 = n5617 ^ n5555;
  assign n5512 = n5499 ^ n5420;
  assign n5513 = n5421 & ~n5512;
  assign n5514 = n5513 ^ n5499;
  assign n5619 = n5618 ^ n5514;
  assign n5509 = n5391 ^ n5388;
  assign n5510 = ~n5501 & ~n5509;
  assign n5511 = n5510 ^ n5500;
  assign n5620 = n5619 ^ n5511;
  assign n5625 = n5624 ^ n5620;
  assign n5733 = ~n5511 & ~n5619;
  assign n5734 = n5511 & n5619;
  assign n5735 = ~n5624 & ~n5734;
  assign n5736 = ~n5733 & ~n5735;
  assign n5720 = ~x23 & n2135;
  assign n5721 = ~x22 & n2139;
  assign n5722 = ~n5720 & ~n5721;
  assign n5723 = x23 & n2142;
  assign n5724 = x22 & n2144;
  assign n5725 = ~n5723 & ~n5724;
  assign n5726 = n5722 & n5725;
  assign n5718 = x15 & x63;
  assign n5711 = x29 & n1204;
  assign n5712 = x28 & n1208;
  assign n5713 = ~n5711 & ~n5712;
  assign n5714 = ~x29 & n1211;
  assign n5715 = ~x28 & n1213;
  assign n5716 = ~n5714 & ~n5715;
  assign n5717 = n5713 & n5716;
  assign n5719 = n5718 ^ n5717;
  assign n5727 = n5726 ^ n5719;
  assign n5707 = n5614 ^ n5605;
  assign n5708 = ~n5607 & ~n5707;
  assign n5709 = n5708 ^ n5606;
  assign n5703 = n5550 ^ n5542;
  assign n5704 = n5550 ^ n5535;
  assign n5705 = n5703 & ~n5704;
  assign n5706 = n5705 ^ n5542;
  assign n5710 = n5709 ^ n5706;
  assign n5728 = n5727 ^ n5710;
  assign n5699 = n5615 ^ n5597;
  assign n5700 = n5598 & ~n5699;
  assign n5701 = n5700 ^ n5615;
  assign n5695 = n5567 ^ n5561;
  assign n5696 = n5564 ^ n5561;
  assign n5697 = ~n5695 & n5696;
  assign n5698 = n5697 ^ n5567;
  assign n5702 = n5701 ^ n5698;
  assign n5729 = n5728 ^ n5702;
  assign n5683 = ~x27 & n1549;
  assign n5684 = ~x26 & n1553;
  assign n5685 = ~n5683 & ~n5684;
  assign n5686 = x27 & n1556;
  assign n5687 = x26 & n1558;
  assign n5688 = ~n5686 & ~n5687;
  assign n5689 = n5685 & n5688;
  assign n5681 = ~n806 & ~n808;
  assign n5674 = ~x31 & n987;
  assign n5675 = ~x30 & n991;
  assign n5676 = ~n5674 & ~n5675;
  assign n5677 = x31 & n994;
  assign n5678 = x30 & n996;
  assign n5679 = ~n5677 & ~n5678;
  assign n5680 = n5676 & n5679;
  assign n5682 = n5681 ^ n5680;
  assign n5690 = n5689 ^ n5682;
  assign n5666 = x25 & n1818;
  assign n5667 = x24 & n1820;
  assign n5668 = ~n5666 & ~n5667;
  assign n5669 = ~x25 & n1811;
  assign n5670 = ~x24 & n1815;
  assign n5671 = ~n5669 & ~n5670;
  assign n5672 = n5668 & n5671;
  assign n5658 = ~x19 & n2770;
  assign n5659 = ~x18 & n2774;
  assign n5660 = ~n5658 & ~n5659;
  assign n5661 = x19 & n2777;
  assign n5662 = x18 & n2779;
  assign n5663 = ~n5661 & ~n5662;
  assign n5664 = n5660 & n5663;
  assign n5651 = ~x17 & n3098;
  assign n5652 = ~x16 & n3102;
  assign n5653 = ~n5651 & ~n5652;
  assign n5654 = x17 & n3105;
  assign n5655 = x16 & n3107;
  assign n5656 = ~n5654 & ~n5655;
  assign n5657 = n5653 & n5656;
  assign n5665 = n5664 ^ n5657;
  assign n5673 = n5672 ^ n5665;
  assign n5691 = n5690 ^ n5673;
  assign n5642 = x21 & n2352;
  assign n5643 = x20 & n2356;
  assign n5644 = ~n5642 & ~n5643;
  assign n5645 = ~x21 & n2359;
  assign n5646 = ~x20 & n2361;
  assign n5647 = ~n5645 & ~n5646;
  assign n5648 = n5644 & n5647;
  assign n5649 = n5648 ^ n5567;
  assign n5639 = n5596 ^ n5581;
  assign n5640 = n5589 & ~n5639;
  assign n5641 = n5640 ^ n5588;
  assign n5650 = n5649 ^ n5641;
  assign n5692 = n5691 ^ n5650;
  assign n5636 = n5528 ^ n5524;
  assign n5637 = n5552 & ~n5636;
  assign n5638 = n5637 ^ n5551;
  assign n5693 = n5692 ^ n5638;
  assign n5633 = n5616 ^ n5569;
  assign n5634 = n5570 & n5633;
  assign n5635 = n5634 ^ n5616;
  assign n5694 = n5693 ^ n5635;
  assign n5730 = n5729 ^ n5694;
  assign n5629 = n5553 ^ n5517;
  assign n5630 = n5521 ^ n5517;
  assign n5631 = n5629 & ~n5630;
  assign n5632 = n5631 ^ n5553;
  assign n5731 = n5730 ^ n5632;
  assign n5626 = n5555 ^ n5514;
  assign n5627 = ~n5618 & n5626;
  assign n5628 = n5627 ^ n5617;
  assign n5732 = n5731 ^ n5628;
  assign n5737 = n5736 ^ n5732;
  assign n5836 = n5628 & n5731;
  assign n5837 = ~n5628 & ~n5731;
  assign n5838 = ~n5736 & ~n5837;
  assign n5839 = ~n5836 & ~n5838;
  assign n5827 = n5689 ^ n5680;
  assign n5828 = ~n5682 & ~n5827;
  assign n5829 = n5828 ^ n5681;
  assign n5824 = n5672 ^ n5657;
  assign n5825 = n5665 & ~n5824;
  assign n5826 = n5825 ^ n5664;
  assign n5830 = n5829 ^ n5826;
  assign n5821 = n5726 ^ n5717;
  assign n5822 = ~n5719 & ~n5821;
  assign n5823 = n5822 ^ n5718;
  assign n5831 = n5830 ^ n5823;
  assign n5817 = n5648 ^ n5641;
  assign n5818 = n5649 & ~n5817;
  assign n5819 = n5818 ^ n5567;
  assign n5814 = n5727 ^ n5709;
  assign n5815 = n5710 & n5814;
  assign n5816 = n5815 ^ n5727;
  assign n5820 = n5819 ^ n5816;
  assign n5832 = n5831 ^ n5820;
  assign n5807 = x49 ^ x31;
  assign n5808 = n990 & n5807;
  assign n5809 = ~n987 & ~n5808;
  assign n5799 = ~x20 & n2770;
  assign n5800 = ~x19 & n2774;
  assign n5801 = ~n5799 & ~n5800;
  assign n5802 = x20 & n2777;
  assign n5803 = x19 & n2779;
  assign n5804 = ~n5802 & ~n5803;
  assign n5805 = n5801 & n5804;
  assign n5792 = ~x22 & n2359;
  assign n5793 = ~x21 & n2361;
  assign n5794 = ~n5792 & ~n5793;
  assign n5795 = x22 & n2352;
  assign n5796 = x21 & n2356;
  assign n5797 = ~n5795 & ~n5796;
  assign n5798 = n5794 & n5797;
  assign n5806 = n5805 ^ n5798;
  assign n5810 = n5809 ^ n5806;
  assign n5783 = x28 & n1556;
  assign n5784 = x27 & n1558;
  assign n5785 = ~n5783 & ~n5784;
  assign n5786 = ~x28 & n1549;
  assign n5787 = ~x27 & n1553;
  assign n5788 = ~n5786 & ~n5787;
  assign n5789 = n5785 & n5788;
  assign n5775 = x24 & n2142;
  assign n5776 = x23 & n2144;
  assign n5777 = ~n5775 & ~n5776;
  assign n5778 = ~x24 & n2135;
  assign n5779 = ~x23 & n2139;
  assign n5780 = ~n5778 & ~n5779;
  assign n5781 = n5777 & n5780;
  assign n5768 = x30 & n1204;
  assign n5769 = x29 & n1208;
  assign n5770 = ~n5768 & ~n5769;
  assign n5771 = ~x30 & n1211;
  assign n5772 = ~x29 & n1213;
  assign n5773 = ~n5771 & ~n5772;
  assign n5774 = n5770 & n5773;
  assign n5782 = n5781 ^ n5774;
  assign n5790 = n5789 ^ n5782;
  assign n5766 = x16 & x63;
  assign n5758 = ~x18 & n3098;
  assign n5759 = ~x17 & n3102;
  assign n5760 = ~n5758 & ~n5759;
  assign n5761 = x18 & n3105;
  assign n5762 = x17 & n3107;
  assign n5763 = ~n5761 & ~n5762;
  assign n5764 = n5760 & n5763;
  assign n5751 = x26 & n1818;
  assign n5752 = x25 & n1820;
  assign n5753 = ~n5751 & ~n5752;
  assign n5754 = ~x26 & n1811;
  assign n5755 = ~x25 & n1815;
  assign n5756 = ~n5754 & ~n5755;
  assign n5757 = n5753 & n5756;
  assign n5765 = n5764 ^ n5757;
  assign n5767 = n5766 ^ n5765;
  assign n5791 = n5790 ^ n5767;
  assign n5811 = n5810 ^ n5791;
  assign n5748 = n5673 ^ n5650;
  assign n5749 = ~n5691 & ~n5748;
  assign n5750 = n5749 ^ n5690;
  assign n5812 = n5811 ^ n5750;
  assign n5745 = n5728 ^ n5701;
  assign n5746 = ~n5702 & ~n5745;
  assign n5747 = n5746 ^ n5728;
  assign n5813 = n5812 ^ n5747;
  assign n5833 = n5832 ^ n5813;
  assign n5741 = n5692 ^ n5635;
  assign n5742 = n5638 ^ n5635;
  assign n5743 = ~n5741 & ~n5742;
  assign n5744 = n5743 ^ n5692;
  assign n5834 = n5833 ^ n5744;
  assign n5738 = n5694 ^ n5632;
  assign n5739 = ~n5730 & n5738;
  assign n5740 = n5739 ^ n5729;
  assign n5835 = n5834 ^ n5740;
  assign n5840 = n5839 ^ n5835;
  assign n5933 = ~n5740 & n5834;
  assign n5934 = n5740 & ~n5834;
  assign n5935 = ~n5839 & ~n5934;
  assign n5936 = ~n5933 & ~n5935;
  assign n5924 = n5766 ^ n5764;
  assign n5925 = ~n5765 & ~n5924;
  assign n5926 = n5925 ^ n5766;
  assign n5927 = n5926 ^ n5809;
  assign n5921 = n5789 ^ n5774;
  assign n5922 = n5782 & ~n5921;
  assign n5923 = n5922 ^ n5781;
  assign n5928 = n5927 ^ n5923;
  assign n5917 = n5809 ^ n5805;
  assign n5918 = ~n5806 & ~n5917;
  assign n5919 = n5918 ^ n5809;
  assign n5914 = n5829 ^ n5823;
  assign n5915 = n5830 & n5914;
  assign n5916 = n5915 ^ n5823;
  assign n5920 = n5919 ^ n5916;
  assign n5929 = n5928 ^ n5920;
  assign n5903 = ~x25 & n2135;
  assign n5904 = ~x24 & n2139;
  assign n5905 = ~n5903 & ~n5904;
  assign n5906 = x25 & n2142;
  assign n5907 = x24 & n2144;
  assign n5908 = ~n5906 & ~n5907;
  assign n5909 = n5905 & n5908;
  assign n5901 = x17 & x63;
  assign n5894 = x19 & n3105;
  assign n5895 = x18 & n3107;
  assign n5896 = ~n5894 & ~n5895;
  assign n5897 = ~x19 & n3098;
  assign n5898 = ~x18 & n3102;
  assign n5899 = ~n5897 & ~n5898;
  assign n5900 = n5896 & n5899;
  assign n5902 = n5901 ^ n5900;
  assign n5910 = n5909 ^ n5902;
  assign n5885 = x21 & n2777;
  assign n5886 = x20 & n2779;
  assign n5887 = ~n5885 & ~n5886;
  assign n5888 = ~x21 & n2770;
  assign n5889 = ~x20 & n2774;
  assign n5890 = ~n5888 & ~n5889;
  assign n5891 = n5887 & n5890;
  assign n5877 = ~x29 & n1549;
  assign n5878 = ~x28 & n1553;
  assign n5879 = ~n5877 & ~n5878;
  assign n5880 = x29 & n1556;
  assign n5881 = x28 & n1558;
  assign n5882 = ~n5880 & ~n5881;
  assign n5883 = n5879 & n5882;
  assign n5870 = ~x23 & n2359;
  assign n5871 = ~x22 & n2361;
  assign n5872 = ~n5870 & ~n5871;
  assign n5873 = x23 & n2352;
  assign n5874 = x22 & n2356;
  assign n5875 = ~n5873 & ~n5874;
  assign n5876 = n5872 & n5875;
  assign n5884 = n5883 ^ n5876;
  assign n5892 = n5891 ^ n5884;
  assign n5862 = ~x27 & n1811;
  assign n5863 = ~x26 & n1815;
  assign n5864 = ~n5862 & ~n5863;
  assign n5865 = x27 & n1818;
  assign n5866 = x26 & n1820;
  assign n5867 = ~n5865 & ~n5866;
  assign n5868 = n5864 & n5867;
  assign n5860 = ~n987 & ~n991;
  assign n5853 = ~x31 & n1211;
  assign n5854 = ~x30 & n1213;
  assign n5855 = ~n5853 & ~n5854;
  assign n5856 = x31 & n1204;
  assign n5857 = x30 & n1208;
  assign n5858 = ~n5856 & ~n5857;
  assign n5859 = n5855 & n5858;
  assign n5861 = n5860 ^ n5859;
  assign n5869 = n5868 ^ n5861;
  assign n5893 = n5892 ^ n5869;
  assign n5911 = n5910 ^ n5893;
  assign n5850 = n5810 ^ n5790;
  assign n5851 = n5791 & ~n5850;
  assign n5852 = n5851 ^ n5810;
  assign n5912 = n5911 ^ n5852;
  assign n5847 = n5831 ^ n5819;
  assign n5848 = n5820 & n5847;
  assign n5849 = n5848 ^ n5831;
  assign n5913 = n5912 ^ n5849;
  assign n5930 = n5929 ^ n5913;
  assign n5844 = n5750 ^ n5747;
  assign n5845 = ~n5812 & n5844;
  assign n5846 = n5845 ^ n5811;
  assign n5931 = n5930 ^ n5846;
  assign n5841 = n5813 ^ n5744;
  assign n5842 = n5833 & ~n5841;
  assign n5843 = n5842 ^ n5832;
  assign n5932 = n5931 ^ n5843;
  assign n5937 = n5936 ^ n5932;
  assign n6026 = n5843 & ~n5931;
  assign n6027 = ~n5843 & n5931;
  assign n6028 = ~n5936 & ~n6027;
  assign n6029 = ~n6026 & ~n6028;
  assign n6012 = ~x22 & n2770;
  assign n6013 = ~x21 & n2774;
  assign n6014 = ~n6012 & ~n6013;
  assign n6015 = x22 & n2777;
  assign n6016 = x21 & n2779;
  assign n6017 = ~n6015 & ~n6016;
  assign n6018 = n6014 & n6017;
  assign n6004 = ~x24 & n2359;
  assign n6005 = ~x23 & n2361;
  assign n6006 = ~n6004 & ~n6005;
  assign n6007 = x24 & n2352;
  assign n6008 = x23 & n2356;
  assign n6009 = ~n6007 & ~n6008;
  assign n6010 = n6006 & n6009;
  assign n5997 = x28 & n1818;
  assign n5998 = x27 & n1820;
  assign n5999 = ~n5997 & ~n5998;
  assign n6000 = ~x28 & n1811;
  assign n6001 = ~x27 & n1815;
  assign n6002 = ~n6000 & ~n6001;
  assign n6003 = n5999 & n6002;
  assign n6011 = n6010 ^ n6003;
  assign n6019 = n6018 ^ n6011;
  assign n5992 = n5909 ^ n5901;
  assign n5993 = n5909 ^ n5900;
  assign n5994 = ~n5992 & ~n5993;
  assign n5995 = n5994 ^ n5901;
  assign n5989 = n5891 ^ n5876;
  assign n5990 = n5884 & ~n5989;
  assign n5991 = n5990 ^ n5883;
  assign n5996 = n5995 ^ n5991;
  assign n6020 = n6019 ^ n5996;
  assign n5986 = n5910 ^ n5869;
  assign n5987 = ~n5893 & ~n5986;
  assign n5988 = n5987 ^ n5892;
  assign n6021 = n6020 ^ n5988;
  assign n5976 = x26 & n2142;
  assign n5977 = x25 & n2144;
  assign n5978 = ~n5976 & ~n5977;
  assign n5979 = ~x26 & n2135;
  assign n5980 = ~x25 & n2139;
  assign n5981 = ~n5979 & ~n5980;
  assign n5982 = n5978 & n5981;
  assign n5974 = x18 & x63;
  assign n5967 = ~x30 & n1549;
  assign n5968 = ~x29 & n1553;
  assign n5969 = ~n5967 & ~n5968;
  assign n5970 = x30 & n1556;
  assign n5971 = x29 & n1558;
  assign n5972 = ~n5970 & ~n5971;
  assign n5973 = n5969 & n5972;
  assign n5975 = n5974 ^ n5973;
  assign n5983 = n5982 ^ n5975;
  assign n5962 = x51 ^ x31;
  assign n5963 = n1207 & n5962;
  assign n5964 = ~n1211 & ~n5963;
  assign n5955 = x20 & n3105;
  assign n5956 = x19 & n3107;
  assign n5957 = ~n5955 & ~n5956;
  assign n5958 = ~x20 & n3098;
  assign n5959 = ~x19 & n3102;
  assign n5960 = ~n5958 & ~n5959;
  assign n5961 = n5957 & n5960;
  assign n5965 = n5964 ^ n5961;
  assign n5951 = n5868 ^ n5860;
  assign n5952 = n5868 ^ n5859;
  assign n5953 = ~n5951 & ~n5952;
  assign n5954 = n5953 ^ n5860;
  assign n5966 = n5965 ^ n5954;
  assign n5984 = n5983 ^ n5966;
  assign n5948 = n5926 ^ n5923;
  assign n5949 = ~n5927 & n5948;
  assign n5950 = n5949 ^ n5809;
  assign n5985 = n5984 ^ n5950;
  assign n6022 = n6021 ^ n5985;
  assign n5944 = n5928 ^ n5919;
  assign n5945 = n5928 ^ n5916;
  assign n5946 = n5944 & ~n5945;
  assign n5947 = n5946 ^ n5919;
  assign n6023 = n6022 ^ n5947;
  assign n5941 = n5852 ^ n5849;
  assign n5942 = ~n5912 & n5941;
  assign n5943 = n5942 ^ n5911;
  assign n6024 = n6023 ^ n5943;
  assign n5938 = n5913 ^ n5846;
  assign n5939 = n5930 & n5938;
  assign n5940 = n5939 ^ n5929;
  assign n6025 = n6024 ^ n5940;
  assign n6030 = n6029 ^ n6025;
  assign n6111 = n5940 & n6024;
  assign n6112 = ~n5940 & ~n6024;
  assign n6113 = ~n6029 & ~n6112;
  assign n6114 = ~n6111 & ~n6113;
  assign n6097 = x23 & n2777;
  assign n6098 = x22 & n2779;
  assign n6099 = ~n6097 & ~n6098;
  assign n6100 = ~x23 & n2770;
  assign n6101 = ~x22 & n2774;
  assign n6102 = ~n6100 & ~n6101;
  assign n6103 = n6099 & n6102;
  assign n6090 = ~x21 & n3098;
  assign n6091 = ~x20 & n3102;
  assign n6092 = ~n6090 & ~n6091;
  assign n6093 = x21 & n3105;
  assign n6094 = x20 & n3107;
  assign n6095 = ~n6093 & ~n6094;
  assign n6096 = n6092 & n6095;
  assign n6104 = n6103 ^ n6096;
  assign n6105 = n6104 ^ n5964;
  assign n6082 = ~x29 & n1811;
  assign n6083 = ~x28 & n1815;
  assign n6084 = ~n6082 & ~n6083;
  assign n6085 = x29 & n1818;
  assign n6086 = x28 & n1820;
  assign n6087 = ~n6085 & ~n6086;
  assign n6088 = n6084 & n6087;
  assign n6080 = x19 & x63;
  assign n6073 = ~x25 & n2359;
  assign n6074 = ~x24 & n2361;
  assign n6075 = ~n6073 & ~n6074;
  assign n6076 = x25 & n2352;
  assign n6077 = x24 & n2356;
  assign n6078 = ~n6076 & ~n6077;
  assign n6079 = n6075 & n6078;
  assign n6081 = n6080 ^ n6079;
  assign n6089 = n6088 ^ n6081;
  assign n6106 = n6105 ^ n6089;
  assign n6070 = n5961 ^ n5954;
  assign n6071 = ~n5965 & n6070;
  assign n6072 = n6071 ^ n5964;
  assign n6107 = n6106 ^ n6072;
  assign n6059 = ~x27 & n2135;
  assign n6060 = ~x26 & n2139;
  assign n6061 = ~n6059 & ~n6060;
  assign n6062 = x27 & n2142;
  assign n6063 = x26 & n2144;
  assign n6064 = ~n6062 & ~n6063;
  assign n6065 = n6061 & n6064;
  assign n6057 = ~n1211 & ~n1213;
  assign n6050 = ~x31 & n1549;
  assign n6051 = ~x30 & n1553;
  assign n6052 = ~n6050 & ~n6051;
  assign n6053 = x31 & n1556;
  assign n6054 = x30 & n1558;
  assign n6055 = ~n6053 & ~n6054;
  assign n6056 = n6052 & n6055;
  assign n6058 = n6057 ^ n6056;
  assign n6066 = n6065 ^ n6058;
  assign n6046 = n5982 ^ n5973;
  assign n6047 = ~n5975 & ~n6046;
  assign n6048 = n6047 ^ n5974;
  assign n6043 = n6018 ^ n6010;
  assign n6044 = ~n6011 & n6043;
  assign n6045 = n6044 ^ n6018;
  assign n6049 = n6048 ^ n6045;
  assign n6067 = n6066 ^ n6049;
  assign n6040 = n6019 ^ n5995;
  assign n6041 = n5996 & ~n6040;
  assign n6042 = n6041 ^ n6019;
  assign n6068 = n6067 ^ n6042;
  assign n6037 = n5966 ^ n5950;
  assign n6038 = ~n5984 & ~n6037;
  assign n6039 = n6038 ^ n5983;
  assign n6069 = n6068 ^ n6039;
  assign n6108 = n6107 ^ n6069;
  assign n6034 = n5988 ^ n5985;
  assign n6035 = ~n6021 & n6034;
  assign n6036 = n6035 ^ n6020;
  assign n6109 = n6108 ^ n6036;
  assign n6031 = n5947 ^ n5943;
  assign n6032 = ~n6023 & n6031;
  assign n6033 = n6032 ^ n6022;
  assign n6110 = n6109 ^ n6033;
  assign n6115 = n6114 ^ n6110;
  assign n6190 = ~n6033 & ~n6109;
  assign n6191 = n6033 & n6109;
  assign n6192 = ~n6114 & ~n6191;
  assign n6193 = ~n6190 & ~n6192;
  assign n6182 = x20 & x63;
  assign n6174 = ~x28 & n2135;
  assign n6175 = ~x27 & n2139;
  assign n6176 = ~n6174 & ~n6175;
  assign n6177 = x28 & n2142;
  assign n6178 = x27 & n2144;
  assign n6179 = ~n6177 & ~n6178;
  assign n6180 = n6176 & n6179;
  assign n6167 = ~x22 & n3098;
  assign n6168 = ~x21 & n3102;
  assign n6169 = ~n6167 & ~n6168;
  assign n6170 = x22 & n3105;
  assign n6171 = x21 & n3107;
  assign n6172 = ~n6170 & ~n6171;
  assign n6173 = n6169 & n6172;
  assign n6181 = n6180 ^ n6173;
  assign n6183 = n6182 ^ n6181;
  assign n6159 = ~x24 & n2770;
  assign n6160 = ~x23 & n2774;
  assign n6161 = ~n6159 & ~n6160;
  assign n6162 = x24 & n2777;
  assign n6163 = x23 & n2779;
  assign n6164 = ~n6162 & ~n6163;
  assign n6165 = n6161 & n6164;
  assign n6151 = ~x30 & n1811;
  assign n6152 = ~x29 & n1815;
  assign n6153 = ~n6151 & ~n6152;
  assign n6154 = x30 & n1818;
  assign n6155 = x29 & n1820;
  assign n6156 = ~n6154 & ~n6155;
  assign n6157 = n6153 & n6156;
  assign n6144 = x26 & n2352;
  assign n6145 = x25 & n2356;
  assign n6146 = ~n6144 & ~n6145;
  assign n6147 = ~x26 & n2359;
  assign n6148 = ~x25 & n2361;
  assign n6149 = ~n6147 & ~n6148;
  assign n6150 = n6146 & n6149;
  assign n6158 = n6157 ^ n6150;
  assign n6166 = n6165 ^ n6158;
  assign n6184 = n6183 ^ n6166;
  assign n6141 = n6103 ^ n5964;
  assign n6142 = ~n6104 & n6141;
  assign n6143 = n6142 ^ n5964;
  assign n6185 = n6184 ^ n6143;
  assign n6135 = x53 ^ x31;
  assign n6136 = n1552 & n6135;
  assign n6137 = ~n1549 & ~n6136;
  assign n6132 = n6065 ^ n6056;
  assign n6133 = ~n6058 & ~n6132;
  assign n6134 = n6133 ^ n6057;
  assign n6138 = n6137 ^ n6134;
  assign n6129 = n6088 ^ n6079;
  assign n6130 = ~n6081 & ~n6129;
  assign n6131 = n6130 ^ n6080;
  assign n6139 = n6138 ^ n6131;
  assign n6126 = n6066 ^ n6048;
  assign n6127 = n6049 & n6126;
  assign n6128 = n6127 ^ n6066;
  assign n6140 = n6139 ^ n6128;
  assign n6186 = n6185 ^ n6140;
  assign n6123 = n6089 ^ n6072;
  assign n6124 = ~n6106 & ~n6123;
  assign n6125 = n6124 ^ n6105;
  assign n6187 = n6186 ^ n6125;
  assign n6120 = n6042 ^ n6039;
  assign n6121 = n6068 & n6120;
  assign n6122 = n6121 ^ n6067;
  assign n6188 = n6187 ^ n6122;
  assign n6116 = n6107 ^ n6036;
  assign n6117 = n6069 ^ n6036;
  assign n6118 = ~n6116 & ~n6117;
  assign n6119 = n6118 ^ n6107;
  assign n6189 = n6188 ^ n6119;
  assign n6194 = n6193 ^ n6189;
  assign n6264 = ~n6119 & n6188;
  assign n6265 = n6119 & ~n6188;
  assign n6266 = ~n6193 & ~n6265;
  assign n6267 = ~n6264 & ~n6266;
  assign n6252 = ~x27 & n2359;
  assign n6253 = ~x26 & n2361;
  assign n6254 = ~n6252 & ~n6253;
  assign n6255 = x27 & n2352;
  assign n6256 = x26 & n2356;
  assign n6257 = ~n6255 & ~n6256;
  assign n6258 = n6254 & n6257;
  assign n6250 = ~n1549 & ~n1553;
  assign n6243 = x31 & n1818;
  assign n6244 = x30 & n1820;
  assign n6245 = ~n6243 & ~n6244;
  assign n6246 = ~x31 & n1811;
  assign n6247 = ~x30 & n1815;
  assign n6248 = ~n6246 & ~n6247;
  assign n6249 = n6245 & n6248;
  assign n6251 = n6250 ^ n6249;
  assign n6259 = n6258 ^ n6251;
  assign n6234 = x23 & n3105;
  assign n6235 = x22 & n3107;
  assign n6236 = ~n6234 & ~n6235;
  assign n6237 = ~x23 & n3098;
  assign n6238 = ~x22 & n3102;
  assign n6239 = ~n6237 & ~n6238;
  assign n6240 = n6236 & n6239;
  assign n6226 = ~x25 & n2770;
  assign n6227 = ~x24 & n2774;
  assign n6228 = ~n6226 & ~n6227;
  assign n6229 = x25 & n2777;
  assign n6230 = x24 & n2779;
  assign n6231 = ~n6229 & ~n6230;
  assign n6232 = n6228 & n6231;
  assign n6219 = x29 & n2142;
  assign n6220 = x28 & n2144;
  assign n6221 = ~n6219 & ~n6220;
  assign n6222 = ~x29 & n2135;
  assign n6223 = ~x28 & n2139;
  assign n6224 = ~n6222 & ~n6223;
  assign n6225 = n6221 & n6224;
  assign n6233 = n6232 ^ n6225;
  assign n6241 = n6240 ^ n6233;
  assign n6216 = n6182 ^ n6180;
  assign n6217 = ~n6181 & ~n6216;
  assign n6218 = n6217 ^ n6182;
  assign n6242 = n6241 ^ n6218;
  assign n6260 = n6259 ^ n6242;
  assign n6211 = x21 & x63;
  assign n6212 = n6211 ^ n6137;
  assign n6208 = n6165 ^ n6150;
  assign n6209 = n6158 & ~n6208;
  assign n6210 = n6209 ^ n6157;
  assign n6213 = n6212 ^ n6210;
  assign n6204 = n6137 ^ n6131;
  assign n6205 = n6134 ^ n6131;
  assign n6206 = n6204 & ~n6205;
  assign n6207 = n6206 ^ n6137;
  assign n6214 = n6213 ^ n6207;
  assign n6201 = n6166 ^ n6143;
  assign n6202 = ~n6184 & ~n6201;
  assign n6203 = n6202 ^ n6183;
  assign n6215 = n6214 ^ n6203;
  assign n6261 = n6260 ^ n6215;
  assign n6198 = n6185 ^ n6139;
  assign n6199 = ~n6140 & n6198;
  assign n6200 = n6199 ^ n6185;
  assign n6262 = n6261 ^ n6200;
  assign n6195 = n6125 ^ n6122;
  assign n6196 = ~n6187 & ~n6195;
  assign n6197 = n6196 ^ n6186;
  assign n6263 = n6262 ^ n6197;
  assign n6268 = n6267 ^ n6263;
  assign n6333 = n6197 & ~n6262;
  assign n6334 = ~n6197 & n6262;
  assign n6335 = ~n6267 & ~n6334;
  assign n6336 = ~n6333 & ~n6335;
  assign n6325 = x55 ^ x31;
  assign n6326 = n1814 & n6325;
  assign n6327 = ~n1811 & ~n6326;
  assign n6317 = x24 & n3105;
  assign n6318 = x23 & n3107;
  assign n6319 = ~n6317 & ~n6318;
  assign n6320 = ~x24 & n3098;
  assign n6321 = ~x23 & n3102;
  assign n6322 = ~n6320 & ~n6321;
  assign n6323 = n6319 & n6322;
  assign n6310 = ~x26 & n2770;
  assign n6311 = ~x25 & n2774;
  assign n6312 = ~n6310 & ~n6311;
  assign n6313 = x26 & n2777;
  assign n6314 = x25 & n2779;
  assign n6315 = ~n6313 & ~n6314;
  assign n6316 = n6312 & n6315;
  assign n6324 = n6323 ^ n6316;
  assign n6328 = n6327 ^ n6324;
  assign n6306 = n6258 ^ n6249;
  assign n6307 = ~n6251 & ~n6306;
  assign n6308 = n6307 ^ n6250;
  assign n6302 = n6240 ^ n6232;
  assign n6303 = n6240 ^ n6225;
  assign n6304 = n6302 & ~n6303;
  assign n6305 = n6304 ^ n6232;
  assign n6309 = n6308 ^ n6305;
  assign n6329 = n6328 ^ n6309;
  assign n6292 = x30 & n2142;
  assign n6293 = x29 & n2144;
  assign n6294 = ~n6292 & ~n6293;
  assign n6295 = ~x30 & n2135;
  assign n6296 = ~x29 & n2139;
  assign n6297 = ~n6295 & ~n6296;
  assign n6298 = n6294 & n6297;
  assign n6290 = x22 & x63;
  assign n6283 = ~x28 & n2359;
  assign n6284 = ~x27 & n2361;
  assign n6285 = ~n6283 & ~n6284;
  assign n6286 = x28 & n2352;
  assign n6287 = x27 & n2356;
  assign n6288 = ~n6286 & ~n6287;
  assign n6289 = n6285 & n6288;
  assign n6291 = n6290 ^ n6289;
  assign n6299 = n6298 ^ n6291;
  assign n6280 = n6210 ^ n6137;
  assign n6281 = ~n6212 & ~n6280;
  assign n6282 = n6281 ^ n6211;
  assign n6300 = n6299 ^ n6282;
  assign n6276 = n6259 ^ n6241;
  assign n6277 = n6259 ^ n6218;
  assign n6278 = ~n6276 & ~n6277;
  assign n6279 = n6278 ^ n6241;
  assign n6301 = n6300 ^ n6279;
  assign n6330 = n6329 ^ n6301;
  assign n6272 = n6213 ^ n6203;
  assign n6273 = n6207 ^ n6203;
  assign n6274 = n6272 & ~n6273;
  assign n6275 = n6274 ^ n6213;
  assign n6331 = n6330 ^ n6275;
  assign n6269 = n6215 ^ n6200;
  assign n6270 = ~n6261 & ~n6269;
  assign n6271 = n6270 ^ n6260;
  assign n6332 = n6331 ^ n6271;
  assign n6337 = n6336 ^ n6332;
  assign n6395 = ~n6271 & n6331;
  assign n6396 = n6271 & ~n6331;
  assign n6397 = ~n6336 & ~n6396;
  assign n6398 = ~n6395 & ~n6397;
  assign n6388 = x23 & x63;
  assign n6380 = x29 & n2352;
  assign n6381 = x28 & n2356;
  assign n6382 = ~n6380 & ~n6381;
  assign n6383 = ~x29 & n2359;
  assign n6384 = ~x28 & n2361;
  assign n6385 = ~n6383 & ~n6384;
  assign n6386 = n6382 & n6385;
  assign n6373 = ~x25 & n3098;
  assign n6374 = ~x24 & n3102;
  assign n6375 = ~n6373 & ~n6374;
  assign n6376 = x25 & n3105;
  assign n6377 = x24 & n3107;
  assign n6378 = ~n6376 & ~n6377;
  assign n6379 = n6375 & n6378;
  assign n6387 = n6386 ^ n6379;
  assign n6389 = n6388 ^ n6387;
  assign n6369 = n6327 ^ n6323;
  assign n6370 = ~n6324 & n6369;
  assign n6371 = n6370 ^ n6327;
  assign n6372 = n6371 ^ n6298;
  assign n6390 = n6389 ^ n6372;
  assign n6360 = ~x27 & n2770;
  assign n6361 = ~x26 & n2774;
  assign n6362 = ~n6360 & ~n6361;
  assign n6363 = x27 & n2777;
  assign n6364 = x26 & n2779;
  assign n6365 = ~n6363 & ~n6364;
  assign n6366 = n6362 & n6365;
  assign n6358 = ~n1811 & ~n1815;
  assign n6351 = ~x31 & n2135;
  assign n6352 = ~x30 & n2139;
  assign n6353 = ~n6351 & ~n6352;
  assign n6354 = x31 & n2142;
  assign n6355 = x30 & n2144;
  assign n6356 = ~n6354 & ~n6355;
  assign n6357 = n6353 & n6356;
  assign n6359 = n6358 ^ n6357;
  assign n6367 = n6366 ^ n6359;
  assign n6347 = n6298 ^ n6290;
  assign n6348 = n6298 ^ n6289;
  assign n6349 = n6347 & n6348;
  assign n6350 = n6349 ^ n6290;
  assign n6368 = n6367 ^ n6350;
  assign n6391 = n6390 ^ n6368;
  assign n6344 = n6328 ^ n6308;
  assign n6345 = n6309 & ~n6344;
  assign n6346 = n6345 ^ n6328;
  assign n6392 = n6391 ^ n6346;
  assign n6341 = n6282 ^ n6279;
  assign n6342 = ~n6300 & n6341;
  assign n6343 = n6342 ^ n6299;
  assign n6393 = n6392 ^ n6343;
  assign n6338 = n6301 ^ n6275;
  assign n6339 = n6330 & ~n6338;
  assign n6340 = n6339 ^ n6329;
  assign n6394 = n6393 ^ n6340;
  assign n6399 = n6398 ^ n6394;
  assign n6450 = n6340 & n6393;
  assign n6451 = ~n6340 & ~n6393;
  assign n6452 = ~n6398 & ~n6451;
  assign n6453 = ~n6450 & ~n6452;
  assign n6437 = ~x30 & n2359;
  assign n6438 = ~x29 & n2361;
  assign n6439 = ~n6437 & ~n6438;
  assign n6440 = x30 & n2352;
  assign n6441 = x29 & n2356;
  assign n6442 = ~n6440 & ~n6441;
  assign n6443 = n6439 & n6442;
  assign n6430 = ~x28 & n2770;
  assign n6431 = ~x27 & n2774;
  assign n6432 = ~n6430 & ~n6431;
  assign n6433 = x28 & n2777;
  assign n6434 = x27 & n2779;
  assign n6435 = ~n6433 & ~n6434;
  assign n6436 = n6432 & n6435;
  assign n6444 = n6443 ^ n6436;
  assign n6427 = n6388 ^ n6386;
  assign n6428 = ~n6387 & ~n6427;
  assign n6429 = n6428 ^ n6388;
  assign n6445 = n6444 ^ n6429;
  assign n6422 = x57 ^ x31;
  assign n6423 = n2138 & n6422;
  assign n6424 = ~n2135 & ~n6423;
  assign n6420 = x24 & x63;
  assign n6413 = x26 & n3105;
  assign n6414 = x25 & n3107;
  assign n6415 = ~n6413 & ~n6414;
  assign n6416 = ~x26 & n3098;
  assign n6417 = ~x25 & n3102;
  assign n6418 = ~n6416 & ~n6417;
  assign n6419 = n6415 & n6418;
  assign n6421 = n6420 ^ n6419;
  assign n6425 = n6424 ^ n6421;
  assign n6410 = n6366 ^ n6357;
  assign n6411 = ~n6359 & ~n6410;
  assign n6412 = n6411 ^ n6358;
  assign n6426 = n6425 ^ n6412;
  assign n6446 = n6445 ^ n6426;
  assign n6406 = n6389 ^ n6298;
  assign n6407 = n6389 ^ n6371;
  assign n6408 = ~n6406 & n6407;
  assign n6409 = n6408 ^ n6298;
  assign n6447 = n6446 ^ n6409;
  assign n6403 = n6390 ^ n6350;
  assign n6404 = n6368 & ~n6403;
  assign n6405 = n6404 ^ n6367;
  assign n6448 = n6447 ^ n6405;
  assign n6400 = n6346 ^ n6343;
  assign n6401 = ~n6392 & ~n6400;
  assign n6402 = n6401 ^ n6391;
  assign n6449 = n6448 ^ n6402;
  assign n6454 = n6453 ^ n6449;
  assign n6500 = n6402 & n6448;
  assign n6501 = ~n6402 & ~n6448;
  assign n6502 = ~n6453 & ~n6501;
  assign n6503 = ~n6500 & ~n6502;
  assign n6493 = x25 & x63;
  assign n6486 = ~x29 & n2770;
  assign n6487 = ~x28 & n2774;
  assign n6488 = ~n6486 & ~n6487;
  assign n6489 = x29 & n2777;
  assign n6490 = x28 & n2779;
  assign n6491 = ~n6489 & ~n6490;
  assign n6492 = n6488 & n6491;
  assign n6494 = n6493 ^ n6492;
  assign n6495 = n6494 ^ n6443;
  assign n6477 = x27 & n3105;
  assign n6478 = x26 & n3107;
  assign n6479 = ~n6477 & ~n6478;
  assign n6480 = ~x27 & n3098;
  assign n6481 = ~x26 & n3102;
  assign n6482 = ~n6480 & ~n6481;
  assign n6483 = n6479 & n6482;
  assign n6475 = ~n2135 & ~n2139;
  assign n6468 = ~x31 & n2359;
  assign n6469 = ~x30 & n2361;
  assign n6470 = ~n6468 & ~n6469;
  assign n6471 = x31 & n2352;
  assign n6472 = x30 & n2356;
  assign n6473 = ~n6471 & ~n6472;
  assign n6474 = n6470 & n6473;
  assign n6476 = n6475 ^ n6474;
  assign n6484 = n6483 ^ n6476;
  assign n6464 = n6424 ^ n6420;
  assign n6465 = n6424 ^ n6419;
  assign n6466 = ~n6464 & ~n6465;
  assign n6467 = n6466 ^ n6420;
  assign n6485 = n6484 ^ n6467;
  assign n6496 = n6495 ^ n6485;
  assign n6461 = n6436 ^ n6429;
  assign n6462 = ~n6444 & n6461;
  assign n6463 = n6462 ^ n6443;
  assign n6497 = n6496 ^ n6463;
  assign n6458 = n6445 ^ n6412;
  assign n6459 = n6426 & n6458;
  assign n6460 = n6459 ^ n6425;
  assign n6498 = n6497 ^ n6460;
  assign n6455 = n6409 ^ n6405;
  assign n6456 = n6447 & n6455;
  assign n6457 = n6456 ^ n6446;
  assign n6499 = n6498 ^ n6457;
  assign n6504 = n6503 ^ n6499;
  assign n6544 = ~n6457 & n6498;
  assign n6545 = n6457 & ~n6498;
  assign n6546 = ~n6503 & ~n6545;
  assign n6547 = ~n6544 & ~n6546;
  assign n6532 = x28 & n3105;
  assign n6533 = x27 & n3107;
  assign n6534 = ~n6532 & ~n6533;
  assign n6535 = ~x28 & n3098;
  assign n6536 = ~x27 & n3102;
  assign n6537 = ~n6535 & ~n6536;
  assign n6538 = n6534 & n6537;
  assign n6530 = x26 & x63;
  assign n6523 = ~x30 & n2770;
  assign n6524 = ~x29 & n2774;
  assign n6525 = ~n6523 & ~n6524;
  assign n6526 = x30 & n2777;
  assign n6527 = x29 & n2779;
  assign n6528 = ~n6526 & ~n6527;
  assign n6529 = n6525 & n6528;
  assign n6531 = n6530 ^ n6529;
  assign n6539 = n6538 ^ n6531;
  assign n6519 = x59 ^ x31;
  assign n6520 = n2355 & n6519;
  assign n6521 = ~n2359 & ~n6520;
  assign n6515 = n6483 ^ n6475;
  assign n6516 = n6483 ^ n6474;
  assign n6517 = ~n6515 & ~n6516;
  assign n6518 = n6517 ^ n6475;
  assign n6522 = n6521 ^ n6518;
  assign n6540 = n6539 ^ n6522;
  assign n6511 = n6493 ^ n6443;
  assign n6512 = n6492 ^ n6443;
  assign n6513 = ~n6511 & ~n6512;
  assign n6514 = n6513 ^ n6493;
  assign n6541 = n6540 ^ n6514;
  assign n6508 = n6495 ^ n6484;
  assign n6509 = ~n6485 & n6508;
  assign n6510 = n6509 ^ n6495;
  assign n6542 = n6541 ^ n6510;
  assign n6505 = n6463 ^ n6460;
  assign n6506 = n6497 & ~n6505;
  assign n6507 = n6506 ^ n6496;
  assign n6543 = n6542 ^ n6507;
  assign n6548 = n6547 ^ n6543;
  assign n6582 = n6507 & n6542;
  assign n6583 = ~n6507 & ~n6542;
  assign n6584 = ~n6547 & ~n6583;
  assign n6585 = ~n6582 & ~n6584;
  assign n6577 = x27 & x63;
  assign n6575 = ~n2359 & ~n2361;
  assign n6568 = x31 & n2777;
  assign n6569 = x30 & n2779;
  assign n6570 = ~n6568 & ~n6569;
  assign n6571 = ~x31 & n2770;
  assign n6572 = ~x30 & n2774;
  assign n6573 = ~n6571 & ~n6572;
  assign n6574 = n6570 & n6573;
  assign n6576 = n6575 ^ n6574;
  assign n6578 = n6577 ^ n6576;
  assign n6559 = ~x29 & n3098;
  assign n6560 = ~x28 & n3102;
  assign n6561 = ~n6559 & ~n6560;
  assign n6562 = x29 & n3105;
  assign n6563 = x28 & n3107;
  assign n6564 = ~n6562 & ~n6563;
  assign n6565 = n6561 & n6564;
  assign n6566 = n6565 ^ n6521;
  assign n6556 = n6538 ^ n6529;
  assign n6557 = ~n6531 & ~n6556;
  assign n6558 = n6557 ^ n6530;
  assign n6567 = n6566 ^ n6558;
  assign n6579 = n6578 ^ n6567;
  assign n6552 = n6539 ^ n6521;
  assign n6553 = n6539 ^ n6518;
  assign n6554 = n6552 & ~n6553;
  assign n6555 = n6554 ^ n6521;
  assign n6580 = n6579 ^ n6555;
  assign n6549 = n6540 ^ n6510;
  assign n6550 = n6541 & ~n6549;
  assign n6551 = n6550 ^ n6514;
  assign n6581 = n6580 ^ n6551;
  assign n6586 = n6585 ^ n6581;
  assign n6612 = n6551 & ~n6580;
  assign n6613 = ~n6551 & n6580;
  assign n6614 = ~n6585 & ~n6613;
  assign n6615 = ~n6612 & ~n6614;
  assign n6605 = x61 ^ x31;
  assign n6606 = n2773 & n6605;
  assign n6607 = ~n2770 & ~n6606;
  assign n6603 = x28 & x63;
  assign n6596 = ~x30 & n3098;
  assign n6597 = ~x29 & n3102;
  assign n6598 = ~n6596 & ~n6597;
  assign n6599 = x30 & n3105;
  assign n6600 = x29 & n3107;
  assign n6601 = ~n6599 & ~n6600;
  assign n6602 = n6598 & n6601;
  assign n6604 = n6603 ^ n6602;
  assign n6608 = n6607 ^ n6604;
  assign n6593 = n6577 ^ n6575;
  assign n6594 = n6576 & n6593;
  assign n6595 = n6594 ^ n6577;
  assign n6609 = n6608 ^ n6595;
  assign n6590 = n6565 ^ n6558;
  assign n6591 = n6566 & n6590;
  assign n6592 = n6591 ^ n6521;
  assign n6610 = n6609 ^ n6592;
  assign n6587 = n6567 ^ n6555;
  assign n6588 = ~n6579 & ~n6587;
  assign n6589 = n6588 ^ n6578;
  assign n6611 = n6610 ^ n6589;
  assign n6616 = n6615 ^ n6611;
  assign n6638 = ~n6589 & n6610;
  assign n6639 = n6589 & ~n6610;
  assign n6640 = ~n6615 & ~n6639;
  assign n6641 = ~n6638 & ~n6640;
  assign n6633 = x29 & x63;
  assign n6631 = ~n2770 & ~n2774;
  assign n6624 = x31 & n3105;
  assign n6625 = x30 & n3107;
  assign n6626 = ~n6624 & ~n6625;
  assign n6627 = ~x31 & n3098;
  assign n6628 = ~x30 & n3102;
  assign n6629 = ~n6627 & ~n6628;
  assign n6630 = n6626 & n6629;
  assign n6632 = n6631 ^ n6630;
  assign n6634 = n6633 ^ n6632;
  assign n6635 = n6634 ^ n6607;
  assign n6620 = n6607 ^ n6603;
  assign n6621 = n6607 ^ n6602;
  assign n6622 = n6620 & n6621;
  assign n6623 = n6622 ^ n6603;
  assign n6636 = n6635 ^ n6623;
  assign n6617 = n6595 ^ n6592;
  assign n6618 = ~n6609 & n6617;
  assign n6619 = n6618 ^ n6608;
  assign n6637 = n6636 ^ n6619;
  assign n6642 = n6641 ^ n6637;
  assign n6656 = ~n6619 & n6636;
  assign n6657 = n6619 & ~n6636;
  assign n6658 = ~n6641 & ~n6657;
  assign n6659 = ~n6656 & ~n6658;
  assign n6652 = x30 & x63;
  assign n6649 = x63 ^ x31;
  assign n6650 = n3101 & n6649;
  assign n6651 = ~n3098 & ~n6650;
  assign n6653 = n6652 ^ n6651;
  assign n6646 = n6633 ^ n6631;
  assign n6647 = n6632 & n6646;
  assign n6648 = n6647 ^ n6633;
  assign n6654 = n6653 ^ n6648;
  assign n6643 = n6634 ^ n6623;
  assign n6644 = n6635 & n6643;
  assign n6645 = n6644 ^ n6607;
  assign n6655 = n6654 ^ n6645;
  assign n6660 = n6659 ^ n6655;
  assign n6668 = ~n3003 & ~n3101;
  assign n6669 = n6668 ^ x31;
  assign n6670 = x63 & ~n6669;
  assign n6671 = n6670 ^ n6652;
  assign n6665 = n6651 ^ n6648;
  assign n6666 = n6653 & n6665;
  assign n6667 = n6666 ^ n6652;
  assign n6672 = n6671 ^ n6667;
  assign n6661 = ~n6645 & n6654;
  assign n6662 = n6645 & ~n6654;
  assign n6663 = ~n6659 & ~n6662;
  assign n6664 = ~n6661 & ~n6663;
  assign n6673 = n6672 ^ n6664;
  assign y0 = n65;
  assign y1 = ~n75;
  assign y2 = ~n85;
  assign y3 = ~n114;
  assign y4 = ~n137;
  assign y5 = n179;
  assign y6 = ~n214;
  assign y7 = n267;
  assign y8 = ~n316;
  assign y9 = ~n382;
  assign y10 = ~n442;
  assign y11 = ~n520;
  assign y12 = ~n591;
  assign y13 = n681;
  assign y14 = n764;
  assign y15 = n866;
  assign y16 = n964;
  assign y17 = n1078;
  assign y18 = ~n1186;
  assign y19 = ~n1312;
  assign y20 = n1435;
  assign y21 = n1574;
  assign y22 = ~n1707;
  assign y23 = ~n1858;
  assign y24 = n2002;
  assign y25 = ~n2167;
  assign y26 = n2326;
  assign y27 = ~n2502;
  assign y28 = ~n2672;
  assign y29 = ~n2860;
  assign y30 = ~n3041;
  assign y31 = n3241;
  assign y32 = n3429;
  assign y33 = ~n3620;
  assign y34 = n3807;
  assign y35 = n3992;
  assign y36 = n4173;
  assign y37 = ~n4348;
  assign y38 = n4512;
  assign y39 = n4672;
  assign y40 = n4825;
  assign y41 = ~n4976;
  assign y42 = ~n5116;
  assign y43 = n5255;
  assign y44 = n5382;
  assign y45 = n5508;
  assign y46 = ~n5625;
  assign y47 = ~n5737;
  assign y48 = n5840;
  assign y49 = n5937;
  assign y50 = ~n6030;
  assign y51 = ~n6115;
  assign y52 = n6194;
  assign y53 = n6268;
  assign y54 = n6337;
  assign y55 = ~n6399;
  assign y56 = ~n6454;
  assign y57 = n6504;
  assign y58 = ~n6548;
  assign y59 = n6586;
  assign y60 = n6616;
  assign y61 = n6642;
  assign y62 = n6660;
  assign y63 = ~n6673;
endmodule
